module top (\CM_rd0[0]_pad , \CM_rd0[10]_pad , \CM_rd0[11]_pad , \CM_rd0[12]_pad , \CM_rd0[13]_pad , \CM_rd0[14]_pad , \CM_rd0[15]_pad , \CM_rd0[16]_pad , \CM_rd0[17]_pad , \CM_rd0[18]_pad , \CM_rd0[19]_pad , \CM_rd0[1]_pad , \CM_rd0[20]_pad , \CM_rd0[21]_pad , \CM_rd0[22]_pad , \CM_rd0[23]_pad , \CM_rd0[2]_pad , \CM_rd0[3]_pad , \CM_rd0[4]_pad , \CM_rd0[5]_pad , \CM_rd0[6]_pad , \CM_rd0[7]_pad , \CM_rd0[8]_pad , \CM_rd0[9]_pad , \CM_rd1[0]_pad , \CM_rd1[10]_pad , \CM_rd1[11]_pad , \CM_rd1[12]_pad , \CM_rd1[13]_pad , \CM_rd1[14]_pad , \CM_rd1[15]_pad , \CM_rd1[16]_pad , \CM_rd1[17]_pad , \CM_rd1[18]_pad , \CM_rd1[19]_pad , \CM_rd1[1]_pad , \CM_rd1[20]_pad , \CM_rd1[21]_pad , \CM_rd1[22]_pad , \CM_rd1[23]_pad , \CM_rd1[2]_pad , \CM_rd1[3]_pad , \CM_rd1[4]_pad , \CM_rd1[5]_pad , \CM_rd1[6]_pad , \CM_rd1[7]_pad , \CM_rd1[8]_pad , \CM_rd1[9]_pad , \CM_rd2[0]_pad , \CM_rd2[10]_pad , \CM_rd2[11]_pad , \CM_rd2[12]_pad , \CM_rd2[13]_pad , \CM_rd2[14]_pad , \CM_rd2[15]_pad , \CM_rd2[16]_pad , \CM_rd2[17]_pad , \CM_rd2[18]_pad , \CM_rd2[19]_pad , \CM_rd2[1]_pad , \CM_rd2[20]_pad , \CM_rd2[21]_pad , \CM_rd2[22]_pad , \CM_rd2[23]_pad , \CM_rd2[2]_pad , \CM_rd2[3]_pad , \CM_rd2[4]_pad , \CM_rd2[5]_pad , \CM_rd2[6]_pad , \CM_rd2[7]_pad , \CM_rd2[8]_pad , \CM_rd2[9]_pad , \CM_rd3[0]_pad , \CM_rd3[10]_pad , \CM_rd3[11]_pad , \CM_rd3[12]_pad , \CM_rd3[13]_pad , \CM_rd3[14]_pad , \CM_rd3[15]_pad , \CM_rd3[16]_pad , \CM_rd3[17]_pad , \CM_rd3[18]_pad , \CM_rd3[19]_pad , \CM_rd3[1]_pad , \CM_rd3[20]_pad , \CM_rd3[21]_pad , \CM_rd3[22]_pad , \CM_rd3[23]_pad , \CM_rd3[2]_pad , \CM_rd3[3]_pad , \CM_rd3[4]_pad , \CM_rd3[5]_pad , \CM_rd3[6]_pad , \CM_rd3[7]_pad , \CM_rd3[8]_pad , \CM_rd3[9]_pad , \CM_rd4[0]_pad , \CM_rd4[10]_pad , \CM_rd4[11]_pad , \CM_rd4[12]_pad , \CM_rd4[13]_pad , \CM_rd4[14]_pad , \CM_rd4[15]_pad , \CM_rd4[16]_pad , \CM_rd4[17]_pad , \CM_rd4[18]_pad , \CM_rd4[19]_pad , \CM_rd4[1]_pad , \CM_rd4[20]_pad , \CM_rd4[21]_pad , \CM_rd4[22]_pad , \CM_rd4[23]_pad , \CM_rd4[2]_pad , \CM_rd4[3]_pad , \CM_rd4[4]_pad , \CM_rd4[5]_pad , \CM_rd4[6]_pad , \CM_rd4[7]_pad , \CM_rd4[8]_pad , \CM_rd4[9]_pad , \CM_rd5[0]_pad , \CM_rd5[10]_pad , \CM_rd5[11]_pad , \CM_rd5[12]_pad , \CM_rd5[13]_pad , \CM_rd5[14]_pad , \CM_rd5[15]_pad , \CM_rd5[16]_pad , \CM_rd5[17]_pad , \CM_rd5[18]_pad , \CM_rd5[19]_pad , \CM_rd5[1]_pad , \CM_rd5[20]_pad , \CM_rd5[21]_pad , \CM_rd5[22]_pad , \CM_rd5[23]_pad , \CM_rd5[2]_pad , \CM_rd5[3]_pad , \CM_rd5[4]_pad , \CM_rd5[5]_pad , \CM_rd5[6]_pad , \CM_rd5[7]_pad , \CM_rd5[8]_pad , \CM_rd5[9]_pad , \CM_rd6[0]_pad , \CM_rd6[10]_pad , \CM_rd6[11]_pad , \CM_rd6[12]_pad , \CM_rd6[13]_pad , \CM_rd6[14]_pad , \CM_rd6[15]_pad , \CM_rd6[16]_pad , \CM_rd6[17]_pad , \CM_rd6[18]_pad , \CM_rd6[19]_pad , \CM_rd6[1]_pad , \CM_rd6[20]_pad , \CM_rd6[21]_pad , \CM_rd6[22]_pad , \CM_rd6[23]_pad , \CM_rd6[2]_pad , \CM_rd6[3]_pad , \CM_rd6[4]_pad , \CM_rd6[5]_pad , \CM_rd6[6]_pad , \CM_rd6[7]_pad , \CM_rd6[8]_pad , \CM_rd6[9]_pad , \CM_rd7[0]_pad , \CM_rd7[10]_pad , \CM_rd7[11]_pad , \CM_rd7[12]_pad , \CM_rd7[13]_pad , \CM_rd7[14]_pad , \CM_rd7[15]_pad , \CM_rd7[16]_pad , \CM_rd7[17]_pad , \CM_rd7[18]_pad , \CM_rd7[19]_pad , \CM_rd7[1]_pad , \CM_rd7[20]_pad , \CM_rd7[21]_pad , \CM_rd7[22]_pad , \CM_rd7[23]_pad , \CM_rd7[2]_pad , \CM_rd7[3]_pad , \CM_rd7[4]_pad , \CM_rd7[5]_pad , \CM_rd7[6]_pad , \CM_rd7[7]_pad , \CM_rd7[8]_pad , \CM_rd7[9]_pad , \CM_rdm[0]_pad , \CM_rdm[10]_pad , \CM_rdm[11]_pad , \CM_rdm[12]_pad , \CM_rdm[13]_pad , \CM_rdm[14]_pad , \CM_rdm[15]_pad , \CM_rdm[16]_pad , \CM_rdm[17]_pad , \CM_rdm[18]_pad , \CM_rdm[19]_pad , \CM_rdm[1]_pad , \CM_rdm[20]_pad , \CM_rdm[21]_pad , \CM_rdm[22]_pad , \CM_rdm[23]_pad , \CM_rdm[2]_pad , \CM_rdm[3]_pad , \CM_rdm[4]_pad , \CM_rdm[5]_pad , \CM_rdm[6]_pad , \CM_rdm[7]_pad , \CM_rdm[8]_pad , \CM_rdm[9]_pad , \DM_rd0[0]_pad , \DM_rd0[10]_pad , \DM_rd0[11]_pad , \DM_rd0[12]_pad , \DM_rd0[13]_pad , \DM_rd0[14]_pad , \DM_rd0[15]_pad , \DM_rd0[1]_pad , \DM_rd0[2]_pad , \DM_rd0[3]_pad , \DM_rd0[4]_pad , \DM_rd0[5]_pad , \DM_rd0[6]_pad , \DM_rd0[7]_pad , \DM_rd0[8]_pad , \DM_rd0[9]_pad , \DM_rd1[0]_pad , \DM_rd1[10]_pad , \DM_rd1[11]_pad , \DM_rd1[12]_pad , \DM_rd1[13]_pad , \DM_rd1[14]_pad , \DM_rd1[15]_pad , \DM_rd1[1]_pad , \DM_rd1[2]_pad , \DM_rd1[3]_pad , \DM_rd1[4]_pad , \DM_rd1[5]_pad , \DM_rd1[6]_pad , \DM_rd1[7]_pad , \DM_rd1[8]_pad , \DM_rd1[9]_pad , \DM_rd2[0]_pad , \DM_rd2[10]_pad , \DM_rd2[11]_pad , \DM_rd2[12]_pad , \DM_rd2[13]_pad , \DM_rd2[14]_pad , \DM_rd2[15]_pad , \DM_rd2[1]_pad , \DM_rd2[2]_pad , \DM_rd2[3]_pad , \DM_rd2[4]_pad , \DM_rd2[5]_pad , \DM_rd2[6]_pad , \DM_rd2[7]_pad , \DM_rd2[8]_pad , \DM_rd2[9]_pad , \DM_rd3[0]_pad , \DM_rd3[10]_pad , \DM_rd3[11]_pad , \DM_rd3[12]_pad , \DM_rd3[13]_pad , \DM_rd3[14]_pad , \DM_rd3[15]_pad , \DM_rd3[1]_pad , \DM_rd3[2]_pad , \DM_rd3[3]_pad , \DM_rd3[4]_pad , \DM_rd3[5]_pad , \DM_rd3[6]_pad , \DM_rd3[7]_pad , \DM_rd3[8]_pad , \DM_rd3[9]_pad , \DM_rd4[0]_pad , \DM_rd4[10]_pad , \DM_rd4[11]_pad , \DM_rd4[12]_pad , \DM_rd4[13]_pad , \DM_rd4[14]_pad , \DM_rd4[15]_pad , \DM_rd4[1]_pad , \DM_rd4[2]_pad , \DM_rd4[3]_pad , \DM_rd4[4]_pad , \DM_rd4[5]_pad , \DM_rd4[6]_pad , \DM_rd4[7]_pad , \DM_rd4[8]_pad , \DM_rd4[9]_pad , \DM_rd5[0]_pad , \DM_rd5[10]_pad , \DM_rd5[11]_pad , \DM_rd5[12]_pad , \DM_rd5[13]_pad , \DM_rd5[14]_pad , \DM_rd5[15]_pad , \DM_rd5[1]_pad , \DM_rd5[2]_pad , \DM_rd5[3]_pad , \DM_rd5[4]_pad , \DM_rd5[5]_pad , \DM_rd5[6]_pad , \DM_rd5[7]_pad , \DM_rd5[8]_pad , \DM_rd5[9]_pad , \DM_rd6[0]_pad , \DM_rd6[10]_pad , \DM_rd6[11]_pad , \DM_rd6[12]_pad , \DM_rd6[13]_pad , \DM_rd6[14]_pad , \DM_rd6[15]_pad , \DM_rd6[1]_pad , \DM_rd6[2]_pad , \DM_rd6[3]_pad , \DM_rd6[4]_pad , \DM_rd6[5]_pad , \DM_rd6[6]_pad , \DM_rd6[7]_pad , \DM_rd6[8]_pad , \DM_rd6[9]_pad , \DM_rd7[0]_pad , \DM_rd7[10]_pad , \DM_rd7[11]_pad , \DM_rd7[12]_pad , \DM_rd7[13]_pad , \DM_rd7[14]_pad , \DM_rd7[15]_pad , \DM_rd7[1]_pad , \DM_rd7[2]_pad , \DM_rd7[3]_pad , \DM_rd7[4]_pad , \DM_rd7[5]_pad , \DM_rd7[6]_pad , \DM_rd7[7]_pad , \DM_rd7[8]_pad , \DM_rd7[9]_pad , \DM_rdm[0]_pad , \DM_rdm[10]_pad , \DM_rdm[11]_pad , \DM_rdm[12]_pad , \DM_rdm[13]_pad , \DM_rdm[14]_pad , \DM_rdm[15]_pad , \DM_rdm[1]_pad , \DM_rdm[2]_pad , \DM_rdm[3]_pad , \DM_rdm[4]_pad , \DM_rdm[5]_pad , \DM_rdm[6]_pad , \DM_rdm[7]_pad , \DM_rdm[8]_pad , \DM_rdm[9]_pad , IACKn_pad, \IRFS0_pad , \IRFS1_pad , \ISCLK0_pad , \ISCLK1_pad , \ITFS0_pad , \ITFS1_pad , \PIO_oe[0]_pad , \PIO_oe[10]_pad , \PIO_oe[11]_pad , \PIO_oe[1]_pad , \PIO_oe[2]_pad , \PIO_oe[3]_pad , \PIO_oe[4]_pad , \PIO_oe[5]_pad , \PIO_oe[6]_pad , \PIO_oe[7]_pad , \PIO_oe[8]_pad , \PIO_oe[9]_pad , \PIO_out[0]_pad , \PIO_out[10]_pad , \PIO_out[11]_pad , \PIO_out[1]_pad , \PIO_out[2]_pad , \PIO_out[3]_pad , \PIO_out[4]_pad , \PIO_out[5]_pad , \PIO_out[6]_pad , \PIO_out[7]_pad , \PIO_out[8]_pad , \PIO_out[9]_pad , PM_bdry_sel_pad, \PM_rd0[0]_pad , \PM_rd0[10]_pad , \PM_rd0[11]_pad , \PM_rd0[12]_pad , \PM_rd0[13]_pad , \PM_rd0[14]_pad , \PM_rd0[15]_pad , \PM_rd0[1]_pad , \PM_rd0[2]_pad , \PM_rd0[3]_pad , \PM_rd0[4]_pad , \PM_rd0[5]_pad , \PM_rd0[6]_pad , \PM_rd0[7]_pad , \PM_rd0[8]_pad , \PM_rd0[9]_pad , \PM_rd1[0]_pad , \PM_rd1[10]_pad , \PM_rd1[11]_pad , \PM_rd1[12]_pad , \PM_rd1[13]_pad , \PM_rd1[14]_pad , \PM_rd1[15]_pad , \PM_rd1[1]_pad , \PM_rd1[2]_pad , \PM_rd1[3]_pad , \PM_rd1[4]_pad , \PM_rd1[5]_pad , \PM_rd1[6]_pad , \PM_rd1[7]_pad , \PM_rd1[8]_pad , \PM_rd1[9]_pad , \PM_rd2[0]_pad , \PM_rd2[10]_pad , \PM_rd2[11]_pad , \PM_rd2[12]_pad , \PM_rd2[13]_pad , \PM_rd2[14]_pad , \PM_rd2[15]_pad , \PM_rd2[1]_pad , \PM_rd2[2]_pad , \PM_rd2[3]_pad , \PM_rd2[4]_pad , \PM_rd2[5]_pad , \PM_rd2[6]_pad , \PM_rd2[7]_pad , \PM_rd2[8]_pad , \PM_rd2[9]_pad , \PM_rd3[0]_pad , \PM_rd3[10]_pad , \PM_rd3[11]_pad , \PM_rd3[12]_pad , \PM_rd3[13]_pad , \PM_rd3[14]_pad , \PM_rd3[15]_pad , \PM_rd3[1]_pad , \PM_rd3[2]_pad , \PM_rd3[3]_pad , \PM_rd3[4]_pad , \PM_rd3[5]_pad , \PM_rd3[6]_pad , \PM_rd3[7]_pad , \PM_rd3[8]_pad , \PM_rd3[9]_pad , \PM_rd4[0]_pad , \PM_rd4[10]_pad , \PM_rd4[11]_pad , \PM_rd4[12]_pad , \PM_rd4[13]_pad , \PM_rd4[14]_pad , \PM_rd4[15]_pad , \PM_rd4[1]_pad , \PM_rd4[2]_pad , \PM_rd4[3]_pad , \PM_rd4[4]_pad , \PM_rd4[5]_pad , \PM_rd4[6]_pad , \PM_rd4[7]_pad , \PM_rd4[8]_pad , \PM_rd4[9]_pad , \PM_rd5[0]_pad , \PM_rd5[10]_pad , \PM_rd5[11]_pad , \PM_rd5[12]_pad , \PM_rd5[13]_pad , \PM_rd5[14]_pad , \PM_rd5[15]_pad , \PM_rd5[1]_pad , \PM_rd5[2]_pad , \PM_rd5[3]_pad , \PM_rd5[4]_pad , \PM_rd5[5]_pad , \PM_rd5[6]_pad , \PM_rd5[7]_pad , \PM_rd5[8]_pad , \PM_rd5[9]_pad , \PM_rd6[0]_pad , \PM_rd6[10]_pad , \PM_rd6[11]_pad , \PM_rd6[12]_pad , \PM_rd6[13]_pad , \PM_rd6[14]_pad , \PM_rd6[15]_pad , \PM_rd6[1]_pad , \PM_rd6[2]_pad , \PM_rd6[3]_pad , \PM_rd6[4]_pad , \PM_rd6[5]_pad , \PM_rd6[6]_pad , \PM_rd6[7]_pad , \PM_rd6[8]_pad , \PM_rd6[9]_pad , \PM_rd7[0]_pad , \PM_rd7[10]_pad , \PM_rd7[11]_pad , \PM_rd7[12]_pad , \PM_rd7[13]_pad , \PM_rd7[14]_pad , \PM_rd7[15]_pad , \PM_rd7[1]_pad , \PM_rd7[2]_pad , \PM_rd7[3]_pad , \PM_rd7[4]_pad , \PM_rd7[5]_pad , \PM_rd7[6]_pad , \PM_rd7[7]_pad , \PM_rd7[8]_pad , \PM_rd7[9]_pad , PWDACK_pad, T_BMODE_pad, T_BRn_pad, T_CLKI_OSC_pad, T_CLKI_PLL_pad, \T_ED[0]_pad , \T_ED[10]_pad , \T_ED[11]_pad , \T_ED[12]_pad , \T_ED[13]_pad , \T_ED[14]_pad , \T_ED[15]_pad , \T_ED[1]_pad , \T_ED[2]_pad , \T_ED[3]_pad , \T_ED[4]_pad , \T_ED[5]_pad , \T_ED[6]_pad , \T_ED[7]_pad , \T_ED[8]_pad , \T_ED[9]_pad , T_ICE_RSTn_pad, T_ID_pad, T_IMS_pad, T_IRDn_pad, \T_IRQ0n_pad , \T_IRQ1n_pad , \T_IRQ2n_pad , \T_IRQE0n_pad , \T_IRQE1n_pad , \T_IRQL1n_pad , T_ISn_pad, T_IWRn_pad, T_MMAP_pad, \T_PIOin[0]_pad , \T_PIOin[10]_pad , \T_PIOin[11]_pad , \T_PIOin[1]_pad , \T_PIOin[2]_pad , \T_PIOin[3]_pad , \T_PIOin[4]_pad , \T_PIOin[5]_pad , \T_PIOin[6]_pad , \T_PIOin[7]_pad , \T_PIOin[8]_pad , \T_PIOin[9]_pad , T_PWDn_pad, \T_RD0_pad , \T_RD1_pad , \T_RFS0_pad , \T_RFS1_pad , T_RSTn_pad, \T_SCLK0_pad , \T_SCLK1_pad , T_Sel_PLL_pad, \T_TFS0_pad , \T_TFS1_pad , \T_TMODE[0]_pad , \T_TMODE[1]_pad , \auctl_BSack_reg/NET0131 , \auctl_DSack_reg/NET0131 , \auctl_R0Sack_reg/NET0131 , \auctl_R1Sack_reg/NET0131 , \auctl_RST_reg/P0001 , \auctl_STEAL_reg/NET0131 , \auctl_T0Sack_reg/NET0131 , \auctl_T1Sack_reg/NET0131 , \bdma_BCTL_reg[0]/NET0131 , \bdma_BCTL_reg[10]/NET0131 , \bdma_BCTL_reg[11]/NET0131 , \bdma_BCTL_reg[12]/NET0131 , \bdma_BCTL_reg[13]/NET0131 , \bdma_BCTL_reg[14]/NET0131 , \bdma_BCTL_reg[15]/NET0131 , \bdma_BCTL_reg[1]/NET0131 , \bdma_BCTL_reg[2]/NET0131 , \bdma_BCTL_reg[3]/NET0131 , \bdma_BCTL_reg[4]/NET0131 , \bdma_BCTL_reg[5]/NET0131 , \bdma_BCTL_reg[6]/NET0131 , \bdma_BCTL_reg[7]/NET0131 , \bdma_BCTL_reg[8]/NET0131 , \bdma_BCTL_reg[9]/NET0131 , \bdma_BDMA_boot_reg/NET0131_reg_syn_10 , \bdma_BDMA_boot_reg/NET0131_reg_syn_2 , \bdma_BDMA_boot_reg/NET0131_reg_syn_8 , \bdma_BDMAmode_reg/NET0131 , \bdma_BEAD_reg[0]/NET0131 , \bdma_BEAD_reg[10]/NET0131 , \bdma_BEAD_reg[11]/NET0131 , \bdma_BEAD_reg[12]/NET0131 , \bdma_BEAD_reg[13]/NET0131 , \bdma_BEAD_reg[1]/NET0131 , \bdma_BEAD_reg[2]/NET0131 , \bdma_BEAD_reg[3]/NET0131 , \bdma_BEAD_reg[4]/NET0131 , \bdma_BEAD_reg[5]/NET0131 , \bdma_BEAD_reg[6]/NET0131 , \bdma_BEAD_reg[7]/NET0131 , \bdma_BEAD_reg[8]/NET0131 , \bdma_BEAD_reg[9]/NET0131 , \bdma_BIAD_reg[0]/NET0131 , \bdma_BIAD_reg[10]/NET0131 , \bdma_BIAD_reg[11]/NET0131 , \bdma_BIAD_reg[12]/NET0131 , \bdma_BIAD_reg[13]/NET0131 , \bdma_BIAD_reg[1]/NET0131 , \bdma_BIAD_reg[2]/NET0131 , \bdma_BIAD_reg[3]/NET0131 , \bdma_BIAD_reg[4]/NET0131 , \bdma_BIAD_reg[5]/NET0131 , \bdma_BIAD_reg[6]/NET0131 , \bdma_BIAD_reg[7]/NET0131 , \bdma_BIAD_reg[8]/NET0131 , \bdma_BIAD_reg[9]/NET0131 , \bdma_BM_cyc_reg/P0001 , \bdma_BMcyc_del_reg/P0001 , \bdma_BOVL_reg[0]/NET0131 , \bdma_BOVL_reg[10]/NET0131 , \bdma_BOVL_reg[11]/NET0131 , \bdma_BOVL_reg[1]/NET0131 , \bdma_BOVL_reg[2]/NET0131 , \bdma_BOVL_reg[3]/NET0131 , \bdma_BOVL_reg[4]/NET0131 , \bdma_BOVL_reg[5]/NET0131 , \bdma_BOVL_reg[6]/NET0131 , \bdma_BOVL_reg[7]/NET0131 , \bdma_BOVL_reg[8]/NET0131 , \bdma_BOVL_reg[9]/NET0131 , \bdma_BRST_s2_reg/NET0131 , \bdma_BRdataBUF_reg[0]/P0001 , \bdma_BRdataBUF_reg[10]/P0001 , \bdma_BRdataBUF_reg[11]/P0001 , \bdma_BRdataBUF_reg[12]/P0001 , \bdma_BRdataBUF_reg[13]/P0001 , \bdma_BRdataBUF_reg[14]/P0001 , \bdma_BRdataBUF_reg[15]/P0001 , \bdma_BRdataBUF_reg[16]/P0001 , \bdma_BRdataBUF_reg[17]/P0001 , \bdma_BRdataBUF_reg[18]/P0001 , \bdma_BRdataBUF_reg[19]/P0001 , \bdma_BRdataBUF_reg[1]/P0001 , \bdma_BRdataBUF_reg[20]/P0001 , \bdma_BRdataBUF_reg[21]/P0001 , \bdma_BRdataBUF_reg[22]/P0001 , \bdma_BRdataBUF_reg[23]/P0001 , \bdma_BRdataBUF_reg[2]/P0001 , \bdma_BRdataBUF_reg[3]/P0001 , \bdma_BRdataBUF_reg[4]/P0001 , \bdma_BRdataBUF_reg[5]/P0001 , \bdma_BRdataBUF_reg[6]/P0001 , \bdma_BRdataBUF_reg[7]/P0001 , \bdma_BRdataBUF_reg[8]/P0001 , \bdma_BRdataBUF_reg[9]/P0001 , \bdma_BSreq_reg/NET0131 , \bdma_BWCOUNT_reg[0]/NET0131 , \bdma_BWCOUNT_reg[10]/NET0131 , \bdma_BWCOUNT_reg[11]/NET0131 , \bdma_BWCOUNT_reg[12]/NET0131 , \bdma_BWCOUNT_reg[13]/NET0131 , \bdma_BWCOUNT_reg[1]/NET0131 , \bdma_BWCOUNT_reg[2]/NET0131 , \bdma_BWCOUNT_reg[3]/NET0131 , \bdma_BWCOUNT_reg[4]/NET0131 , \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_2 , \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_8 , \bdma_BWCOUNT_reg[6]/NET0131 , \bdma_BWCOUNT_reg[7]/NET0131 , \bdma_BWCOUNT_reg[8]/NET0131 , \bdma_BWCOUNT_reg[9]/NET0131 , \bdma_BWRn_reg/NET0131 , \bdma_BWcnt_reg[0]/NET0131 , \bdma_BWcnt_reg[1]/NET0131 , \bdma_BWcnt_reg[2]/NET0131 , \bdma_BWcnt_reg[3]/NET0131 , \bdma_BWcnt_reg[4]/NET0131 , \bdma_BWdataBUF_h_reg[0]/P0001 , \bdma_BWdataBUF_h_reg[10]/P0001 , \bdma_BWdataBUF_h_reg[11]/P0001 , \bdma_BWdataBUF_h_reg[12]/P0001 , \bdma_BWdataBUF_h_reg[13]/P0001 , \bdma_BWdataBUF_h_reg[14]/P0001 , \bdma_BWdataBUF_h_reg[15]/P0001 , \bdma_BWdataBUF_h_reg[16]/P0001 , \bdma_BWdataBUF_h_reg[17]/P0001 , \bdma_BWdataBUF_h_reg[18]/P0001 , \bdma_BWdataBUF_h_reg[19]/P0001 , \bdma_BWdataBUF_h_reg[1]/P0001 , \bdma_BWdataBUF_h_reg[20]/P0001 , \bdma_BWdataBUF_h_reg[21]/P0001 , \bdma_BWdataBUF_h_reg[22]/P0001 , \bdma_BWdataBUF_h_reg[23]/P0001 , \bdma_BWdataBUF_h_reg[2]/P0001 , \bdma_BWdataBUF_h_reg[3]/P0001 , \bdma_BWdataBUF_h_reg[4]/P0001 , \bdma_BWdataBUF_h_reg[5]/P0001 , \bdma_BWdataBUF_h_reg[6]/P0001 , \bdma_BWdataBUF_h_reg[7]/P0001 , \bdma_BWdataBUF_h_reg[8]/P0001 , \bdma_BWdataBUF_h_reg[9]/P0001 , \bdma_BWdataBUF_reg[0]/P0001 , \bdma_BWdataBUF_reg[1]/P0001 , \bdma_BWdataBUF_reg[2]/P0001 , \bdma_BWdataBUF_reg[3]/P0001 , \bdma_BWdataBUF_reg[4]/P0001 , \bdma_BWdataBUF_reg[5]/P0001 , \bdma_BWdataBUF_reg[6]/P0001 , \bdma_BWdataBUF_reg[7]/P0001 , \bdma_CMcnt_reg[0]/NET0131 , \bdma_CMcnt_reg[1]/NET0131 , \bdma_DM_2nd_reg/NET0131 , \bdma_RST_pin_reg/P0001 , \bdma_WRlat_reg/P0001 , \clkc_Awake_reg/NET0131 , \clkc_CLKOUT_reg/NET0131 , \clkc_CTR_cnt_reg[0]/NET0131 , \clkc_CTR_cnt_reg[1]/NET0131 , \clkc_Cnt128_reg/NET0131 , \clkc_Cnt4096_reg/NET0131 , \clkc_Cnt4096_s1_reg/NET0131 , \clkc_Cnt4096_s2_reg/NET0131 , \clkc_DSPoff_reg/NET0131 , \clkc_OSCoff_reg/NET0131 , \clkc_OSCoff_set_reg/P0001 , \clkc_OUTcnt_reg[0]/NET0131 , \clkc_OUTcnt_reg[1]/NET0131 , \clkc_OUTcnt_reg[2]/NET0131 , \clkc_OUTcnt_reg[3]/NET0131 , \clkc_OUTcnt_reg[4]/NET0131 , \clkc_OUTcnt_reg[5]/NET0131 , \clkc_OUTcnt_reg[6]/NET0131 , \clkc_RSTtext_reg/P0001 , \clkc_SIDLE_s1_reg/NET0131 , \clkc_SIDLE_s2_reg/NET0131 , \clkc_SLEEP_reg/NET0131 , \clkc_STBY_reg/NET0131 , \clkc_STDcnt_reg[0]/NET0131 , \clkc_STDcnt_reg[10]/NET0131 , \clkc_STDcnt_reg[1]/NET0131 , \clkc_STDcnt_reg[2]/NET0131 , \clkc_STDcnt_reg[3]/NET0131 , \clkc_STDcnt_reg[4]/NET0131 , \clkc_STDcnt_reg[5]/NET0131 , \clkc_STDcnt_reg[6]/NET0131 , \clkc_STDcnt_reg[7]/NET0131 , \clkc_STDcnt_reg[8]/NET0131 , \clkc_STDcnt_reg[9]/NET0131 , \clkc_SlowDn_reg/NET0131 , \clkc_SlowDn_s1_reg/P0001 , \clkc_SlowDn_s2_reg/P0001 , \clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131 , \clkc_ckr_reg_DO_reg[0]/NET0131 , \clkc_ckr_reg_DO_reg[10]/NET0131 , \clkc_ckr_reg_DO_reg[11]/NET0131 , \clkc_ckr_reg_DO_reg[12]/NET0131 , \clkc_ckr_reg_DO_reg[13]/NET0131 , \clkc_ckr_reg_DO_reg[14]/NET0131 , \clkc_ckr_reg_DO_reg[15]/NET0131 , \clkc_ckr_reg_DO_reg[1]/NET0131 , \clkc_ckr_reg_DO_reg[2]/NET0131 , \clkc_ckr_reg_DO_reg[3]/NET0131 , \clkc_ckr_reg_DO_reg[4]/NET0131 , \clkc_ckr_reg_DO_reg[5]/NET0131 , \clkc_ckr_reg_DO_reg[6]/NET0131 , \clkc_ckr_reg_DO_reg[7]/NET0131 , \clkc_ckr_reg_DO_reg[8]/NET0131 , \clkc_ckr_reg_DO_reg[9]/NET0131 , \clkc_oscntr_reg_DO_reg[0]/NET0131 , \clkc_oscntr_reg_DO_reg[10]/NET0131 , \clkc_oscntr_reg_DO_reg[11]/NET0131 , \clkc_oscntr_reg_DO_reg[1]/NET0131 , \clkc_oscntr_reg_DO_reg[2]/NET0131 , \clkc_oscntr_reg_DO_reg[3]/NET0131 , \clkc_oscntr_reg_DO_reg[4]/NET0131 , \clkc_oscntr_reg_DO_reg[5]/NET0131 , \clkc_oscntr_reg_DO_reg[6]/NET0131 , \clkc_oscntr_reg_DO_reg[7]/NET0131 , \clkc_oscntr_reg_DO_reg[8]/NET0131 , \clkc_oscntr_reg_DO_reg[9]/NET0131 , \core_c_dec_ALUop_E_reg/P0001 , \core_c_dec_BR_Ed_reg/P0001 , \core_c_dec_Call_Ed_reg/P0001 , \core_c_dec_DIVQ_E_reg/P0001 , \core_c_dec_DIVS_E_reg/P0001 , \core_c_dec_DU_Eg_reg/P0001 , \core_c_dec_Double_E_reg/P0001 , \core_c_dec_Dummy_E_reg/NET0131 , \core_c_dec_EXIT_E_reg/P0001 , \core_c_dec_IDLE_Eg_reg/P0001 , \core_c_dec_IRE_reg[0]/NET0131 , \core_c_dec_IRE_reg[10]/NET0131 , \core_c_dec_IRE_reg[11]/NET0131 , \core_c_dec_IRE_reg[12]/NET0131 , \core_c_dec_IRE_reg[13]/NET0131 , \core_c_dec_IRE_reg[14]/NET0131 , \core_c_dec_IRE_reg[15]/NET0131 , \core_c_dec_IRE_reg[16]/NET0131 , \core_c_dec_IRE_reg[17]/NET0131 , \core_c_dec_IRE_reg[18]/NET0131 , \core_c_dec_IRE_reg[19]/NET0131 , \core_c_dec_IRE_reg[1]/NET0131 , \core_c_dec_IRE_reg[2]/NET0131 , \core_c_dec_IRE_reg[3]/NET0131 , \core_c_dec_IRE_reg[4]/NET0131 , \core_c_dec_IRE_reg[5]/NET0131 , \core_c_dec_IRE_reg[6]/NET0131 , \core_c_dec_IRE_reg[7]/NET0131 , \core_c_dec_IRE_reg[8]/NET0131 , \core_c_dec_IRE_reg[9]/NET0131 , \core_c_dec_IR_reg[0]/NET0131 , \core_c_dec_IR_reg[10]/NET0131 , \core_c_dec_IR_reg[11]/NET0131 , \core_c_dec_IR_reg[12]/NET0131 , \core_c_dec_IR_reg[13]/NET0131 , \core_c_dec_IR_reg[14]/NET0131 , \core_c_dec_IR_reg[15]/NET0131 , \core_c_dec_IR_reg[16]/NET0131 , \core_c_dec_IR_reg[17]/NET0131 , \core_c_dec_IR_reg[18]/NET0131 , \core_c_dec_IR_reg[19]/NET0131 , \core_c_dec_IR_reg[1]/NET0131 , \core_c_dec_IR_reg[20]/NET0131 , \core_c_dec_IR_reg[21]/NET0131 , \core_c_dec_IR_reg[22]/NET0131 , \core_c_dec_IR_reg[23]/NET0131 , \core_c_dec_IR_reg[2]/NET0131 , \core_c_dec_IR_reg[3]/NET0131 , \core_c_dec_IR_reg[4]/NET0131 , \core_c_dec_IR_reg[5]/NET0131 , \core_c_dec_IR_reg[6]/NET0131 , \core_c_dec_IR_reg[7]/NET0131 , \core_c_dec_IR_reg[8]/NET0131 , \core_c_dec_IR_reg[9]/NET0131 , \core_c_dec_Long_Cg_reg/P0001 , \core_c_dec_Long_Eg_reg/P0001 , \core_c_dec_MACdep_Eg_reg/P0001 , \core_c_dec_MACop_E_reg/P0001 , \core_c_dec_MFALU_Ei_reg/NET0131 , \core_c_dec_MFAR_E_reg/P0001 , \core_c_dec_MFASTAT_E_reg/P0001 , \core_c_dec_MFAX0_E_reg/P0001 , \core_c_dec_MFAX1_E_reg/P0001 , \core_c_dec_MFAY0_E_reg/P0001 , \core_c_dec_MFAY1_E_reg/P0001 , \core_c_dec_MFCNTR_E_reg/P0001 , \core_c_dec_MFDAG1_Ei_reg/NET0131 , \core_c_dec_MFDAG2_Ei_reg/NET0131 , \core_c_dec_MFDMOVL_E_reg/P0001 , \core_c_dec_MFICNTL_E_reg/P0001 , \core_c_dec_MFIDR_E_reg/P0001 , \core_c_dec_MFIMASK_E_reg/P0001 , \core_c_dec_MFIreg_E_reg[0]/P0001 , \core_c_dec_MFIreg_E_reg[1]/P0001 , \core_c_dec_MFIreg_E_reg[2]/P0001 , \core_c_dec_MFIreg_E_reg[3]/P0001 , \core_c_dec_MFIreg_E_reg[4]/P0001 , \core_c_dec_MFIreg_E_reg[5]/P0001 , \core_c_dec_MFIreg_E_reg[6]/P0001 , \core_c_dec_MFIreg_E_reg[7]/P0001 , \core_c_dec_MFLreg_E_reg[0]/P0001 , \core_c_dec_MFLreg_E_reg[1]/P0001 , \core_c_dec_MFLreg_E_reg[2]/P0001 , \core_c_dec_MFLreg_E_reg[3]/P0001 , \core_c_dec_MFLreg_E_reg[4]/P0001 , \core_c_dec_MFLreg_E_reg[5]/P0001 , \core_c_dec_MFLreg_E_reg[6]/P0001 , \core_c_dec_MFLreg_E_reg[7]/P0001 , \core_c_dec_MFMAC_Ei_reg/NET0131 , \core_c_dec_MFMR0_E_reg/P0001 , \core_c_dec_MFMR1_E_reg/P0001 , \core_c_dec_MFMR2_E_reg/P0001 , \core_c_dec_MFMSTAT_E_reg/P0001 , \core_c_dec_MFMX0_E_reg/P0001 , \core_c_dec_MFMX1_E_reg/P0001 , \core_c_dec_MFMY0_E_reg/P0001 , \core_c_dec_MFMY1_E_reg/P0001 , \core_c_dec_MFMreg_E_reg[0]/P0001 , \core_c_dec_MFMreg_E_reg[1]/P0001 , \core_c_dec_MFMreg_E_reg[2]/P0001 , \core_c_dec_MFMreg_E_reg[3]/P0001 , \core_c_dec_MFMreg_E_reg[4]/P0001 , \core_c_dec_MFMreg_E_reg[5]/P0001 , \core_c_dec_MFMreg_E_reg[6]/P0001 , \core_c_dec_MFMreg_E_reg[7]/P0001 , \core_c_dec_MFPMOVL_E_reg/P0001 , \core_c_dec_MFPSQ_Ei_reg/NET0131 , \core_c_dec_MFRX0_E_reg/P0001 , \core_c_dec_MFRX1_E_reg/P0001 , \core_c_dec_MFSB_E_reg/P0001 , \core_c_dec_MFSE_E_reg/P0001 , \core_c_dec_MFSHT_Ei_reg/NET0131 , \core_c_dec_MFSI_E_reg/P0001 , \core_c_dec_MFSPT_Ei_reg/NET0131 , \core_c_dec_MFSR0_E_reg/P0001 , \core_c_dec_MFSR1_E_reg/P0001 , \core_c_dec_MFSSTAT_E_reg/P0001 , \core_c_dec_MFTX0_E_reg/P0001 , \core_c_dec_MFTX1_E_reg/P0001 , \core_c_dec_MFtoppcs_Eg_reg/P0001 , \core_c_dec_MTAR_E_reg/P0001 , \core_c_dec_MTASTAT_E_reg/P0001 , \core_c_dec_MTAX0_E_reg/P0001 , \core_c_dec_MTAX1_E_reg/P0001 , \core_c_dec_MTAY0_E_reg/P0001 , \core_c_dec_MTAY1_E_reg/P0001 , \core_c_dec_MTCNTR_Eg_reg/P0001 , \core_c_dec_MTDMOVL_E_reg/P0001 , \core_c_dec_MTICNTL_Eg_reg/P0001 , \core_c_dec_MTIDR_E_reg/P0001 , \core_c_dec_MTIFC_Eg_reg/P0001 , \core_c_dec_MTIMASK_Eg_reg/P0001 , \core_c_dec_MTIreg_E_reg[0]/P0001 , \core_c_dec_MTIreg_E_reg[1]/P0001 , \core_c_dec_MTIreg_E_reg[2]/P0001 , \core_c_dec_MTIreg_E_reg[3]/P0001 , \core_c_dec_MTIreg_E_reg[4]/P0001 , \core_c_dec_MTIreg_E_reg[5]/P0001 , \core_c_dec_MTIreg_E_reg[6]/P0001 , \core_c_dec_MTIreg_E_reg[7]/P0001 , \core_c_dec_MTLreg_E_reg[0]/P0001 , \core_c_dec_MTLreg_E_reg[1]/P0001 , \core_c_dec_MTLreg_E_reg[2]/P0001 , \core_c_dec_MTLreg_E_reg[3]/P0001 , \core_c_dec_MTLreg_E_reg[4]/P0001 , \core_c_dec_MTLreg_E_reg[5]/P0001 , \core_c_dec_MTLreg_E_reg[6]/P0001 , \core_c_dec_MTLreg_E_reg[7]/P0001 , \core_c_dec_MTMR0_E_reg/P0001 , \core_c_dec_MTMR1_E_reg/P0001 , \core_c_dec_MTMR2_E_reg/P0001 , \core_c_dec_MTMSTAT_Eg_reg/P0001 , \core_c_dec_MTMX0_E_reg/P0001 , \core_c_dec_MTMX1_E_reg/P0001 , \core_c_dec_MTMY0_E_reg/P0001 , \core_c_dec_MTMY1_E_reg/P0001 , \core_c_dec_MTMreg_E_reg[0]/P0001 , \core_c_dec_MTMreg_E_reg[1]/P0001 , \core_c_dec_MTMreg_E_reg[2]/P0001 , \core_c_dec_MTMreg_E_reg[3]/P0001 , \core_c_dec_MTMreg_E_reg[4]/P0001 , \core_c_dec_MTMreg_E_reg[5]/P0001 , \core_c_dec_MTMreg_E_reg[6]/P0001 , \core_c_dec_MTMreg_E_reg[7]/P0001 , \core_c_dec_MTOWRCNTR_Eg_reg/P0001 , \core_c_dec_MTPMOVL_E_reg/P0001 , \core_c_dec_MTRX0_E_reg/P0001 , \core_c_dec_MTRX1_E_reg/P0001 , \core_c_dec_MTSB_E_reg/P0001 , \core_c_dec_MTSE_E_reg/P0001 , \core_c_dec_MTSI_E_reg/P0001 , \core_c_dec_MTSR0_E_reg/P0001 , \core_c_dec_MTSR1_E_reg/P0001 , \core_c_dec_MTTX0_E_reg/P0001 , \core_c_dec_MTTX1_E_reg/P0001 , \core_c_dec_MTtoppcs_Eg_reg/P0001 , \core_c_dec_Modctl_Eg_reg/P0001 , \core_c_dec_MpopLP_Eg_reg/P0001 , \core_c_dec_NOP_E_reg/P0001 , \core_c_dec_Nrti_Ed_reg/P0001 , \core_c_dec_Nseq_Ed_reg/P0001 , \core_c_dec_PPclr_reg/P0001 , \core_c_dec_Post1_E_reg/P0001 , \core_c_dec_Post2_E_reg/P0001 , \core_c_dec_Prderr_Cg_reg/NET0131 , \core_c_dec_RET_Ed_reg/P0001 , \core_c_dec_RTI_Ed_reg/P0001 , \core_c_dec_SHTop_E_reg/P0001 , \core_c_dec_Stkctl_Eg_reg/P0001 , \core_c_dec_Usecond_E_reg/P0001 , \core_c_dec_accCM_E_reg/NET0131 , \core_c_dec_accPM_E_reg/P0001 , \core_c_dec_cdAM_E_reg/P0001 , \core_c_dec_imSHT_E_reg/P0001 , \core_c_dec_imm14_E_reg/P0001 , \core_c_dec_imm16_E_reg/P0001 , \core_c_dec_pMFALU_Ei_reg/NET0131 , \core_c_dec_pMFMAC_Ei_reg/NET0131 , \core_c_dec_pMFSHT_Ei_reg/NET0131 , \core_c_dec_rdCM_E_reg/NET0131 , \core_c_dec_satMR_E_reg/P0001 , \core_c_dec_updAF_E_reg/P0001 , \core_c_dec_updAR_E_reg/P0001 , \core_c_dec_updMF_E_reg/P0001 , \core_c_dec_updMR_E_reg/P0001 , \core_c_dec_updSR_E_reg/P0001 , \core_c_psq_CE_reg/NET0131 , \core_c_psq_CNTR_reg_DO_reg[0]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[10]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[11]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[12]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[13]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[1]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[2]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[3]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[4]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[5]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[6]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[7]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[8]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[9]/NET0131 , \core_c_psq_CNTRval_reg/NET0131 , \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 , \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 , \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 , \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 , \core_c_psq_DRA_reg[0]/P0001 , \core_c_psq_DRA_reg[10]/P0001 , \core_c_psq_DRA_reg[11]/P0001 , \core_c_psq_DRA_reg[12]/P0001 , \core_c_psq_DRA_reg[13]/P0001 , \core_c_psq_DRA_reg[1]/P0001 , \core_c_psq_DRA_reg[2]/P0001 , \core_c_psq_DRA_reg[3]/P0001 , \core_c_psq_DRA_reg[4]/P0001 , \core_c_psq_DRA_reg[5]/P0001 , \core_c_psq_DRA_reg[6]/P0001 , \core_c_psq_DRA_reg[7]/P0001 , \core_c_psq_DRA_reg[8]/P0001 , \core_c_psq_DRA_reg[9]/P0001 , \core_c_psq_ECYC_reg/P0001 , \core_c_psq_EXA_reg[0]/P0001 , \core_c_psq_EXA_reg[10]/P0001 , \core_c_psq_EXA_reg[11]/P0001 , \core_c_psq_EXA_reg[12]/P0001 , \core_c_psq_EXA_reg[13]/P0001 , \core_c_psq_EXA_reg[1]/P0001 , \core_c_psq_EXA_reg[2]/P0001 , \core_c_psq_EXA_reg[3]/P0001 , \core_c_psq_EXA_reg[4]/P0001 , \core_c_psq_EXA_reg[5]/P0001 , \core_c_psq_EXA_reg[6]/P0001 , \core_c_psq_EXA_reg[7]/P0001 , \core_c_psq_EXA_reg[8]/P0001 , \core_c_psq_EXA_reg[9]/P0001 , \core_c_psq_Eqend_D_reg/P0001 , \core_c_psq_Eqend_Ed_reg/P0001 , \core_c_psq_ICNTL_reg_DO_reg[0]/NET0131 , \core_c_psq_ICNTL_reg_DO_reg[1]/NET0131 , \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 , \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 , \core_c_psq_IFA_reg[0]/P0001 , \core_c_psq_IFA_reg[10]/P0001 , \core_c_psq_IFA_reg[11]/P0001 , \core_c_psq_IFA_reg[12]/P0001 , \core_c_psq_IFA_reg[13]/P0001 , \core_c_psq_IFA_reg[1]/P0001 , \core_c_psq_IFA_reg[2]/P0001 , \core_c_psq_IFA_reg[3]/P0001 , \core_c_psq_IFA_reg[4]/P0001 , \core_c_psq_IFA_reg[5]/P0001 , \core_c_psq_IFA_reg[6]/P0001 , \core_c_psq_IFA_reg[7]/P0001 , \core_c_psq_IFA_reg[8]/P0001 , \core_c_psq_IFA_reg[9]/P0001 , \core_c_psq_IFC_reg[0]/NET0131 , \core_c_psq_IFC_reg[10]/NET0131 , \core_c_psq_IFC_reg[11]/NET0131 , \core_c_psq_IFC_reg[12]/NET0131 , \core_c_psq_IFC_reg[13]/NET0131 , \core_c_psq_IFC_reg[14]/NET0131 , \core_c_psq_IFC_reg[15]/NET0131 , \core_c_psq_IFC_reg[1]/NET0131 , \core_c_psq_IFC_reg[2]/NET0131 , \core_c_psq_IFC_reg[3]/NET0131 , \core_c_psq_IFC_reg[4]/NET0131 , \core_c_psq_IFC_reg[5]/NET0131 , \core_c_psq_IFC_reg[6]/NET0131 , \core_c_psq_IFC_reg[7]/NET0131 , \core_c_psq_IFC_reg[8]/NET0131 , \core_c_psq_IFC_reg[9]/NET0131 , \core_c_psq_IMASK_reg[0]/NET0131 , \core_c_psq_IMASK_reg[1]/NET0131 , \core_c_psq_IMASK_reg[2]/NET0131 , \core_c_psq_IMASK_reg[3]/NET0131 , \core_c_psq_IMASK_reg[4]/NET0131 , \core_c_psq_IMASK_reg[5]/NET0131 , \core_c_psq_IMASK_reg[6]/NET0131 , \core_c_psq_IMASK_reg[7]/NET0131 , \core_c_psq_IMASK_reg[8]/NET0131 , \core_c_psq_IMASK_reg[9]/NET0131 , \core_c_psq_INT_en_reg/NET0131 , \core_c_psq_Iact_E_reg[0]/NET0131 , \core_c_psq_Iact_E_reg[10]/NET0131 , \core_c_psq_Iact_E_reg[1]/NET0131 , \core_c_psq_Iact_E_reg[2]/NET0131 , \core_c_psq_Iact_E_reg[3]/NET0131 , \core_c_psq_Iact_E_reg[4]/NET0131 , \core_c_psq_Iact_E_reg[5]/NET0131 , \core_c_psq_Iact_E_reg[6]/NET0131 , \core_c_psq_Iact_E_reg[7]/NET0131 , \core_c_psq_Iact_E_reg[8]/NET0131 , \core_c_psq_Iact_E_reg[9]/NET0131 , \core_c_psq_Iflag_reg[0]/NET0131 , \core_c_psq_Iflag_reg[10]/NET0131 , \core_c_psq_Iflag_reg[11]/NET0131 , \core_c_psq_Iflag_reg[12]/NET0131 , \core_c_psq_Iflag_reg[1]/NET0131 , \core_c_psq_Iflag_reg[2]/NET0131 , \core_c_psq_Iflag_reg[3]/NET0131 , \core_c_psq_Iflag_reg[4]/NET0131 , \core_c_psq_Iflag_reg[5]/NET0131 , \core_c_psq_Iflag_reg[6]/NET0131 , \core_c_psq_Iflag_reg[7]/NET0131 , \core_c_psq_Iflag_reg[8]/NET0131 , \core_c_psq_Iflag_reg[9]/NET0131 , \core_c_psq_MGNT_reg/NET0131 , \core_c_psq_MREQ_reg/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[0]/P0002 , \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 , \core_c_psq_PCS2or3_reg/NET0131 , \core_c_psq_PCS_reg[0]/NET0131 , \core_c_psq_PCS_reg[10]/NET0131 , \core_c_psq_PCS_reg[11]/NET0131 , \core_c_psq_PCS_reg[12]/NET0131 , \core_c_psq_PCS_reg[13]/NET0131 , \core_c_psq_PCS_reg[14]/NET0131 , \core_c_psq_PCS_reg[15]/NET0131 , \core_c_psq_PCS_reg[1]/NET0131 , \core_c_psq_PCS_reg[2]/NET0131 , \core_c_psq_PCS_reg[3]/NET0131 , \core_c_psq_PCS_reg[4]/NET0131 , \core_c_psq_PCS_reg[5]/NET0131 , \core_c_psq_PCS_reg[6]/NET0131 , \core_c_psq_PCS_reg[7]/NET0131 , \core_c_psq_PCS_reg[8]/NET0131 , \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 , \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 , \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 , \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 , \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 , \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 , \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 , \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 , \core_c_psq_SRST_reg/P0001 , \core_c_psq_SSTAT_reg[0]/NET0131 , \core_c_psq_SSTAT_reg[1]/NET0131 , \core_c_psq_SSTAT_reg[2]/NET0131 , \core_c_psq_SSTAT_reg[3]/NET0131 , \core_c_psq_SSTAT_reg[4]/NET0131 , \core_c_psq_SSTAT_reg[5]/NET0131 , \core_c_psq_SSTAT_reg[6]/NET0131 , \core_c_psq_SSTAT_reg[7]/NET0131 , \core_c_psq_TRAP_Eg_reg/NET0131 , \core_c_psq_TRAP_R_L_reg/NET0131 , \core_c_psq_T_IRQ0_s1_reg/P0001 , \core_c_psq_T_IRQ0p_reg/P0001 , \core_c_psq_T_IRQ1_s1_reg/P0001 , \core_c_psq_T_IRQ1p_reg/P0001 , \core_c_psq_T_IRQ2_s1_reg/P0001 , \core_c_psq_T_IRQ2p_reg/P0001 , \core_c_psq_T_IRQE0_reg/P0001 , \core_c_psq_T_IRQE0_s1_reg/P0001 , \core_c_psq_T_IRQE1_reg/P0001 , \core_c_psq_T_IRQE1_s1_reg/P0001 , \core_c_psq_T_IRQL0p_reg/P0001 , \core_c_psq_T_IRQL1p_reg/P0001 , \core_c_psq_T_PWRDN_reg/P0001 , \core_c_psq_T_PWRDN_s1_reg/P0001 , \core_c_psq_Taddr_Eb_reg[0]/P0001 , \core_c_psq_Taddr_Eb_reg[10]/P0001 , \core_c_psq_Taddr_Eb_reg[11]/P0001 , \core_c_psq_Taddr_Eb_reg[12]/P0001 , \core_c_psq_Taddr_Eb_reg[13]/P0001 , \core_c_psq_Taddr_Eb_reg[1]/P0001 , \core_c_psq_Taddr_Eb_reg[2]/P0001 , \core_c_psq_Taddr_Eb_reg[3]/P0001 , \core_c_psq_Taddr_Eb_reg[4]/P0001 , \core_c_psq_Taddr_Eb_reg[5]/P0001 , \core_c_psq_Taddr_Eb_reg[6]/P0001 , \core_c_psq_Taddr_Eb_reg[7]/P0001 , \core_c_psq_Taddr_Eb_reg[8]/P0001 , \core_c_psq_Taddr_Eb_reg[9]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001 , \core_c_psq_cntstk_ptr_reg[0]/NET0131 , \core_c_psq_cntstk_ptr_reg[1]/NET0131 , \core_c_psq_cntstk_ptr_reg[2]/NET0131 , \core_c_psq_irq0_de_IN_syn_reg/P0001 , \core_c_psq_irq0_de_OUT_reg/P0001 , \core_c_psq_irq1_de_IN_syn_reg/P0001 , \core_c_psq_irq1_de_OUT_reg/P0001 , \core_c_psq_irq2_de_IN_syn_reg/P0001 , \core_c_psq_irq2_de_OUT_reg/P0001 , \core_c_psq_irql0_de_IN_syn_reg/P0001 , \core_c_psq_irql0_de_OUT_reg/P0001 , \core_c_psq_irql1_de_IN_syn_reg/P0001 , \core_c_psq_irql1_de_OUT_reg/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001 , \core_c_psq_lpstk_ptr_reg[0]/NET0131 , \core_c_psq_lpstk_ptr_reg[1]/NET0131 , \core_c_psq_lpstk_ptr_reg[2]/NET0131 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001 , \core_c_psq_pcstk_ptr_reg[0]/NET0131 , \core_c_psq_pcstk_ptr_reg[1]/NET0131 , \core_c_psq_pcstk_ptr_reg[2]/NET0131 , \core_c_psq_pcstk_ptr_reg[3]/NET0131 , \core_c_psq_pcstk_ptr_reg[4]/NET0131 , \core_c_psq_ststk_ptr_reg[0]/NET0131 , \core_c_psq_ststk_ptr_reg[1]/NET0131 , \core_c_psq_ststk_ptr_reg[2]/NET0131 , \core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001 , \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I_reg[0]/NET0131 , \core_dag_ilm1reg_I_reg[10]/NET0131 , \core_dag_ilm1reg_I_reg[11]/NET0131 , \core_dag_ilm1reg_I_reg[12]/NET0131 , \core_dag_ilm1reg_I_reg[13]/NET0131 , \core_dag_ilm1reg_I_reg[1]/NET0131 , \core_dag_ilm1reg_I_reg[2]/NET0131 , \core_dag_ilm1reg_I_reg[3]/NET0131 , \core_dag_ilm1reg_I_reg[4]/NET0131 , \core_dag_ilm1reg_I_reg[5]/NET0131 , \core_dag_ilm1reg_I_reg[6]/NET0131 , \core_dag_ilm1reg_I_reg[7]/NET0131 , \core_dag_ilm1reg_I_reg[8]/NET0131 , \core_dag_ilm1reg_I_reg[9]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_L_reg[0]/NET0131 , \core_dag_ilm1reg_L_reg[10]/NET0131 , \core_dag_ilm1reg_L_reg[11]/NET0131 , \core_dag_ilm1reg_L_reg[12]/NET0131 , \core_dag_ilm1reg_L_reg[13]/NET0131 , \core_dag_ilm1reg_L_reg[1]/NET0131 , \core_dag_ilm1reg_L_reg[2]/NET0131 , \core_dag_ilm1reg_L_reg[3]/NET0131 , \core_dag_ilm1reg_L_reg[4]/NET0131 , \core_dag_ilm1reg_L_reg[5]/NET0131 , \core_dag_ilm1reg_L_reg[6]/NET0131 , \core_dag_ilm1reg_L_reg[7]/NET0131 , \core_dag_ilm1reg_L_reg[8]/NET0131 , \core_dag_ilm1reg_L_reg[9]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_M_reg[0]/NET0131 , \core_dag_ilm1reg_M_reg[10]/NET0131 , \core_dag_ilm1reg_M_reg[11]/NET0131 , \core_dag_ilm1reg_M_reg[12]/NET0131 , \core_dag_ilm1reg_M_reg[13]/NET0131 , \core_dag_ilm1reg_M_reg[1]/NET0131 , \core_dag_ilm1reg_M_reg[2]/NET0131 , \core_dag_ilm1reg_M_reg[3]/NET0131 , \core_dag_ilm1reg_M_reg[4]/NET0131 , \core_dag_ilm1reg_M_reg[5]/NET0131 , \core_dag_ilm1reg_M_reg[6]/NET0131 , \core_dag_ilm1reg_M_reg[7]/NET0131 , \core_dag_ilm1reg_M_reg[8]/NET0131 , \core_dag_ilm1reg_M_reg[9]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[0]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[1]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[2]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[3]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[4]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131 , \core_dag_ilm1reg_STEALI_E_reg[0]/P0001 , \core_dag_ilm1reg_STEALI_E_reg[1]/P0001 , \core_dag_ilm1reg_STEALI_E_reg[2]/P0001 , \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_IL_E_reg[0]/P0001 , \core_dag_ilm2reg_IL_E_reg[1]/P0001 , \core_dag_ilm2reg_I_reg[0]/NET0131 , \core_dag_ilm2reg_I_reg[10]/NET0131 , \core_dag_ilm2reg_I_reg[11]/NET0131 , \core_dag_ilm2reg_I_reg[12]/NET0131 , \core_dag_ilm2reg_I_reg[13]/NET0131 , \core_dag_ilm2reg_I_reg[1]/NET0131 , \core_dag_ilm2reg_I_reg[2]/NET0131 , \core_dag_ilm2reg_I_reg[3]/NET0131 , \core_dag_ilm2reg_I_reg[4]/NET0131 , \core_dag_ilm2reg_I_reg[5]/NET0131 , \core_dag_ilm2reg_I_reg[6]/NET0131 , \core_dag_ilm2reg_I_reg[7]/NET0131 , \core_dag_ilm2reg_I_reg[8]/NET0131 , \core_dag_ilm2reg_I_reg[9]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_L_reg[0]/NET0131 , \core_dag_ilm2reg_L_reg[10]/NET0131 , \core_dag_ilm2reg_L_reg[11]/NET0131 , \core_dag_ilm2reg_L_reg[12]/NET0131 , \core_dag_ilm2reg_L_reg[13]/NET0131 , \core_dag_ilm2reg_L_reg[1]/NET0131 , \core_dag_ilm2reg_L_reg[2]/NET0131 , \core_dag_ilm2reg_L_reg[3]/NET0131 , \core_dag_ilm2reg_L_reg[4]/NET0131 , \core_dag_ilm2reg_L_reg[5]/NET0131 , \core_dag_ilm2reg_L_reg[6]/NET0131 , \core_dag_ilm2reg_L_reg[7]/NET0131 , \core_dag_ilm2reg_L_reg[8]/NET0131 , \core_dag_ilm2reg_L_reg[9]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_M_E_reg[0]/NET0131 , \core_dag_ilm2reg_M_E_reg[1]/NET0131 , \core_dag_ilm2reg_M_reg[0]/NET0131 , \core_dag_ilm2reg_M_reg[10]/NET0131 , \core_dag_ilm2reg_M_reg[11]/NET0131 , \core_dag_ilm2reg_M_reg[12]/NET0131 , \core_dag_ilm2reg_M_reg[13]/NET0131 , \core_dag_ilm2reg_M_reg[1]/NET0131 , \core_dag_ilm2reg_M_reg[2]/NET0131 , \core_dag_ilm2reg_M_reg[3]/NET0131 , \core_dag_ilm2reg_M_reg[4]/NET0131 , \core_dag_ilm2reg_M_reg[5]/NET0131 , \core_dag_ilm2reg_M_reg[6]/NET0131 , \core_dag_ilm2reg_M_reg[7]/NET0131 , \core_dag_ilm2reg_M_reg[8]/NET0131 , \core_dag_ilm2reg_M_reg[9]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 , \core_dag_modulo1_R0wrap_reg/P0001 , \core_dag_modulo1_R1wrap_reg/P0001 , \core_dag_modulo1_T0wrap_reg/P0001 , \core_dag_modulo1_T1wrap_reg/P0001 , \core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 , \core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 , \core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 , \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 , \core_eu_ea_alu_ea_dec_AMF_E_reg[4]/NET0131 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001 , \core_eu_ec_cun_AC_reg/P0001 , \core_eu_ec_cun_AN_reg/P0001 , \core_eu_ec_cun_AQ_reg/P0001 , \core_eu_ec_cun_AS_reg/P0001 , \core_eu_ec_cun_AV_reg/P0001 , \core_eu_ec_cun_AZ_reg/P0001 , \core_eu_ec_cun_COND_E_reg[0]/P0001 , \core_eu_ec_cun_COND_E_reg[1]/P0001 , \core_eu_ec_cun_COND_E_reg[2]/P0001 , \core_eu_ec_cun_COND_E_reg[3]/P0001 , \core_eu_ec_cun_MV_reg/P0000_reg_syn_2 , \core_eu_ec_cun_MVi_pre_C_reg/P0001 , \core_eu_ec_cun_SS_reg/P0001 , \core_eu_ec_cun_TERM_E_reg[0]/P0001 , \core_eu_ec_cun_TERM_E_reg[1]/P0001 , \core_eu_ec_cun_TERM_E_reg[2]/P0001 , \core_eu_ec_cun_TERM_E_reg[3]/P0001 , \core_eu_ec_cun_condOK_CE_reg/P0001 , \core_eu_ec_cun_mven_FFout_reg/NET0131 , \core_eu_ec_cun_termOK_CE_reg/P0001 , \core_eu_ec_cun_updateMV_C_reg/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_Sq_E_reg/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 , \core_eu_em_mac_em_reg_s1_reg/P0000_reg_syn_2 , \core_eu_em_mac_em_reg_s2_reg/P0000_reg_syn_2 , \core_eu_es_sht_es_reg_SBr_reg[0]/P0001 , \core_eu_es_sht_es_reg_SBr_reg[1]/P0001 , \core_eu_es_sht_es_reg_SBr_reg[2]/P0001 , \core_eu_es_sht_es_reg_SBr_reg[3]/P0001 , \core_eu_es_sht_es_reg_SBr_reg[4]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[0]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[1]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[2]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[3]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[4]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001 , \emc_DMDoe_reg/NET0131 , \emc_DMDreg_reg[0]/P0001 , \emc_DMDreg_reg[10]/P0001 , \emc_DMDreg_reg[11]/P0001 , \emc_DMDreg_reg[12]/P0001 , \emc_DMDreg_reg[13]/P0001 , \emc_DMDreg_reg[14]/P0001 , \emc_DMDreg_reg[15]/P0001 , \emc_DMDreg_reg[1]/P0001 , \emc_DMDreg_reg[2]/P0001 , \emc_DMDreg_reg[3]/P0001 , \emc_DMDreg_reg[4]/P0001 , \emc_DMDreg_reg[5]/P0001 , \emc_DMDreg_reg[6]/P0001 , \emc_DMDreg_reg[7]/P0001 , \emc_DMDreg_reg[8]/P0001 , \emc_DMDreg_reg[9]/P0001 , \emc_DMcst_reg/NET0131 , \emc_ECMA_reg[0]/P0001 , \emc_ECMA_reg[10]/P0001 , \emc_ECMA_reg[11]/P0001 , \emc_ECMA_reg[12]/P0001 , \emc_ECMA_reg[1]/P0001 , \emc_ECMA_reg[2]/P0001 , \emc_ECMA_reg[3]/P0001 , \emc_ECMA_reg[4]/P0001 , \emc_ECMA_reg[5]/P0001 , \emc_ECMA_reg[6]/P0001 , \emc_ECMA_reg[7]/P0001 , \emc_ECMA_reg[8]/P0001 , \emc_ECMA_reg[9]/P0001 , \emc_ECMDreg_reg[0]/P0001 , \emc_ECMDreg_reg[10]/P0001 , \emc_ECMDreg_reg[11]/P0001 , \emc_ECMDreg_reg[12]/P0001 , \emc_ECMDreg_reg[13]/P0001 , \emc_ECMDreg_reg[14]/P0001 , \emc_ECMDreg_reg[15]/P0001 , \emc_ECMDreg_reg[16]/P0001 , \emc_ECMDreg_reg[17]/P0001 , \emc_ECMDreg_reg[18]/P0001 , \emc_ECMDreg_reg[19]/P0001 , \emc_ECMDreg_reg[1]/P0001 , \emc_ECMDreg_reg[20]/P0001 , \emc_ECMDreg_reg[21]/P0001 , \emc_ECMDreg_reg[22]/P0001 , \emc_ECMDreg_reg[23]/P0001 , \emc_ECMDreg_reg[2]/P0001 , \emc_ECMDreg_reg[3]/P0001 , \emc_ECMDreg_reg[4]/P0001 , \emc_ECMDreg_reg[5]/P0001 , \emc_ECMDreg_reg[6]/P0001 , \emc_ECMDreg_reg[7]/P0001 , \emc_ECMDreg_reg[8]/P0001 , \emc_ECMDreg_reg[9]/P0001 , \emc_ECMcs_reg/NET0131 , \emc_ECS_reg[0]/NET0131 , \emc_ECS_reg[1]/NET0131 , \emc_ECS_reg[2]/NET0131 , \emc_ECS_reg[3]/NET0131 , \emc_ED_oei_reg/P0001 , \emc_EXTC_Eg_syn_reg/P0001 , \emc_IOcst_reg/NET0131 , \emc_PMDoe_reg/NET0131 , \emc_PMDreg_reg[0]/P0001 , \emc_PMDreg_reg[10]/P0001 , \emc_PMDreg_reg[11]/P0001 , \emc_PMDreg_reg[12]/P0001 , \emc_PMDreg_reg[13]/P0001 , \emc_PMDreg_reg[14]/P0001 , \emc_PMDreg_reg[15]/P0001 , \emc_PMDreg_reg[1]/P0001 , \emc_PMDreg_reg[2]/P0001 , \emc_PMDreg_reg[3]/P0001 , \emc_PMDreg_reg[4]/P0001 , \emc_PMDreg_reg[5]/P0001 , \emc_PMDreg_reg[6]/P0001 , \emc_PMDreg_reg[7]/P0001 , \emc_PMDreg_reg[8]/P0001 , \emc_PMDreg_reg[9]/P0001 , \emc_PMcst_reg/NET0131 , \emc_RWcnt_reg[0]/P0001 , \emc_RWcnt_reg[1]/P0001 , \emc_RWcnt_reg[2]/P0001 , \emc_RWcnt_reg[3]/P0001 , \emc_RWcnt_reg[4]/P0001 , \emc_RWcnt_reg[5]/P0001 , \emc_WRn_h_reg/P0001 , \emc_WSCRext_reg_DO_reg[0]/NET0131 , \emc_WSCRext_reg_DO_reg[1]/NET0131 , \emc_WSCRext_reg_DO_reg[2]/NET0131 , \emc_WSCRext_reg_DO_reg[3]/NET0131 , \emc_WSCRext_reg_DO_reg[4]/NET0131 , \emc_WSCRext_reg_DO_reg[5]/NET0131 , \emc_WSCRext_reg_DO_reg[6]/NET0131 , \emc_WSCRext_reg_DO_reg[7]/NET0131 , \emc_WSCRreg_DO_reg[0]/NET0131 , \emc_WSCRreg_DO_reg[10]/NET0131 , \emc_WSCRreg_DO_reg[11]/NET0131 , \emc_WSCRreg_DO_reg[12]/NET0131 , \emc_WSCRreg_DO_reg[13]/NET0131 , \emc_WSCRreg_DO_reg[14]/NET0131 , \emc_WSCRreg_DO_reg[1]/NET0131 , \emc_WSCRreg_DO_reg[2]/NET0131 , \emc_WSCRreg_DO_reg[3]/NET0131 , \emc_WSCRreg_DO_reg[4]/NET0131 , \emc_WSCRreg_DO_reg[5]/NET0131 , \emc_WSCRreg_DO_reg[6]/NET0131 , \emc_WSCRreg_DO_reg[7]/NET0131 , \emc_WSCRreg_DO_reg[8]/NET0131 , \emc_WSCRreg_DO_reg[9]/NET0131 , \emc_eRDY_reg/NET0131 , \emc_selDMDi_reg/P0001 , \emc_selPMDi_reg/P0001 , \idma_CM_oe_reg/P0001 , \idma_CMo_oe0_reg/P0001 , \idma_CMo_oe1_reg/P0001 , \idma_CMo_oe2_reg/P0001 , \idma_CMo_oe3_reg/P0001 , \idma_CMo_oe4_reg/P0001 , \idma_CMo_oe5_reg/P0001 , \idma_CMo_oe6_reg/P0001 , \idma_CMo_oe7_reg/P0001 , \idma_DCTL_reg[0]/NET0131 , \idma_DCTL_reg[10]/NET0131 , \idma_DCTL_reg[11]/NET0131 , \idma_DCTL_reg[12]/NET0131 , \idma_DCTL_reg[13]/NET0131 , \idma_DCTL_reg[14]/NET0131 , \idma_DCTL_reg[1]/NET0131 , \idma_DCTL_reg[2]/NET0131 , \idma_DCTL_reg[3]/NET0131 , \idma_DCTL_reg[4]/NET0131 , \idma_DCTL_reg[5]/NET0131 , \idma_DCTL_reg[6]/NET0131 , \idma_DCTL_reg[7]/NET0131 , \idma_DCTL_reg[8]/NET0131 , \idma_DCTL_reg[9]/NET0131 , \idma_DOVL_reg[0]/NET0131 , \idma_DOVL_reg[10]/NET0131 , \idma_DOVL_reg[11]/NET0131 , \idma_DOVL_reg[1]/NET0131 , \idma_DOVL_reg[2]/NET0131 , \idma_DOVL_reg[3]/NET0131 , \idma_DOVL_reg[4]/NET0131 , \idma_DOVL_reg[5]/NET0131 , \idma_DOVL_reg[6]/NET0131 , \idma_DOVL_reg[7]/NET0131 , \idma_DOVL_reg[8]/NET0131 , \idma_DOVL_reg[9]/NET0131 , \idma_DSreq_reg/NET0131 , \idma_DTMP_H_reg[0]/P0001 , \idma_DTMP_H_reg[10]/P0001 , \idma_DTMP_H_reg[11]/P0001 , \idma_DTMP_H_reg[12]/P0001 , \idma_DTMP_H_reg[13]/P0001 , \idma_DTMP_H_reg[14]/P0001 , \idma_DTMP_H_reg[15]/P0001 , \idma_DTMP_H_reg[1]/P0001 , \idma_DTMP_H_reg[2]/P0001 , \idma_DTMP_H_reg[3]/P0001 , \idma_DTMP_H_reg[4]/P0001 , \idma_DTMP_H_reg[5]/P0001 , \idma_DTMP_H_reg[6]/P0001 , \idma_DTMP_H_reg[7]/P0001 , \idma_DTMP_H_reg[8]/P0001 , \idma_DTMP_H_reg[9]/P0001 , \idma_DTMP_L_reg[0]/P0001 , \idma_DTMP_L_reg[1]/P0001 , \idma_DTMP_L_reg[2]/P0001 , \idma_DTMP_L_reg[3]/P0001 , \idma_DTMP_L_reg[4]/P0001 , \idma_DTMP_L_reg[5]/P0001 , \idma_DTMP_L_reg[6]/P0001 , \idma_DTMP_L_reg[7]/P0001 , \idma_IADi_reg[0]/P0001 , \idma_IADi_reg[10]/P0001 , \idma_IADi_reg[11]/P0001 , \idma_IADi_reg[12]/P0001 , \idma_IADi_reg[13]/P0001 , \idma_IADi_reg[14]/P0001 , \idma_IADi_reg[15]/P0001 , \idma_IADi_reg[1]/P0001 , \idma_IADi_reg[2]/P0001 , \idma_IADi_reg[3]/P0001 , \idma_IADi_reg[4]/P0001 , \idma_IADi_reg[5]/P0001 , \idma_IADi_reg[6]/P0001 , \idma_IADi_reg[7]/P0001 , \idma_IADi_reg[8]/P0001 , \idma_IADi_reg[9]/P0001 , \idma_IAL_reg/P0001 , \idma_IDMA_boot_reg/NET0131_reg_syn_10 , \idma_IDMA_boot_reg/NET0131_reg_syn_2 , \idma_IDMA_boot_reg/NET0131_reg_syn_8 , \idma_IRDn_reg/P0001 , \idma_ISn_reg/P0001 , \idma_IWRn_reg/P0001 , \idma_PCrd_1st_reg/NET0131 , \idma_PM_1st_reg/NET0131 , \idma_RDCMD_d1_reg/P0001 , \idma_RDCMD_reg/P0001 , \idma_RDcnt_reg[0]/NET0131 , \idma_RDcnt_reg[1]/NET0131 , \idma_RDcnt_reg[2]/NET0131 , \idma_RDcyc_reg/NET0131 , \idma_WRCMD_d1_reg/P0001 , \idma_WRCMD_reg/P0001 , \idma_WRcnt_reg[0]/NET0131 , \idma_WRcnt_reg[1]/NET0131 , \idma_WRcnt_reg[2]/NET0131 , \idma_WRcyc_reg/NET0131 , \idma_WRtrue_reg/NET0131 , \memc_DM_oe_reg/P0001 , \memc_DMo_oe0_reg/P0001 , \memc_DMo_oe1_reg/P0001 , \memc_DMo_oe2_reg/P0001 , \memc_DMo_oe3_reg/P0001 , \memc_DMo_oe4_reg/P0001 , \memc_DMo_oe5_reg/P0001 , \memc_DMo_oe6_reg/P0001 , \memc_DMo_oe7_reg/P0001 , \memc_Dread_E_reg/NET0131 , \memc_Dwrite_C_reg/NET0131 , \memc_Dwrite_E_reg/NET0131 , \memc_EXTC_E_reg/NET0131 , \memc_EXTC_Eg_reg/NET0131_reg_syn_10 , \memc_EXTC_Eg_reg/NET0131_reg_syn_2 , \memc_EXTC_Eg_reg/NET0131_reg_syn_8 , \memc_IOcmd_E_reg/NET0131 , \memc_LDaST_Eg_reg/NET0131 , \memc_MMR_web_reg/NET0131 , \memc_PMo_oe0_reg/P0001 , \memc_PMo_oe1_reg/P0001 , \memc_PMo_oe2_reg/P0001 , \memc_PMo_oe3_reg/P0001 , \memc_PMo_oe4_reg/P0001 , \memc_PMo_oe5_reg/P0001 , \memc_PMo_oe6_reg/P0001 , \memc_PMo_oe7_reg/P0001 , \memc_Pread_E_reg/NET0131 , \memc_Pwrite_C_reg/NET0131 , \memc_Pwrite_E_reg/NET0131 , \memc_STI_Cg_reg/NET0131 , \memc_accDM_E_reg/NET0131 , \memc_accPM_E_reg/NET0131 , \memc_ldSREG_E_reg/NET0131 , \memc_selMIO_E_reg/P0001 , \memc_usysr_DO_reg[0]/NET0131 , \memc_usysr_DO_reg[10]/NET0131 , \memc_usysr_DO_reg[11]/NET0131 , \memc_usysr_DO_reg[12]/NET0131 , \memc_usysr_DO_reg[13]/NET0131 , \memc_usysr_DO_reg[14]/NET0131 , \memc_usysr_DO_reg[15]/NET0131 , \memc_usysr_DO_reg[1]/NET0131 , \memc_usysr_DO_reg[2]/NET0131 , \memc_usysr_DO_reg[3]/NET0131 , \memc_usysr_DO_reg[4]/NET0131 , \memc_usysr_DO_reg[5]/NET0131 , \memc_usysr_DO_reg[6]/NET0131 , \memc_usysr_DO_reg[7]/NET0131 , \memc_usysr_DO_reg[8]/NET0131 , \memc_usysr_DO_reg[9]/NET0131 , \pio_PINT_reg[0]/NET0131 , \pio_PINT_reg[10]/NET0131 , \pio_PINT_reg[11]/NET0131 , \pio_PINT_reg[1]/NET0131 , \pio_PINT_reg[2]/NET0131 , \pio_PINT_reg[3]/NET0131 , \pio_PINT_reg[4]/NET0131 , \pio_PINT_reg[5]/NET0131 , \pio_PINT_reg[6]/NET0131 , \pio_PINT_reg[7]/NET0131 , \pio_PINT_reg[8]/NET0131 , \pio_PINT_reg[9]/NET0131 , \pio_PIO_IN_P_reg[0]/P0001 , \pio_PIO_IN_P_reg[10]/P0001 , \pio_PIO_IN_P_reg[11]/P0001 , \pio_PIO_IN_P_reg[1]/P0001 , \pio_PIO_IN_P_reg[2]/P0001 , \pio_PIO_IN_P_reg[3]/P0001 , \pio_PIO_IN_P_reg[4]/P0001 , \pio_PIO_IN_P_reg[5]/P0001 , \pio_PIO_IN_P_reg[6]/P0001 , \pio_PIO_IN_P_reg[7]/P0001 , \pio_PIO_IN_P_reg[8]/P0001 , \pio_PIO_IN_P_reg[9]/P0001 , \pio_PIO_RES_OUT_reg[0]/P0001 , \pio_PIO_RES_OUT_reg[10]/P0001 , \pio_PIO_RES_OUT_reg[11]/P0001 , \pio_PIO_RES_OUT_reg[1]/P0001 , \pio_PIO_RES_OUT_reg[2]/P0001 , \pio_PIO_RES_OUT_reg[3]/P0001 , \pio_PIO_RES_OUT_reg[4]/P0001 , \pio_PIO_RES_OUT_reg[5]/P0001 , \pio_PIO_RES_OUT_reg[6]/P0001 , \pio_PIO_RES_OUT_reg[7]/P0001 , \pio_PIO_RES_OUT_reg[8]/P0001 , \pio_PIO_RES_OUT_reg[9]/P0001 , \pio_PIO_RES_reg[0]/NET0131 , \pio_PIO_RES_reg[10]/NET0131 , \pio_PIO_RES_reg[11]/NET0131 , \pio_PIO_RES_reg[1]/NET0131 , \pio_PIO_RES_reg[2]/NET0131 , \pio_PIO_RES_reg[3]/NET0131 , \pio_PIO_RES_reg[4]/NET0131 , \pio_PIO_RES_reg[5]/NET0131 , \pio_PIO_RES_reg[6]/NET0131 , \pio_PIO_RES_reg[7]/NET0131 , \pio_PIO_RES_reg[8]/NET0131 , \pio_PIO_RES_reg[9]/NET0131 , \pio_pmask_reg_DO_reg[0]/NET0131 , \pio_pmask_reg_DO_reg[10]/NET0131 , \pio_pmask_reg_DO_reg[11]/NET0131 , \pio_pmask_reg_DO_reg[1]/NET0131 , \pio_pmask_reg_DO_reg[2]/NET0131 , \pio_pmask_reg_DO_reg[3]/NET0131 , \pio_pmask_reg_DO_reg[4]/NET0131 , \pio_pmask_reg_DO_reg[5]/NET0131 , \pio_pmask_reg_DO_reg[6]/NET0131 , \pio_pmask_reg_DO_reg[7]/NET0131 , \pio_pmask_reg_DO_reg[8]/NET0131 , \pio_pmask_reg_DO_reg[9]/NET0131 , \regout_STD_C_reg[0]/P0001 , \regout_STD_C_reg[10]/P0001 , \regout_STD_C_reg[11]/P0001 , \regout_STD_C_reg[12]/P0001 , \regout_STD_C_reg[13]/P0001 , \regout_STD_C_reg[14]/P0001 , \regout_STD_C_reg[15]/P0001 , \regout_STD_C_reg[1]/P0001 , \regout_STD_C_reg[2]/P0001 , \regout_STD_C_reg[3]/P0001 , \regout_STD_C_reg[4]/P0001 , \regout_STD_C_reg[5]/P0001 , \regout_STD_C_reg[6]/P0001 , \regout_STD_C_reg[7]/P0001 , \regout_STD_C_reg[8]/P0001 , \regout_STD_C_reg[9]/P0001 , \sice_CLR_I_reg/NET0131 , \sice_CLR_M_reg/NET0131 , \sice_CMRW_reg/NET0131 , \sice_DBR1_reg[0]/P0001 , \sice_DBR1_reg[10]/P0001 , \sice_DBR1_reg[11]/P0001 , \sice_DBR1_reg[12]/P0001 , \sice_DBR1_reg[13]/P0001 , \sice_DBR1_reg[14]/P0001 , \sice_DBR1_reg[15]/P0001 , \sice_DBR1_reg[16]/P0001 , \sice_DBR1_reg[17]/P0001 , \sice_DBR1_reg[18]/P0001 , \sice_DBR1_reg[1]/P0001 , \sice_DBR1_reg[2]/P0001 , \sice_DBR1_reg[3]/P0001 , \sice_DBR1_reg[4]/P0001 , \sice_DBR1_reg[5]/P0001 , \sice_DBR1_reg[6]/P0001 , \sice_DBR1_reg[7]/P0001 , \sice_DBR1_reg[8]/P0001 , \sice_DBR1_reg[9]/P0001 , \sice_DBR2_reg[0]/P0001 , \sice_DBR2_reg[10]/P0001 , \sice_DBR2_reg[11]/P0001 , \sice_DBR2_reg[12]/P0001 , \sice_DBR2_reg[13]/P0001 , \sice_DBR2_reg[14]/P0001 , \sice_DBR2_reg[15]/P0001 , \sice_DBR2_reg[16]/P0001 , \sice_DBR2_reg[17]/P0001 , \sice_DBR2_reg[18]/P0001 , \sice_DBR2_reg[1]/P0001 , \sice_DBR2_reg[2]/P0001 , \sice_DBR2_reg[3]/P0001 , \sice_DBR2_reg[4]/P0001 , \sice_DBR2_reg[5]/P0001 , \sice_DBR2_reg[6]/P0001 , \sice_DBR2_reg[7]/P0001 , \sice_DBR2_reg[8]/P0001 , \sice_DBR2_reg[9]/P0001 , \sice_DMR1_reg[0]/NET0131 , \sice_DMR1_reg[10]/NET0131 , \sice_DMR1_reg[11]/NET0131 , \sice_DMR1_reg[12]/NET0131 , \sice_DMR1_reg[13]/NET0131 , \sice_DMR1_reg[14]/NET0131 , \sice_DMR1_reg[15]/NET0131 , \sice_DMR1_reg[16]/NET0131 , \sice_DMR1_reg[17]/NET0131 , \sice_DMR1_reg[1]/NET0131 , \sice_DMR1_reg[2]/NET0131 , \sice_DMR1_reg[3]/NET0131 , \sice_DMR1_reg[4]/NET0131 , \sice_DMR1_reg[5]/NET0131 , \sice_DMR1_reg[6]/NET0131 , \sice_DMR1_reg[7]/NET0131 , \sice_DMR1_reg[8]/NET0131 , \sice_DMR1_reg[9]/NET0131 , \sice_DMR2_reg[0]/NET0131 , \sice_DMR2_reg[10]/NET0131 , \sice_DMR2_reg[11]/NET0131 , \sice_DMR2_reg[12]/NET0131 , \sice_DMR2_reg[13]/NET0131 , \sice_DMR2_reg[14]/NET0131 , \sice_DMR2_reg[15]/NET0131 , \sice_DMR2_reg[16]/NET0131 , \sice_DMR2_reg[17]/NET0131 , \sice_DMR2_reg[1]/NET0131 , \sice_DMR2_reg[2]/NET0131 , \sice_DMR2_reg[3]/NET0131 , \sice_DMR2_reg[4]/NET0131 , \sice_DMR2_reg[5]/NET0131 , \sice_DMR2_reg[6]/NET0131 , \sice_DMR2_reg[7]/NET0131 , \sice_DMR2_reg[8]/NET0131 , \sice_DMR2_reg[9]/NET0131 , \sice_GOICE_1_reg/NET0131 , \sice_GOICE_2_reg/NET0131 , \sice_GOICE_s1_reg/NET0131 , \sice_GOICE_syn_reg/P0001 , \sice_GO_NX_reg/NET0131 , \sice_GO_NXi_reg/NET0131 , \sice_HALT_E_reg/P0001 , \sice_IAR_reg[0]/NET0131 , \sice_IAR_reg[1]/NET0131 , \sice_IAR_reg[2]/NET0131 , \sice_IAR_reg[3]/NET0131 , \sice_IBR1_reg[0]/P0001 , \sice_IBR1_reg[10]/P0001 , \sice_IBR1_reg[11]/P0001 , \sice_IBR1_reg[12]/P0001 , \sice_IBR1_reg[13]/P0001 , \sice_IBR1_reg[14]/P0001 , \sice_IBR1_reg[15]/P0001 , \sice_IBR1_reg[16]/P0001 , \sice_IBR1_reg[17]/P0001 , \sice_IBR1_reg[1]/P0001 , \sice_IBR1_reg[2]/P0001 , \sice_IBR1_reg[3]/P0001 , \sice_IBR1_reg[4]/P0001 , \sice_IBR1_reg[5]/P0001 , \sice_IBR1_reg[6]/P0001 , \sice_IBR1_reg[7]/P0001 , \sice_IBR1_reg[8]/P0001 , \sice_IBR1_reg[9]/P0001 , \sice_IBR2_reg[0]/P0001 , \sice_IBR2_reg[10]/P0001 , \sice_IBR2_reg[11]/P0001 , \sice_IBR2_reg[12]/P0001 , \sice_IBR2_reg[13]/P0001 , \sice_IBR2_reg[14]/P0001 , \sice_IBR2_reg[15]/P0001 , \sice_IBR2_reg[16]/P0001 , \sice_IBR2_reg[17]/P0001 , \sice_IBR2_reg[1]/P0001 , \sice_IBR2_reg[2]/P0001 , \sice_IBR2_reg[3]/P0001 , \sice_IBR2_reg[4]/P0001 , \sice_IBR2_reg[5]/P0001 , \sice_IBR2_reg[6]/P0001 , \sice_IBR2_reg[7]/P0001 , \sice_IBR2_reg[8]/P0001 , \sice_IBR2_reg[9]/P0001 , \sice_ICS_reg[0]/NET0131 , \sice_ICS_reg[1]/NET0131 , \sice_ICS_reg[2]/NET0131 , \sice_ICYC_clr_reg/NET0131 , \sice_ICYC_en_reg/NET0131 , \sice_ICYC_en_syn_reg/P0001 , \sice_ICYC_reg[0]/NET0131 , \sice_ICYC_reg[10]/NET0131 , \sice_ICYC_reg[11]/NET0131 , \sice_ICYC_reg[12]/NET0131 , \sice_ICYC_reg[13]/NET0131 , \sice_ICYC_reg[14]/NET0131 , \sice_ICYC_reg[15]/NET0131 , \sice_ICYC_reg[16]/NET0131 , \sice_ICYC_reg[17]/NET0131 , \sice_ICYC_reg[18]/NET0131 , \sice_ICYC_reg[19]/NET0131 , \sice_ICYC_reg[1]/NET0131 , \sice_ICYC_reg[20]/NET0131 , \sice_ICYC_reg[21]/NET0131 , \sice_ICYC_reg[22]/NET0131 , \sice_ICYC_reg[23]/NET0131 , \sice_ICYC_reg[2]/NET0131 , \sice_ICYC_reg[3]/NET0131 , \sice_ICYC_reg[4]/NET0131 , \sice_ICYC_reg[5]/NET0131 , \sice_ICYC_reg[6]/NET0131 , \sice_ICYC_reg[7]/NET0131 , \sice_ICYC_reg[8]/NET0131 , \sice_ICYC_reg[9]/NET0131 , \sice_IDONE_reg/NET0131 , \sice_IIRC_reg[0]/NET0131 , \sice_IIRC_reg[10]/NET0131 , \sice_IIRC_reg[11]/NET0131 , \sice_IIRC_reg[12]/NET0131 , \sice_IIRC_reg[13]/NET0131 , \sice_IIRC_reg[14]/NET0131 , \sice_IIRC_reg[15]/NET0131 , \sice_IIRC_reg[16]/NET0131 , \sice_IIRC_reg[17]/NET0131 , \sice_IIRC_reg[18]/NET0131 , \sice_IIRC_reg[19]/NET0131 , \sice_IIRC_reg[1]/NET0131 , \sice_IIRC_reg[20]/NET0131 , \sice_IIRC_reg[21]/NET0131 , \sice_IIRC_reg[22]/NET0131 , \sice_IIRC_reg[23]/NET0131 , \sice_IIRC_reg[2]/NET0131 , \sice_IIRC_reg[3]/NET0131 , \sice_IIRC_reg[4]/NET0131 , \sice_IIRC_reg[5]/NET0131 , \sice_IIRC_reg[6]/NET0131 , \sice_IIRC_reg[7]/NET0131 , \sice_IIRC_reg[8]/NET0131 , \sice_IIRC_reg[9]/NET0131 , \sice_IMR1_reg[0]/NET0131 , \sice_IMR1_reg[10]/NET0131 , \sice_IMR1_reg[11]/NET0131 , \sice_IMR1_reg[12]/NET0131 , \sice_IMR1_reg[13]/NET0131 , \sice_IMR1_reg[14]/NET0131 , \sice_IMR1_reg[15]/NET0131 , \sice_IMR1_reg[16]/NET0131 , \sice_IMR1_reg[17]/NET0131 , \sice_IMR1_reg[1]/NET0131 , \sice_IMR1_reg[2]/NET0131 , \sice_IMR1_reg[3]/NET0131 , \sice_IMR1_reg[4]/NET0131 , \sice_IMR1_reg[5]/NET0131 , \sice_IMR1_reg[6]/NET0131 , \sice_IMR1_reg[7]/NET0131 , \sice_IMR1_reg[8]/NET0131 , \sice_IMR1_reg[9]/NET0131 , \sice_IMR2_reg[0]/NET0131 , \sice_IMR2_reg[10]/NET0131 , \sice_IMR2_reg[11]/NET0131 , \sice_IMR2_reg[12]/NET0131 , \sice_IMR2_reg[13]/NET0131 , \sice_IMR2_reg[14]/NET0131 , \sice_IMR2_reg[15]/NET0131 , \sice_IMR2_reg[16]/NET0131 , \sice_IMR2_reg[17]/NET0131 , \sice_IMR2_reg[1]/NET0131 , \sice_IMR2_reg[2]/NET0131 , \sice_IMR2_reg[3]/NET0131 , \sice_IMR2_reg[4]/NET0131 , \sice_IMR2_reg[5]/NET0131 , \sice_IMR2_reg[6]/NET0131 , \sice_IMR2_reg[7]/NET0131 , \sice_IMR2_reg[8]/NET0131 , \sice_IMR2_reg[9]/NET0131 , \sice_IRR_reg[0]/P0001 , \sice_IRR_reg[10]/P0001 , \sice_IRR_reg[11]/P0001 , \sice_IRR_reg[12]/P0001 , \sice_IRR_reg[13]/P0001 , \sice_IRR_reg[1]/P0001 , \sice_IRR_reg[2]/P0001 , \sice_IRR_reg[3]/P0001 , \sice_IRR_reg[4]/P0001 , \sice_IRR_reg[5]/P0001 , \sice_IRR_reg[6]/P0001 , \sice_IRR_reg[7]/P0001 , \sice_IRR_reg[8]/P0001 , \sice_IRR_reg[9]/P0001 , \sice_IRST_reg/NET0131 , \sice_IRST_syn_reg/P0001 , \sice_ITR_reg[0]/NET0131 , \sice_ITR_reg[1]/NET0131 , \sice_ITR_reg[2]/NET0131 , \sice_OE_reg/P0001 , \sice_RCS_reg[0]/NET0131 , \sice_RCS_reg[1]/NET0131 , \sice_RST_req_reg/NET0131 , \sice_SPC_reg[0]/P0001 , \sice_SPC_reg[10]/P0001 , \sice_SPC_reg[11]/P0001 , \sice_SPC_reg[12]/P0001 , \sice_SPC_reg[13]/P0001 , \sice_SPC_reg[14]/P0001 , \sice_SPC_reg[15]/P0001 , \sice_SPC_reg[16]/P0001 , \sice_SPC_reg[17]/P0001 , \sice_SPC_reg[18]/P0001 , \sice_SPC_reg[19]/P0001 , \sice_SPC_reg[1]/P0001 , \sice_SPC_reg[20]/P0001 , \sice_SPC_reg[21]/P0001 , \sice_SPC_reg[22]/P0001 , \sice_SPC_reg[23]/P0001 , \sice_SPC_reg[2]/P0001 , \sice_SPC_reg[3]/P0001 , \sice_SPC_reg[4]/P0001 , \sice_SPC_reg[5]/P0001 , \sice_SPC_reg[6]/P0001 , \sice_SPC_reg[7]/P0001 , \sice_SPC_reg[8]/P0001 , \sice_SPC_reg[9]/P0001 , \sice_UpdDR_sd1_reg/P0001 , \sice_UpdDR_sd2_reg/P0001 , \sice_idr0_reg_DO_reg[0]/P0001 , \sice_idr0_reg_DO_reg[10]/P0001 , \sice_idr0_reg_DO_reg[11]/P0001 , \sice_idr0_reg_DO_reg[1]/P0001 , \sice_idr0_reg_DO_reg[2]/P0001 , \sice_idr0_reg_DO_reg[3]/P0001 , \sice_idr0_reg_DO_reg[4]/P0001 , \sice_idr0_reg_DO_reg[5]/P0001 , \sice_idr0_reg_DO_reg[6]/P0001 , \sice_idr0_reg_DO_reg[7]/P0001 , \sice_idr0_reg_DO_reg[8]/P0001 , \sice_idr0_reg_DO_reg[9]/P0001 , \sice_idr1_reg_DO_reg[0]/P0001 , \sice_idr1_reg_DO_reg[10]/P0001 , \sice_idr1_reg_DO_reg[11]/P0001 , \sice_idr1_reg_DO_reg[1]/P0001 , \sice_idr1_reg_DO_reg[2]/P0001 , \sice_idr1_reg_DO_reg[3]/P0001 , \sice_idr1_reg_DO_reg[4]/P0001 , \sice_idr1_reg_DO_reg[5]/P0001 , \sice_idr1_reg_DO_reg[6]/P0001 , \sice_idr1_reg_DO_reg[7]/P0001 , \sice_idr1_reg_DO_reg[8]/P0001 , \sice_idr1_reg_DO_reg[9]/P0001 , \sport0_cfg_FSi_cnt_reg[0]/NET0131 , \sport0_cfg_FSi_cnt_reg[10]/NET0131 , \sport0_cfg_FSi_cnt_reg[11]/NET0131 , \sport0_cfg_FSi_cnt_reg[12]/NET0131 , \sport0_cfg_FSi_cnt_reg[13]/NET0131 , \sport0_cfg_FSi_cnt_reg[14]/NET0131 , \sport0_cfg_FSi_cnt_reg[15]/NET0131 , \sport0_cfg_FSi_cnt_reg[1]/NET0131 , \sport0_cfg_FSi_cnt_reg[2]/NET0131 , \sport0_cfg_FSi_cnt_reg[3]/NET0131 , \sport0_cfg_FSi_cnt_reg[4]/NET0131 , \sport0_cfg_FSi_cnt_reg[5]/NET0131 , \sport0_cfg_FSi_cnt_reg[6]/NET0131 , \sport0_cfg_FSi_cnt_reg[7]/NET0131 , \sport0_cfg_FSi_cnt_reg[8]/NET0131 , \sport0_cfg_FSi_cnt_reg[9]/NET0131 , \sport0_cfg_FSi_reg/NET0131 , \sport0_cfg_RFSg_d1_reg/NET0131 , \sport0_cfg_RFSg_d2_reg/NET0131 , \sport0_cfg_RFSg_d3_reg/NET0131 , \sport0_cfg_RFSgi_d_reg/NET0131 , \sport0_cfg_SCLKi_cnt_reg[0]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[10]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[11]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[12]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[13]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[14]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[15]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[1]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[2]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[3]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[4]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[5]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[6]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[7]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[8]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[9]/NET0131 , \sport0_cfg_SCLKi_h_reg/NET0131 , \sport0_cfg_SP_ENg_D1_reg/P0001 , \sport0_cfg_SP_ENg_reg/NET0131 , \sport0_cfg_TFSg_d1_reg/NET0131 , \sport0_cfg_TFSg_d2_reg/NET0131 , \sport0_cfg_TFSg_d3_reg/NET0131 , \sport0_cfg_TFSgi_d_reg/NET0131 , \sport0_regs_AUTO_a_reg[12]/NET0131 , \sport0_regs_AUTO_a_reg[13]/NET0131 , \sport0_regs_AUTO_a_reg[14]/NET0131 , \sport0_regs_AUTO_a_reg[15]/NET0131 , \sport0_regs_AUTOreg_DO_reg[0]/NET0131 , \sport0_regs_AUTOreg_DO_reg[10]/NET0131 , \sport0_regs_AUTOreg_DO_reg[11]/NET0131 , \sport0_regs_AUTOreg_DO_reg[1]/NET0131 , \sport0_regs_AUTOreg_DO_reg[2]/NET0131 , \sport0_regs_AUTOreg_DO_reg[3]/NET0131 , \sport0_regs_AUTOreg_DO_reg[4]/NET0131 , \sport0_regs_AUTOreg_DO_reg[5]/NET0131 , \sport0_regs_AUTOreg_DO_reg[6]/NET0131 , \sport0_regs_AUTOreg_DO_reg[7]/NET0131 , \sport0_regs_AUTOreg_DO_reg[8]/NET0131 , \sport0_regs_AUTOreg_DO_reg[9]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[0]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[10]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[11]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[12]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[13]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[14]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[15]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[1]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[2]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[3]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[4]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[5]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[6]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[7]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[8]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[9]/NET0131 , \sport0_regs_MWORDreg_DO_reg[0]/NET0131 , \sport0_regs_MWORDreg_DO_reg[10]/NET0131 , \sport0_regs_MWORDreg_DO_reg[1]/NET0131 , \sport0_regs_MWORDreg_DO_reg[2]/NET0131 , \sport0_regs_MWORDreg_DO_reg[3]/NET0131 , \sport0_regs_MWORDreg_DO_reg[4]/NET0131 , \sport0_regs_MWORDreg_DO_reg[5]/NET0131 , \sport0_regs_MWORDreg_DO_reg[6]/NET0131 , \sport0_regs_MWORDreg_DO_reg[7]/NET0131 , \sport0_regs_MWORDreg_DO_reg[8]/NET0131 , \sport0_regs_MWORDreg_DO_reg[9]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 , \sport0_regs_SCTLreg_DO_reg[0]/NET0131 , \sport0_regs_SCTLreg_DO_reg[10]/NET0131 , \sport0_regs_SCTLreg_DO_reg[11]/NET0131 , \sport0_regs_SCTLreg_DO_reg[12]/NET0131 , \sport0_regs_SCTLreg_DO_reg[13]/NET0131 , \sport0_regs_SCTLreg_DO_reg[15]/NET0131 , \sport0_regs_SCTLreg_DO_reg[1]/NET0131 , \sport0_regs_SCTLreg_DO_reg[2]/NET0131 , \sport0_regs_SCTLreg_DO_reg[3]/NET0131 , \sport0_regs_SCTLreg_DO_reg[4]/NET0131 , \sport0_regs_SCTLreg_DO_reg[5]/NET0131 , \sport0_regs_SCTLreg_DO_reg[6]/NET0131 , \sport0_regs_SCTLreg_DO_reg[7]/NET0131 , \sport0_rxctl_Bcnt_reg[0]/NET0131 , \sport0_rxctl_Bcnt_reg[1]/NET0131 , \sport0_rxctl_Bcnt_reg[2]/NET0131 , \sport0_rxctl_Bcnt_reg[3]/NET0131 , \sport0_rxctl_Bcnt_reg[4]/NET0131 , \sport0_rxctl_ISRa_reg/P0001 , \sport0_rxctl_LMcnt_reg[0]/NET0131 , \sport0_rxctl_LMcnt_reg[1]/NET0131 , \sport0_rxctl_LMcnt_reg[2]/NET0131 , \sport0_rxctl_LMcnt_reg[3]/NET0131 , \sport0_rxctl_LMcnt_reg[4]/NET0131 , \sport0_rxctl_RCS_reg[0]/NET0131 , \sport0_rxctl_RCS_reg[1]/NET0131 , \sport0_rxctl_RCS_reg[2]/NET0131 , \sport0_rxctl_RSreq_reg/NET0131 , \sport0_rxctl_RXSHT_reg[0]/P0001 , \sport0_rxctl_RXSHT_reg[10]/P0001 , \sport0_rxctl_RXSHT_reg[11]/P0001 , \sport0_rxctl_RXSHT_reg[12]/P0001 , \sport0_rxctl_RXSHT_reg[13]/P0001 , \sport0_rxctl_RXSHT_reg[14]/P0001 , \sport0_rxctl_RXSHT_reg[15]/P0001 , \sport0_rxctl_RXSHT_reg[1]/P0001 , \sport0_rxctl_RXSHT_reg[2]/P0001 , \sport0_rxctl_RXSHT_reg[3]/P0001 , \sport0_rxctl_RXSHT_reg[4]/P0001 , \sport0_rxctl_RXSHT_reg[5]/P0001 , \sport0_rxctl_RXSHT_reg[6]/P0001 , \sport0_rxctl_RXSHT_reg[7]/P0001 , \sport0_rxctl_RXSHT_reg[8]/P0001 , \sport0_rxctl_RXSHT_reg[9]/P0001 , \sport0_rxctl_RX_reg[0]/P0001 , \sport0_rxctl_RX_reg[10]/P0001 , \sport0_rxctl_RX_reg[11]/P0001 , \sport0_rxctl_RX_reg[12]/P0001 , \sport0_rxctl_RX_reg[13]/P0001 , \sport0_rxctl_RX_reg[14]/P0001 , \sport0_rxctl_RX_reg[15]/P0001 , \sport0_rxctl_RX_reg[1]/P0001 , \sport0_rxctl_RX_reg[2]/P0001 , \sport0_rxctl_RX_reg[3]/P0001 , \sport0_rxctl_RX_reg[4]/P0001 , \sport0_rxctl_RX_reg[5]/P0001 , \sport0_rxctl_RX_reg[6]/P0001 , \sport0_rxctl_RX_reg[7]/P0001 , \sport0_rxctl_RX_reg[8]/P0001 , \sport0_rxctl_RX_reg[9]/P0001 , \sport0_rxctl_SLOT1_EXT_reg[2]/NET0131 , \sport0_rxctl_SLOT1_EXT_reg[3]/NET0131 , \sport0_rxctl_TAG_SLOT_reg/P0001 , \sport0_rxctl_Wcnt_reg[0]/NET0131 , \sport0_rxctl_Wcnt_reg[1]/NET0131 , \sport0_rxctl_Wcnt_reg[2]/NET0131 , \sport0_rxctl_Wcnt_reg[3]/NET0131 , \sport0_rxctl_Wcnt_reg[4]/NET0131 , \sport0_rxctl_Wcnt_reg[5]/NET0131 , \sport0_rxctl_Wcnt_reg[6]/NET0131 , \sport0_rxctl_Wcnt_reg[7]/NET0131 , \sport0_rxctl_a_sync1_reg/P0001 , \sport0_rxctl_a_sync2_reg/P0001 , \sport0_rxctl_ldRX_cmp_reg/P0001 , \sport0_rxctl_sht2nd_reg/P0001 , \sport0_txctl_Bcnt_reg[0]/NET0131 , \sport0_txctl_Bcnt_reg[1]/NET0131 , \sport0_txctl_Bcnt_reg[2]/NET0131 , \sport0_txctl_Bcnt_reg[3]/NET0131 , \sport0_txctl_Bcnt_reg[4]/NET0131 , \sport0_txctl_SP_EN_D1_reg/P0001 , \sport0_txctl_TCS_reg[0]/NET0131 , \sport0_txctl_TCS_reg[1]/NET0131 , \sport0_txctl_TCS_reg[2]/NET0131 , \sport0_txctl_TSreq_reg/NET0131 , \sport0_txctl_TSreqi_reg/NET0131 , \sport0_txctl_TXSHT_reg[0]/P0001 , \sport0_txctl_TXSHT_reg[10]/P0001 , \sport0_txctl_TXSHT_reg[11]/P0001 , \sport0_txctl_TXSHT_reg[12]/P0001 , \sport0_txctl_TXSHT_reg[13]/P0001 , \sport0_txctl_TXSHT_reg[14]/P0001 , \sport0_txctl_TXSHT_reg[15]/P0001 , \sport0_txctl_TXSHT_reg[1]/P0001 , \sport0_txctl_TXSHT_reg[2]/P0001 , \sport0_txctl_TXSHT_reg[3]/P0001 , \sport0_txctl_TXSHT_reg[4]/P0001 , \sport0_txctl_TXSHT_reg[5]/P0001 , \sport0_txctl_TXSHT_reg[6]/P0001 , \sport0_txctl_TXSHT_reg[7]/P0001 , \sport0_txctl_TXSHT_reg[8]/P0001 , \sport0_txctl_TXSHT_reg[9]/P0001 , \sport0_txctl_TX_reg[0]/P0001 , \sport0_txctl_TX_reg[10]/P0001 , \sport0_txctl_TX_reg[11]/P0001 , \sport0_txctl_TX_reg[12]/P0001 , \sport0_txctl_TX_reg[13]/P0001 , \sport0_txctl_TX_reg[14]/P0001 , \sport0_txctl_TX_reg[15]/P0001 , \sport0_txctl_TX_reg[1]/P0001 , \sport0_txctl_TX_reg[2]/P0001 , \sport0_txctl_TX_reg[3]/P0001 , \sport0_txctl_TX_reg[4]/P0001 , \sport0_txctl_TX_reg[5]/P0001 , \sport0_txctl_TX_reg[6]/P0001 , \sport0_txctl_TX_reg[7]/P0001 , \sport0_txctl_TX_reg[8]/P0001 , \sport0_txctl_TX_reg[9]/P0001 , \sport0_txctl_Wcnt_reg[0]/NET0131 , \sport0_txctl_Wcnt_reg[1]/NET0131 , \sport0_txctl_Wcnt_reg[2]/NET0131 , \sport0_txctl_Wcnt_reg[3]/NET0131 , \sport0_txctl_Wcnt_reg[4]/NET0131 , \sport0_txctl_Wcnt_reg[5]/NET0131 , \sport0_txctl_Wcnt_reg[6]/NET0131 , \sport0_txctl_Wcnt_reg[7]/NET0131 , \sport0_txctl_b_sync1_reg/P0001 , \sport0_txctl_c_sync1_reg/P0001 , \sport0_txctl_c_sync2_reg/P0001 , \sport0_txctl_ldTX_cmp_reg/P0001 , \sport1_cfg_FSi_cnt_reg[0]/NET0131 , \sport1_cfg_FSi_cnt_reg[10]/NET0131 , \sport1_cfg_FSi_cnt_reg[11]/NET0131 , \sport1_cfg_FSi_cnt_reg[12]/NET0131 , \sport1_cfg_FSi_cnt_reg[13]/NET0131 , \sport1_cfg_FSi_cnt_reg[14]/NET0131 , \sport1_cfg_FSi_cnt_reg[15]/NET0131 , \sport1_cfg_FSi_cnt_reg[1]/NET0131 , \sport1_cfg_FSi_cnt_reg[2]/NET0131 , \sport1_cfg_FSi_cnt_reg[3]/NET0131 , \sport1_cfg_FSi_cnt_reg[4]/NET0131 , \sport1_cfg_FSi_cnt_reg[5]/NET0131 , \sport1_cfg_FSi_cnt_reg[6]/NET0131 , \sport1_cfg_FSi_cnt_reg[7]/NET0131 , \sport1_cfg_FSi_cnt_reg[8]/NET0131 , \sport1_cfg_FSi_cnt_reg[9]/NET0131 , \sport1_cfg_FSi_reg/NET0131 , \sport1_cfg_RFSg_d1_reg/NET0131 , \sport1_cfg_RFSg_d2_reg/NET0131 , \sport1_cfg_RFSg_d3_reg/NET0131 , \sport1_cfg_RFSgi_d_reg/NET0131 , \sport1_cfg_SCLKi_cnt_reg[0]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[10]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[11]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[12]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[13]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[14]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[15]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[1]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[2]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[3]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[4]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[5]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[6]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[7]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[8]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[9]/NET0131 , \sport1_cfg_SCLKi_h_reg/NET0131 , \sport1_cfg_SP_ENg_D1_reg/P0001 , \sport1_cfg_SP_ENg_reg/NET0131 , \sport1_cfg_TFSg_d1_reg/NET0131 , \sport1_cfg_TFSg_d2_reg/NET0131 , \sport1_cfg_TFSg_d3_reg/NET0131 , \sport1_cfg_TFSgi_d_reg/NET0131 , \sport1_regs_AUTOreg_DO_reg[0]/NET0131 , \sport1_regs_AUTOreg_DO_reg[10]/NET0131 , \sport1_regs_AUTOreg_DO_reg[11]/NET0131 , \sport1_regs_AUTOreg_DO_reg[1]/NET0131 , \sport1_regs_AUTOreg_DO_reg[2]/NET0131 , \sport1_regs_AUTOreg_DO_reg[3]/NET0131 , \sport1_regs_AUTOreg_DO_reg[4]/NET0131 , \sport1_regs_AUTOreg_DO_reg[5]/NET0131 , \sport1_regs_AUTOreg_DO_reg[6]/NET0131 , \sport1_regs_AUTOreg_DO_reg[7]/NET0131 , \sport1_regs_AUTOreg_DO_reg[8]/NET0131 , \sport1_regs_AUTOreg_DO_reg[9]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[0]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[10]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[11]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[12]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[13]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[14]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[15]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[1]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[2]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[3]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[4]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[5]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[6]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[7]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[8]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[9]/NET0131 , \sport1_regs_MWORDreg_DO_reg[0]/NET0131 , \sport1_regs_MWORDreg_DO_reg[10]/NET0131 , \sport1_regs_MWORDreg_DO_reg[1]/NET0131 , \sport1_regs_MWORDreg_DO_reg[2]/NET0131 , \sport1_regs_MWORDreg_DO_reg[3]/NET0131 , \sport1_regs_MWORDreg_DO_reg[4]/NET0131 , \sport1_regs_MWORDreg_DO_reg[5]/NET0131 , \sport1_regs_MWORDreg_DO_reg[6]/NET0131 , \sport1_regs_MWORDreg_DO_reg[7]/NET0131 , \sport1_regs_MWORDreg_DO_reg[8]/NET0131 , \sport1_regs_MWORDreg_DO_reg[9]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 , \sport1_regs_SCTLreg_DO_reg[0]/NET0131 , \sport1_regs_SCTLreg_DO_reg[10]/NET0131 , \sport1_regs_SCTLreg_DO_reg[11]/NET0131 , \sport1_regs_SCTLreg_DO_reg[12]/NET0131 , \sport1_regs_SCTLreg_DO_reg[13]/NET0131 , \sport1_regs_SCTLreg_DO_reg[15]/NET0131 , \sport1_regs_SCTLreg_DO_reg[1]/NET0131 , \sport1_regs_SCTLreg_DO_reg[2]/NET0131 , \sport1_regs_SCTLreg_DO_reg[3]/NET0131 , \sport1_regs_SCTLreg_DO_reg[4]/NET0131 , \sport1_regs_SCTLreg_DO_reg[5]/NET0131 , \sport1_regs_SCTLreg_DO_reg[6]/NET0131 , \sport1_regs_SCTLreg_DO_reg[7]/NET0131 , \sport1_rxctl_Bcnt_reg[0]/NET0131 , \sport1_rxctl_Bcnt_reg[1]/NET0131 , \sport1_rxctl_Bcnt_reg[2]/NET0131 , \sport1_rxctl_Bcnt_reg[3]/NET0131 , \sport1_rxctl_Bcnt_reg[4]/NET0131 , \sport1_rxctl_ISRa_reg/P0001 , \sport1_rxctl_LMcnt_reg[0]/NET0131 , \sport1_rxctl_LMcnt_reg[1]/NET0131 , \sport1_rxctl_LMcnt_reg[2]/NET0131 , \sport1_rxctl_LMcnt_reg[3]/NET0131 , \sport1_rxctl_LMcnt_reg[4]/NET0131 , \sport1_rxctl_RCS_reg[0]/NET0131 , \sport1_rxctl_RCS_reg[1]/NET0131 , \sport1_rxctl_RCS_reg[2]/NET0131 , \sport1_rxctl_RSreq_reg/NET0131 , \sport1_rxctl_RXSHT_reg[0]/P0001 , \sport1_rxctl_RXSHT_reg[10]/P0001 , \sport1_rxctl_RXSHT_reg[11]/P0001 , \sport1_rxctl_RXSHT_reg[12]/P0001 , \sport1_rxctl_RXSHT_reg[13]/P0001 , \sport1_rxctl_RXSHT_reg[14]/P0001 , \sport1_rxctl_RXSHT_reg[15]/P0001 , \sport1_rxctl_RXSHT_reg[1]/P0001 , \sport1_rxctl_RXSHT_reg[2]/P0001 , \sport1_rxctl_RXSHT_reg[3]/P0001 , \sport1_rxctl_RXSHT_reg[4]/P0001 , \sport1_rxctl_RXSHT_reg[5]/P0001 , \sport1_rxctl_RXSHT_reg[6]/P0001 , \sport1_rxctl_RXSHT_reg[7]/P0001 , \sport1_rxctl_RXSHT_reg[8]/P0001 , \sport1_rxctl_RXSHT_reg[9]/P0001 , \sport1_rxctl_RX_reg[0]/P0001 , \sport1_rxctl_RX_reg[10]/P0001 , \sport1_rxctl_RX_reg[11]/P0001 , \sport1_rxctl_RX_reg[12]/P0001 , \sport1_rxctl_RX_reg[13]/P0001 , \sport1_rxctl_RX_reg[14]/P0001 , \sport1_rxctl_RX_reg[15]/P0001 , \sport1_rxctl_RX_reg[1]/P0001 , \sport1_rxctl_RX_reg[2]/P0001 , \sport1_rxctl_RX_reg[3]/P0001 , \sport1_rxctl_RX_reg[4]/P0001 , \sport1_rxctl_RX_reg[5]/P0001 , \sport1_rxctl_RX_reg[6]/P0001 , \sport1_rxctl_RX_reg[7]/P0001 , \sport1_rxctl_RX_reg[8]/P0001 , \sport1_rxctl_RX_reg[9]/P0001 , \sport1_rxctl_SLOT1_EXT_reg[2]/NET0131 , \sport1_rxctl_SLOT1_EXT_reg[3]/NET0131 , \sport1_rxctl_TAG_SLOT_reg/P0001 , \sport1_rxctl_Wcnt_reg[0]/NET0131 , \sport1_rxctl_Wcnt_reg[1]/NET0131 , \sport1_rxctl_Wcnt_reg[2]/NET0131 , \sport1_rxctl_Wcnt_reg[3]/NET0131 , \sport1_rxctl_Wcnt_reg[4]/NET0131 , \sport1_rxctl_Wcnt_reg[5]/NET0131 , \sport1_rxctl_Wcnt_reg[6]/NET0131 , \sport1_rxctl_Wcnt_reg[7]/NET0131 , \sport1_rxctl_a_sync1_reg/P0001 , \sport1_rxctl_a_sync2_reg/P0001 , \sport1_rxctl_sht2nd_reg/P0001 , \sport1_txctl_Bcnt_reg[0]/NET0131 , \sport1_txctl_Bcnt_reg[1]/NET0131 , \sport1_txctl_Bcnt_reg[2]/NET0131 , \sport1_txctl_Bcnt_reg[3]/NET0131 , \sport1_txctl_Bcnt_reg[4]/NET0131 , \sport1_txctl_SP_EN_D1_reg/P0001 , \sport1_txctl_TCS_reg[0]/NET0131 , \sport1_txctl_TCS_reg[1]/NET0131 , \sport1_txctl_TCS_reg[2]/NET0131 , \sport1_txctl_TSreq_reg/NET0131 , \sport1_txctl_TSreqi_reg/NET0131 , \sport1_txctl_TXSHT_reg[0]/P0001 , \sport1_txctl_TXSHT_reg[10]/P0001 , \sport1_txctl_TXSHT_reg[11]/P0001 , \sport1_txctl_TXSHT_reg[12]/P0001 , \sport1_txctl_TXSHT_reg[13]/P0001 , \sport1_txctl_TXSHT_reg[14]/P0001 , \sport1_txctl_TXSHT_reg[15]/P0001 , \sport1_txctl_TXSHT_reg[1]/P0001 , \sport1_txctl_TXSHT_reg[2]/P0001 , \sport1_txctl_TXSHT_reg[3]/P0001 , \sport1_txctl_TXSHT_reg[4]/P0001 , \sport1_txctl_TXSHT_reg[5]/P0001 , \sport1_txctl_TXSHT_reg[6]/P0001 , \sport1_txctl_TXSHT_reg[7]/P0001 , \sport1_txctl_TXSHT_reg[8]/P0001 , \sport1_txctl_TXSHT_reg[9]/P0001 , \sport1_txctl_TX_reg[0]/P0001 , \sport1_txctl_TX_reg[10]/P0001 , \sport1_txctl_TX_reg[11]/P0001 , \sport1_txctl_TX_reg[12]/P0001 , \sport1_txctl_TX_reg[13]/P0001 , \sport1_txctl_TX_reg[14]/P0001 , \sport1_txctl_TX_reg[15]/P0001 , \sport1_txctl_TX_reg[1]/P0001 , \sport1_txctl_TX_reg[2]/P0001 , \sport1_txctl_TX_reg[3]/P0001 , \sport1_txctl_TX_reg[4]/P0001 , \sport1_txctl_TX_reg[5]/P0001 , \sport1_txctl_TX_reg[6]/P0001 , \sport1_txctl_TX_reg[7]/P0001 , \sport1_txctl_TX_reg[8]/P0001 , \sport1_txctl_TX_reg[9]/P0001 , \sport1_txctl_Wcnt_reg[0]/NET0131 , \sport1_txctl_Wcnt_reg[1]/NET0131 , \sport1_txctl_Wcnt_reg[2]/NET0131 , \sport1_txctl_Wcnt_reg[3]/NET0131 , \sport1_txctl_Wcnt_reg[4]/NET0131 , \sport1_txctl_Wcnt_reg[5]/NET0131 , \sport1_txctl_Wcnt_reg[6]/NET0131 , \sport1_txctl_Wcnt_reg[7]/NET0131 , \sport1_txctl_c_sync1_reg/P0001 , \sport1_txctl_c_sync2_reg/P0001 , \tm_MSTAT5_syn_reg/NET0131 , \tm_TCR_TMP_reg[0]/NET0131 , \tm_TCR_TMP_reg[10]/NET0131 , \tm_TCR_TMP_reg[11]/NET0131 , \tm_TCR_TMP_reg[12]/NET0131 , \tm_TCR_TMP_reg[13]/NET0131 , \tm_TCR_TMP_reg[14]/NET0131 , \tm_TCR_TMP_reg[15]/NET0131 , \tm_TCR_TMP_reg[1]/NET0131 , \tm_TCR_TMP_reg[2]/NET0131 , \tm_TCR_TMP_reg[3]/NET0131 , \tm_TCR_TMP_reg[4]/NET0131 , \tm_TCR_TMP_reg[5]/NET0131 , \tm_TCR_TMP_reg[6]/NET0131 , \tm_TCR_TMP_reg[7]/NET0131 , \tm_TCR_TMP_reg[8]/NET0131 , \tm_TCR_TMP_reg[9]/NET0131 , \tm_TINT_GEN1_reg/NET0131 , \tm_TINT_GEN2_reg/NET0131 , \tm_TSR_TMP_reg[0]/NET0131 , \tm_TSR_TMP_reg[1]/NET0131 , \tm_TSR_TMP_reg[2]/NET0131 , \tm_TSR_TMP_reg[3]/NET0131 , \tm_TSR_TMP_reg[4]/NET0131 , \tm_TSR_TMP_reg[5]/NET0131 , \tm_TSR_TMP_reg[6]/NET0131 , \tm_TSR_TMP_reg[7]/NET0131 , \tm_WR_TCR_KEEP_TO_TMCLK_p_reg/NET0131 , \tm_WR_TCR_TMP_GEN1_reg/P0001 , \tm_WR_TCR_TMP_GEN2_reg/P0001 , \tm_WR_TCR_p_reg/P0001 , \tm_WR_TSR_KEEP_TO_TMCLK_p_reg/NET0131 , \tm_WR_TSR_TMP_GEN1_reg/P0001 , \tm_WR_TSR_TMP_GEN2_reg/P0001 , \tm_WR_TSR_p_reg/P0001 , \tm_tcr_reg_DO_reg[0]/NET0131 , \tm_tcr_reg_DO_reg[10]/NET0131 , \tm_tcr_reg_DO_reg[11]/NET0131 , \tm_tcr_reg_DO_reg[12]/NET0131 , \tm_tcr_reg_DO_reg[13]/NET0131 , \tm_tcr_reg_DO_reg[14]/NET0131 , \tm_tcr_reg_DO_reg[15]/NET0131 , \tm_tcr_reg_DO_reg[1]/NET0131 , \tm_tcr_reg_DO_reg[2]/NET0131 , \tm_tcr_reg_DO_reg[3]/NET0131 , \tm_tcr_reg_DO_reg[4]/NET0131 , \tm_tcr_reg_DO_reg[5]/NET0131 , \tm_tcr_reg_DO_reg[6]/NET0131 , \tm_tcr_reg_DO_reg[7]/NET0131 , \tm_tcr_reg_DO_reg[8]/NET0131 , \tm_tcr_reg_DO_reg[9]/NET0131 , \tm_tpr_reg_DO_reg[0]/NET0131 , \tm_tpr_reg_DO_reg[10]/NET0131 , \tm_tpr_reg_DO_reg[11]/NET0131 , \tm_tpr_reg_DO_reg[12]/NET0131 , \tm_tpr_reg_DO_reg[13]/NET0131 , \tm_tpr_reg_DO_reg[14]/NET0131 , \tm_tpr_reg_DO_reg[15]/NET0131 , \tm_tpr_reg_DO_reg[1]/NET0131 , \tm_tpr_reg_DO_reg[2]/NET0131 , \tm_tpr_reg_DO_reg[3]/NET0131 , \tm_tpr_reg_DO_reg[4]/NET0131 , \tm_tpr_reg_DO_reg[5]/NET0131 , \tm_tpr_reg_DO_reg[6]/NET0131 , \tm_tpr_reg_DO_reg[7]/NET0131 , \tm_tpr_reg_DO_reg[8]/NET0131 , \tm_tpr_reg_DO_reg[9]/NET0131 , \tm_tsr_reg_DO_reg[0]/NET0131 , \tm_tsr_reg_DO_reg[1]/NET0131 , \tm_tsr_reg_DO_reg[2]/NET0131 , \tm_tsr_reg_DO_reg[3]/NET0131 , \tm_tsr_reg_DO_reg[4]/NET0131 , \tm_tsr_reg_DO_reg[5]/NET0131 , \tm_tsr_reg_DO_reg[6]/NET0131 , \tm_tsr_reg_DO_reg[7]/NET0131 , \tm_tsr_reg_DO_reg[8]/NET0131 , CLKO_pad, \CMAinx[0]_pad , \CMAinx[10]_pad , \CMAinx[11]_pad , \CMAinx[1]_pad , \CMAinx[2]_pad , \CMAinx[3]_pad , \CMAinx[4]_pad , \CMAinx[5]_pad , \CMAinx[6]_pad , \CMAinx[7]_pad , \CMAinx[8]_pad , \CMAinx[9]_pad , CMSn_pad, CM_cs_pad, \CM_wd[0]_pad , \CM_wd[10]_pad , \CM_wd[11]_pad , \CM_wd[12]_pad , \CM_wd[13]_pad , \CM_wd[14]_pad , \CM_wd[15]_pad , \CM_wd[16]_pad , \CM_wd[17]_pad , \CM_wd[18]_pad , \CM_wd[19]_pad , \CM_wd[1]_pad , \CM_wd[20]_pad , \CM_wd[21]_pad , \CM_wd[22]_pad , \CM_wd[23]_pad , \CM_wd[2]_pad , \CM_wd[3]_pad , \CM_wd[4]_pad , \CM_wd[5]_pad , \CM_wd[6]_pad , \CM_wd[7]_pad , \CM_wd[8]_pad , \CM_wd[9]_pad , CM_web_pad, \CMo_cs0_pad , \CMo_cs1_pad , \CMo_cs2_pad , \CMo_cs3_pad , \CMo_cs4_pad , \CMo_cs5_pad , \CMo_cs6_pad , \CMo_cs7_pad , \DMAinx[0]_pad , \DMAinx[10]_pad , \DMAinx[11]_pad , \DMAinx[12]_pad , \DMAinx[13]_pad , \DMAinx[1]_pad , \DMAinx[2]_pad , \DMAinx[3]_pad , \DMAinx[4]_pad , \DMAinx[5]_pad , \DMAinx[6]_pad , \DMAinx[7]_pad , \DMAinx[8]_pad , \DMAinx[9]_pad , DMSn_pad, DM_cs_pad, \DM_wd[0]_pad , \DM_wd[10]_pad , \DM_wd[11]_pad , \DM_wd[12]_pad , \DM_wd[13]_pad , \DM_wd[14]_pad , \DM_wd[15]_pad , \DM_wd[1]_pad , \DM_wd[2]_pad , \DM_wd[3]_pad , \DM_wd[4]_pad , \DM_wd[5]_pad , \DM_wd[6]_pad , \DM_wd[7]_pad , \DM_wd[8]_pad , \DM_wd[9]_pad , \DMo_cs0_pad , \DMo_cs1_pad , \DMo_cs2_pad , \DMo_cs3_pad , \DMo_cs4_pad , \DMo_cs5_pad , \DMo_cs6_pad , \DMo_cs7_pad , \DSPCLK_cm1_pad , \EA_do[0]_pad , \EA_do[10]_pad , \EA_do[12]_pad , \EA_do[13]_pad , \EA_do[14]_pad , \EA_do[1]_pad , \EA_do[2]_pad , \EA_do[3]_pad , \EA_do[4]_pad , \EA_do[5]_pad , \EA_do[6]_pad , \EA_do[7]_pad , \EA_do[8]_pad , \EA_do[9]_pad , EA_oe_pad, \ED_do[0]_pad , \ED_do[10]_pad , \ED_do[11]_pad , \ED_do[12]_pad , \ED_do[13]_pad , \ED_do[14]_pad , \ED_do[15]_pad , \ED_do[1]_pad , \ED_do[2]_pad , \ED_do[3]_pad , \ED_do[4]_pad , \ED_do[5]_pad , \ED_do[6]_pad , \ED_do[7]_pad , \ED_do[8]_pad , \ED_do[9]_pad , \ED_oe_14_8_pad , \ED_oe_7_0_pad , \IAD_do[0]_pad , \IAD_do[10]_pad , \IAD_do[11]_pad , \IAD_do[12]_pad , \IAD_do[13]_pad , \IAD_do[14]_pad , \IAD_do[15]_pad , \IAD_do[1]_pad , \IAD_do[2]_pad , \IAD_do[3]_pad , \IAD_do[4]_pad , \IAD_do[5]_pad , \IAD_do[6]_pad , \IAD_do[7]_pad , \IAD_do[8]_pad , \IAD_do[9]_pad , IAD_oe_pad, IDoe_pad, IOSn_pad, \PMAinx[0]_pad , \PMAinx[10]_pad , \PMAinx[11]_pad , \PMAinx[1]_pad , \PMAinx[2]_pad , \PMAinx[3]_pad , \PMAinx[4]_pad , \PMAinx[5]_pad , \PMAinx[6]_pad , \PMAinx[7]_pad , \PMAinx[8]_pad , \PMAinx[9]_pad , \PM_wd[0]_pad , \PM_wd[10]_pad , \PM_wd[11]_pad , \PM_wd[12]_pad , \PM_wd[13]_pad , \PM_wd[14]_pad , \PM_wd[15]_pad , \PM_wd[1]_pad , \PM_wd[2]_pad , \PM_wd[3]_pad , \PM_wd[4]_pad , \PM_wd[5]_pad , \PM_wd[6]_pad , \PM_wd[7]_pad , \PM_wd[8]_pad , \PM_wd[9]_pad , \PMo_cs0_pad , \PMo_cs1_pad , \PMo_cs2_pad , \PMo_cs3_pad , \PMo_cs4_pad , \PMo_cs5_pad , \PMo_cs6_pad , \PMo_cs7_pad , \PMo_oe0_pad , \RFS0_pad , \RFS1_pad , \SCLK0_pad , \SCLK1_pad , \TD0_pad , \TD1_pad , \TFS0_pad , \TFS1_pad , \T_ISn_syn_2 , WRn_pad, XTALoffn_pad, \_al_n0 , \bdma_BDMA_boot_reg/NET0131_reg_syn_3 , \bdma_BDMA_boot_reg/n0 , \bdma_BM_cyc_reg/P0000 , \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_3 , \core_c_psq_MGNT_reg/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001_reg_syn_3 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001_reg_syn_3 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001_reg_syn_3 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001_reg_syn_3 , \core_eu_ec_cun_MVi_pre_C_reg/P0001_reg_syn_3 , \core_eu_em_mac_em_reg_Sq_E_reg/P0001_reg_syn_3 , \emc_DMDreg_reg[8]/P0001_reg_syn_3 , \emc_DMDreg_reg[9]/P0001_reg_syn_3 , \emc_ECMcs_reg/P0001 , \emc_PMDreg_reg[8]/P0001_reg_syn_3 , \emc_PMDreg_reg[9]/P0001_reg_syn_3 , \g10/_0_ , \g1000/_0_ , \g10000/_0_ , \g10001/_0_ , \g10002/_0_ , \g10003/_0_ , \g10004/_0_ , \g10005/_0_ , \g10007/_0_ , \g10008/_0_ , \g10009/_0_ , \g1001/_3_ , \g10010/_0_ , \g10011/_0_ , \g10012/_0_ , \g10013/_0_ , \g10014/_0_ , \g10015/_0_ , \g10016/_0_ , \g10017/_0_ , \g10018/_0_ , \g10019/_0_ , \g1002/_3_ , \g10020/_0_ , \g10021/_0_ , \g10022/_0_ , \g10023/_0_ , \g10024/_0_ , \g10025/_0_ , \g10026/_0_ , \g10027/_0_ , \g10028/_0_ , \g10029/_0_ , \g1003/_0_ , \g10030/_0_ , \g10031/_0_ , \g10032/_0_ , \g10033/_0_ , \g10034/_0_ , \g10035/_0_ , \g10036/_0_ , \g10037/_0_ , \g10038/_0_ , \g10039/_0_ , \g10040/_0_ , \g10041/_0_ , \g10042/_0_ , \g10043/_0_ , \g10044/_0_ , \g10045/_0_ , \g10046/_0_ , \g10047/_0_ , \g10048/_0_ , \g10049/_0_ , \g10050/_0_ , \g10051/_0_ , \g10052/_0_ , \g10053/_0_ , \g10054/_0_ , \g10055/_0_ , \g10056/_0_ , \g10057/_0_ , \g10058/_0_ , \g10059/_0_ , \g10060/_0_ , \g10061/_0_ , \g10062/_0_ , \g10063/_0_ , \g10064/_0_ , \g10065/_0_ , \g10066/_0_ , \g10067/_0_ , \g10068/_0_ , \g10069/_0_ , \g10070/_0_ , \g10071/_0_ , \g10072/_0_ , \g10073/_0_ , \g10074/_0_ , \g10075/_0_ , \g10076/_0_ , \g10077/_0_ , \g10078/_0_ , \g10080/_0_ , \g10081/_0_ , \g10083/_0_ , \g10089/_0_ , \g1009/_0_ , \g10090/_0_ , \g10091/_0_ , \g10092/_0_ , \g10093/_0_ , \g10094/_0_ , \g1010/_0_ , \g10108/_3_ , \g1011/_0_ , \g10110/_0_ , \g10111/_0_ , \g10113/_3_ , \g10115/_3_ , \g1013/_0_ , \g1014/_0_ , \g10152/_0_ , \g10153/_0_ , \g10154/_0_ , \g10155/_0_ , \g10156/_0_ , \g10157/_0_ , \g10158/_0_ , \g10159/_0_ , \g1016/_0_ , \g10160/_0_ , \g10161/_0_ , \g10162/_0_ , \g10163/_0_ , \g10164/_0_ , \g10165/_0_ , \g1017/_0_ , \g10170/_3_ , \g1018/_0_ , \g10190/_3_ , \g10194/_3_ , \g10198/_0_ , \g10199/_0_ , \g102/_0_ , \g103/_0_ , \g104/_0_ , \g105/_0_ , \g10598/_0_ , \g106/_0_ , \g10667/_0_ , \g10683/_0_ , \g10685/_0_ , \g107/_0_ , \g10721/_0_ , \g10758/_0_ , \g10765/_0_ , \g10778/_0_ , \g10791/_0_ , \g108/_0_ , \g10887/_0_ , \g1089/_0_ , \g109/_0_ , \g1090/_0_ , \g1091/_0_ , \g1092/_0_ , \g10923/_0_ , \g1093/_0_ , \g10930/_0_ , \g10931/_0_ , \g10936/_0_ , \g1097/_0_ , \g11/_0_ , \g110/_0_ , \g1101/_0_ , \g11013/_0_ , \g1102/_0_ , \g1103/_0_ , \g11032/_0_ , \g1104/_0_ , \g1105/_0_ , \g1107/_0_ , \g11074/_0_ , \g11077/_0_ , \g1108/_0_ , \g1109/_0_ , \g11112/_0_ , \g11115/_0_ , \g11116/_0_ , \g11119/_0_ , \g11120/_0_ , \g1113/_0_ , \g1115/_0_ , \g1116/_0_ , \g1117/_0_ , \g11267/_0_ , \g11281/_0_ , \g11287/_0_ , \g11300/_0_ , \g11323/_0_ , \g11325/_2__syn_2 , \g11345/_2_ , \g11470/_0_ , \g11471/_0_ , \g11472/_0_ , \g11473/_0_ , \g11474/_0_ , \g11476/_0_ , \g11477/_0_ , \g11496/_0_ , \g11497/_0_ , \g11498/_0_ , \g11499/_0_ , \g11500/_0_ , \g11501/_0_ , \g11502/_0_ , \g11503/_0_ , \g11504/_0_ , \g11505/_0_ , \g11506/_0_ , \g11507/_0_ , \g11509/_0_ , \g11510/_0_ , \g11515/_0_ , \g11516/_0_ , \g11520/_0_ , \g11521/_0_ , \g11576/_0_ , \g11577/_0_ , \g11578/_0_ , \g11579/_0_ , \g11580/_0_ , \g11581/_0_ , \g11582/_0_ , \g11583/_0_ , \g11584/_0_ , \g11585/_0_ , \g11586/_0_ , \g11587/_0_ , \g11588/_0_ , \g11589/_0_ , \g11591/_0_ , \g11593/_0_ , \g11595/_0_ , \g11596/_0_ , \g11597/_0_ , \g11605/_0_ , \g11606/_0_ , \g11607/_0_ , \g11608/_0_ , \g11609/_0_ , \g11610/_0_ , \g11611/_0_ , \g11612/_0_ , \g11613/_0_ , \g11615/_0_ , \g11616/_0_ , \g11617/_0_ , \g11651/_3_ , \g11704/_0_ , \g11705/_0_ , \g11709/_0_ , \g11722/_0_ , \g11723/_0_ , \g119/_0_ , \g1192/_0_ , \g11994/_0_ , \g120/_0_ , \g1200/_0_ , \g12003/_0_ , \g1201/_0_ , \g12019/_0_ , \g1203/_3_ , \g1204/_3_ , \g1207/_0_ , \g1208/_0_ , \g12092/_0_ , \g1210/_0_ , \g1211/_0_ , \g1212/_0_ , \g1213/_0_ , \g12145/_0_ , \g12155/_0_ , \g12186/_0_ , \g12187/_0_ , \g12192/_0_ , \g12201/_0_ , \g12202/_0_ , \g12203/_0_ , \g12204/_0_ , \g12207/_0_ , \g12229/_3_ , \g12267/_0_ , \g12276/_0_ , \g12278/_0_ , \g12279/_0_ , \g12280/_0_ , \g12302/_0_ , \g12316/_0_ , \g12317/_0_ , \g12319/_0_ , \g12328/_3_ , \g1233/_0_ , \g12348/_0_ , \g12351/_0_ , \g12352/_0_ , \g12353/_0_ , \g12354/_0_ , \g12355/_0_ , \g1237/_0_ , \g124/_0_ , \g12444/_0_ , \g125/_0_ , \g12637/_0_ , \g12639/_0_ , \g12658/_0_ , \g12659/_0_ , \g12660/_0_ , \g12663/_0_ , \g12664/_0_ , \g12665/_0_ , \g12672/_3_ , \g12673/_3_ , \g12674/_3_ , \g12675/_3_ , \g12676/_3_ , \g12677/_3_ , \g12678/_0_ , \g12679/_3_ , \g12697/_3_ , \g12701/_3_ , \g12711/_2_ , \g12713/_2_ , \g12715/_2_ , \g12717/_2_ , \g12718/_2__syn_2 , \g1272/_0_ , \g12728/_1__syn_2 , \g12730/_3_ , \g12741/_1__syn_2 , \g12746/_0__syn_2 , \g12748/_0_ , \g12749/_0_ , \g12759/_1__syn_2 , \g12760/_0_ , \g12762/_0_ , \g12763/_0_ , \g12764/_0_ , \g12765/_0_ , \g12766/_0_ , \g12767/_0_ , \g12768/_0_ , \g12769/_0_ , \g12770/_0_ , \g12771/_0_ , \g12772/_0_ , \g12773/_0_ , \g12774/_0_ , \g12775/_0_ , \g12776/_0_ , \g12777/_0_ , \g12778/_0_ , \g12779/_0_ , \g1278/_0_ , \g12780/_0_ , \g12781/_0_ , \g12782/_0_ , \g12783/_0_ , \g12784/_0_ , \g12785/_0_ , \g12786/_0_ , \g12787/_0_ , \g12788/_0_ , \g12789/_0_ , \g12790/_0_ , \g12791/_0_ , \g12792/_0_ , \g12793/_0_ , \g12794/_0_ , \g12795/_0_ , \g12796/_0_ , \g12797/_0_ , \g12798/_0_ , \g12799/_0_ , \g12800/_0_ , \g12801/_0_ , \g12802/_0_ , \g12803/_0_ , \g12804/_0_ , \g12805/_0_ , \g12806/_0_ , \g12807/_0_ , \g12808/_0_ , \g12809/_0_ , \g1281/_0_ , \g12810/_0_ , \g12811/_0_ , \g12812/_0_ , \g12813/_0_ , \g12814/_0_ , \g12815/_0_ , \g12816/_0_ , \g12817/_0_ , \g12818/_0_ , \g12819/_0_ , \g1282/_0_ , \g12820/_0_ , \g12821/_0_ , \g12822/_0_ , \g12823/_0_ , \g12824/_0_ , \g12825/_0_ , \g12826/_0_ , \g12827/_0_ , \g12828/_0_ , \g12829/_0_ , \g12830/_0_ , \g12831/_0_ , \g12832/_0_ , \g12833/_0_ , \g12835/_0_ , \g12836/_0_ , \g12838/_0_ , \g12848/_0_ , \g12849/_0_ , \g1285/_0_ , \g12850/_0_ , \g12857/_0_ , \g12858/_0_ , \g12859/_0_ , \g12861/_0_ , \g12862/_0_ , \g12868/_0_ , \g12869/_0_ , \g1287/_0_ , \g12870/_0_ , \g12871/_0_ , \g12872/_0_ , \g12873/_0_ , \g12874/_0_ , \g12875/_0_ , \g12876/_0_ , \g12877/_0_ , \g12878/_0_ , \g12879/_0_ , \g12880/_0_ , \g12881/_0_ , \g12882/_0_ , \g12883/_0_ , \g12884/_0_ , \g12885/_0_ , \g12886/_0_ , \g12887/_0_ , \g12888/_0_ , \g12889/_0_ , \g1289/_0_ , \g12890/_0_ , \g12891/_0_ , \g12894/_0_ , \g12898/_0_ , \g12899/_0_ , \g12900/_0_ , \g12901/_0_ , \g12902/_0_ , \g12903/_0_ , \g12906/_0_ , \g12907/_0_ , \g12908/_0_ , \g12912/_0_ , \g12913/_0_ , \g12914/_0_ , \g12915/_0_ , \g12916/_0_ , \g12917/_0_ , \g12918/_0_ , \g12919/_0_ , \g12920/_0_ , \g12921/_0_ , \g12922/_0_ , \g12923/_0_ , \g12924/_0_ , \g12925/_0_ , \g12926/_0_ , \g12932/_0_ , \g12933/_0_ , \g12936/_0_ , \g12955/_0_ , \g13015/_0_ , \g13016/_0_ , \g13017/_0_ , \g13018/_0_ , \g13019/_0_ , \g13020/_0_ , \g13021/_0_ , \g13024/_0_ , \g13025/_0_ , \g13027/_0_ , \g13028/_0_ , \g13030/_0_ , \g13031/_0_ , \g13033/_0_ , \g13047/_0_ , \g13060/_0_ , \g13062/_0_ , \g13063/_0_ , \g13064/_0_ , \g13067/_0_ , \g13068/_0_ , \g13069/_0_ , \g13070/_0_ , \g13072/_0_ , \g13094/_0_ , \g13104/_0_ , \g13110/_0_ , \g13114/_0_ , \g13115/_0_ , \g13116/_0_ , \g13117/_0_ , \g13118/_0_ , \g13119/_0_ , \g13120/_0_ , \g13121/_0_ , \g13124/_0_ , \g13125/_0_ , \g13127/_0_ , \g13128/_0_ , \g13129/_0_ , \g13130/_0_ , \g13131/_0_ , \g13132/_0_ , \g13133/_0_ , \g13134/_0_ , \g13138/_0_ , \g13139/_0_ , \g13140/_0_ , \g13141/_0_ , \g13142/_0_ , \g13143/_0_ , \g13144/_0_ , \g13146/_0_ , \g13150/_0_ , \g13152/_0_ , \g13154/_0_ , \g13155/_0_ , \g13156/_0_ , \g13157/_0_ , \g13158/_0_ , \g1320/_3_ , \g13266/_0_ , \g13269/_0_ , \g13274/_0_ , \g13277/_0_ , \g13280/_0_ , \g13283/_0_ , \g13294/_0_ , \g13330/_0_ , \g13333/_0_ , \g13334/_0_ , \g13335/_0_ , \g13336/_0_ , \g13337/_0_ , \g13338/_0_ , \g13345/_0_ , \g13346/_0_ , \g13347/_0_ , \g13348/_0_ , \g13349/_0_ , \g13350/_0_ , \g13351/_0_ , \g13352/_0_ , \g13486/_0_ , \g13488/_0_ , \g13508/_0_ , \g13509/_0_ , \g13510/_0_ , \g13511/_0_ , \g13512/_0_ , \g13513/_0_ , \g13514/_0_ , \g13515/_0_ , \g13516/_0_ , \g13517/_0_ , \g13518/_0_ , \g13519/_0_ , \g13520/_0_ , \g13521/_0_ , \g13540/_0_ , \g13541/_0_ , \g13542/_0_ , \g13543/_0_ , \g13544/_0_ , \g13545/_0_ , \g13546/_0_ , \g13547/_0_ , \g13548/_0_ , \g13549/_0_ , \g13550/_0_ , \g13551/_0_ , \g13552/_0_ , \g13553/_0_ , \g13554/_0_ , \g13555/_0_ , \g13556/_0_ , \g13557/_0_ , \g13558/_0_ , \g13559/_0_ , \g13560/_0_ , \g13561/_0_ , \g13562/_0_ , \g13563/_0_ , \g13564/_0_ , \g13565/_0_ , \g13566/_0_ , \g13567/_0_ , \g13568/_0_ , \g13569/_0_ , \g13570/_0_ , \g13571/_0_ , \g13572/_0_ , \g137/_3_ , \g1387/_3_ , \g1388/_3_ , \g1389/_0_ , \g139/_0_ , \g1390/_0_ , \g1393/_0_ , \g140/_0_ , \g141/_0_ , \g14173/_0_ , \g14176/_0_ , \g142/_3_ , \g14273/_1__syn_2 , \g14274/_0_ , \g14280/_0_ , \g14281/_0_ , \g143/_3_ , \g14354/_3__syn_2 , \g14370/_0_ , \g14385/_0_ , \g14386/_0_ , \g144/_3_ , \g14407/_0_ , \g14412/_0_ , \g14435/_0_ , \g14439/_0_ , \g145/_0_ , \g14522/_0_ , \g14528/_0_ , \g14533/_0_ , \g14581/_1_ , \g14582/_0_ , \g146/_3_ , \g14671/_0_ , \g14672/_0_ , \g147/_0_ , \g1473/_0_ , \g148/_0_ , \g14826/_0_ , \g149/_0_ , \g14908/_0_ , \g14911/_0_ , \g14936/_2_ , \g1494/_0_ , \g1495/_0_ , \g14950/_2_ , \g14953/_2_ , \g15003/_0_ , \g15004/_0_ , \g15006/_0_ , \g15007/_0_ , \g15008/_0_ , \g15009/_0_ , \g15010/_0_ , \g15011/_0_ , \g15012/_0_ , \g15013/_0_ , \g15014/_0_ , \g15015/_0_ , \g15016/_0_ , \g15017/_0_ , \g15018/_0_ , \g15019/_0_ , \g15035/_0_ , \g15036/_0_ , \g15038/_0_ , \g15039/_0_ , \g15040/_0_ , \g15041/_0_ , \g15042/_0_ , \g15043/_0_ , \g15044/_0_ , \g15045/_0_ , \g15046/_0_ , \g15056/_00_ , \g151/_0_ , \g15193/_0_ , \g152/_0_ , \g15256/_0_ , \g153/_0_ , \g15393/_0_ , \g15394/_0_ , \g15395/_0_ , \g15396/_0_ , \g15397/_0_ , \g15398/_0_ , \g15399/_0_ , \g154/_0_ , \g15400/_0_ , \g15401/_0_ , \g15402/_0_ , \g15403/_0_ , \g15404/_0_ , \g15405/_0_ , \g15406/_0_ , \g15407/_0_ , \g15408/_0_ , \g15473/_0_ , \g15650/_0_ , \g15651/_0_ , \g15652/_0_ , \g15653/_0_ , \g15662/_0_ , \g15663/_0_ , \g15664/_0_ , \g15665/_0_ , \g15666/_0_ , \g15667/_0_ , \g15668/_0_ , \g15669/_0_ , \g15670/_0_ , \g15671/_0_ , \g15672/_0_ , \g15673/_0_ , \g15674/_0_ , \g15675/_0_ , \g1569/_0_ , \g1570/_0_ , \g1575/_0_ , \g1576/_0_ , \g15922/_1_ , \g15970/_0_ , \g16059/_0_ , \g1606/_3_ , \g16124/_0_ , \g16144/_0_ , \g16202/_0_ , \g16214/_0_ , \g16247/_0_ , \g16257/_0_ , \g16274/_1_ , \g16324/_0_ , \g16343/_1__syn_2 , \g16381/_0_ , \g16383/_0_ , \g16386/_0_ , \g16414/_1__syn_2 , \g16416/_0__syn_2 , \g16448/_0_ , \g16460/_1_ , \g16625/_3_ , \g16662/_0_ , \g16668/_1__syn_2 , \g16692/_0_ , \g16721/_0_ , \g16723/_0_ , \g16725/_0_ , \g16726/_0_ , \g16727/_0_ , \g16728/_0_ , \g16729/_0_ , \g16730/_0_ , \g16731/_0_ , \g16732/_0_ , \g16733/_0_ , \g16734/_0_ , \g16735/_0_ , \g16736/_0_ , \g16737/_0_ , \g16738/_0_ , \g16739/_0_ , \g16740/_0_ , \g16741/_0_ , \g16742/_0_ , \g16743/_0_ , \g16747/_0_ , \g16748/_0_ , \g16749/_0_ , \g16750/_0_ , \g16753/_0_ , \g16754/_0_ , \g16755/_0_ , \g16756/_0_ , \g16757/_0_ , \g16758/_0_ , \g16761/_0_ , \g16765/_0_ , \g16766/_0_ , \g16767/_0_ , \g16768/_0_ , \g16769/_0_ , \g16772/_0_ , \g16785/_0_ , \g16786/_0_ , \g16787/_0_ , \g16788/_0_ , \g16789/_0_ , \g16790/_0_ , \g16791/_0_ , \g16804/_0_ , \g16805/_0_ , \g16806/_0_ , \g16807/_0_ , \g16808/_0_ , \g16809/_0_ , \g16810/_0_ , \g16811/_0_ , \g16812/_0_ , \g16813/_0_ , \g16814/_0_ , \g16815/_0_ , \g16816/_0_ , \g16817/_0_ , \g16819/_0_ , \g16822/_0_ , \g16823/_0_ , \g16824/_0_ , \g16825/_0_ , \g16828/_0_ , \g16829/_0_ , \g16830/_0_ , \g16831/_0_ , \g16832/_0_ , \g16833/_0_ , \g16834/_0_ , \g16835/_0_ , \g16836/_0_ , \g16837/_0_ , \g16840/_0_ , \g16841/_0_ , \g16842/_0_ , \g16843/_0_ , \g16846/_0_ , \g16847/_0_ , \g16848/_0_ , \g16849/_0_ , \g16850/_0_ , \g16851/_0_ , \g16852/_0_ , \g16853/_0_ , \g16854/_0_ , \g16855/_0_ , \g16856/_0_ , \g16857/_0_ , \g16859/_0_ , \g16862/_0_ , \g16865/_0_ , \g16866/_0_ , \g16867/_0_ , \g16868/_0_ , \g16869/_0_ , \g16870/_0_ , \g16871/_0_ , \g16872/_0_ , \g16873/_0_ , \g16874/_0_ , \g16875/_0_ , \g16876/_0_ , \g16877/_0_ , \g16878/_0_ , \g16879/_0_ , \g16880/_0_ , \g16881/_0_ , \g16882/_0_ , \g16884/_0_ , \g16887/_0_ , \g16891/_0_ , \g16892/_0_ , \g16893/_0_ , \g16894/_0_ , \g16895/_0_ , \g16897/_0_ , \g16898/_0_ , \g16899/_0_ , \g16900/_0_ , \g16901/_0_ , \g16902/_0_ , \g16903/_0_ , \g16904/_0_ , \g16905/_0_ , \g16906/_0_ , \g16907/_0_ , \g16908/_0_ , \g16909/_0_ , \g16910/_0_ , \g16912/_0_ , \g16914/_0_ , \g16915/_0_ , \g16950/_0_ , \g16951/_0_ , \g16952/_0_ , \g16953/_0_ , \g16954/_0_ , \g16955/_0_ , \g16956/_0_ , \g16957/_0_ , \g16958/_0_ , \g16959/_0_ , \g16960/_0_ , \g16961/_0_ , \g16962/_0_ , \g16963/_0_ , \g16964/_0_ , \g16965/_0_ , \g16966/_0_ , \g16967/_0_ , \g16968/_0_ , \g16970/_0_ , \g17102/_3_ , \g17106/_0_ , \g17107/_0_ , \g17109/_0_ , \g17110/_0_ , \g17111/_0_ , \g17112/_0_ , \g17115/_0_ , \g17116/_0_ , \g17119/_0_ , \g17120/_0_ , \g17122/_0_ , \g17123/_0_ , \g17124/_0_ , \g17125/_0_ , \g17126/_0_ , \g17127/_0_ , \g17128/_0_ , \g17130/_0_ , \g17131/_0_ , \g17132/_0_ , \g17133/_0_ , \g17134/_0_ , \g17135/_0_ , \g17136/_0_ , \g17137/_0_ , \g17138/_0_ , \g17140/_0_ , \g17141/_0_ , \g17142/_0_ , \g17143/_0_ , \g17144/_0_ , \g17145/_0_ , \g17146/_0_ , \g17147/_0_ , \g17148/_0_ , \g17149/_0_ , \g17150/_0_ , \g17151/_0_ , \g17152/_0_ , \g17153/_0_ , \g17154/_0_ , \g17155/_0_ , \g17157/_0_ , \g17159/_0_ , \g17160/_0_ , \g17161/_0_ , \g17162/_0_ , \g17163/_0_ , \g17164/_0_ , \g17165/_0_ , \g17166/_0_ , \g17168/_0_ , \g17171/_0_ , \g17173/_0_ , \g17177/_0_ , \g17178/_0_ , \g17179/_0_ , \g17180/_0_ , \g17182/_0_ , \g17183/_0_ , \g17184/_0_ , \g17185/_0_ , \g17186/_0_ , \g17188/_0_ , \g17189/_0_ , \g17190/_0_ , \g17191/_0_ , \g17193/_0_ , \g17194/_0_ , \g17195/_0_ , \g17196/_0_ , \g17197/_0_ , \g17198/_0_ , \g17199/_0_ , \g17200/_0_ , \g17201/_0_ , \g17202/_0_ , \g17203/_0_ , \g17204/_0_ , \g17205/_0_ , \g17206/_0_ , \g17207/_0_ , \g17208/_0_ , \g17209/_0_ , \g17210/_0_ , \g17211/_0_ , \g17212/_0_ , \g17213/_0_ , \g17214/_0_ , \g17215/_0_ , \g17216/_0_ , \g17217/_0_ , \g17218/_0_ , \g17219/_0_ , \g17223/_0_ , \g17224/_0_ , \g17225/_0_ , \g17226/_0_ , \g17227/_0_ , \g17228/_0_ , \g17229/_0_ , \g17231/_0_ , \g17232/_0_ , \g17233/_0_ , \g17234/_0_ , \g17237/_0_ , \g17239/_0_ , \g17240/_0_ , \g17243/_0_ , \g17246/_0_ , \g17247/_0_ , \g17248/_0_ , \g17249/_0_ , \g17250/_0_ , \g17251/_0_ , \g17252/_0_ , \g17253/_0_ , \g17254/_0_ , \g17258/_0_ , \g17261/_0_ , \g17262/_0_ , \g17269/_0_ , \g17271/_0_ , \g17274/_0_ , \g17275/_0_ , \g17276/_0_ , \g17277/_0_ , \g17278/_0_ , \g17279/_0_ , \g17280/_0_ , \g17281/_0_ , \g17282/_0_ , \g17283/_0_ , \g17285/_0_ , \g17290/_0_ , \g17292/_0_ , \g17293/_0_ , \g17296/_0_ , \g17297/_0_ , \g17298/_0_ , \g173/_0_ , \g17303/_0_ , \g17304/_0_ , \g17305/_0_ , \g17306/_0_ , \g17307/_0_ , \g17308/_0_ , \g17309/_0_ , \g17310/_0_ , \g17311/_0_ , \g17312/_0_ , \g17314/_0_ , \g17315/_0_ , \g17316/_0_ , \g17317/_0_ , \g17318/_0_ , \g17319/_0_ , \g17320/_0_ , \g17321/_0_ , \g17322/_0_ , \g17323/_0_ , \g17324/_0_ , \g17325/_0_ , \g17326/_0_ , \g17327/_0_ , \g17328/_0_ , \g17329/_0_ , \g17330/_0_ , \g17331/_0_ , \g17332/_0_ , \g17333/_0_ , \g17335/_0_ , \g17336/_0_ , \g17337/_0_ , \g17338/_0_ , \g17339/_0_ , \g17340/_0_ , \g17342/_0_ , \g17343/_0_ , \g17347/_0_ , \g17350/_0_ , \g17354/_0_ , \g17356/_0_ , \g17357/_0_ , \g17358/_0_ , \g17359/_0_ , \g17360/_0_ , \g17415/_0_ , \g17441/_0_ , \g17442/_0_ , \g17451/_0_ , \g17457/_0_ , \g17458/_0_ , \g17459/_0_ , \g17460/_0_ , \g17461/_0_ , \g17462/_0_ , \g17463/_0_ , \g17464/_0_ , \g17465/_0_ , \g17466/_0_ , \g17467/_0_ , \g17468/_0_ , \g17469/_0_ , \g17470/_0_ , \g17471/_0_ , \g17472/_0_ , \g175/_3_ , \g1750/_0_ , \g176/_3_ , \g17619/_0_ , \g17620/_0_ , \g1763/_3_ , \g1764/_3_ , \g1768/_0_ , \g1769/_0_ , \g177/_3_ , \g17737/_0_ , \g17747/_0_ , \g178/_3_ , \g17814/_1_ , \g17815/_0_ , \g17821/_1_ , \g17821/_1__syn_2 , \g17872/_0_ , \g179/_3_ , \g17902/_0_ , \g180/_3_ , \g18020/_1_ , \g18057/_0_ , \g18096/_0_ , \g18099/_0_ , \g18107/_0_ , \g18133/_0_ , \g18140/_1_ , \g18153/_0_ , \g182/_0_ , \g18218/_0_ , \g18244/_0_ , \g18262/_0_ , \g18267/_0_ , \g18387/_1__syn_2 , \g184/_0_ , \g18478/_1_ , \g18585/_3_ , \g18608/_0_ , \g18609/_0_ , \g18613/_0_ , \g18618/_0_ , \g18647/_0_ , \g18687/_2_ , \g18707/_0_ , \g18748/_0_ , \g18753/_0_ , \g18758/_0_ , \g18759/_0_ , \g18760/_0_ , \g18761/_0_ , \g18762/_0_ , \g18763/_0_ , \g18764/_0_ , \g18765/_0_ , \g18766/_0_ , \g18767/_0_ , \g18768/_0_ , \g18770/_0_ , \g18771/_0_ , \g18788/_0_ , \g18796/_0_ , \g18800/_0_ , \g18801/_0_ , \g18802/_0_ , \g18803/_0_ , \g18804/_0_ , \g18805/_0_ , \g18807/_0_ , \g18840/_0_ , \g18843/_0_ , \g18844/_0_ , \g18846/_0_ , \g18847/_0_ , \g18848/_0_ , \g18849/_0_ , \g18850/_0_ , \g18851/_0_ , \g18852/_0_ , \g18853/_0_ , \g18854/_0_ , \g18855/_0_ , \g18856/_0_ , \g18858/_0_ , \g18860/_0_ , \g18861/_0_ , \g18863/_0_ , \g18864/_0_ , \g18866/_0_ , \g18867/_0_ , \g18868/_0_ , \g18869/_0_ , \g18870/_0_ , \g18871/_0_ , \g18872/_0_ , \g18873/_0_ , \g18874/_0_ , \g18875/_0_ , \g18876/_0_ , \g18877/_0_ , \g18878/_0_ , \g18879/_0_ , \g18880/_0_ , \g18881/_0_ , \g18882/_0_ , \g18883/_0_ , \g18888/_0_ , \g18892/_0_ , \g18895/_0_ , \g18896/_0_ , \g18897/_0_ , \g18905/_0_ , \g18908/_0_ , \g18909/_0_ , \g18912/_0_ , \g18918/_0_ , \g18919/_0_ , \g18920/_0_ , \g18921/_0_ , \g18922/_0_ , \g18924/_0_ , \g18925/_0_ , \g18927/_0_ , \g18930/_0_ , \g18966/_0_ , \g18968/_0_ , \g18970/_0_ , \g18974/_0_ , \g18975/_0_ , \g18977/_0_ , \g18981/_0_ , \g18983/_0_ , \g18985/_0_ , \g18987/_0_ , \g18989/_0_ , \g18991/_0_ , \g18992/_0_ , \g18993/_0_ , \g18994/_0_ , \g18995/_0_ , \g18996/_0_ , \g18997/_0_ , \g18998/_0_ , \g18999/_0_ , \g19001/_0_ , \g19003/_0_ , \g19005/_0_ , \g19006/_0_ , \g19014/_0_ , \g19016/_0_ , \g19018/_0_ , \g19020/_0_ , \g19022/_0_ , \g19056/_3_ , \g19058/_3_ , \g19060/_3_ , \g19062/_3_ , \g1910/_0_ , \g19186/_0_ , \g19188/_0_ , \g19235/_0_ , \g19239/_0_ , \g19244/_0_ , \g19253/_0_ , \g19254/_0_ , \g19259/_0_ , \g19261/_0_ , \g19267/_0_ , \g19277/_0_ , \g19278/_0_ , \g19280/_0_ , \g19281/_0_ , \g19282/_0_ , \g19283/_0_ , \g19284/_0_ , \g19285/_0_ , \g19286/_0_ , \g19287/_0_ , \g19288/_0_ , \g19289/_0_ , \g19290/_0_ , \g19291/_0_ , \g19292/_0_ , \g19293/_0_ , \g19294/_0_ , \g19295/_0_ , \g19296/_0_ , \g19297/_0_ , \g19298/_0_ , \g19299/_0_ , \g19300/_0_ , \g19301/_0_ , \g19302/_0_ , \g19303/_0_ , \g19304/_0_ , \g19305/_0_ , \g19306/_0_ , \g19307/_0_ , \g19308/_0_ , \g19315/_0_ , \g19316/_0_ , \g19317/_0_ , \g19318/_0_ , \g19319/_0_ , \g19320/_0_ , \g19321/_0_ , \g19322/_0_ , \g19323/_0_ , \g19325/_3_ , \g19326/_3_ , \g19333/_3_ , \g19341/_3_ , \g19347/_3_ , \g19377/_3_ , \g19381/_3_ , \g19393/_0_ , \g19401/_0_ , \g19402/_0_ , \g195/_2_ , \g19513/_0_ , \g19514/_0_ , \g19515/_0_ , \g19516/_0_ , \g1952/_3_ , \g19529/_0_ , \g19530/_0_ , \g19531/_0_ , \g19532/_0_ , \g19533/_0_ , \g19534/_0_ , \g19535/_0_ , \g19536/_0_ , \g19537/_0_ , \g19539/_0_ , \g19546/_0_ , \g19552/_0_ , \g19553/_0_ , \g19562/_0_ , \g19563/_0_ , \g19564/_0_ , \g19572/_0_ , \g19575/_0_ , \g19615/_0_ , \g19686/_0_ , \g19688/_0_ , \g197/_0_ , \g19729/_0_ , \g19774/_0_ , \g19777/_0_ , \g19791/_0_ , \g19818/_0_ , \g19819/_0_ , \g19828/_0_ , \g19852/_1_ , \g19860/_0_ , \g19861/_0_ , \g19864/_0_ , \g19886/_0_ , \g19887/_0_ , \g199/_0_ , \g19908/_0_ , \g19918/_0_ , \g19927/_0_ , \g19933/_0_ , \g200/_0_ , \g20019/_0_ , \g20046/_0_ , \g20068/_1_ , \g20080/_1_ , \g201/_0_ , \g20137/_0_ , \g20139/_0_ , \g20141/_0_ , \g20152/_1_ , \g20154/_00_ , \g202/_0_ , \g20206/_0_ , \g20211/_2_ , \g20217/_2_ , \g20239/_0_ , \g20265/_2_ , \g20266/_0_ , \g20272/_2_ , \g20278/_2_ , \g20283/_0_ , \g20285/_2_ , \g20288/_2__syn_2 , \g20293/_0_ , \g20295/_2_ , \g203/_0_ , \g20302/_2_ , \g20303/_2_ , \g20304/_2_ , \g20311/_2_ , \g20326/_0_ , \g20330/_0_ , \g2034/_0_ , \g20345/_0_ , \g20346/_0_ , \g2035/_0_ , \g20363/_0_ , \g20364/_0_ , \g204/_0_ , \g2047/_0_ , \g20483/_0_ , \g20493/_00_ , \g205/_0_ , \g20569/_0_ , \g20570/_0_ , \g20571/_0_ , \g206/_0_ , \g20613/_0_ , \g20615/_0_ , \g20657/_1__syn_2 , \g20660/_0_ , \g20685/_0_ , \g207/_0_ , \g20713/_1_ , \g20747/_1_ , \g20784/_0_ , \g20820/_1_ , \g20859/_0_ , \g20873/_2_ , \g20886/_0_ , \g20887/_0_ , \g20891/_2__syn_2 , \g20907/_2_ , \g20936/_2__syn_2 , \g20937/_1_ , \g20955/_0_ , \g20959/_2__syn_2 , \g20967/_0_ , \g20971/_2__syn_2 , \g20974/_1__syn_2 , \g21015/_1_ , \g21051/_2_ , \g21079/_1_ , \g21081/_1_ , \g21087/_2__syn_2 , \g21114/_1_ , \g21116/_1_ , \g21120/_2__syn_2 , \g21147/_0_ , \g21179/_1_ , \g21185/_1_ , \g21223/_0_ , \g21242/_0_ , \g21253/_0_ , \g21257/_0_ , \g21323/_1_ , \g21324/_1_ , \g21366/_0_ , \g21385/_2_ , \g21464/_0_ , \g21475/_3_ , \g21481/_0_ , \g21482/_0_ , \g21494/_3_ , \g21500/_3_ , \g21507/_3_ , \g21511/_3_ , \g21537/_1_ , \g21568/_0_ , \g21591/_0_ , \g21604/_0_ , \g21605/_3_ , \g21606/_0_ , \g21607/_0_ , \g21608/_0_ , \g21609/_0_ , \g21610/_0_ , \g21611/_0_ , \g21612/_0_ , \g21613/_0_ , \g21614/_0_ , \g21615/_0_ , \g21616/_0_ , \g21617/_0_ , \g21618/_0_ , \g21621/_0_ , \g21640/_0_ , \g21678/_0_ , \g21679/_0_ , \g21686/_0_ , \g21692/_3_ , \g21696/_0_ , \g21698/_0_ , \g21702/_3_ , \g21707/_0_ , \g21709/_0_ , \g21728/_0_ , \g21729/_0_ , \g21731/_0_ , \g21732/_0_ , \g21733/_0_ , \g21736/_0_ , \g21744/_3_ , \g21753/_0_ , \g21754/_0_ , \g21755/_0_ , \g21756/_0_ , \g21757/_0_ , \g21759/_0_ , \g21761/_0_ , \g21763/_0_ , \g21764/_0_ , \g21766/_0_ , \g2180/_0_ , \g21853/_3_ , \g21861/_3_ , \g21863/_3_ , \g21869/_3_ , \g2187/_0_ , \g21875/_3_ , \g21877/_3_ , \g21879/_3_ , \g2188/_0_ , \g21900/_0_ , \g22080/_0_ , \g22082/_0_ , \g22135/_0_ , \g22145/_1_ , \g22225/_0_ , \g223/_0_ , \g22354/_0_ , \g224/_0_ , \g22412/_0_ , \g22415/_1__syn_2 , \g225/_0_ , \g2257/_0_ , \g226/_3_ , \g22624/_0_ , \g227/_3_ , \g22702/_0_ , \g22919/_1__syn_2 , \g22933/_0_ , \g22954/_0_ , \g22989/_1_ , \g23529/_0_ , \g23539/_0_ , \g2362/_2_ , \g23766/_0_ , \g24/_3_ , \g24018/_0_ , \g2416/_0_ , \g2420/_0_ , \g24213/_0_ , \g24301/_0_ , \g2479/_0_ , \g248/_3_ , \g2480/_0_ , \g2481/_0_ , \g2482/_0_ , \g2483/_0_ , \g2484/_0_ , \g2485/_0_ , \g2486/_0_ , \g2487/_0_ , \g2488/_0_ , \g249/_3_ , \g2490/_0_ , \g2491/_0_ , \g2492/_0_ , \g2493/_0_ , \g2494/_0_ , \g2495/_0_ , \g2496/_0_ , \g2497/_0_ , \g2507/_0_ , \g2508/_0_ , \g2509/_0_ , \g2510/_0_ , \g2511/_0_ , \g2512/_0_ , \g2513/_0_ , \g2514/_0_ , \g2515/_0_ , \g2516/_0_ , \g25237/_0_ , \g2558/_0_ , \g2562/_0_ , \g2563/_0_ , \g2564/_0_ , \g2565/_0_ , \g2566/_0_ , \g2567/_0_ , \g2699/_0_ , \g27/_2_ , \g271/_0_ , \g272/_3_ , \g273/_3_ , \g274/_3_ , \g275/_3_ , \g276/_3_ , \g277/_3_ , \g2787/_3_ , \g2788/_3_ , \g279/_0_ , \g2795/_0_ , \g2796/_0_ , \g280/_0_ , \g2842/_3_ , \g29/_1_ , \g2927/_0_ , \g2978/_0_ , \g2979/_0_ , \g2980/_0_ , \g2981/_0_ , \g2982/_0_ , \g2983/_0_ , \g2984/_0_ , \g2985/_0_ , \g3021/_3_ , \g3022/_3_ , \g3023/_3_ , \g3024/_3_ , \g3025/_3_ , \g3026/_3_ , \g3027/_3_ , \g3028/_3_ , \g3029/_3_ , \g3030/_3_ , \g3031/_3_ , \g3032/_3_ , \g3033/_3_ , \g3034/_3_ , \g3035/_3_ , \g3036/_3_ , \g3037/_3_ , \g3038/_3_ , \g3039/_3_ , \g3040/_3_ , \g3041/_3_ , \g3042/_3_ , \g3049/_0_ , \g3050/_0_ , \g3051/_0_ , \g3052/_0_ , \g3053/_0_ , \g3054/_0_ , \g3058/_0_ , \g3059/_0_ , \g3088/_0_ , \g3089/_0_ , \g3090/_0_ , \g3091/_0_ , \g3092/_0_ , \g3093/_0_ , \g3094/_0_ , \g3095/_0_ , \g314/_0_ , \g3147/_3_ , \g3148/_3_ , \g3189/_0_ , \g3190/_0_ , \g3191/_0_ , \g3192/_0_ , \g3193/_0_ , \g3194/_0_ , \g3195/_0_ , \g3196/_0_ , \g3197/_0_ , \g3198/_0_ , \g3199/_0_ , \g32/_0_ , \g320/_3_ , \g3200/_0_ , \g3201/_0_ , \g3202/_0_ , \g3203/_0_ , \g3204/_0_ , \g321/_3_ , \g325/_3_ , \g3271/_2_ , \g33/_0_ , \g3363/_0_ , \g3413/_0_ , \g3414/_0_ , \g352/_0_ , \g355/_0_ , \g356/_3_ , \g357/_3_ , \g35_dup/_1_ , \g36/_3_ , \g365/_3_ , \g366/_3_ , \g367/_3_ , \g368/_3_ , \g3687/_0_ , \g369/_3_ , \g37/_3_ , \g370/_3_ , \g372/_3_ , \g374/_3_ , \g3740/_0_ , \g375/_3_ , \g376/_3_ , \g3878/_0_ , \g3879/_0_ , \g388/_3_ , \g3880/_0_ , \g3881/_0_ , \g3882/_0_ , \g389/_3_ , \g3894/_0_ , \g3895/_0_ , \g3896/_0_ , \g3897/_0_ , \g3898/_0_ , \g392/_3_ , \g393/_3_ , \g394/_3_ , \g395/_3_ , \g396/_3_ , \g397/_3_ , \g398/_3_ , \g399/_3_ , \g401/_3_ , \g402/_3_ , \g404/_3_ , \g4048/_0_ , \g405/_3_ , \g4050/_0_ , \g406/_3_ , \g407/_3_ , \g410/_3_ , \g411/_3_ , \g412/_3_ , \g413/_3_ , \g415/_3_ , \g416/_3_ , \g42/_0_ , \g4216/_3_ , \g4217/_3_ , \g4218/_3_ , \g4219/_3_ , \g4296/_0_ , \g4297/_0_ , \g4298/_0_ , \g4299/_0_ , \g43/_0_ , \g4300/_0_ , \g4301/_0_ , \g4302/_0_ , \g4303/_0_ , \g4304/_0_ , \g4305/_0_ , \g4306/_0_ , \g4307/_0_ , \g4308/_0_ , \g4309/_0_ , \g4310/_0_ , \g4311/_0_ , \g4312/_0_ , \g4313/_0_ , \g4314/_0_ , \g4315/_0_ , \g4316/_0_ , \g4317/_0_ , \g4318/_0_ , \g4319/_0_ , \g4320/_0_ , \g4321/_0_ , \g4322/_0_ , \g4323/_0_ , \g436/_0_ , \g44/_0_ , \g448/_3_ , \g45/_0_ , \g4587/_0_ , \g4588/_0_ , \g46/_0_ , \g4601/_0_ , \g4602/_0_ , \g4613/_3_ , \g4614/_3_ , \g4615/_3_ , \g463/_0_ , \g465/_0_ , \g4653/_0_ , \g4654/_0_ , \g4655/_0_ , \g4656/_0_ , \g4659/_0_ , \g466/_0_ , \g468/_3_ , \g469/_3_ , \g4697/_0_ , \g47/_3_ , \g470/_0_ , \g471/_0_ , \g4755/_0_ , \g476/_0_ , \g48/_3_ , \g480/_00_ , \g4839/_0_ , \g4840/_0_ , \g485/_3_ , \g4854/_0_ , \g4855/_0_ , \g4859/_0_ , \g486/_3_ , \g4860/_0_ , \g4880/_0_ , \g4881/_0_ , \g4882/_0_ , \g4883/_0_ , \g4884/_0_ , \g4885/_0_ , \g4886/_0_ , \g4887/_0_ , \g4888/_0_ , \g49/_0_ , \g494/_0_ , \g499/_1_ , \g50/_0_ , \g5002/_0_ , \g5003/_0_ , \g5009/_0_ , \g5010/_0_ , \g5011/_0_ , \g5014/_0_ , \g51/_0_ , \g5105/_0_ , \g5129/_2_ , \g5132/_0_ , \g5135/_0_ , \g5168/_0_ , \g5169/_0_ , \g5173/_0_ , \g5224/_0_ , \g5225/_0_ , \g5226/_0_ , \g5227/_0_ , \g5334/_0_ , \g5335/_0_ , \g5336/_0_ , \g5337/_0_ , \g5338/_0_ , \g5339/_0_ , \g5340/_0_ , \g5341/_0_ , \g5342/_0_ , \g5343/_0_ , \g5344/_0_ , \g5345/_0_ , \g5346/_0_ , \g5347/_0_ , \g5348/_0_ , \g5349/_0_ , \g5395/_0_ , \g54/_0_ , \g5434/_0_ , \g5447/_0_ , \g5450/_0_ , \g5451/_0_ , \g5452/_0_ , \g5453/_0_ , \g5454/_0_ , \g5461/_0_ , \g5483/_0_ , \g5484/_0_ , \g5492/_0_ , \g5493/_0_ , \g5496/_3_ , \g5497/_3_ , \g55/_0_ , \g5500/_0_ , \g5502/_0_ , \g5503/_0_ , \g5506/_0_ , \g5511/_0_ , \g5518/_0_ , \g5519/_0_ , \g5520/_0_ , \g5522/_0_ , \g5523/_0_ , \g5524/_0_ , \g5525/_0_ , \g5532/_0_ , \g5533/_0_ , \g5534/_0_ , \g5535/_0_ , \g5536/_0_ , \g5537/_0_ , \g5538/_0_ , \g5546/_0_ , \g5555/_00_ , \g5593/_0_ , \g5614/_2_ , \g567/_0_ , \g5677/_0_ , \g5678/_0_ , \g5682/_0_ , \g5683/_0_ , \g5684/_0_ , \g5686/_0_ , \g5687/_0_ , \g5689/_0_ , \g5690/_0_ , \g5691/_0_ , \g5692/_0_ , \g5698/_0_ , \g5699/_0_ , \g5700/_0_ , \g5701/_0_ , \g5702/_0_ , \g5703/_0_ , \g5704/_0_ , \g5709/_0_ , \g5711/_0_ , \g5714/_0_ , \g572/_0_ , \g5723/_0_ , \g5724/_0_ , \g5725/_0_ , \g573/_0_ , \g5739/_0_ , \g5740/_0_ , \g575/_0_ , \g5756/_0_ , \g5757/_0_ , \g5758/_0_ , \g5759/_0_ , \g576/_0_ , \g5760/_0_ , \g5761/_0_ , \g5762/_0_ , \g5763/_0_ , \g577/_0_ , \g5772/_0_ , \g5773/_0_ , \g5774/_0_ , \g5775/_0_ , \g5776/_0_ , \g5777/_0_ , \g578/_0_ , \g5781/_0_ , \g5783/_0_ , \g5784/_0_ , \g5785/_0_ , \g5786/_0_ , \g5787/_0_ , \g5788/_0_ , \g5789/_0_ , \g579/_0_ , \g5790/_0_ , \g5791/_0_ , \g5792/_0_ , \g5794/_0_ , \g5795/_0_ , \g5796/_0_ , \g580/_0_ , \g5801/_0_ , \g5802/_0_ , \g5803/_0_ , \g5804/_0_ , \g5805/_0_ , \g581/_0_ , \g5814/_0_ , \g582/_0_ , \g583/_0_ , \g5849/_3_ , \g585/_0_ , \g586/_0_ , \g587/_0_ , \g588/_0_ , \g589/_0_ , \g590/_0_ , \g591/_0_ , \g592/_0_ , \g593/_0_ , \g594/_0_ , \g595/_0_ , \g596/_0_ , \g597/_0_ , \g5971/_0_ , \g5972/_0_ , \g5976/_0_ , \g598/_0_ , \g5989/_0_ , \g599/_0_ , \g600/_0_ , \g601/_0_ , \g602/_0_ , \g603/_0_ , \g604/_0_ , \g605/_0_ , \g6092/_0_ , \g6093/_2_ , \g6094/_0_ , \g6114/_0_ , \g614/_3_ , \g6148/_0_ , \g6149/_0_ , \g6171/_0_ , \g6172/_0_ , \g6173/_0_ , \g6174/_0_ , \g6175/_0_ , \g6176/_0_ , \g6177/_0_ , \g6178/_0_ , \g6179/_0_ , \g6180/_0_ , \g6181/_0_ , \g6182/_0_ , \g6183/_0_ , \g6184/_0_ , \g6185/_0_ , \g6186/_0_ , \g6187/_0_ , \g6193/_0_ , \g6196/_0_ , \g6197/_0_ , \g6198/_3_ , \g6200/_2_ , \g6202/_2_ , \g6203/_3_ , \g6204/_3_ , \g6209/_0_ , \g6211/_0_ , \g6215/_0_ , \g6217/_0_ , \g6219/_0_ , \g6220/_0_ , \g6222/_0_ , \g6224/_0_ , \g6228/_0_ , \g6238/_0_ , \g6239/_0_ , \g6240/_0_ , \g6242/_0_ , \g6243/_0_ , \g6244/_0_ , \g6245/_0_ , \g6246/_0_ , \g6248/_0_ , \g6249/_0_ , \g6259/_0_ , \g6260/_0_ , \g6261/_0_ , \g6262/_0_ , \g6263/_0_ , \g6264/_0_ , \g6265/_0_ , \g6266/_0_ , \g6267/_0_ , \g6268/_0_ , \g6269/_0_ , \g6270/_0_ , \g6271/_0_ , \g6272/_0_ , \g6277/_0_ , \g6318/_0_ , \g6326/_0_ , \g6329/_0_ , \g6330/_0_ , \g6331/_0_ , \g6332/_0_ , \g6333/_0_ , \g6334/_0_ , \g6335/_0_ , \g6336/_0_ , \g6337/_0_ , \g6338/_0_ , \g6339/_0_ , \g6340/_0_ , \g6341/_0_ , \g6342/_0_ , \g6343/_0_ , \g6344/_0_ , \g6345/_0_ , \g6346/_0_ , \g6347/_0_ , \g6348/_0_ , \g6349/_0_ , \g6350/_0_ , \g6351/_0_ , \g6352/_0_ , \g6353/_0_ , \g6354/_0_ , \g6355/_0_ , \g6361/_0_ , \g637/_0_ , \g638/_0_ , \g639/_3_ , \g64/_3_ , \g640/_3_ , \g6419/_0_ , \g6442/_0_ , \g6442/_1_ , \g6489/_0_ , \g6490/_0_ , \g65/_3_ , \g6513/_0_ , \g6515/_0_ , \g6571/_0_ , \g6588/_0_ , \g6589/_0_ , \g6638/_0_ , \g6639/_0_ , \g6653/_0_ , \g6654/_3_ , \g6655/_0_ , \g6656/_0_ , \g6657/_0_ , \g6687/_0_ , \g6688/_0_ , \g6689/_0_ , \g6690/_0_ , \g6691/_0_ , \g6692/_0_ , \g6693/_0_ , \g6694/_0_ , \g6701/_0_ , \g6706/_0_ , \g6711/_0_ , \g6727/_0_ , \g6728/_0_ , \g6736/_0_ , \g6739/_0_ , \g6742/_0_ , \g6746/_0_ , \g6752/_0_ , \g6771/_0_ , \g684/_0_ , \g685/_0_ , \g686/_0_ , \g687/_0_ , \g688/_0_ , \g689/_0_ , \g690/_0_ , \g691/_0_ , \g692/_0_ , \g693/_0_ , \g696/_3_ , \g697/_3_ , \g699/_0_ , \g7/_0_ , \g700/_0_ , \g7005/_0_ , \g7056/_0_ , \g7057/_0_ , \g7058/_0_ , \g7060/_0_ , \g7075/_0_ , \g7086/_0_ , \g7087/_0_ , \g7089/_0_ , \g7108/_0_ , \g7109/_0_ , \g7112/_0_ , \g7172/_2_ , \g7210/_2_ , \g7211/_0_ , \g7212/_0_ , \g7213/_0_ , \g7214/_0_ , \g7215/_0_ , \g7216/_0_ , \g7217/_3_ , \g7218/_0_ , \g7219/_0_ , \g7220/_0_ , \g7222/_0_ , \g7227/_2_ , \g723/_3_ , \g7234/_0_ , \g7237/_3_ , \g7238/_3_ , \g7239/_3_ , \g724/_3_ , \g7240/_3_ , \g7241/_3_ , \g7242/_3_ , \g7243/_3_ , \g7244/_0_ , \g7245/_0_ , \g7246/_0_ , \g7247/_0_ , \g7248/_0_ , \g7249/_0_ , \g7250/_0_ , \g7251/_0_ , \g7253/_0_ , \g7254/_0_ , \g7255/_0_ , \g7256/_0_ , \g7257/_0_ , \g7258/_0_ , \g7261/_0_ , \g7264/_0_ , \g7265/_0_ , \g7266/_0_ , \g7267/_0_ , \g7268/_0_ , \g7269/_0_ , \g7278/_0_ , \g7279/_0_ , \g7280/_0_ , \g7281/_0_ , \g7282/_0_ , \g7283/_0_ , \g7284/_0_ , \g7285/_0_ , \g7286/_3_ , \g7288/_3_ , \g7291/_0_ , \g7296/_3_ , \g73/_0_ , \g7302/_3_ , \g7306/_3_ , \g7310/_3_ , \g7311/_3_ , \g7312/_3_ , \g7313/_3_ , \g7314/_3_ , \g7315/_3_ , \g7316/_3_ , \g7317/_3_ , \g7323/_3_ , \g7324/_3_ , \g7325/_3_ , \g7327/_0_ , \g7362/_0_ , \g74/_0_ , \g75/_0_ , \g7512/_0_ , \g7513/_0_ , \g7514/_0_ , \g7515/_0_ , \g7516/_0_ , \g7518/_0_ , \g7528/_0_ , \g7529/_0_ , \g7548/_0_ , \g7549/_0_ , \g7550/_0_ , \g7575/_0_ , \g7576/_0_ , \g7577/_0_ , \g7578/_0_ , \g7579/_0_ , \g7580/_0_ , \g7581/_0_ , \g7582/_0_ , \g7583/_0_ , \g7584/_0_ , \g7585/_0_ , \g7586/_0_ , \g7587/_0_ , \g7588/_0_ , \g7589/_0_ , \g7590/_0_ , \g7591/_0_ , \g7592/_0_ , \g7593/_0_ , \g7594/_0_ , \g7595/_0_ , \g7596/_0_ , \g7597/_0_ , \g7598/_0_ , \g7599/_0_ , \g76/_0_ , \g7600/_0_ , \g7601/_0_ , \g7602/_0_ , \g7603/_0_ , \g7604/_0_ , \g7614/_0_ , \g7618/_0_ , \g762/_0_ , \g7634/_0_ , \g766/_0_ , \g767/_0_ , \g768/_0_ , \g769/_0_ , \g77/_0_ , \g770/_3_ , \g771/_3_ , \g7715/_0_ , \g774/_0_ , \g7746/_0_ , \g7753/_0_ , \g7754/_0_ , \g7755/_0_ , \g7756/_0_ , \g7757/_0_ , \g7758/_0_ , \g7759/_0_ , \g7760/_0_ , \g7761/_0_ , \g7762/_0_ , \g7763/_0_ , \g7764/_0_ , \g7765/_0_ , \g7766/_0_ , \g7778/_0_ , \g7779/_0_ , \g7780/_0_ , \g7781/_0_ , \g7782/_0_ , \g7784/_0_ , \g78/_0_ , \g7800/_0_ , \g7823/_3_ , \g7837/_0_ , \g7841/_0_ , \g7842/_0_ , \g7843/_0_ , \g7844/_0_ , \g7845/_0_ , \g7846/_0_ , \g7847/_0_ , \g7849/_0_ , \g7850/_0_ , \g7852/_0_ , \g7854/_0_ , \g7855/_0_ , \g7857/_0_ , \g7858/_0_ , \g7859/_0_ , \g7860/_0_ , \g7861/_0_ , \g7862/_0_ , \g7863/_0_ , \g7864/_0_ , \g7865/_0_ , \g7866/_0_ , \g7867/_0_ , \g7868/_0_ , \g7869/_0_ , \g7870/_0_ , \g7871/_0_ , \g79211/_3_ , \g79258/_3_ , \g79299/_3_ , \g79316/_2_ , \g79342/_3_ , \g79401/_3_ , \g79452/_3_ , \g79457/_3_ , \g7951/_0_ , \g79541/_3_ , \g7958/_0_ , \g79598/_3_ , \g79654/_3_ , \g79675/_3_ , \g7971/_0_ , \g7972/_0_ , \g7973/_3_ , \g79753/_3_ , \g7976/_3_ , \g79855/_3_ , \g79858/_3_ , \g79997/_3_ , \g8/_0_ , \g80008/_3_ , \g80011/_0_ , \g80104/_0_ , \g80172/_1_ , \g80195/_3_ , \g80238/_3_ , \g80290/_2_ , \g80294/_0_ , \g80302/_0_ , \g80327/_0_ , \g80360/_3_ , \g80373/_0_ , \g80401/_0_ , \g80410/_0_ , \g80475/_0_ , \g80476/_0_ , \g80516/_3_ , \g80536/_0_ , \g80537/_0_ , \g80572/_0_ , \g80573/_0_ , \g80609/_2_ , \g80610/_2_ , \g80676/_0_ , \g80798/_0_ , \g80807/_0_ , \g80890/_2_ , \g80904/_0_ , \g81719/_2_ , \g81746/_0_ , \g81775/_0_ , \g81872/_0_ , \g81961/_0_ , \g81968/_0_ , \g82096/_0_ , \g82123/_0_ , \g82147/_0_ , \g82147/_1_ , \g82335/_0_ , \g82338/_2_ , \g82368/_0_ , \g82460/_2_ , \g82469/_0_ , \g82481/_0_ , \g82625/_1_ , \g82711/_0_ , \g82772/_0_ , \g82946/_0_ , \g82947/_0_ , \g82956/_0_ , \g83003/_0_ , \g83006/_1_ , \g83415/_0_ , \g83498/_0_ , \g837/_0_ , \g838/_0_ , \g83863/_0_ , \g839/_0_ , \g84049/_3_ , \g84050/_3_ , \g84077/_2_ , \g842/_0_ , \g84245/_0_ , \g843/_0_ , \g844/_0_ , \g84448/_0_ , \g84478/_3_ , \g845/_0_ , \g846/_0_ , \g847/_0_ , \g848/_0_ , \g8487/_0_ , \g8488/_0_ , \g8489/_0_ , \g849/_0_ , \g8490/_0_ , \g84904/_0_ , \g8491/_0_ , \g8492/_0_ , \g8493/_0_ , \g8494/_0_ , \g8496/_0_ , \g8517/_0_ , \g8534/_0_ , \g8538/_0_ , \g8540/_0_ , \g8576/_2_ , \g8597/_0_ , \g8598/_0_ , \g8599/_0_ , \g8600/_0_ , \g8601/_0_ , \g8602/_0_ , \g8603/_0_ , \g8605/_0_ , \g8606/_0_ , \g8607/_0_ , \g8608/_0_ , \g8609/_0_ , \g8610/_0_ , \g8611/_0_ , \g8612/_0_ , \g8613/_0_ , \g8614/_0_ , \g8615/_0_ , \g8617/_0_ , \g8643/_0_ , \g8644/_0_ , \g8645/_0_ , \g8646/_0_ , \g8647/_0_ , \g8648/_0_ , \g8650/_0_ , \g8651/_0_ , \g8652/_0_ , \g8653/_0_ , \g8654/_0_ , \g8655/_0_ , \g8656/_0_ , \g8657/_0_ , \g8658/_0_ , \g8659/_0_ , \g8660/_0_ , \g8665/_00_ , \g8666/_00_ , \g8667/_00_ , \g8668/_00_ , \g8669/_00_ , \g86715/_0_ , \g86745/_3_ , \g8691/_0_ , \g8700/_0_ , \g8701/_0_ , \g8702/_0_ , \g8703/_0_ , \g8704/_0_ , \g8705/_0_ , \g87063/_0_ , \g87114/_0_ , \g8712/_0_ , \g8713/_0_ , \g8714/_0_ , \g87171/_1_ , \g87252/_1_ , \g87298/_0_ , \g8730/_0_ , \g8741/_0_ , \g8747/_0_ , \g87480/_0_ , \g87484/_2_ , \g87488/_1__syn_2 , \g8761/_0_ , \g8762/_0_ , \g8763/_0_ , \g8764/_0_ , \g8765/_0_ , \g8775/_0_ , \g8776/_0_ , \g8777/_0_ , \g8778/_0_ , \g8784/_0_ , \g8804/_0_ , \g8807/_0_ , \g8808/_0_ , \g8809/_0_ , \g8810/_0_ , \g8811/_0_ , \g8812/_0_ , \g8813/_0_ , \g8814/_0_ , \g8815/_0_ , \g8816/_0_ , \g8817/_0_ , \g8818/_0_ , \g8819/_0_ , \g8820/_0_ , \g8821/_0_ , \g8822/_0_ , \g8823/_0_ , \g8824/_0_ , \g8825/_0_ , \g8826/_0_ , \g8827/_0_ , \g8828/_0_ , \g8829/_0_ , \g8830/_0_ , \g8831/_0_ , \g8832/_0_ , \g8833/_0_ , \g8834/_0_ , \g8835/_0_ , \g8836/_0_ , \g8837/_0_ , \g8838/_0_ , \g8839/_0_ , \g8840/_0_ , \g8842/_0_ , \g8843/_0_ , \g8846/_0_ , \g8848/_0_ , \g8857/_0_ , \g8895/_0_ , \g8902/_3_ , \g8903/_3_ , \g8904/_3_ , \g8905/_3_ , \g8906/_3_ , \g8909/_0_ , \g8910/_0_ , \g8911/_0_ , \g8924/_3_ , \g8926/_3_ , \g8927/_3_ , \g8943/_0_ , \g8944/_0_ , \g8958/_3_ , \g8960/_00_ , \g8961/_3_ , \g8965/_0_ , \g8966/_0_ , \g8967/_0_ , \g8968/_0_ , \g9/_0_ , \g9123/_0_ , \g9125/_0_ , \g9126/_0_ , \g913/_0_ , \g915/_0_ , \g916/_0_ , \g917/_0_ , \g918/_0_ , \g919/_0_ , \g920/_3_ , \g921/_3_ , \g925/_0_ , \g926/_0_ , \g927/_0_ , \g928/_0_ , \g929/_0_ , \g930/_0_ , \g9336/_0_ , \g9337/_0_ , \g939/_3_ , \g9396/_0_ , \g9397/_0_ , \g9399/_0_ , \g9400/_0_ , \g9401/_0_ , \g9402/_0_ , \g9403/_0_ , \g9404/_0_ , \g9415/_0_ , \g9418/_0_ , \g9419/_0_ , \g9420/_0_ , \g9446/_0_ , \g9465/_0_ , \g9493/_0_ , \g9536/_0_ , \g9537/_0_ , \g9538/_0_ , \g9539/_0_ , \g9540/_0_ , \g9541/_0_ , \g9542/_0_ , \g955/_2_ , \g9561/_0_ , \g9562/_0_ , \g9563/_0_ , \g9564/_0_ , \g9565/_0_ , \g9566/_0_ , \g9567/_0_ , \g9568/_0_ , \g9569/_0_ , \g9570/_0_ , \g9571/_0_ , \g9572/_0_ , \g9573/_0_ , \g9574/_0_ , \g9575/_0_ , \g9576/_0_ , \g9577/_0_ , \g9578/_0_ , \g9579/_0_ , \g9580/_0_ , \g9581/_0_ , \g9582/_0_ , \g9583/_0_ , \g9584/_0_ , \g9585/_0_ , \g9586/_0_ , \g9587/_0_ , \g9588/_0_ , \g9589/_0_ , \g9590/_0_ , \g9591/_0_ , \g9592/_0_ , \g9593/_0_ , \g9594/_0_ , \g9595/_0_ , \g9596/_0_ , \g9597/_0_ , \g9598/_0_ , \g9599/_0_ , \g9600/_0_ , \g9601/_0_ , \g9602/_0_ , \g9603/_0_ , \g9604/_0_ , \g9605/_0_ , \g9606/_0_ , \g9607/_0_ , \g9608/_0_ , \g9609/_0_ , \g9610/_0_ , \g9611/_0_ , \g9612/_0_ , \g9613/_0_ , \g9614/_0_ , \g9615/_0_ , \g9616/_0_ , \g9617/_0_ , \g9618/_0_ , \g9619/_0_ , \g9620/_0_ , \g9621/_0_ , \g9622/_0_ , \g9623/_0_ , \g9624/_0_ , \g9625/_0_ , \g9626/_0_ , \g9627/_0_ , \g9628/_0_ , \g9629/_0_ , \g9630/_0_ , \g9631/_0_ , \g9632/_0_ , \g9633/_0_ , \g9634/_0_ , \g9635/_0_ , \g9636/_0_ , \g9637/_0_ , \g9638/_0_ , \g9639/_0_ , \g9640/_0_ , \g9641/_0_ , \g9642/_0_ , \g9643/_0_ , \g9644/_0_ , \g9645/_0_ , \g9646/_0_ , \g9647/_0_ , \g9648/_0_ , \g9649/_0_ , \g9650/_0_ , \g9651/_0_ , \g9652/_0_ , \g9653/_0_ , \g9654/_0_ , \g9655/_0_ , \g9656/_0_ , \g9657/_0_ , \g9658/_0_ , \g9659/_0_ , \g9660/_0_ , \g9661/_0_ , \g9662/_0_ , \g9663/_0_ , \g9664/_0_ , \g9665/_0_ , \g9666/_0_ , \g9667/_0_ , \g9668/_0_ , \g9669/_0_ , \g9670/_0_ , \g9671/_0_ , \g9672/_0_ , \g9673/_0_ , \g9674/_0_ , \g9675/_0_ , \g9676/_0_ , \g9677/_0_ , \g9678/_0_ , \g9681/_0_ , \g9683/_0_ , \g9689/_0_ , \g9692/_0_ , \g9694/_0_ , \g9695/_0_ , \g9701/_0_ , \g9702/_0_ , \g9703/_0_ , \g9704/_0_ , \g9709/_0_ , \g9710/_0_ , \g9711/_0_ , \g9712/_0_ , \g9720/_0_ , \g9721/_0_ , \g9722/_0_ , \g9726/_0_ , \g9733/_0_ , \g9734/_0_ , \g9735/_0_ , \g9736/_0_ , \g9737/_0_ , \g9738/_0_ , \g9739/_0_ , \g9740/_0_ , \g9741/_0_ , \g9742/_0_ , \g9743/_0_ , \g9744/_0_ , \g9745/_0_ , \g9746/_0_ , \g9747/_0_ , \g9748/_0_ , \g9749/_0_ , \g9750/_0_ , \g9751/_0_ , \g9752/_0_ , \g9753/_0_ , \g9754/_0_ , \g9755/_0_ , \g9756/_0_ , \g9757/_0_ , \g9758/_0_ , \g9759/_0_ , \g9760/_0_ , \g9761/_0_ , \g9762/_0_ , \g9763/_0_ , \g9764/_0_ , \g9765/_0_ , \g9766/_0_ , \g9767/_0_ , \g9768/_0_ , \g9769/_0_ , \g9770/_0_ , \g9771/_0_ , \g9772/_0_ , \g9773/_0_ , \g9774/_0_ , \g9775/_0_ , \g9776/_0_ , \g9777/_0_ , \g9778/_0_ , \g9779/_0_ , \g9780/_0_ , \g9781/_0_ , \g9782/_0_ , \g9783/_0_ , \g9784/_0_ , \g9785/_0_ , \g9786/_0_ , \g9787/_0_ , \g9788/_0_ , \g9789/_0_ , \g9790/_0_ , \g9791/_0_ , \g9792/_0_ , \g9793/_0_ , \g9794/_0_ , \g9795/_0_ , \g9796/_0_ , \g9797/_0_ , \g9798/_0_ , \g9799/_0_ , \g9800/_0_ , \g9801/_0_ , \g9802/_0_ , \g9803/_0_ , \g9804/_0_ , \g9805/_0_ , \g9806/_0_ , \g9807/_0_ , \g9808/_0_ , \g9809/_0_ , \g9810/_0_ , \g9811/_0_ , \g9812/_0_ , \g9813/_0_ , \g9814/_0_ , \g9815/_0_ , \g9816/_0_ , \g9817/_0_ , \g9818/_0_ , \g9819/_0_ , \g9820/_0_ , \g9821/_0_ , \g9822/_0_ , \g9823/_0_ , \g9824/_0_ , \g9825/_0_ , \g9826/_0_ , \g9827/_0_ , \g9828/_0_ , \g9829/_0_ , \g9830/_0_ , \g9831/_0_ , \g9832/_0_ , \g9833/_0_ , \g9835/_0_ , \g9836/_0_ , \g9837/_0_ , \g9838/_0_ , \g9839/_0_ , \g9840/_0_ , \g9841/_0_ , \g9842/_0_ , \g9844/_0_ , \g9845/_0_ , \g9846/_0_ , \g9848/_0_ , \g9849/_0_ , \g9850/_0_ , \g9851/_0_ , \g9853/_0_ , \g9854/_0_ , \g9855/_0_ , \g9856/_0_ , \g9857/_0_ , \g9858/_0_ , \g9859/_0_ , \g9860/_0_ , \g9862/_0_ , \g9863/_0_ , \g9864/_0_ , \g9865/_0_ , \g9867/_0_ , \g9868/_0_ , \g9876/_0_ , \g9877/_0_ , \g9878/_0_ , \g9879/_0_ , \g9880/_0_ , \g9881/_0_ , \g9898/_0_ , \g9900/_0_ , \g9901/_0_ , \g9902/_0_ , \g9903/_0_ , \g9904/_0_ , \g9905/_0_ , \g9906/_0_ , \g9907/_0_ , \g9908/_0_ , \g9909/_0_ , \g9910/_0_ , \g9911/_0_ , \g9912/_0_ , \g9913/_0_ , \g9914/_0_ , \g9915/_0_ , \g9916/_0_ , \g9917/_0_ , \g9918/_0_ , \g9919/_0_ , \g992/_0_ , \g9920/_0_ , \g9921/_0_ , \g9922/_0_ , \g9923/_0_ , \g9924/_0_ , \g9925/_0_ , \g9926/_0_ , \g9927/_0_ , \g9928/_0_ , \g9929/_0_ , \g9930/_0_ , \g9931/_0_ , \g9932/_0_ , \g9933/_0_ , \g9934/_0_ , \g9935/_0_ , \g9936/_0_ , \g9937/_0_ , \g9938/_0_ , \g9939/_0_ , \g9940/_0_ , \g9941/_0_ , \g9942/_0_ , \g9943/_0_ , \g9944/_0_ , \g9945/_0_ , \g9946/_0_ , \g9947/_0_ , \g9948/_0_ , \g9949/_0_ , \g9950/_0_ , \g9951/_0_ , \g9952/_0_ , \g9953/_0_ , \g9954/_0_ , \g9955/_0_ , \g9956/_0_ , \g9957/_0_ , \g9958/_0_ , \g9959/_0_ , \g9960/_0_ , \g9961/_0_ , \g9962/_0_ , \g9963/_0_ , \g9964/_0_ , \g9965/_0_ , \g9966/_0_ , \g9967/_0_ , \g9968/_0_ , \g9969/_0_ , \g9970/_0_ , \g9971/_0_ , \g9972/_0_ , \g9973/_0_ , \g9974/_0_ , \g9975/_0_ , \g9976/_0_ , \g9977/_0_ , \g9978/_0_ , \g9979/_0_ , \g9980/_0_ , \g9981/_0_ , \g9982/_0_ , \g9983/_0_ , \g9984/_0_ , \g9985/_0_ , \g9987/_0_ , \g9988/_0_ , \g9989/_0_ , \g999/_0_ , \g9990/_0_ , \g9991/_0_ , \g9992/_0_ , \g9993/_0_ , \g9994/_0_ , \g9995/_0_ , \g9996/_0_ , \g9997/_0_ , \g9998/_0_ , \g9999/_0_ , \idma_IDMA_boot_reg/NET0131_reg_syn_3 , \memc_EXTC_Eg_reg/NET0131 , \memc_EXTC_Eg_reg/NET0131_reg_syn_3 , \memc_EXTC_Eg_reg/n0 , \pio_PIO_IN_P_reg[0]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[10]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[11]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[1]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[2]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[3]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[4]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[5]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[6]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[7]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[8]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[9]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[0]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[10]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[2]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[4]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[6]/P0001_reg_syn_3 , \sice_GO_NXi_reg/NET0131_reg_syn_3 , \sport0_rxctl_RXSHT_reg[0]/P0001_reg_syn_3 , \sport0_rxctl_RXSHT_reg[1]/P0001_reg_syn_3 , \sport1_rxctl_RXSHT_reg[0]/P0001_reg_syn_3 , \sport1_rxctl_RXSHT_reg[1]/P0001_reg_syn_3 );
	input \CM_rd0[0]_pad  ;
	input \CM_rd0[10]_pad  ;
	input \CM_rd0[11]_pad  ;
	input \CM_rd0[12]_pad  ;
	input \CM_rd0[13]_pad  ;
	input \CM_rd0[14]_pad  ;
	input \CM_rd0[15]_pad  ;
	input \CM_rd0[16]_pad  ;
	input \CM_rd0[17]_pad  ;
	input \CM_rd0[18]_pad  ;
	input \CM_rd0[19]_pad  ;
	input \CM_rd0[1]_pad  ;
	input \CM_rd0[20]_pad  ;
	input \CM_rd0[21]_pad  ;
	input \CM_rd0[22]_pad  ;
	input \CM_rd0[23]_pad  ;
	input \CM_rd0[2]_pad  ;
	input \CM_rd0[3]_pad  ;
	input \CM_rd0[4]_pad  ;
	input \CM_rd0[5]_pad  ;
	input \CM_rd0[6]_pad  ;
	input \CM_rd0[7]_pad  ;
	input \CM_rd0[8]_pad  ;
	input \CM_rd0[9]_pad  ;
	input \CM_rd1[0]_pad  ;
	input \CM_rd1[10]_pad  ;
	input \CM_rd1[11]_pad  ;
	input \CM_rd1[12]_pad  ;
	input \CM_rd1[13]_pad  ;
	input \CM_rd1[14]_pad  ;
	input \CM_rd1[15]_pad  ;
	input \CM_rd1[16]_pad  ;
	input \CM_rd1[17]_pad  ;
	input \CM_rd1[18]_pad  ;
	input \CM_rd1[19]_pad  ;
	input \CM_rd1[1]_pad  ;
	input \CM_rd1[20]_pad  ;
	input \CM_rd1[21]_pad  ;
	input \CM_rd1[22]_pad  ;
	input \CM_rd1[23]_pad  ;
	input \CM_rd1[2]_pad  ;
	input \CM_rd1[3]_pad  ;
	input \CM_rd1[4]_pad  ;
	input \CM_rd1[5]_pad  ;
	input \CM_rd1[6]_pad  ;
	input \CM_rd1[7]_pad  ;
	input \CM_rd1[8]_pad  ;
	input \CM_rd1[9]_pad  ;
	input \CM_rd2[0]_pad  ;
	input \CM_rd2[10]_pad  ;
	input \CM_rd2[11]_pad  ;
	input \CM_rd2[12]_pad  ;
	input \CM_rd2[13]_pad  ;
	input \CM_rd2[14]_pad  ;
	input \CM_rd2[15]_pad  ;
	input \CM_rd2[16]_pad  ;
	input \CM_rd2[17]_pad  ;
	input \CM_rd2[18]_pad  ;
	input \CM_rd2[19]_pad  ;
	input \CM_rd2[1]_pad  ;
	input \CM_rd2[20]_pad  ;
	input \CM_rd2[21]_pad  ;
	input \CM_rd2[22]_pad  ;
	input \CM_rd2[23]_pad  ;
	input \CM_rd2[2]_pad  ;
	input \CM_rd2[3]_pad  ;
	input \CM_rd2[4]_pad  ;
	input \CM_rd2[5]_pad  ;
	input \CM_rd2[6]_pad  ;
	input \CM_rd2[7]_pad  ;
	input \CM_rd2[8]_pad  ;
	input \CM_rd2[9]_pad  ;
	input \CM_rd3[0]_pad  ;
	input \CM_rd3[10]_pad  ;
	input \CM_rd3[11]_pad  ;
	input \CM_rd3[12]_pad  ;
	input \CM_rd3[13]_pad  ;
	input \CM_rd3[14]_pad  ;
	input \CM_rd3[15]_pad  ;
	input \CM_rd3[16]_pad  ;
	input \CM_rd3[17]_pad  ;
	input \CM_rd3[18]_pad  ;
	input \CM_rd3[19]_pad  ;
	input \CM_rd3[1]_pad  ;
	input \CM_rd3[20]_pad  ;
	input \CM_rd3[21]_pad  ;
	input \CM_rd3[22]_pad  ;
	input \CM_rd3[23]_pad  ;
	input \CM_rd3[2]_pad  ;
	input \CM_rd3[3]_pad  ;
	input \CM_rd3[4]_pad  ;
	input \CM_rd3[5]_pad  ;
	input \CM_rd3[6]_pad  ;
	input \CM_rd3[7]_pad  ;
	input \CM_rd3[8]_pad  ;
	input \CM_rd3[9]_pad  ;
	input \CM_rd4[0]_pad  ;
	input \CM_rd4[10]_pad  ;
	input \CM_rd4[11]_pad  ;
	input \CM_rd4[12]_pad  ;
	input \CM_rd4[13]_pad  ;
	input \CM_rd4[14]_pad  ;
	input \CM_rd4[15]_pad  ;
	input \CM_rd4[16]_pad  ;
	input \CM_rd4[17]_pad  ;
	input \CM_rd4[18]_pad  ;
	input \CM_rd4[19]_pad  ;
	input \CM_rd4[1]_pad  ;
	input \CM_rd4[20]_pad  ;
	input \CM_rd4[21]_pad  ;
	input \CM_rd4[22]_pad  ;
	input \CM_rd4[23]_pad  ;
	input \CM_rd4[2]_pad  ;
	input \CM_rd4[3]_pad  ;
	input \CM_rd4[4]_pad  ;
	input \CM_rd4[5]_pad  ;
	input \CM_rd4[6]_pad  ;
	input \CM_rd4[7]_pad  ;
	input \CM_rd4[8]_pad  ;
	input \CM_rd4[9]_pad  ;
	input \CM_rd5[0]_pad  ;
	input \CM_rd5[10]_pad  ;
	input \CM_rd5[11]_pad  ;
	input \CM_rd5[12]_pad  ;
	input \CM_rd5[13]_pad  ;
	input \CM_rd5[14]_pad  ;
	input \CM_rd5[15]_pad  ;
	input \CM_rd5[16]_pad  ;
	input \CM_rd5[17]_pad  ;
	input \CM_rd5[18]_pad  ;
	input \CM_rd5[19]_pad  ;
	input \CM_rd5[1]_pad  ;
	input \CM_rd5[20]_pad  ;
	input \CM_rd5[21]_pad  ;
	input \CM_rd5[22]_pad  ;
	input \CM_rd5[23]_pad  ;
	input \CM_rd5[2]_pad  ;
	input \CM_rd5[3]_pad  ;
	input \CM_rd5[4]_pad  ;
	input \CM_rd5[5]_pad  ;
	input \CM_rd5[6]_pad  ;
	input \CM_rd5[7]_pad  ;
	input \CM_rd5[8]_pad  ;
	input \CM_rd5[9]_pad  ;
	input \CM_rd6[0]_pad  ;
	input \CM_rd6[10]_pad  ;
	input \CM_rd6[11]_pad  ;
	input \CM_rd6[12]_pad  ;
	input \CM_rd6[13]_pad  ;
	input \CM_rd6[14]_pad  ;
	input \CM_rd6[15]_pad  ;
	input \CM_rd6[16]_pad  ;
	input \CM_rd6[17]_pad  ;
	input \CM_rd6[18]_pad  ;
	input \CM_rd6[19]_pad  ;
	input \CM_rd6[1]_pad  ;
	input \CM_rd6[20]_pad  ;
	input \CM_rd6[21]_pad  ;
	input \CM_rd6[22]_pad  ;
	input \CM_rd6[23]_pad  ;
	input \CM_rd6[2]_pad  ;
	input \CM_rd6[3]_pad  ;
	input \CM_rd6[4]_pad  ;
	input \CM_rd6[5]_pad  ;
	input \CM_rd6[6]_pad  ;
	input \CM_rd6[7]_pad  ;
	input \CM_rd6[8]_pad  ;
	input \CM_rd6[9]_pad  ;
	input \CM_rd7[0]_pad  ;
	input \CM_rd7[10]_pad  ;
	input \CM_rd7[11]_pad  ;
	input \CM_rd7[12]_pad  ;
	input \CM_rd7[13]_pad  ;
	input \CM_rd7[14]_pad  ;
	input \CM_rd7[15]_pad  ;
	input \CM_rd7[16]_pad  ;
	input \CM_rd7[17]_pad  ;
	input \CM_rd7[18]_pad  ;
	input \CM_rd7[19]_pad  ;
	input \CM_rd7[1]_pad  ;
	input \CM_rd7[20]_pad  ;
	input \CM_rd7[21]_pad  ;
	input \CM_rd7[22]_pad  ;
	input \CM_rd7[23]_pad  ;
	input \CM_rd7[2]_pad  ;
	input \CM_rd7[3]_pad  ;
	input \CM_rd7[4]_pad  ;
	input \CM_rd7[5]_pad  ;
	input \CM_rd7[6]_pad  ;
	input \CM_rd7[7]_pad  ;
	input \CM_rd7[8]_pad  ;
	input \CM_rd7[9]_pad  ;
	input \CM_rdm[0]_pad  ;
	input \CM_rdm[10]_pad  ;
	input \CM_rdm[11]_pad  ;
	input \CM_rdm[12]_pad  ;
	input \CM_rdm[13]_pad  ;
	input \CM_rdm[14]_pad  ;
	input \CM_rdm[15]_pad  ;
	input \CM_rdm[16]_pad  ;
	input \CM_rdm[17]_pad  ;
	input \CM_rdm[18]_pad  ;
	input \CM_rdm[19]_pad  ;
	input \CM_rdm[1]_pad  ;
	input \CM_rdm[20]_pad  ;
	input \CM_rdm[21]_pad  ;
	input \CM_rdm[22]_pad  ;
	input \CM_rdm[23]_pad  ;
	input \CM_rdm[2]_pad  ;
	input \CM_rdm[3]_pad  ;
	input \CM_rdm[4]_pad  ;
	input \CM_rdm[5]_pad  ;
	input \CM_rdm[6]_pad  ;
	input \CM_rdm[7]_pad  ;
	input \CM_rdm[8]_pad  ;
	input \CM_rdm[9]_pad  ;
	input \DM_rd0[0]_pad  ;
	input \DM_rd0[10]_pad  ;
	input \DM_rd0[11]_pad  ;
	input \DM_rd0[12]_pad  ;
	input \DM_rd0[13]_pad  ;
	input \DM_rd0[14]_pad  ;
	input \DM_rd0[15]_pad  ;
	input \DM_rd0[1]_pad  ;
	input \DM_rd0[2]_pad  ;
	input \DM_rd0[3]_pad  ;
	input \DM_rd0[4]_pad  ;
	input \DM_rd0[5]_pad  ;
	input \DM_rd0[6]_pad  ;
	input \DM_rd0[7]_pad  ;
	input \DM_rd0[8]_pad  ;
	input \DM_rd0[9]_pad  ;
	input \DM_rd1[0]_pad  ;
	input \DM_rd1[10]_pad  ;
	input \DM_rd1[11]_pad  ;
	input \DM_rd1[12]_pad  ;
	input \DM_rd1[13]_pad  ;
	input \DM_rd1[14]_pad  ;
	input \DM_rd1[15]_pad  ;
	input \DM_rd1[1]_pad  ;
	input \DM_rd1[2]_pad  ;
	input \DM_rd1[3]_pad  ;
	input \DM_rd1[4]_pad  ;
	input \DM_rd1[5]_pad  ;
	input \DM_rd1[6]_pad  ;
	input \DM_rd1[7]_pad  ;
	input \DM_rd1[8]_pad  ;
	input \DM_rd1[9]_pad  ;
	input \DM_rd2[0]_pad  ;
	input \DM_rd2[10]_pad  ;
	input \DM_rd2[11]_pad  ;
	input \DM_rd2[12]_pad  ;
	input \DM_rd2[13]_pad  ;
	input \DM_rd2[14]_pad  ;
	input \DM_rd2[15]_pad  ;
	input \DM_rd2[1]_pad  ;
	input \DM_rd2[2]_pad  ;
	input \DM_rd2[3]_pad  ;
	input \DM_rd2[4]_pad  ;
	input \DM_rd2[5]_pad  ;
	input \DM_rd2[6]_pad  ;
	input \DM_rd2[7]_pad  ;
	input \DM_rd2[8]_pad  ;
	input \DM_rd2[9]_pad  ;
	input \DM_rd3[0]_pad  ;
	input \DM_rd3[10]_pad  ;
	input \DM_rd3[11]_pad  ;
	input \DM_rd3[12]_pad  ;
	input \DM_rd3[13]_pad  ;
	input \DM_rd3[14]_pad  ;
	input \DM_rd3[15]_pad  ;
	input \DM_rd3[1]_pad  ;
	input \DM_rd3[2]_pad  ;
	input \DM_rd3[3]_pad  ;
	input \DM_rd3[4]_pad  ;
	input \DM_rd3[5]_pad  ;
	input \DM_rd3[6]_pad  ;
	input \DM_rd3[7]_pad  ;
	input \DM_rd3[8]_pad  ;
	input \DM_rd3[9]_pad  ;
	input \DM_rd4[0]_pad  ;
	input \DM_rd4[10]_pad  ;
	input \DM_rd4[11]_pad  ;
	input \DM_rd4[12]_pad  ;
	input \DM_rd4[13]_pad  ;
	input \DM_rd4[14]_pad  ;
	input \DM_rd4[15]_pad  ;
	input \DM_rd4[1]_pad  ;
	input \DM_rd4[2]_pad  ;
	input \DM_rd4[3]_pad  ;
	input \DM_rd4[4]_pad  ;
	input \DM_rd4[5]_pad  ;
	input \DM_rd4[6]_pad  ;
	input \DM_rd4[7]_pad  ;
	input \DM_rd4[8]_pad  ;
	input \DM_rd4[9]_pad  ;
	input \DM_rd5[0]_pad  ;
	input \DM_rd5[10]_pad  ;
	input \DM_rd5[11]_pad  ;
	input \DM_rd5[12]_pad  ;
	input \DM_rd5[13]_pad  ;
	input \DM_rd5[14]_pad  ;
	input \DM_rd5[15]_pad  ;
	input \DM_rd5[1]_pad  ;
	input \DM_rd5[2]_pad  ;
	input \DM_rd5[3]_pad  ;
	input \DM_rd5[4]_pad  ;
	input \DM_rd5[5]_pad  ;
	input \DM_rd5[6]_pad  ;
	input \DM_rd5[7]_pad  ;
	input \DM_rd5[8]_pad  ;
	input \DM_rd5[9]_pad  ;
	input \DM_rd6[0]_pad  ;
	input \DM_rd6[10]_pad  ;
	input \DM_rd6[11]_pad  ;
	input \DM_rd6[12]_pad  ;
	input \DM_rd6[13]_pad  ;
	input \DM_rd6[14]_pad  ;
	input \DM_rd6[15]_pad  ;
	input \DM_rd6[1]_pad  ;
	input \DM_rd6[2]_pad  ;
	input \DM_rd6[3]_pad  ;
	input \DM_rd6[4]_pad  ;
	input \DM_rd6[5]_pad  ;
	input \DM_rd6[6]_pad  ;
	input \DM_rd6[7]_pad  ;
	input \DM_rd6[8]_pad  ;
	input \DM_rd6[9]_pad  ;
	input \DM_rd7[0]_pad  ;
	input \DM_rd7[10]_pad  ;
	input \DM_rd7[11]_pad  ;
	input \DM_rd7[12]_pad  ;
	input \DM_rd7[13]_pad  ;
	input \DM_rd7[14]_pad  ;
	input \DM_rd7[15]_pad  ;
	input \DM_rd7[1]_pad  ;
	input \DM_rd7[2]_pad  ;
	input \DM_rd7[3]_pad  ;
	input \DM_rd7[4]_pad  ;
	input \DM_rd7[5]_pad  ;
	input \DM_rd7[6]_pad  ;
	input \DM_rd7[7]_pad  ;
	input \DM_rd7[8]_pad  ;
	input \DM_rd7[9]_pad  ;
	input \DM_rdm[0]_pad  ;
	input \DM_rdm[10]_pad  ;
	input \DM_rdm[11]_pad  ;
	input \DM_rdm[12]_pad  ;
	input \DM_rdm[13]_pad  ;
	input \DM_rdm[14]_pad  ;
	input \DM_rdm[15]_pad  ;
	input \DM_rdm[1]_pad  ;
	input \DM_rdm[2]_pad  ;
	input \DM_rdm[3]_pad  ;
	input \DM_rdm[4]_pad  ;
	input \DM_rdm[5]_pad  ;
	input \DM_rdm[6]_pad  ;
	input \DM_rdm[7]_pad  ;
	input \DM_rdm[8]_pad  ;
	input \DM_rdm[9]_pad  ;
	input IACKn_pad ;
	input \IRFS0_pad  ;
	input \IRFS1_pad  ;
	input \ISCLK0_pad  ;
	input \ISCLK1_pad  ;
	input \ITFS0_pad  ;
	input \ITFS1_pad  ;
	input \PIO_oe[0]_pad  ;
	input \PIO_oe[10]_pad  ;
	input \PIO_oe[11]_pad  ;
	input \PIO_oe[1]_pad  ;
	input \PIO_oe[2]_pad  ;
	input \PIO_oe[3]_pad  ;
	input \PIO_oe[4]_pad  ;
	input \PIO_oe[5]_pad  ;
	input \PIO_oe[6]_pad  ;
	input \PIO_oe[7]_pad  ;
	input \PIO_oe[8]_pad  ;
	input \PIO_oe[9]_pad  ;
	input \PIO_out[0]_pad  ;
	input \PIO_out[10]_pad  ;
	input \PIO_out[11]_pad  ;
	input \PIO_out[1]_pad  ;
	input \PIO_out[2]_pad  ;
	input \PIO_out[3]_pad  ;
	input \PIO_out[4]_pad  ;
	input \PIO_out[5]_pad  ;
	input \PIO_out[6]_pad  ;
	input \PIO_out[7]_pad  ;
	input \PIO_out[8]_pad  ;
	input \PIO_out[9]_pad  ;
	input PM_bdry_sel_pad ;
	input \PM_rd0[0]_pad  ;
	input \PM_rd0[10]_pad  ;
	input \PM_rd0[11]_pad  ;
	input \PM_rd0[12]_pad  ;
	input \PM_rd0[13]_pad  ;
	input \PM_rd0[14]_pad  ;
	input \PM_rd0[15]_pad  ;
	input \PM_rd0[1]_pad  ;
	input \PM_rd0[2]_pad  ;
	input \PM_rd0[3]_pad  ;
	input \PM_rd0[4]_pad  ;
	input \PM_rd0[5]_pad  ;
	input \PM_rd0[6]_pad  ;
	input \PM_rd0[7]_pad  ;
	input \PM_rd0[8]_pad  ;
	input \PM_rd0[9]_pad  ;
	input \PM_rd1[0]_pad  ;
	input \PM_rd1[10]_pad  ;
	input \PM_rd1[11]_pad  ;
	input \PM_rd1[12]_pad  ;
	input \PM_rd1[13]_pad  ;
	input \PM_rd1[14]_pad  ;
	input \PM_rd1[15]_pad  ;
	input \PM_rd1[1]_pad  ;
	input \PM_rd1[2]_pad  ;
	input \PM_rd1[3]_pad  ;
	input \PM_rd1[4]_pad  ;
	input \PM_rd1[5]_pad  ;
	input \PM_rd1[6]_pad  ;
	input \PM_rd1[7]_pad  ;
	input \PM_rd1[8]_pad  ;
	input \PM_rd1[9]_pad  ;
	input \PM_rd2[0]_pad  ;
	input \PM_rd2[10]_pad  ;
	input \PM_rd2[11]_pad  ;
	input \PM_rd2[12]_pad  ;
	input \PM_rd2[13]_pad  ;
	input \PM_rd2[14]_pad  ;
	input \PM_rd2[15]_pad  ;
	input \PM_rd2[1]_pad  ;
	input \PM_rd2[2]_pad  ;
	input \PM_rd2[3]_pad  ;
	input \PM_rd2[4]_pad  ;
	input \PM_rd2[5]_pad  ;
	input \PM_rd2[6]_pad  ;
	input \PM_rd2[7]_pad  ;
	input \PM_rd2[8]_pad  ;
	input \PM_rd2[9]_pad  ;
	input \PM_rd3[0]_pad  ;
	input \PM_rd3[10]_pad  ;
	input \PM_rd3[11]_pad  ;
	input \PM_rd3[12]_pad  ;
	input \PM_rd3[13]_pad  ;
	input \PM_rd3[14]_pad  ;
	input \PM_rd3[15]_pad  ;
	input \PM_rd3[1]_pad  ;
	input \PM_rd3[2]_pad  ;
	input \PM_rd3[3]_pad  ;
	input \PM_rd3[4]_pad  ;
	input \PM_rd3[5]_pad  ;
	input \PM_rd3[6]_pad  ;
	input \PM_rd3[7]_pad  ;
	input \PM_rd3[8]_pad  ;
	input \PM_rd3[9]_pad  ;
	input \PM_rd4[0]_pad  ;
	input \PM_rd4[10]_pad  ;
	input \PM_rd4[11]_pad  ;
	input \PM_rd4[12]_pad  ;
	input \PM_rd4[13]_pad  ;
	input \PM_rd4[14]_pad  ;
	input \PM_rd4[15]_pad  ;
	input \PM_rd4[1]_pad  ;
	input \PM_rd4[2]_pad  ;
	input \PM_rd4[3]_pad  ;
	input \PM_rd4[4]_pad  ;
	input \PM_rd4[5]_pad  ;
	input \PM_rd4[6]_pad  ;
	input \PM_rd4[7]_pad  ;
	input \PM_rd4[8]_pad  ;
	input \PM_rd4[9]_pad  ;
	input \PM_rd5[0]_pad  ;
	input \PM_rd5[10]_pad  ;
	input \PM_rd5[11]_pad  ;
	input \PM_rd5[12]_pad  ;
	input \PM_rd5[13]_pad  ;
	input \PM_rd5[14]_pad  ;
	input \PM_rd5[15]_pad  ;
	input \PM_rd5[1]_pad  ;
	input \PM_rd5[2]_pad  ;
	input \PM_rd5[3]_pad  ;
	input \PM_rd5[4]_pad  ;
	input \PM_rd5[5]_pad  ;
	input \PM_rd5[6]_pad  ;
	input \PM_rd5[7]_pad  ;
	input \PM_rd5[8]_pad  ;
	input \PM_rd5[9]_pad  ;
	input \PM_rd6[0]_pad  ;
	input \PM_rd6[10]_pad  ;
	input \PM_rd6[11]_pad  ;
	input \PM_rd6[12]_pad  ;
	input \PM_rd6[13]_pad  ;
	input \PM_rd6[14]_pad  ;
	input \PM_rd6[15]_pad  ;
	input \PM_rd6[1]_pad  ;
	input \PM_rd6[2]_pad  ;
	input \PM_rd6[3]_pad  ;
	input \PM_rd6[4]_pad  ;
	input \PM_rd6[5]_pad  ;
	input \PM_rd6[6]_pad  ;
	input \PM_rd6[7]_pad  ;
	input \PM_rd6[8]_pad  ;
	input \PM_rd6[9]_pad  ;
	input \PM_rd7[0]_pad  ;
	input \PM_rd7[10]_pad  ;
	input \PM_rd7[11]_pad  ;
	input \PM_rd7[12]_pad  ;
	input \PM_rd7[13]_pad  ;
	input \PM_rd7[14]_pad  ;
	input \PM_rd7[15]_pad  ;
	input \PM_rd7[1]_pad  ;
	input \PM_rd7[2]_pad  ;
	input \PM_rd7[3]_pad  ;
	input \PM_rd7[4]_pad  ;
	input \PM_rd7[5]_pad  ;
	input \PM_rd7[6]_pad  ;
	input \PM_rd7[7]_pad  ;
	input \PM_rd7[8]_pad  ;
	input \PM_rd7[9]_pad  ;
	input PWDACK_pad ;
	input T_BMODE_pad ;
	input T_BRn_pad ;
	input T_CLKI_OSC_pad ;
	input T_CLKI_PLL_pad ;
	input \T_ED[0]_pad  ;
	input \T_ED[10]_pad  ;
	input \T_ED[11]_pad  ;
	input \T_ED[12]_pad  ;
	input \T_ED[13]_pad  ;
	input \T_ED[14]_pad  ;
	input \T_ED[15]_pad  ;
	input \T_ED[1]_pad  ;
	input \T_ED[2]_pad  ;
	input \T_ED[3]_pad  ;
	input \T_ED[4]_pad  ;
	input \T_ED[5]_pad  ;
	input \T_ED[6]_pad  ;
	input \T_ED[7]_pad  ;
	input \T_ED[8]_pad  ;
	input \T_ED[9]_pad  ;
	input T_ICE_RSTn_pad ;
	input T_ID_pad ;
	input T_IMS_pad ;
	input T_IRDn_pad ;
	input \T_IRQ0n_pad  ;
	input \T_IRQ1n_pad  ;
	input \T_IRQ2n_pad  ;
	input \T_IRQE0n_pad  ;
	input \T_IRQE1n_pad  ;
	input \T_IRQL1n_pad  ;
	input T_ISn_pad ;
	input T_IWRn_pad ;
	input T_MMAP_pad ;
	input \T_PIOin[0]_pad  ;
	input \T_PIOin[10]_pad  ;
	input \T_PIOin[11]_pad  ;
	input \T_PIOin[1]_pad  ;
	input \T_PIOin[2]_pad  ;
	input \T_PIOin[3]_pad  ;
	input \T_PIOin[4]_pad  ;
	input \T_PIOin[5]_pad  ;
	input \T_PIOin[6]_pad  ;
	input \T_PIOin[7]_pad  ;
	input \T_PIOin[8]_pad  ;
	input \T_PIOin[9]_pad  ;
	input T_PWDn_pad ;
	input \T_RD0_pad  ;
	input \T_RD1_pad  ;
	input \T_RFS0_pad  ;
	input \T_RFS1_pad  ;
	input T_RSTn_pad ;
	input \T_SCLK0_pad  ;
	input \T_SCLK1_pad  ;
	input T_Sel_PLL_pad ;
	input \T_TFS0_pad  ;
	input \T_TFS1_pad  ;
	input \T_TMODE[0]_pad  ;
	input \T_TMODE[1]_pad  ;
	input \auctl_BSack_reg/NET0131  ;
	input \auctl_DSack_reg/NET0131  ;
	input \auctl_R0Sack_reg/NET0131  ;
	input \auctl_R1Sack_reg/NET0131  ;
	input \auctl_RST_reg/P0001  ;
	input \auctl_STEAL_reg/NET0131  ;
	input \auctl_T0Sack_reg/NET0131  ;
	input \auctl_T1Sack_reg/NET0131  ;
	input \bdma_BCTL_reg[0]/NET0131  ;
	input \bdma_BCTL_reg[10]/NET0131  ;
	input \bdma_BCTL_reg[11]/NET0131  ;
	input \bdma_BCTL_reg[12]/NET0131  ;
	input \bdma_BCTL_reg[13]/NET0131  ;
	input \bdma_BCTL_reg[14]/NET0131  ;
	input \bdma_BCTL_reg[15]/NET0131  ;
	input \bdma_BCTL_reg[1]/NET0131  ;
	input \bdma_BCTL_reg[2]/NET0131  ;
	input \bdma_BCTL_reg[3]/NET0131  ;
	input \bdma_BCTL_reg[4]/NET0131  ;
	input \bdma_BCTL_reg[5]/NET0131  ;
	input \bdma_BCTL_reg[6]/NET0131  ;
	input \bdma_BCTL_reg[7]/NET0131  ;
	input \bdma_BCTL_reg[8]/NET0131  ;
	input \bdma_BCTL_reg[9]/NET0131  ;
	input \bdma_BDMA_boot_reg/NET0131_reg_syn_10  ;
	input \bdma_BDMA_boot_reg/NET0131_reg_syn_2  ;
	input \bdma_BDMA_boot_reg/NET0131_reg_syn_8  ;
	input \bdma_BDMAmode_reg/NET0131  ;
	input \bdma_BEAD_reg[0]/NET0131  ;
	input \bdma_BEAD_reg[10]/NET0131  ;
	input \bdma_BEAD_reg[11]/NET0131  ;
	input \bdma_BEAD_reg[12]/NET0131  ;
	input \bdma_BEAD_reg[13]/NET0131  ;
	input \bdma_BEAD_reg[1]/NET0131  ;
	input \bdma_BEAD_reg[2]/NET0131  ;
	input \bdma_BEAD_reg[3]/NET0131  ;
	input \bdma_BEAD_reg[4]/NET0131  ;
	input \bdma_BEAD_reg[5]/NET0131  ;
	input \bdma_BEAD_reg[6]/NET0131  ;
	input \bdma_BEAD_reg[7]/NET0131  ;
	input \bdma_BEAD_reg[8]/NET0131  ;
	input \bdma_BEAD_reg[9]/NET0131  ;
	input \bdma_BIAD_reg[0]/NET0131  ;
	input \bdma_BIAD_reg[10]/NET0131  ;
	input \bdma_BIAD_reg[11]/NET0131  ;
	input \bdma_BIAD_reg[12]/NET0131  ;
	input \bdma_BIAD_reg[13]/NET0131  ;
	input \bdma_BIAD_reg[1]/NET0131  ;
	input \bdma_BIAD_reg[2]/NET0131  ;
	input \bdma_BIAD_reg[3]/NET0131  ;
	input \bdma_BIAD_reg[4]/NET0131  ;
	input \bdma_BIAD_reg[5]/NET0131  ;
	input \bdma_BIAD_reg[6]/NET0131  ;
	input \bdma_BIAD_reg[7]/NET0131  ;
	input \bdma_BIAD_reg[8]/NET0131  ;
	input \bdma_BIAD_reg[9]/NET0131  ;
	input \bdma_BM_cyc_reg/P0001  ;
	input \bdma_BMcyc_del_reg/P0001  ;
	input \bdma_BOVL_reg[0]/NET0131  ;
	input \bdma_BOVL_reg[10]/NET0131  ;
	input \bdma_BOVL_reg[11]/NET0131  ;
	input \bdma_BOVL_reg[1]/NET0131  ;
	input \bdma_BOVL_reg[2]/NET0131  ;
	input \bdma_BOVL_reg[3]/NET0131  ;
	input \bdma_BOVL_reg[4]/NET0131  ;
	input \bdma_BOVL_reg[5]/NET0131  ;
	input \bdma_BOVL_reg[6]/NET0131  ;
	input \bdma_BOVL_reg[7]/NET0131  ;
	input \bdma_BOVL_reg[8]/NET0131  ;
	input \bdma_BOVL_reg[9]/NET0131  ;
	input \bdma_BRST_s2_reg/NET0131  ;
	input \bdma_BRdataBUF_reg[0]/P0001  ;
	input \bdma_BRdataBUF_reg[10]/P0001  ;
	input \bdma_BRdataBUF_reg[11]/P0001  ;
	input \bdma_BRdataBUF_reg[12]/P0001  ;
	input \bdma_BRdataBUF_reg[13]/P0001  ;
	input \bdma_BRdataBUF_reg[14]/P0001  ;
	input \bdma_BRdataBUF_reg[15]/P0001  ;
	input \bdma_BRdataBUF_reg[16]/P0001  ;
	input \bdma_BRdataBUF_reg[17]/P0001  ;
	input \bdma_BRdataBUF_reg[18]/P0001  ;
	input \bdma_BRdataBUF_reg[19]/P0001  ;
	input \bdma_BRdataBUF_reg[1]/P0001  ;
	input \bdma_BRdataBUF_reg[20]/P0001  ;
	input \bdma_BRdataBUF_reg[21]/P0001  ;
	input \bdma_BRdataBUF_reg[22]/P0001  ;
	input \bdma_BRdataBUF_reg[23]/P0001  ;
	input \bdma_BRdataBUF_reg[2]/P0001  ;
	input \bdma_BRdataBUF_reg[3]/P0001  ;
	input \bdma_BRdataBUF_reg[4]/P0001  ;
	input \bdma_BRdataBUF_reg[5]/P0001  ;
	input \bdma_BRdataBUF_reg[6]/P0001  ;
	input \bdma_BRdataBUF_reg[7]/P0001  ;
	input \bdma_BRdataBUF_reg[8]/P0001  ;
	input \bdma_BRdataBUF_reg[9]/P0001  ;
	input \bdma_BSreq_reg/NET0131  ;
	input \bdma_BWCOUNT_reg[0]/NET0131  ;
	input \bdma_BWCOUNT_reg[10]/NET0131  ;
	input \bdma_BWCOUNT_reg[11]/NET0131  ;
	input \bdma_BWCOUNT_reg[12]/NET0131  ;
	input \bdma_BWCOUNT_reg[13]/NET0131  ;
	input \bdma_BWCOUNT_reg[1]/NET0131  ;
	input \bdma_BWCOUNT_reg[2]/NET0131  ;
	input \bdma_BWCOUNT_reg[3]/NET0131  ;
	input \bdma_BWCOUNT_reg[4]/NET0131  ;
	input \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_2  ;
	input \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_8  ;
	input \bdma_BWCOUNT_reg[6]/NET0131  ;
	input \bdma_BWCOUNT_reg[7]/NET0131  ;
	input \bdma_BWCOUNT_reg[8]/NET0131  ;
	input \bdma_BWCOUNT_reg[9]/NET0131  ;
	input \bdma_BWRn_reg/NET0131  ;
	input \bdma_BWcnt_reg[0]/NET0131  ;
	input \bdma_BWcnt_reg[1]/NET0131  ;
	input \bdma_BWcnt_reg[2]/NET0131  ;
	input \bdma_BWcnt_reg[3]/NET0131  ;
	input \bdma_BWcnt_reg[4]/NET0131  ;
	input \bdma_BWdataBUF_h_reg[0]/P0001  ;
	input \bdma_BWdataBUF_h_reg[10]/P0001  ;
	input \bdma_BWdataBUF_h_reg[11]/P0001  ;
	input \bdma_BWdataBUF_h_reg[12]/P0001  ;
	input \bdma_BWdataBUF_h_reg[13]/P0001  ;
	input \bdma_BWdataBUF_h_reg[14]/P0001  ;
	input \bdma_BWdataBUF_h_reg[15]/P0001  ;
	input \bdma_BWdataBUF_h_reg[16]/P0001  ;
	input \bdma_BWdataBUF_h_reg[17]/P0001  ;
	input \bdma_BWdataBUF_h_reg[18]/P0001  ;
	input \bdma_BWdataBUF_h_reg[19]/P0001  ;
	input \bdma_BWdataBUF_h_reg[1]/P0001  ;
	input \bdma_BWdataBUF_h_reg[20]/P0001  ;
	input \bdma_BWdataBUF_h_reg[21]/P0001  ;
	input \bdma_BWdataBUF_h_reg[22]/P0001  ;
	input \bdma_BWdataBUF_h_reg[23]/P0001  ;
	input \bdma_BWdataBUF_h_reg[2]/P0001  ;
	input \bdma_BWdataBUF_h_reg[3]/P0001  ;
	input \bdma_BWdataBUF_h_reg[4]/P0001  ;
	input \bdma_BWdataBUF_h_reg[5]/P0001  ;
	input \bdma_BWdataBUF_h_reg[6]/P0001  ;
	input \bdma_BWdataBUF_h_reg[7]/P0001  ;
	input \bdma_BWdataBUF_h_reg[8]/P0001  ;
	input \bdma_BWdataBUF_h_reg[9]/P0001  ;
	input \bdma_BWdataBUF_reg[0]/P0001  ;
	input \bdma_BWdataBUF_reg[1]/P0001  ;
	input \bdma_BWdataBUF_reg[2]/P0001  ;
	input \bdma_BWdataBUF_reg[3]/P0001  ;
	input \bdma_BWdataBUF_reg[4]/P0001  ;
	input \bdma_BWdataBUF_reg[5]/P0001  ;
	input \bdma_BWdataBUF_reg[6]/P0001  ;
	input \bdma_BWdataBUF_reg[7]/P0001  ;
	input \bdma_CMcnt_reg[0]/NET0131  ;
	input \bdma_CMcnt_reg[1]/NET0131  ;
	input \bdma_DM_2nd_reg/NET0131  ;
	input \bdma_RST_pin_reg/P0001  ;
	input \bdma_WRlat_reg/P0001  ;
	input \clkc_Awake_reg/NET0131  ;
	input \clkc_CLKOUT_reg/NET0131  ;
	input \clkc_CTR_cnt_reg[0]/NET0131  ;
	input \clkc_CTR_cnt_reg[1]/NET0131  ;
	input \clkc_Cnt128_reg/NET0131  ;
	input \clkc_Cnt4096_reg/NET0131  ;
	input \clkc_Cnt4096_s1_reg/NET0131  ;
	input \clkc_Cnt4096_s2_reg/NET0131  ;
	input \clkc_DSPoff_reg/NET0131  ;
	input \clkc_OSCoff_reg/NET0131  ;
	input \clkc_OSCoff_set_reg/P0001  ;
	input \clkc_OUTcnt_reg[0]/NET0131  ;
	input \clkc_OUTcnt_reg[1]/NET0131  ;
	input \clkc_OUTcnt_reg[2]/NET0131  ;
	input \clkc_OUTcnt_reg[3]/NET0131  ;
	input \clkc_OUTcnt_reg[4]/NET0131  ;
	input \clkc_OUTcnt_reg[5]/NET0131  ;
	input \clkc_OUTcnt_reg[6]/NET0131  ;
	input \clkc_RSTtext_reg/P0001  ;
	input \clkc_SIDLE_s1_reg/NET0131  ;
	input \clkc_SIDLE_s2_reg/NET0131  ;
	input \clkc_SLEEP_reg/NET0131  ;
	input \clkc_STBY_reg/NET0131  ;
	input \clkc_STDcnt_reg[0]/NET0131  ;
	input \clkc_STDcnt_reg[10]/NET0131  ;
	input \clkc_STDcnt_reg[1]/NET0131  ;
	input \clkc_STDcnt_reg[2]/NET0131  ;
	input \clkc_STDcnt_reg[3]/NET0131  ;
	input \clkc_STDcnt_reg[4]/NET0131  ;
	input \clkc_STDcnt_reg[5]/NET0131  ;
	input \clkc_STDcnt_reg[6]/NET0131  ;
	input \clkc_STDcnt_reg[7]/NET0131  ;
	input \clkc_STDcnt_reg[8]/NET0131  ;
	input \clkc_STDcnt_reg[9]/NET0131  ;
	input \clkc_SlowDn_reg/NET0131  ;
	input \clkc_SlowDn_s1_reg/P0001  ;
	input \clkc_SlowDn_s2_reg/P0001  ;
	input \clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131  ;
	input \clkc_ckr_reg_DO_reg[0]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[10]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[11]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[12]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[13]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[14]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[15]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[1]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[2]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[3]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[4]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[5]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[6]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[7]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[8]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[9]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[0]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[10]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[11]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[1]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[2]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[3]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[4]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[5]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[6]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[7]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[8]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[9]/NET0131  ;
	input \core_c_dec_ALUop_E_reg/P0001  ;
	input \core_c_dec_BR_Ed_reg/P0001  ;
	input \core_c_dec_Call_Ed_reg/P0001  ;
	input \core_c_dec_DIVQ_E_reg/P0001  ;
	input \core_c_dec_DIVS_E_reg/P0001  ;
	input \core_c_dec_DU_Eg_reg/P0001  ;
	input \core_c_dec_Double_E_reg/P0001  ;
	input \core_c_dec_Dummy_E_reg/NET0131  ;
	input \core_c_dec_EXIT_E_reg/P0001  ;
	input \core_c_dec_IDLE_Eg_reg/P0001  ;
	input \core_c_dec_IRE_reg[0]/NET0131  ;
	input \core_c_dec_IRE_reg[10]/NET0131  ;
	input \core_c_dec_IRE_reg[11]/NET0131  ;
	input \core_c_dec_IRE_reg[12]/NET0131  ;
	input \core_c_dec_IRE_reg[13]/NET0131  ;
	input \core_c_dec_IRE_reg[14]/NET0131  ;
	input \core_c_dec_IRE_reg[15]/NET0131  ;
	input \core_c_dec_IRE_reg[16]/NET0131  ;
	input \core_c_dec_IRE_reg[17]/NET0131  ;
	input \core_c_dec_IRE_reg[18]/NET0131  ;
	input \core_c_dec_IRE_reg[19]/NET0131  ;
	input \core_c_dec_IRE_reg[1]/NET0131  ;
	input \core_c_dec_IRE_reg[2]/NET0131  ;
	input \core_c_dec_IRE_reg[3]/NET0131  ;
	input \core_c_dec_IRE_reg[4]/NET0131  ;
	input \core_c_dec_IRE_reg[5]/NET0131  ;
	input \core_c_dec_IRE_reg[6]/NET0131  ;
	input \core_c_dec_IRE_reg[7]/NET0131  ;
	input \core_c_dec_IRE_reg[8]/NET0131  ;
	input \core_c_dec_IRE_reg[9]/NET0131  ;
	input \core_c_dec_IR_reg[0]/NET0131  ;
	input \core_c_dec_IR_reg[10]/NET0131  ;
	input \core_c_dec_IR_reg[11]/NET0131  ;
	input \core_c_dec_IR_reg[12]/NET0131  ;
	input \core_c_dec_IR_reg[13]/NET0131  ;
	input \core_c_dec_IR_reg[14]/NET0131  ;
	input \core_c_dec_IR_reg[15]/NET0131  ;
	input \core_c_dec_IR_reg[16]/NET0131  ;
	input \core_c_dec_IR_reg[17]/NET0131  ;
	input \core_c_dec_IR_reg[18]/NET0131  ;
	input \core_c_dec_IR_reg[19]/NET0131  ;
	input \core_c_dec_IR_reg[1]/NET0131  ;
	input \core_c_dec_IR_reg[20]/NET0131  ;
	input \core_c_dec_IR_reg[21]/NET0131  ;
	input \core_c_dec_IR_reg[22]/NET0131  ;
	input \core_c_dec_IR_reg[23]/NET0131  ;
	input \core_c_dec_IR_reg[2]/NET0131  ;
	input \core_c_dec_IR_reg[3]/NET0131  ;
	input \core_c_dec_IR_reg[4]/NET0131  ;
	input \core_c_dec_IR_reg[5]/NET0131  ;
	input \core_c_dec_IR_reg[6]/NET0131  ;
	input \core_c_dec_IR_reg[7]/NET0131  ;
	input \core_c_dec_IR_reg[8]/NET0131  ;
	input \core_c_dec_IR_reg[9]/NET0131  ;
	input \core_c_dec_Long_Cg_reg/P0001  ;
	input \core_c_dec_Long_Eg_reg/P0001  ;
	input \core_c_dec_MACdep_Eg_reg/P0001  ;
	input \core_c_dec_MACop_E_reg/P0001  ;
	input \core_c_dec_MFALU_Ei_reg/NET0131  ;
	input \core_c_dec_MFAR_E_reg/P0001  ;
	input \core_c_dec_MFASTAT_E_reg/P0001  ;
	input \core_c_dec_MFAX0_E_reg/P0001  ;
	input \core_c_dec_MFAX1_E_reg/P0001  ;
	input \core_c_dec_MFAY0_E_reg/P0001  ;
	input \core_c_dec_MFAY1_E_reg/P0001  ;
	input \core_c_dec_MFCNTR_E_reg/P0001  ;
	input \core_c_dec_MFDAG1_Ei_reg/NET0131  ;
	input \core_c_dec_MFDAG2_Ei_reg/NET0131  ;
	input \core_c_dec_MFDMOVL_E_reg/P0001  ;
	input \core_c_dec_MFICNTL_E_reg/P0001  ;
	input \core_c_dec_MFIDR_E_reg/P0001  ;
	input \core_c_dec_MFIMASK_E_reg/P0001  ;
	input \core_c_dec_MFIreg_E_reg[0]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[1]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[2]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[3]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[4]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[5]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[6]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[7]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[0]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[1]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[2]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[3]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[4]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[5]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[6]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[7]/P0001  ;
	input \core_c_dec_MFMAC_Ei_reg/NET0131  ;
	input \core_c_dec_MFMR0_E_reg/P0001  ;
	input \core_c_dec_MFMR1_E_reg/P0001  ;
	input \core_c_dec_MFMR2_E_reg/P0001  ;
	input \core_c_dec_MFMSTAT_E_reg/P0001  ;
	input \core_c_dec_MFMX0_E_reg/P0001  ;
	input \core_c_dec_MFMX1_E_reg/P0001  ;
	input \core_c_dec_MFMY0_E_reg/P0001  ;
	input \core_c_dec_MFMY1_E_reg/P0001  ;
	input \core_c_dec_MFMreg_E_reg[0]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[1]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[2]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[3]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[4]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[5]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[6]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[7]/P0001  ;
	input \core_c_dec_MFPMOVL_E_reg/P0001  ;
	input \core_c_dec_MFPSQ_Ei_reg/NET0131  ;
	input \core_c_dec_MFRX0_E_reg/P0001  ;
	input \core_c_dec_MFRX1_E_reg/P0001  ;
	input \core_c_dec_MFSB_E_reg/P0001  ;
	input \core_c_dec_MFSE_E_reg/P0001  ;
	input \core_c_dec_MFSHT_Ei_reg/NET0131  ;
	input \core_c_dec_MFSI_E_reg/P0001  ;
	input \core_c_dec_MFSPT_Ei_reg/NET0131  ;
	input \core_c_dec_MFSR0_E_reg/P0001  ;
	input \core_c_dec_MFSR1_E_reg/P0001  ;
	input \core_c_dec_MFSSTAT_E_reg/P0001  ;
	input \core_c_dec_MFTX0_E_reg/P0001  ;
	input \core_c_dec_MFTX1_E_reg/P0001  ;
	input \core_c_dec_MFtoppcs_Eg_reg/P0001  ;
	input \core_c_dec_MTAR_E_reg/P0001  ;
	input \core_c_dec_MTASTAT_E_reg/P0001  ;
	input \core_c_dec_MTAX0_E_reg/P0001  ;
	input \core_c_dec_MTAX1_E_reg/P0001  ;
	input \core_c_dec_MTAY0_E_reg/P0001  ;
	input \core_c_dec_MTAY1_E_reg/P0001  ;
	input \core_c_dec_MTCNTR_Eg_reg/P0001  ;
	input \core_c_dec_MTDMOVL_E_reg/P0001  ;
	input \core_c_dec_MTICNTL_Eg_reg/P0001  ;
	input \core_c_dec_MTIDR_E_reg/P0001  ;
	input \core_c_dec_MTIFC_Eg_reg/P0001  ;
	input \core_c_dec_MTIMASK_Eg_reg/P0001  ;
	input \core_c_dec_MTIreg_E_reg[0]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[1]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[2]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[3]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[4]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[5]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[6]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[7]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[0]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[1]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[2]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[3]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[4]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[5]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[6]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[7]/P0001  ;
	input \core_c_dec_MTMR0_E_reg/P0001  ;
	input \core_c_dec_MTMR1_E_reg/P0001  ;
	input \core_c_dec_MTMR2_E_reg/P0001  ;
	input \core_c_dec_MTMSTAT_Eg_reg/P0001  ;
	input \core_c_dec_MTMX0_E_reg/P0001  ;
	input \core_c_dec_MTMX1_E_reg/P0001  ;
	input \core_c_dec_MTMY0_E_reg/P0001  ;
	input \core_c_dec_MTMY1_E_reg/P0001  ;
	input \core_c_dec_MTMreg_E_reg[0]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[1]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[2]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[3]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[4]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[5]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[6]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[7]/P0001  ;
	input \core_c_dec_MTOWRCNTR_Eg_reg/P0001  ;
	input \core_c_dec_MTPMOVL_E_reg/P0001  ;
	input \core_c_dec_MTRX0_E_reg/P0001  ;
	input \core_c_dec_MTRX1_E_reg/P0001  ;
	input \core_c_dec_MTSB_E_reg/P0001  ;
	input \core_c_dec_MTSE_E_reg/P0001  ;
	input \core_c_dec_MTSI_E_reg/P0001  ;
	input \core_c_dec_MTSR0_E_reg/P0001  ;
	input \core_c_dec_MTSR1_E_reg/P0001  ;
	input \core_c_dec_MTTX0_E_reg/P0001  ;
	input \core_c_dec_MTTX1_E_reg/P0001  ;
	input \core_c_dec_MTtoppcs_Eg_reg/P0001  ;
	input \core_c_dec_Modctl_Eg_reg/P0001  ;
	input \core_c_dec_MpopLP_Eg_reg/P0001  ;
	input \core_c_dec_NOP_E_reg/P0001  ;
	input \core_c_dec_Nrti_Ed_reg/P0001  ;
	input \core_c_dec_Nseq_Ed_reg/P0001  ;
	input \core_c_dec_PPclr_reg/P0001  ;
	input \core_c_dec_Post1_E_reg/P0001  ;
	input \core_c_dec_Post2_E_reg/P0001  ;
	input \core_c_dec_Prderr_Cg_reg/NET0131  ;
	input \core_c_dec_RET_Ed_reg/P0001  ;
	input \core_c_dec_RTI_Ed_reg/P0001  ;
	input \core_c_dec_SHTop_E_reg/P0001  ;
	input \core_c_dec_Stkctl_Eg_reg/P0001  ;
	input \core_c_dec_Usecond_E_reg/P0001  ;
	input \core_c_dec_accCM_E_reg/NET0131  ;
	input \core_c_dec_accPM_E_reg/P0001  ;
	input \core_c_dec_cdAM_E_reg/P0001  ;
	input \core_c_dec_imSHT_E_reg/P0001  ;
	input \core_c_dec_imm14_E_reg/P0001  ;
	input \core_c_dec_imm16_E_reg/P0001  ;
	input \core_c_dec_pMFALU_Ei_reg/NET0131  ;
	input \core_c_dec_pMFMAC_Ei_reg/NET0131  ;
	input \core_c_dec_pMFSHT_Ei_reg/NET0131  ;
	input \core_c_dec_rdCM_E_reg/NET0131  ;
	input \core_c_dec_satMR_E_reg/P0001  ;
	input \core_c_dec_updAF_E_reg/P0001  ;
	input \core_c_dec_updAR_E_reg/P0001  ;
	input \core_c_dec_updMF_E_reg/P0001  ;
	input \core_c_dec_updMR_E_reg/P0001  ;
	input \core_c_dec_updSR_E_reg/P0001  ;
	input \core_c_psq_CE_reg/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  ;
	input \core_c_psq_CNTRval_reg/NET0131  ;
	input \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  ;
	input \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  ;
	input \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  ;
	input \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  ;
	input \core_c_psq_DRA_reg[0]/P0001  ;
	input \core_c_psq_DRA_reg[10]/P0001  ;
	input \core_c_psq_DRA_reg[11]/P0001  ;
	input \core_c_psq_DRA_reg[12]/P0001  ;
	input \core_c_psq_DRA_reg[13]/P0001  ;
	input \core_c_psq_DRA_reg[1]/P0001  ;
	input \core_c_psq_DRA_reg[2]/P0001  ;
	input \core_c_psq_DRA_reg[3]/P0001  ;
	input \core_c_psq_DRA_reg[4]/P0001  ;
	input \core_c_psq_DRA_reg[5]/P0001  ;
	input \core_c_psq_DRA_reg[6]/P0001  ;
	input \core_c_psq_DRA_reg[7]/P0001  ;
	input \core_c_psq_DRA_reg[8]/P0001  ;
	input \core_c_psq_DRA_reg[9]/P0001  ;
	input \core_c_psq_ECYC_reg/P0001  ;
	input \core_c_psq_EXA_reg[0]/P0001  ;
	input \core_c_psq_EXA_reg[10]/P0001  ;
	input \core_c_psq_EXA_reg[11]/P0001  ;
	input \core_c_psq_EXA_reg[12]/P0001  ;
	input \core_c_psq_EXA_reg[13]/P0001  ;
	input \core_c_psq_EXA_reg[1]/P0001  ;
	input \core_c_psq_EXA_reg[2]/P0001  ;
	input \core_c_psq_EXA_reg[3]/P0001  ;
	input \core_c_psq_EXA_reg[4]/P0001  ;
	input \core_c_psq_EXA_reg[5]/P0001  ;
	input \core_c_psq_EXA_reg[6]/P0001  ;
	input \core_c_psq_EXA_reg[7]/P0001  ;
	input \core_c_psq_EXA_reg[8]/P0001  ;
	input \core_c_psq_EXA_reg[9]/P0001  ;
	input \core_c_psq_Eqend_D_reg/P0001  ;
	input \core_c_psq_Eqend_Ed_reg/P0001  ;
	input \core_c_psq_ICNTL_reg_DO_reg[0]/NET0131  ;
	input \core_c_psq_ICNTL_reg_DO_reg[1]/NET0131  ;
	input \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131  ;
	input \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  ;
	input \core_c_psq_IFA_reg[0]/P0001  ;
	input \core_c_psq_IFA_reg[10]/P0001  ;
	input \core_c_psq_IFA_reg[11]/P0001  ;
	input \core_c_psq_IFA_reg[12]/P0001  ;
	input \core_c_psq_IFA_reg[13]/P0001  ;
	input \core_c_psq_IFA_reg[1]/P0001  ;
	input \core_c_psq_IFA_reg[2]/P0001  ;
	input \core_c_psq_IFA_reg[3]/P0001  ;
	input \core_c_psq_IFA_reg[4]/P0001  ;
	input \core_c_psq_IFA_reg[5]/P0001  ;
	input \core_c_psq_IFA_reg[6]/P0001  ;
	input \core_c_psq_IFA_reg[7]/P0001  ;
	input \core_c_psq_IFA_reg[8]/P0001  ;
	input \core_c_psq_IFA_reg[9]/P0001  ;
	input \core_c_psq_IFC_reg[0]/NET0131  ;
	input \core_c_psq_IFC_reg[10]/NET0131  ;
	input \core_c_psq_IFC_reg[11]/NET0131  ;
	input \core_c_psq_IFC_reg[12]/NET0131  ;
	input \core_c_psq_IFC_reg[13]/NET0131  ;
	input \core_c_psq_IFC_reg[14]/NET0131  ;
	input \core_c_psq_IFC_reg[15]/NET0131  ;
	input \core_c_psq_IFC_reg[1]/NET0131  ;
	input \core_c_psq_IFC_reg[2]/NET0131  ;
	input \core_c_psq_IFC_reg[3]/NET0131  ;
	input \core_c_psq_IFC_reg[4]/NET0131  ;
	input \core_c_psq_IFC_reg[5]/NET0131  ;
	input \core_c_psq_IFC_reg[6]/NET0131  ;
	input \core_c_psq_IFC_reg[7]/NET0131  ;
	input \core_c_psq_IFC_reg[8]/NET0131  ;
	input \core_c_psq_IFC_reg[9]/NET0131  ;
	input \core_c_psq_IMASK_reg[0]/NET0131  ;
	input \core_c_psq_IMASK_reg[1]/NET0131  ;
	input \core_c_psq_IMASK_reg[2]/NET0131  ;
	input \core_c_psq_IMASK_reg[3]/NET0131  ;
	input \core_c_psq_IMASK_reg[4]/NET0131  ;
	input \core_c_psq_IMASK_reg[5]/NET0131  ;
	input \core_c_psq_IMASK_reg[6]/NET0131  ;
	input \core_c_psq_IMASK_reg[7]/NET0131  ;
	input \core_c_psq_IMASK_reg[8]/NET0131  ;
	input \core_c_psq_IMASK_reg[9]/NET0131  ;
	input \core_c_psq_INT_en_reg/NET0131  ;
	input \core_c_psq_Iact_E_reg[0]/NET0131  ;
	input \core_c_psq_Iact_E_reg[10]/NET0131  ;
	input \core_c_psq_Iact_E_reg[1]/NET0131  ;
	input \core_c_psq_Iact_E_reg[2]/NET0131  ;
	input \core_c_psq_Iact_E_reg[3]/NET0131  ;
	input \core_c_psq_Iact_E_reg[4]/NET0131  ;
	input \core_c_psq_Iact_E_reg[5]/NET0131  ;
	input \core_c_psq_Iact_E_reg[6]/NET0131  ;
	input \core_c_psq_Iact_E_reg[7]/NET0131  ;
	input \core_c_psq_Iact_E_reg[8]/NET0131  ;
	input \core_c_psq_Iact_E_reg[9]/NET0131  ;
	input \core_c_psq_Iflag_reg[0]/NET0131  ;
	input \core_c_psq_Iflag_reg[10]/NET0131  ;
	input \core_c_psq_Iflag_reg[11]/NET0131  ;
	input \core_c_psq_Iflag_reg[12]/NET0131  ;
	input \core_c_psq_Iflag_reg[1]/NET0131  ;
	input \core_c_psq_Iflag_reg[2]/NET0131  ;
	input \core_c_psq_Iflag_reg[3]/NET0131  ;
	input \core_c_psq_Iflag_reg[4]/NET0131  ;
	input \core_c_psq_Iflag_reg[5]/NET0131  ;
	input \core_c_psq_Iflag_reg[6]/NET0131  ;
	input \core_c_psq_Iflag_reg[7]/NET0131  ;
	input \core_c_psq_Iflag_reg[8]/NET0131  ;
	input \core_c_psq_Iflag_reg[9]/NET0131  ;
	input \core_c_psq_MGNT_reg/NET0131  ;
	input \core_c_psq_MREQ_reg/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  ;
	input \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  ;
	input \core_c_psq_PCS2or3_reg/NET0131  ;
	input \core_c_psq_PCS_reg[0]/NET0131  ;
	input \core_c_psq_PCS_reg[10]/NET0131  ;
	input \core_c_psq_PCS_reg[11]/NET0131  ;
	input \core_c_psq_PCS_reg[12]/NET0131  ;
	input \core_c_psq_PCS_reg[13]/NET0131  ;
	input \core_c_psq_PCS_reg[14]/NET0131  ;
	input \core_c_psq_PCS_reg[15]/NET0131  ;
	input \core_c_psq_PCS_reg[1]/NET0131  ;
	input \core_c_psq_PCS_reg[2]/NET0131  ;
	input \core_c_psq_PCS_reg[3]/NET0131  ;
	input \core_c_psq_PCS_reg[4]/NET0131  ;
	input \core_c_psq_PCS_reg[5]/NET0131  ;
	input \core_c_psq_PCS_reg[6]/NET0131  ;
	input \core_c_psq_PCS_reg[7]/NET0131  ;
	input \core_c_psq_PCS_reg[8]/NET0131  ;
	input \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  ;
	input \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  ;
	input \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  ;
	input \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  ;
	input \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  ;
	input \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  ;
	input \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  ;
	input \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  ;
	input \core_c_psq_SRST_reg/P0001  ;
	input \core_c_psq_SSTAT_reg[0]/NET0131  ;
	input \core_c_psq_SSTAT_reg[1]/NET0131  ;
	input \core_c_psq_SSTAT_reg[2]/NET0131  ;
	input \core_c_psq_SSTAT_reg[3]/NET0131  ;
	input \core_c_psq_SSTAT_reg[4]/NET0131  ;
	input \core_c_psq_SSTAT_reg[5]/NET0131  ;
	input \core_c_psq_SSTAT_reg[6]/NET0131  ;
	input \core_c_psq_SSTAT_reg[7]/NET0131  ;
	input \core_c_psq_TRAP_Eg_reg/NET0131  ;
	input \core_c_psq_TRAP_R_L_reg/NET0131  ;
	input \core_c_psq_T_IRQ0_s1_reg/P0001  ;
	input \core_c_psq_T_IRQ0p_reg/P0001  ;
	input \core_c_psq_T_IRQ1_s1_reg/P0001  ;
	input \core_c_psq_T_IRQ1p_reg/P0001  ;
	input \core_c_psq_T_IRQ2_s1_reg/P0001  ;
	input \core_c_psq_T_IRQ2p_reg/P0001  ;
	input \core_c_psq_T_IRQE0_reg/P0001  ;
	input \core_c_psq_T_IRQE0_s1_reg/P0001  ;
	input \core_c_psq_T_IRQE1_reg/P0001  ;
	input \core_c_psq_T_IRQE1_s1_reg/P0001  ;
	input \core_c_psq_T_IRQL0p_reg/P0001  ;
	input \core_c_psq_T_IRQL1p_reg/P0001  ;
	input \core_c_psq_T_PWRDN_reg/P0001  ;
	input \core_c_psq_T_PWRDN_s1_reg/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[0]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[10]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[11]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[12]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[13]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[1]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[2]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[3]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[4]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[5]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[6]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[7]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[8]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[9]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001  ;
	input \core_c_psq_cntstk_ptr_reg[0]/NET0131  ;
	input \core_c_psq_cntstk_ptr_reg[1]/NET0131  ;
	input \core_c_psq_cntstk_ptr_reg[2]/NET0131  ;
	input \core_c_psq_irq0_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irq0_de_OUT_reg/P0001  ;
	input \core_c_psq_irq1_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irq1_de_OUT_reg/P0001  ;
	input \core_c_psq_irq2_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irq2_de_OUT_reg/P0001  ;
	input \core_c_psq_irql0_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irql0_de_OUT_reg/P0001  ;
	input \core_c_psq_irql1_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irql1_de_OUT_reg/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001  ;
	input \core_c_psq_lpstk_ptr_reg[0]/NET0131  ;
	input \core_c_psq_lpstk_ptr_reg[1]/NET0131  ;
	input \core_c_psq_lpstk_ptr_reg[2]/NET0131  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001  ;
	input \core_c_psq_pcstk_ptr_reg[0]/NET0131  ;
	input \core_c_psq_pcstk_ptr_reg[1]/NET0131  ;
	input \core_c_psq_pcstk_ptr_reg[2]/NET0131  ;
	input \core_c_psq_pcstk_ptr_reg[3]/NET0131  ;
	input \core_c_psq_pcstk_ptr_reg[4]/NET0131  ;
	input \core_c_psq_ststk_ptr_reg[0]/NET0131  ;
	input \core_c_psq_ststk_ptr_reg[1]/NET0131  ;
	input \core_c_psq_ststk_ptr_reg[2]/NET0131  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_STEALI_E_reg[0]/P0001  ;
	input \core_dag_ilm1reg_STEALI_E_reg[1]/P0001  ;
	input \core_dag_ilm1reg_STEALI_E_reg[2]/P0001  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_IL_E_reg[0]/P0001  ;
	input \core_dag_ilm2reg_IL_E_reg[1]/P0001  ;
	input \core_dag_ilm2reg_I_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M_E_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M_E_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  ;
	input \core_dag_modulo1_R0wrap_reg/P0001  ;
	input \core_dag_modulo1_R1wrap_reg/P0001  ;
	input \core_dag_modulo1_T0wrap_reg/P0001  ;
	input \core_dag_modulo1_T1wrap_reg/P0001  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[4]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001  ;
	input \core_eu_ec_cun_AC_reg/P0001  ;
	input \core_eu_ec_cun_AN_reg/P0001  ;
	input \core_eu_ec_cun_AQ_reg/P0001  ;
	input \core_eu_ec_cun_AS_reg/P0001  ;
	input \core_eu_ec_cun_AV_reg/P0001  ;
	input \core_eu_ec_cun_AZ_reg/P0001  ;
	input \core_eu_ec_cun_COND_E_reg[0]/P0001  ;
	input \core_eu_ec_cun_COND_E_reg[1]/P0001  ;
	input \core_eu_ec_cun_COND_E_reg[2]/P0001  ;
	input \core_eu_ec_cun_COND_E_reg[3]/P0001  ;
	input \core_eu_ec_cun_MV_reg/P0000_reg_syn_2  ;
	input \core_eu_ec_cun_MVi_pre_C_reg/P0001  ;
	input \core_eu_ec_cun_SS_reg/P0001  ;
	input \core_eu_ec_cun_TERM_E_reg[0]/P0001  ;
	input \core_eu_ec_cun_TERM_E_reg[1]/P0001  ;
	input \core_eu_ec_cun_TERM_E_reg[2]/P0001  ;
	input \core_eu_ec_cun_TERM_E_reg[3]/P0001  ;
	input \core_eu_ec_cun_condOK_CE_reg/P0001  ;
	input \core_eu_ec_cun_mven_FFout_reg/NET0131  ;
	input \core_eu_ec_cun_termOK_CE_reg/P0001  ;
	input \core_eu_ec_cun_updateMV_C_reg/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_Sq_E_reg/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2  ;
	input \core_eu_em_mac_em_reg_s1_reg/P0000_reg_syn_2  ;
	input \core_eu_em_mac_em_reg_s2_reg/P0000_reg_syn_2  ;
	input \core_eu_es_sht_es_reg_SBr_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_SBr_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_SBr_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_SBr_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_SBr_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001  ;
	input \emc_DMDoe_reg/NET0131  ;
	input \emc_DMDreg_reg[0]/P0001  ;
	input \emc_DMDreg_reg[10]/P0001  ;
	input \emc_DMDreg_reg[11]/P0001  ;
	input \emc_DMDreg_reg[12]/P0001  ;
	input \emc_DMDreg_reg[13]/P0001  ;
	input \emc_DMDreg_reg[14]/P0001  ;
	input \emc_DMDreg_reg[15]/P0001  ;
	input \emc_DMDreg_reg[1]/P0001  ;
	input \emc_DMDreg_reg[2]/P0001  ;
	input \emc_DMDreg_reg[3]/P0001  ;
	input \emc_DMDreg_reg[4]/P0001  ;
	input \emc_DMDreg_reg[5]/P0001  ;
	input \emc_DMDreg_reg[6]/P0001  ;
	input \emc_DMDreg_reg[7]/P0001  ;
	input \emc_DMDreg_reg[8]/P0001  ;
	input \emc_DMDreg_reg[9]/P0001  ;
	input \emc_DMcst_reg/NET0131  ;
	input \emc_ECMA_reg[0]/P0001  ;
	input \emc_ECMA_reg[10]/P0001  ;
	input \emc_ECMA_reg[11]/P0001  ;
	input \emc_ECMA_reg[12]/P0001  ;
	input \emc_ECMA_reg[1]/P0001  ;
	input \emc_ECMA_reg[2]/P0001  ;
	input \emc_ECMA_reg[3]/P0001  ;
	input \emc_ECMA_reg[4]/P0001  ;
	input \emc_ECMA_reg[5]/P0001  ;
	input \emc_ECMA_reg[6]/P0001  ;
	input \emc_ECMA_reg[7]/P0001  ;
	input \emc_ECMA_reg[8]/P0001  ;
	input \emc_ECMA_reg[9]/P0001  ;
	input \emc_ECMDreg_reg[0]/P0001  ;
	input \emc_ECMDreg_reg[10]/P0001  ;
	input \emc_ECMDreg_reg[11]/P0001  ;
	input \emc_ECMDreg_reg[12]/P0001  ;
	input \emc_ECMDreg_reg[13]/P0001  ;
	input \emc_ECMDreg_reg[14]/P0001  ;
	input \emc_ECMDreg_reg[15]/P0001  ;
	input \emc_ECMDreg_reg[16]/P0001  ;
	input \emc_ECMDreg_reg[17]/P0001  ;
	input \emc_ECMDreg_reg[18]/P0001  ;
	input \emc_ECMDreg_reg[19]/P0001  ;
	input \emc_ECMDreg_reg[1]/P0001  ;
	input \emc_ECMDreg_reg[20]/P0001  ;
	input \emc_ECMDreg_reg[21]/P0001  ;
	input \emc_ECMDreg_reg[22]/P0001  ;
	input \emc_ECMDreg_reg[23]/P0001  ;
	input \emc_ECMDreg_reg[2]/P0001  ;
	input \emc_ECMDreg_reg[3]/P0001  ;
	input \emc_ECMDreg_reg[4]/P0001  ;
	input \emc_ECMDreg_reg[5]/P0001  ;
	input \emc_ECMDreg_reg[6]/P0001  ;
	input \emc_ECMDreg_reg[7]/P0001  ;
	input \emc_ECMDreg_reg[8]/P0001  ;
	input \emc_ECMDreg_reg[9]/P0001  ;
	input \emc_ECMcs_reg/NET0131  ;
	input \emc_ECS_reg[0]/NET0131  ;
	input \emc_ECS_reg[1]/NET0131  ;
	input \emc_ECS_reg[2]/NET0131  ;
	input \emc_ECS_reg[3]/NET0131  ;
	input \emc_ED_oei_reg/P0001  ;
	input \emc_EXTC_Eg_syn_reg/P0001  ;
	input \emc_IOcst_reg/NET0131  ;
	input \emc_PMDoe_reg/NET0131  ;
	input \emc_PMDreg_reg[0]/P0001  ;
	input \emc_PMDreg_reg[10]/P0001  ;
	input \emc_PMDreg_reg[11]/P0001  ;
	input \emc_PMDreg_reg[12]/P0001  ;
	input \emc_PMDreg_reg[13]/P0001  ;
	input \emc_PMDreg_reg[14]/P0001  ;
	input \emc_PMDreg_reg[15]/P0001  ;
	input \emc_PMDreg_reg[1]/P0001  ;
	input \emc_PMDreg_reg[2]/P0001  ;
	input \emc_PMDreg_reg[3]/P0001  ;
	input \emc_PMDreg_reg[4]/P0001  ;
	input \emc_PMDreg_reg[5]/P0001  ;
	input \emc_PMDreg_reg[6]/P0001  ;
	input \emc_PMDreg_reg[7]/P0001  ;
	input \emc_PMDreg_reg[8]/P0001  ;
	input \emc_PMDreg_reg[9]/P0001  ;
	input \emc_PMcst_reg/NET0131  ;
	input \emc_RWcnt_reg[0]/P0001  ;
	input \emc_RWcnt_reg[1]/P0001  ;
	input \emc_RWcnt_reg[2]/P0001  ;
	input \emc_RWcnt_reg[3]/P0001  ;
	input \emc_RWcnt_reg[4]/P0001  ;
	input \emc_RWcnt_reg[5]/P0001  ;
	input \emc_WRn_h_reg/P0001  ;
	input \emc_WSCRext_reg_DO_reg[0]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[1]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[2]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[3]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[4]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[5]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[6]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[7]/NET0131  ;
	input \emc_WSCRreg_DO_reg[0]/NET0131  ;
	input \emc_WSCRreg_DO_reg[10]/NET0131  ;
	input \emc_WSCRreg_DO_reg[11]/NET0131  ;
	input \emc_WSCRreg_DO_reg[12]/NET0131  ;
	input \emc_WSCRreg_DO_reg[13]/NET0131  ;
	input \emc_WSCRreg_DO_reg[14]/NET0131  ;
	input \emc_WSCRreg_DO_reg[1]/NET0131  ;
	input \emc_WSCRreg_DO_reg[2]/NET0131  ;
	input \emc_WSCRreg_DO_reg[3]/NET0131  ;
	input \emc_WSCRreg_DO_reg[4]/NET0131  ;
	input \emc_WSCRreg_DO_reg[5]/NET0131  ;
	input \emc_WSCRreg_DO_reg[6]/NET0131  ;
	input \emc_WSCRreg_DO_reg[7]/NET0131  ;
	input \emc_WSCRreg_DO_reg[8]/NET0131  ;
	input \emc_WSCRreg_DO_reg[9]/NET0131  ;
	input \emc_eRDY_reg/NET0131  ;
	input \emc_selDMDi_reg/P0001  ;
	input \emc_selPMDi_reg/P0001  ;
	input \idma_CM_oe_reg/P0001  ;
	input \idma_CMo_oe0_reg/P0001  ;
	input \idma_CMo_oe1_reg/P0001  ;
	input \idma_CMo_oe2_reg/P0001  ;
	input \idma_CMo_oe3_reg/P0001  ;
	input \idma_CMo_oe4_reg/P0001  ;
	input \idma_CMo_oe5_reg/P0001  ;
	input \idma_CMo_oe6_reg/P0001  ;
	input \idma_CMo_oe7_reg/P0001  ;
	input \idma_DCTL_reg[0]/NET0131  ;
	input \idma_DCTL_reg[10]/NET0131  ;
	input \idma_DCTL_reg[11]/NET0131  ;
	input \idma_DCTL_reg[12]/NET0131  ;
	input \idma_DCTL_reg[13]/NET0131  ;
	input \idma_DCTL_reg[14]/NET0131  ;
	input \idma_DCTL_reg[1]/NET0131  ;
	input \idma_DCTL_reg[2]/NET0131  ;
	input \idma_DCTL_reg[3]/NET0131  ;
	input \idma_DCTL_reg[4]/NET0131  ;
	input \idma_DCTL_reg[5]/NET0131  ;
	input \idma_DCTL_reg[6]/NET0131  ;
	input \idma_DCTL_reg[7]/NET0131  ;
	input \idma_DCTL_reg[8]/NET0131  ;
	input \idma_DCTL_reg[9]/NET0131  ;
	input \idma_DOVL_reg[0]/NET0131  ;
	input \idma_DOVL_reg[10]/NET0131  ;
	input \idma_DOVL_reg[11]/NET0131  ;
	input \idma_DOVL_reg[1]/NET0131  ;
	input \idma_DOVL_reg[2]/NET0131  ;
	input \idma_DOVL_reg[3]/NET0131  ;
	input \idma_DOVL_reg[4]/NET0131  ;
	input \idma_DOVL_reg[5]/NET0131  ;
	input \idma_DOVL_reg[6]/NET0131  ;
	input \idma_DOVL_reg[7]/NET0131  ;
	input \idma_DOVL_reg[8]/NET0131  ;
	input \idma_DOVL_reg[9]/NET0131  ;
	input \idma_DSreq_reg/NET0131  ;
	input \idma_DTMP_H_reg[0]/P0001  ;
	input \idma_DTMP_H_reg[10]/P0001  ;
	input \idma_DTMP_H_reg[11]/P0001  ;
	input \idma_DTMP_H_reg[12]/P0001  ;
	input \idma_DTMP_H_reg[13]/P0001  ;
	input \idma_DTMP_H_reg[14]/P0001  ;
	input \idma_DTMP_H_reg[15]/P0001  ;
	input \idma_DTMP_H_reg[1]/P0001  ;
	input \idma_DTMP_H_reg[2]/P0001  ;
	input \idma_DTMP_H_reg[3]/P0001  ;
	input \idma_DTMP_H_reg[4]/P0001  ;
	input \idma_DTMP_H_reg[5]/P0001  ;
	input \idma_DTMP_H_reg[6]/P0001  ;
	input \idma_DTMP_H_reg[7]/P0001  ;
	input \idma_DTMP_H_reg[8]/P0001  ;
	input \idma_DTMP_H_reg[9]/P0001  ;
	input \idma_DTMP_L_reg[0]/P0001  ;
	input \idma_DTMP_L_reg[1]/P0001  ;
	input \idma_DTMP_L_reg[2]/P0001  ;
	input \idma_DTMP_L_reg[3]/P0001  ;
	input \idma_DTMP_L_reg[4]/P0001  ;
	input \idma_DTMP_L_reg[5]/P0001  ;
	input \idma_DTMP_L_reg[6]/P0001  ;
	input \idma_DTMP_L_reg[7]/P0001  ;
	input \idma_IADi_reg[0]/P0001  ;
	input \idma_IADi_reg[10]/P0001  ;
	input \idma_IADi_reg[11]/P0001  ;
	input \idma_IADi_reg[12]/P0001  ;
	input \idma_IADi_reg[13]/P0001  ;
	input \idma_IADi_reg[14]/P0001  ;
	input \idma_IADi_reg[15]/P0001  ;
	input \idma_IADi_reg[1]/P0001  ;
	input \idma_IADi_reg[2]/P0001  ;
	input \idma_IADi_reg[3]/P0001  ;
	input \idma_IADi_reg[4]/P0001  ;
	input \idma_IADi_reg[5]/P0001  ;
	input \idma_IADi_reg[6]/P0001  ;
	input \idma_IADi_reg[7]/P0001  ;
	input \idma_IADi_reg[8]/P0001  ;
	input \idma_IADi_reg[9]/P0001  ;
	input \idma_IAL_reg/P0001  ;
	input \idma_IDMA_boot_reg/NET0131_reg_syn_10  ;
	input \idma_IDMA_boot_reg/NET0131_reg_syn_2  ;
	input \idma_IDMA_boot_reg/NET0131_reg_syn_8  ;
	input \idma_IRDn_reg/P0001  ;
	input \idma_ISn_reg/P0001  ;
	input \idma_IWRn_reg/P0001  ;
	input \idma_PCrd_1st_reg/NET0131  ;
	input \idma_PM_1st_reg/NET0131  ;
	input \idma_RDCMD_d1_reg/P0001  ;
	input \idma_RDCMD_reg/P0001  ;
	input \idma_RDcnt_reg[0]/NET0131  ;
	input \idma_RDcnt_reg[1]/NET0131  ;
	input \idma_RDcnt_reg[2]/NET0131  ;
	input \idma_RDcyc_reg/NET0131  ;
	input \idma_WRCMD_d1_reg/P0001  ;
	input \idma_WRCMD_reg/P0001  ;
	input \idma_WRcnt_reg[0]/NET0131  ;
	input \idma_WRcnt_reg[1]/NET0131  ;
	input \idma_WRcnt_reg[2]/NET0131  ;
	input \idma_WRcyc_reg/NET0131  ;
	input \idma_WRtrue_reg/NET0131  ;
	input \memc_DM_oe_reg/P0001  ;
	input \memc_DMo_oe0_reg/P0001  ;
	input \memc_DMo_oe1_reg/P0001  ;
	input \memc_DMo_oe2_reg/P0001  ;
	input \memc_DMo_oe3_reg/P0001  ;
	input \memc_DMo_oe4_reg/P0001  ;
	input \memc_DMo_oe5_reg/P0001  ;
	input \memc_DMo_oe6_reg/P0001  ;
	input \memc_DMo_oe7_reg/P0001  ;
	input \memc_Dread_E_reg/NET0131  ;
	input \memc_Dwrite_C_reg/NET0131  ;
	input \memc_Dwrite_E_reg/NET0131  ;
	input \memc_EXTC_E_reg/NET0131  ;
	input \memc_EXTC_Eg_reg/NET0131_reg_syn_10  ;
	input \memc_EXTC_Eg_reg/NET0131_reg_syn_2  ;
	input \memc_EXTC_Eg_reg/NET0131_reg_syn_8  ;
	input \memc_IOcmd_E_reg/NET0131  ;
	input \memc_LDaST_Eg_reg/NET0131  ;
	input \memc_MMR_web_reg/NET0131  ;
	input \memc_PMo_oe0_reg/P0001  ;
	input \memc_PMo_oe1_reg/P0001  ;
	input \memc_PMo_oe2_reg/P0001  ;
	input \memc_PMo_oe3_reg/P0001  ;
	input \memc_PMo_oe4_reg/P0001  ;
	input \memc_PMo_oe5_reg/P0001  ;
	input \memc_PMo_oe6_reg/P0001  ;
	input \memc_PMo_oe7_reg/P0001  ;
	input \memc_Pread_E_reg/NET0131  ;
	input \memc_Pwrite_C_reg/NET0131  ;
	input \memc_Pwrite_E_reg/NET0131  ;
	input \memc_STI_Cg_reg/NET0131  ;
	input \memc_accDM_E_reg/NET0131  ;
	input \memc_accPM_E_reg/NET0131  ;
	input \memc_ldSREG_E_reg/NET0131  ;
	input \memc_selMIO_E_reg/P0001  ;
	input \memc_usysr_DO_reg[0]/NET0131  ;
	input \memc_usysr_DO_reg[10]/NET0131  ;
	input \memc_usysr_DO_reg[11]/NET0131  ;
	input \memc_usysr_DO_reg[12]/NET0131  ;
	input \memc_usysr_DO_reg[13]/NET0131  ;
	input \memc_usysr_DO_reg[14]/NET0131  ;
	input \memc_usysr_DO_reg[15]/NET0131  ;
	input \memc_usysr_DO_reg[1]/NET0131  ;
	input \memc_usysr_DO_reg[2]/NET0131  ;
	input \memc_usysr_DO_reg[3]/NET0131  ;
	input \memc_usysr_DO_reg[4]/NET0131  ;
	input \memc_usysr_DO_reg[5]/NET0131  ;
	input \memc_usysr_DO_reg[6]/NET0131  ;
	input \memc_usysr_DO_reg[7]/NET0131  ;
	input \memc_usysr_DO_reg[8]/NET0131  ;
	input \memc_usysr_DO_reg[9]/NET0131  ;
	input \pio_PINT_reg[0]/NET0131  ;
	input \pio_PINT_reg[10]/NET0131  ;
	input \pio_PINT_reg[11]/NET0131  ;
	input \pio_PINT_reg[1]/NET0131  ;
	input \pio_PINT_reg[2]/NET0131  ;
	input \pio_PINT_reg[3]/NET0131  ;
	input \pio_PINT_reg[4]/NET0131  ;
	input \pio_PINT_reg[5]/NET0131  ;
	input \pio_PINT_reg[6]/NET0131  ;
	input \pio_PINT_reg[7]/NET0131  ;
	input \pio_PINT_reg[8]/NET0131  ;
	input \pio_PINT_reg[9]/NET0131  ;
	input \pio_PIO_IN_P_reg[0]/P0001  ;
	input \pio_PIO_IN_P_reg[10]/P0001  ;
	input \pio_PIO_IN_P_reg[11]/P0001  ;
	input \pio_PIO_IN_P_reg[1]/P0001  ;
	input \pio_PIO_IN_P_reg[2]/P0001  ;
	input \pio_PIO_IN_P_reg[3]/P0001  ;
	input \pio_PIO_IN_P_reg[4]/P0001  ;
	input \pio_PIO_IN_P_reg[5]/P0001  ;
	input \pio_PIO_IN_P_reg[6]/P0001  ;
	input \pio_PIO_IN_P_reg[7]/P0001  ;
	input \pio_PIO_IN_P_reg[8]/P0001  ;
	input \pio_PIO_IN_P_reg[9]/P0001  ;
	input \pio_PIO_RES_OUT_reg[0]/P0001  ;
	input \pio_PIO_RES_OUT_reg[10]/P0001  ;
	input \pio_PIO_RES_OUT_reg[11]/P0001  ;
	input \pio_PIO_RES_OUT_reg[1]/P0001  ;
	input \pio_PIO_RES_OUT_reg[2]/P0001  ;
	input \pio_PIO_RES_OUT_reg[3]/P0001  ;
	input \pio_PIO_RES_OUT_reg[4]/P0001  ;
	input \pio_PIO_RES_OUT_reg[5]/P0001  ;
	input \pio_PIO_RES_OUT_reg[6]/P0001  ;
	input \pio_PIO_RES_OUT_reg[7]/P0001  ;
	input \pio_PIO_RES_OUT_reg[8]/P0001  ;
	input \pio_PIO_RES_OUT_reg[9]/P0001  ;
	input \pio_PIO_RES_reg[0]/NET0131  ;
	input \pio_PIO_RES_reg[10]/NET0131  ;
	input \pio_PIO_RES_reg[11]/NET0131  ;
	input \pio_PIO_RES_reg[1]/NET0131  ;
	input \pio_PIO_RES_reg[2]/NET0131  ;
	input \pio_PIO_RES_reg[3]/NET0131  ;
	input \pio_PIO_RES_reg[4]/NET0131  ;
	input \pio_PIO_RES_reg[5]/NET0131  ;
	input \pio_PIO_RES_reg[6]/NET0131  ;
	input \pio_PIO_RES_reg[7]/NET0131  ;
	input \pio_PIO_RES_reg[8]/NET0131  ;
	input \pio_PIO_RES_reg[9]/NET0131  ;
	input \pio_pmask_reg_DO_reg[0]/NET0131  ;
	input \pio_pmask_reg_DO_reg[10]/NET0131  ;
	input \pio_pmask_reg_DO_reg[11]/NET0131  ;
	input \pio_pmask_reg_DO_reg[1]/NET0131  ;
	input \pio_pmask_reg_DO_reg[2]/NET0131  ;
	input \pio_pmask_reg_DO_reg[3]/NET0131  ;
	input \pio_pmask_reg_DO_reg[4]/NET0131  ;
	input \pio_pmask_reg_DO_reg[5]/NET0131  ;
	input \pio_pmask_reg_DO_reg[6]/NET0131  ;
	input \pio_pmask_reg_DO_reg[7]/NET0131  ;
	input \pio_pmask_reg_DO_reg[8]/NET0131  ;
	input \pio_pmask_reg_DO_reg[9]/NET0131  ;
	input \regout_STD_C_reg[0]/P0001  ;
	input \regout_STD_C_reg[10]/P0001  ;
	input \regout_STD_C_reg[11]/P0001  ;
	input \regout_STD_C_reg[12]/P0001  ;
	input \regout_STD_C_reg[13]/P0001  ;
	input \regout_STD_C_reg[14]/P0001  ;
	input \regout_STD_C_reg[15]/P0001  ;
	input \regout_STD_C_reg[1]/P0001  ;
	input \regout_STD_C_reg[2]/P0001  ;
	input \regout_STD_C_reg[3]/P0001  ;
	input \regout_STD_C_reg[4]/P0001  ;
	input \regout_STD_C_reg[5]/P0001  ;
	input \regout_STD_C_reg[6]/P0001  ;
	input \regout_STD_C_reg[7]/P0001  ;
	input \regout_STD_C_reg[8]/P0001  ;
	input \regout_STD_C_reg[9]/P0001  ;
	input \sice_CLR_I_reg/NET0131  ;
	input \sice_CLR_M_reg/NET0131  ;
	input \sice_CMRW_reg/NET0131  ;
	input \sice_DBR1_reg[0]/P0001  ;
	input \sice_DBR1_reg[10]/P0001  ;
	input \sice_DBR1_reg[11]/P0001  ;
	input \sice_DBR1_reg[12]/P0001  ;
	input \sice_DBR1_reg[13]/P0001  ;
	input \sice_DBR1_reg[14]/P0001  ;
	input \sice_DBR1_reg[15]/P0001  ;
	input \sice_DBR1_reg[16]/P0001  ;
	input \sice_DBR1_reg[17]/P0001  ;
	input \sice_DBR1_reg[18]/P0001  ;
	input \sice_DBR1_reg[1]/P0001  ;
	input \sice_DBR1_reg[2]/P0001  ;
	input \sice_DBR1_reg[3]/P0001  ;
	input \sice_DBR1_reg[4]/P0001  ;
	input \sice_DBR1_reg[5]/P0001  ;
	input \sice_DBR1_reg[6]/P0001  ;
	input \sice_DBR1_reg[7]/P0001  ;
	input \sice_DBR1_reg[8]/P0001  ;
	input \sice_DBR1_reg[9]/P0001  ;
	input \sice_DBR2_reg[0]/P0001  ;
	input \sice_DBR2_reg[10]/P0001  ;
	input \sice_DBR2_reg[11]/P0001  ;
	input \sice_DBR2_reg[12]/P0001  ;
	input \sice_DBR2_reg[13]/P0001  ;
	input \sice_DBR2_reg[14]/P0001  ;
	input \sice_DBR2_reg[15]/P0001  ;
	input \sice_DBR2_reg[16]/P0001  ;
	input \sice_DBR2_reg[17]/P0001  ;
	input \sice_DBR2_reg[18]/P0001  ;
	input \sice_DBR2_reg[1]/P0001  ;
	input \sice_DBR2_reg[2]/P0001  ;
	input \sice_DBR2_reg[3]/P0001  ;
	input \sice_DBR2_reg[4]/P0001  ;
	input \sice_DBR2_reg[5]/P0001  ;
	input \sice_DBR2_reg[6]/P0001  ;
	input \sice_DBR2_reg[7]/P0001  ;
	input \sice_DBR2_reg[8]/P0001  ;
	input \sice_DBR2_reg[9]/P0001  ;
	input \sice_DMR1_reg[0]/NET0131  ;
	input \sice_DMR1_reg[10]/NET0131  ;
	input \sice_DMR1_reg[11]/NET0131  ;
	input \sice_DMR1_reg[12]/NET0131  ;
	input \sice_DMR1_reg[13]/NET0131  ;
	input \sice_DMR1_reg[14]/NET0131  ;
	input \sice_DMR1_reg[15]/NET0131  ;
	input \sice_DMR1_reg[16]/NET0131  ;
	input \sice_DMR1_reg[17]/NET0131  ;
	input \sice_DMR1_reg[1]/NET0131  ;
	input \sice_DMR1_reg[2]/NET0131  ;
	input \sice_DMR1_reg[3]/NET0131  ;
	input \sice_DMR1_reg[4]/NET0131  ;
	input \sice_DMR1_reg[5]/NET0131  ;
	input \sice_DMR1_reg[6]/NET0131  ;
	input \sice_DMR1_reg[7]/NET0131  ;
	input \sice_DMR1_reg[8]/NET0131  ;
	input \sice_DMR1_reg[9]/NET0131  ;
	input \sice_DMR2_reg[0]/NET0131  ;
	input \sice_DMR2_reg[10]/NET0131  ;
	input \sice_DMR2_reg[11]/NET0131  ;
	input \sice_DMR2_reg[12]/NET0131  ;
	input \sice_DMR2_reg[13]/NET0131  ;
	input \sice_DMR2_reg[14]/NET0131  ;
	input \sice_DMR2_reg[15]/NET0131  ;
	input \sice_DMR2_reg[16]/NET0131  ;
	input \sice_DMR2_reg[17]/NET0131  ;
	input \sice_DMR2_reg[1]/NET0131  ;
	input \sice_DMR2_reg[2]/NET0131  ;
	input \sice_DMR2_reg[3]/NET0131  ;
	input \sice_DMR2_reg[4]/NET0131  ;
	input \sice_DMR2_reg[5]/NET0131  ;
	input \sice_DMR2_reg[6]/NET0131  ;
	input \sice_DMR2_reg[7]/NET0131  ;
	input \sice_DMR2_reg[8]/NET0131  ;
	input \sice_DMR2_reg[9]/NET0131  ;
	input \sice_GOICE_1_reg/NET0131  ;
	input \sice_GOICE_2_reg/NET0131  ;
	input \sice_GOICE_s1_reg/NET0131  ;
	input \sice_GOICE_syn_reg/P0001  ;
	input \sice_GO_NX_reg/NET0131  ;
	input \sice_GO_NXi_reg/NET0131  ;
	input \sice_HALT_E_reg/P0001  ;
	input \sice_IAR_reg[0]/NET0131  ;
	input \sice_IAR_reg[1]/NET0131  ;
	input \sice_IAR_reg[2]/NET0131  ;
	input \sice_IAR_reg[3]/NET0131  ;
	input \sice_IBR1_reg[0]/P0001  ;
	input \sice_IBR1_reg[10]/P0001  ;
	input \sice_IBR1_reg[11]/P0001  ;
	input \sice_IBR1_reg[12]/P0001  ;
	input \sice_IBR1_reg[13]/P0001  ;
	input \sice_IBR1_reg[14]/P0001  ;
	input \sice_IBR1_reg[15]/P0001  ;
	input \sice_IBR1_reg[16]/P0001  ;
	input \sice_IBR1_reg[17]/P0001  ;
	input \sice_IBR1_reg[1]/P0001  ;
	input \sice_IBR1_reg[2]/P0001  ;
	input \sice_IBR1_reg[3]/P0001  ;
	input \sice_IBR1_reg[4]/P0001  ;
	input \sice_IBR1_reg[5]/P0001  ;
	input \sice_IBR1_reg[6]/P0001  ;
	input \sice_IBR1_reg[7]/P0001  ;
	input \sice_IBR1_reg[8]/P0001  ;
	input \sice_IBR1_reg[9]/P0001  ;
	input \sice_IBR2_reg[0]/P0001  ;
	input \sice_IBR2_reg[10]/P0001  ;
	input \sice_IBR2_reg[11]/P0001  ;
	input \sice_IBR2_reg[12]/P0001  ;
	input \sice_IBR2_reg[13]/P0001  ;
	input \sice_IBR2_reg[14]/P0001  ;
	input \sice_IBR2_reg[15]/P0001  ;
	input \sice_IBR2_reg[16]/P0001  ;
	input \sice_IBR2_reg[17]/P0001  ;
	input \sice_IBR2_reg[1]/P0001  ;
	input \sice_IBR2_reg[2]/P0001  ;
	input \sice_IBR2_reg[3]/P0001  ;
	input \sice_IBR2_reg[4]/P0001  ;
	input \sice_IBR2_reg[5]/P0001  ;
	input \sice_IBR2_reg[6]/P0001  ;
	input \sice_IBR2_reg[7]/P0001  ;
	input \sice_IBR2_reg[8]/P0001  ;
	input \sice_IBR2_reg[9]/P0001  ;
	input \sice_ICS_reg[0]/NET0131  ;
	input \sice_ICS_reg[1]/NET0131  ;
	input \sice_ICS_reg[2]/NET0131  ;
	input \sice_ICYC_clr_reg/NET0131  ;
	input \sice_ICYC_en_reg/NET0131  ;
	input \sice_ICYC_en_syn_reg/P0001  ;
	input \sice_ICYC_reg[0]/NET0131  ;
	input \sice_ICYC_reg[10]/NET0131  ;
	input \sice_ICYC_reg[11]/NET0131  ;
	input \sice_ICYC_reg[12]/NET0131  ;
	input \sice_ICYC_reg[13]/NET0131  ;
	input \sice_ICYC_reg[14]/NET0131  ;
	input \sice_ICYC_reg[15]/NET0131  ;
	input \sice_ICYC_reg[16]/NET0131  ;
	input \sice_ICYC_reg[17]/NET0131  ;
	input \sice_ICYC_reg[18]/NET0131  ;
	input \sice_ICYC_reg[19]/NET0131  ;
	input \sice_ICYC_reg[1]/NET0131  ;
	input \sice_ICYC_reg[20]/NET0131  ;
	input \sice_ICYC_reg[21]/NET0131  ;
	input \sice_ICYC_reg[22]/NET0131  ;
	input \sice_ICYC_reg[23]/NET0131  ;
	input \sice_ICYC_reg[2]/NET0131  ;
	input \sice_ICYC_reg[3]/NET0131  ;
	input \sice_ICYC_reg[4]/NET0131  ;
	input \sice_ICYC_reg[5]/NET0131  ;
	input \sice_ICYC_reg[6]/NET0131  ;
	input \sice_ICYC_reg[7]/NET0131  ;
	input \sice_ICYC_reg[8]/NET0131  ;
	input \sice_ICYC_reg[9]/NET0131  ;
	input \sice_IDONE_reg/NET0131  ;
	input \sice_IIRC_reg[0]/NET0131  ;
	input \sice_IIRC_reg[10]/NET0131  ;
	input \sice_IIRC_reg[11]/NET0131  ;
	input \sice_IIRC_reg[12]/NET0131  ;
	input \sice_IIRC_reg[13]/NET0131  ;
	input \sice_IIRC_reg[14]/NET0131  ;
	input \sice_IIRC_reg[15]/NET0131  ;
	input \sice_IIRC_reg[16]/NET0131  ;
	input \sice_IIRC_reg[17]/NET0131  ;
	input \sice_IIRC_reg[18]/NET0131  ;
	input \sice_IIRC_reg[19]/NET0131  ;
	input \sice_IIRC_reg[1]/NET0131  ;
	input \sice_IIRC_reg[20]/NET0131  ;
	input \sice_IIRC_reg[21]/NET0131  ;
	input \sice_IIRC_reg[22]/NET0131  ;
	input \sice_IIRC_reg[23]/NET0131  ;
	input \sice_IIRC_reg[2]/NET0131  ;
	input \sice_IIRC_reg[3]/NET0131  ;
	input \sice_IIRC_reg[4]/NET0131  ;
	input \sice_IIRC_reg[5]/NET0131  ;
	input \sice_IIRC_reg[6]/NET0131  ;
	input \sice_IIRC_reg[7]/NET0131  ;
	input \sice_IIRC_reg[8]/NET0131  ;
	input \sice_IIRC_reg[9]/NET0131  ;
	input \sice_IMR1_reg[0]/NET0131  ;
	input \sice_IMR1_reg[10]/NET0131  ;
	input \sice_IMR1_reg[11]/NET0131  ;
	input \sice_IMR1_reg[12]/NET0131  ;
	input \sice_IMR1_reg[13]/NET0131  ;
	input \sice_IMR1_reg[14]/NET0131  ;
	input \sice_IMR1_reg[15]/NET0131  ;
	input \sice_IMR1_reg[16]/NET0131  ;
	input \sice_IMR1_reg[17]/NET0131  ;
	input \sice_IMR1_reg[1]/NET0131  ;
	input \sice_IMR1_reg[2]/NET0131  ;
	input \sice_IMR1_reg[3]/NET0131  ;
	input \sice_IMR1_reg[4]/NET0131  ;
	input \sice_IMR1_reg[5]/NET0131  ;
	input \sice_IMR1_reg[6]/NET0131  ;
	input \sice_IMR1_reg[7]/NET0131  ;
	input \sice_IMR1_reg[8]/NET0131  ;
	input \sice_IMR1_reg[9]/NET0131  ;
	input \sice_IMR2_reg[0]/NET0131  ;
	input \sice_IMR2_reg[10]/NET0131  ;
	input \sice_IMR2_reg[11]/NET0131  ;
	input \sice_IMR2_reg[12]/NET0131  ;
	input \sice_IMR2_reg[13]/NET0131  ;
	input \sice_IMR2_reg[14]/NET0131  ;
	input \sice_IMR2_reg[15]/NET0131  ;
	input \sice_IMR2_reg[16]/NET0131  ;
	input \sice_IMR2_reg[17]/NET0131  ;
	input \sice_IMR2_reg[1]/NET0131  ;
	input \sice_IMR2_reg[2]/NET0131  ;
	input \sice_IMR2_reg[3]/NET0131  ;
	input \sice_IMR2_reg[4]/NET0131  ;
	input \sice_IMR2_reg[5]/NET0131  ;
	input \sice_IMR2_reg[6]/NET0131  ;
	input \sice_IMR2_reg[7]/NET0131  ;
	input \sice_IMR2_reg[8]/NET0131  ;
	input \sice_IMR2_reg[9]/NET0131  ;
	input \sice_IRR_reg[0]/P0001  ;
	input \sice_IRR_reg[10]/P0001  ;
	input \sice_IRR_reg[11]/P0001  ;
	input \sice_IRR_reg[12]/P0001  ;
	input \sice_IRR_reg[13]/P0001  ;
	input \sice_IRR_reg[1]/P0001  ;
	input \sice_IRR_reg[2]/P0001  ;
	input \sice_IRR_reg[3]/P0001  ;
	input \sice_IRR_reg[4]/P0001  ;
	input \sice_IRR_reg[5]/P0001  ;
	input \sice_IRR_reg[6]/P0001  ;
	input \sice_IRR_reg[7]/P0001  ;
	input \sice_IRR_reg[8]/P0001  ;
	input \sice_IRR_reg[9]/P0001  ;
	input \sice_IRST_reg/NET0131  ;
	input \sice_IRST_syn_reg/P0001  ;
	input \sice_ITR_reg[0]/NET0131  ;
	input \sice_ITR_reg[1]/NET0131  ;
	input \sice_ITR_reg[2]/NET0131  ;
	input \sice_OE_reg/P0001  ;
	input \sice_RCS_reg[0]/NET0131  ;
	input \sice_RCS_reg[1]/NET0131  ;
	input \sice_RST_req_reg/NET0131  ;
	input \sice_SPC_reg[0]/P0001  ;
	input \sice_SPC_reg[10]/P0001  ;
	input \sice_SPC_reg[11]/P0001  ;
	input \sice_SPC_reg[12]/P0001  ;
	input \sice_SPC_reg[13]/P0001  ;
	input \sice_SPC_reg[14]/P0001  ;
	input \sice_SPC_reg[15]/P0001  ;
	input \sice_SPC_reg[16]/P0001  ;
	input \sice_SPC_reg[17]/P0001  ;
	input \sice_SPC_reg[18]/P0001  ;
	input \sice_SPC_reg[19]/P0001  ;
	input \sice_SPC_reg[1]/P0001  ;
	input \sice_SPC_reg[20]/P0001  ;
	input \sice_SPC_reg[21]/P0001  ;
	input \sice_SPC_reg[22]/P0001  ;
	input \sice_SPC_reg[23]/P0001  ;
	input \sice_SPC_reg[2]/P0001  ;
	input \sice_SPC_reg[3]/P0001  ;
	input \sice_SPC_reg[4]/P0001  ;
	input \sice_SPC_reg[5]/P0001  ;
	input \sice_SPC_reg[6]/P0001  ;
	input \sice_SPC_reg[7]/P0001  ;
	input \sice_SPC_reg[8]/P0001  ;
	input \sice_SPC_reg[9]/P0001  ;
	input \sice_UpdDR_sd1_reg/P0001  ;
	input \sice_UpdDR_sd2_reg/P0001  ;
	input \sice_idr0_reg_DO_reg[0]/P0001  ;
	input \sice_idr0_reg_DO_reg[10]/P0001  ;
	input \sice_idr0_reg_DO_reg[11]/P0001  ;
	input \sice_idr0_reg_DO_reg[1]/P0001  ;
	input \sice_idr0_reg_DO_reg[2]/P0001  ;
	input \sice_idr0_reg_DO_reg[3]/P0001  ;
	input \sice_idr0_reg_DO_reg[4]/P0001  ;
	input \sice_idr0_reg_DO_reg[5]/P0001  ;
	input \sice_idr0_reg_DO_reg[6]/P0001  ;
	input \sice_idr0_reg_DO_reg[7]/P0001  ;
	input \sice_idr0_reg_DO_reg[8]/P0001  ;
	input \sice_idr0_reg_DO_reg[9]/P0001  ;
	input \sice_idr1_reg_DO_reg[0]/P0001  ;
	input \sice_idr1_reg_DO_reg[10]/P0001  ;
	input \sice_idr1_reg_DO_reg[11]/P0001  ;
	input \sice_idr1_reg_DO_reg[1]/P0001  ;
	input \sice_idr1_reg_DO_reg[2]/P0001  ;
	input \sice_idr1_reg_DO_reg[3]/P0001  ;
	input \sice_idr1_reg_DO_reg[4]/P0001  ;
	input \sice_idr1_reg_DO_reg[5]/P0001  ;
	input \sice_idr1_reg_DO_reg[6]/P0001  ;
	input \sice_idr1_reg_DO_reg[7]/P0001  ;
	input \sice_idr1_reg_DO_reg[8]/P0001  ;
	input \sice_idr1_reg_DO_reg[9]/P0001  ;
	input \sport0_cfg_FSi_cnt_reg[0]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[10]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[11]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[12]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[13]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[14]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[15]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[1]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[2]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[3]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[4]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[5]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[6]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[7]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[8]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[9]/NET0131  ;
	input \sport0_cfg_FSi_reg/NET0131  ;
	input \sport0_cfg_RFSg_d1_reg/NET0131  ;
	input \sport0_cfg_RFSg_d2_reg/NET0131  ;
	input \sport0_cfg_RFSg_d3_reg/NET0131  ;
	input \sport0_cfg_RFSgi_d_reg/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[0]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[10]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[11]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[12]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[13]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[14]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[15]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[1]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[2]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[3]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[4]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[5]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[6]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[7]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[8]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[9]/NET0131  ;
	input \sport0_cfg_SCLKi_h_reg/NET0131  ;
	input \sport0_cfg_SP_ENg_D1_reg/P0001  ;
	input \sport0_cfg_SP_ENg_reg/NET0131  ;
	input \sport0_cfg_TFSg_d1_reg/NET0131  ;
	input \sport0_cfg_TFSg_d2_reg/NET0131  ;
	input \sport0_cfg_TFSg_d3_reg/NET0131  ;
	input \sport0_cfg_TFSgi_d_reg/NET0131  ;
	input \sport0_regs_AUTO_a_reg[12]/NET0131  ;
	input \sport0_regs_AUTO_a_reg[13]/NET0131  ;
	input \sport0_regs_AUTO_a_reg[14]/NET0131  ;
	input \sport0_regs_AUTO_a_reg[15]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[11]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[7]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[8]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[9]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[11]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[12]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[13]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[14]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[15]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[7]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[8]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[9]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[7]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[8]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[9]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[11]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[12]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[13]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[15]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[7]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[0]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[1]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[2]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[3]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[4]/NET0131  ;
	input \sport0_rxctl_ISRa_reg/P0001  ;
	input \sport0_rxctl_LMcnt_reg[0]/NET0131  ;
	input \sport0_rxctl_LMcnt_reg[1]/NET0131  ;
	input \sport0_rxctl_LMcnt_reg[2]/NET0131  ;
	input \sport0_rxctl_LMcnt_reg[3]/NET0131  ;
	input \sport0_rxctl_LMcnt_reg[4]/NET0131  ;
	input \sport0_rxctl_RCS_reg[0]/NET0131  ;
	input \sport0_rxctl_RCS_reg[1]/NET0131  ;
	input \sport0_rxctl_RCS_reg[2]/NET0131  ;
	input \sport0_rxctl_RSreq_reg/NET0131  ;
	input \sport0_rxctl_RXSHT_reg[0]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[10]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[11]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[12]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[13]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[14]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[15]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[1]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[2]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[3]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[4]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[5]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[6]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[7]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[8]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[9]/P0001  ;
	input \sport0_rxctl_RX_reg[0]/P0001  ;
	input \sport0_rxctl_RX_reg[10]/P0001  ;
	input \sport0_rxctl_RX_reg[11]/P0001  ;
	input \sport0_rxctl_RX_reg[12]/P0001  ;
	input \sport0_rxctl_RX_reg[13]/P0001  ;
	input \sport0_rxctl_RX_reg[14]/P0001  ;
	input \sport0_rxctl_RX_reg[15]/P0001  ;
	input \sport0_rxctl_RX_reg[1]/P0001  ;
	input \sport0_rxctl_RX_reg[2]/P0001  ;
	input \sport0_rxctl_RX_reg[3]/P0001  ;
	input \sport0_rxctl_RX_reg[4]/P0001  ;
	input \sport0_rxctl_RX_reg[5]/P0001  ;
	input \sport0_rxctl_RX_reg[6]/P0001  ;
	input \sport0_rxctl_RX_reg[7]/P0001  ;
	input \sport0_rxctl_RX_reg[8]/P0001  ;
	input \sport0_rxctl_RX_reg[9]/P0001  ;
	input \sport0_rxctl_SLOT1_EXT_reg[2]/NET0131  ;
	input \sport0_rxctl_SLOT1_EXT_reg[3]/NET0131  ;
	input \sport0_rxctl_TAG_SLOT_reg/P0001  ;
	input \sport0_rxctl_Wcnt_reg[0]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[1]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[2]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[3]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[4]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[5]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[6]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[7]/NET0131  ;
	input \sport0_rxctl_a_sync1_reg/P0001  ;
	input \sport0_rxctl_a_sync2_reg/P0001  ;
	input \sport0_rxctl_ldRX_cmp_reg/P0001  ;
	input \sport0_rxctl_sht2nd_reg/P0001  ;
	input \sport0_txctl_Bcnt_reg[0]/NET0131  ;
	input \sport0_txctl_Bcnt_reg[1]/NET0131  ;
	input \sport0_txctl_Bcnt_reg[2]/NET0131  ;
	input \sport0_txctl_Bcnt_reg[3]/NET0131  ;
	input \sport0_txctl_Bcnt_reg[4]/NET0131  ;
	input \sport0_txctl_SP_EN_D1_reg/P0001  ;
	input \sport0_txctl_TCS_reg[0]/NET0131  ;
	input \sport0_txctl_TCS_reg[1]/NET0131  ;
	input \sport0_txctl_TCS_reg[2]/NET0131  ;
	input \sport0_txctl_TSreq_reg/NET0131  ;
	input \sport0_txctl_TSreqi_reg/NET0131  ;
	input \sport0_txctl_TXSHT_reg[0]/P0001  ;
	input \sport0_txctl_TXSHT_reg[10]/P0001  ;
	input \sport0_txctl_TXSHT_reg[11]/P0001  ;
	input \sport0_txctl_TXSHT_reg[12]/P0001  ;
	input \sport0_txctl_TXSHT_reg[13]/P0001  ;
	input \sport0_txctl_TXSHT_reg[14]/P0001  ;
	input \sport0_txctl_TXSHT_reg[15]/P0001  ;
	input \sport0_txctl_TXSHT_reg[1]/P0001  ;
	input \sport0_txctl_TXSHT_reg[2]/P0001  ;
	input \sport0_txctl_TXSHT_reg[3]/P0001  ;
	input \sport0_txctl_TXSHT_reg[4]/P0001  ;
	input \sport0_txctl_TXSHT_reg[5]/P0001  ;
	input \sport0_txctl_TXSHT_reg[6]/P0001  ;
	input \sport0_txctl_TXSHT_reg[7]/P0001  ;
	input \sport0_txctl_TXSHT_reg[8]/P0001  ;
	input \sport0_txctl_TXSHT_reg[9]/P0001  ;
	input \sport0_txctl_TX_reg[0]/P0001  ;
	input \sport0_txctl_TX_reg[10]/P0001  ;
	input \sport0_txctl_TX_reg[11]/P0001  ;
	input \sport0_txctl_TX_reg[12]/P0001  ;
	input \sport0_txctl_TX_reg[13]/P0001  ;
	input \sport0_txctl_TX_reg[14]/P0001  ;
	input \sport0_txctl_TX_reg[15]/P0001  ;
	input \sport0_txctl_TX_reg[1]/P0001  ;
	input \sport0_txctl_TX_reg[2]/P0001  ;
	input \sport0_txctl_TX_reg[3]/P0001  ;
	input \sport0_txctl_TX_reg[4]/P0001  ;
	input \sport0_txctl_TX_reg[5]/P0001  ;
	input \sport0_txctl_TX_reg[6]/P0001  ;
	input \sport0_txctl_TX_reg[7]/P0001  ;
	input \sport0_txctl_TX_reg[8]/P0001  ;
	input \sport0_txctl_TX_reg[9]/P0001  ;
	input \sport0_txctl_Wcnt_reg[0]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[1]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[2]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[3]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[4]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[5]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[6]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[7]/NET0131  ;
	input \sport0_txctl_b_sync1_reg/P0001  ;
	input \sport0_txctl_c_sync1_reg/P0001  ;
	input \sport0_txctl_c_sync2_reg/P0001  ;
	input \sport0_txctl_ldTX_cmp_reg/P0001  ;
	input \sport1_cfg_FSi_cnt_reg[0]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[10]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[11]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[12]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[13]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[14]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[15]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[1]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[2]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[3]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[4]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[5]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[6]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[7]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[8]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[9]/NET0131  ;
	input \sport1_cfg_FSi_reg/NET0131  ;
	input \sport1_cfg_RFSg_d1_reg/NET0131  ;
	input \sport1_cfg_RFSg_d2_reg/NET0131  ;
	input \sport1_cfg_RFSg_d3_reg/NET0131  ;
	input \sport1_cfg_RFSgi_d_reg/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[0]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[10]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[11]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[12]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[13]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[14]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[15]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[1]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[2]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[3]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[4]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[5]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[6]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[7]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[8]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[9]/NET0131  ;
	input \sport1_cfg_SCLKi_h_reg/NET0131  ;
	input \sport1_cfg_SP_ENg_D1_reg/P0001  ;
	input \sport1_cfg_SP_ENg_reg/NET0131  ;
	input \sport1_cfg_TFSg_d1_reg/NET0131  ;
	input \sport1_cfg_TFSg_d2_reg/NET0131  ;
	input \sport1_cfg_TFSg_d3_reg/NET0131  ;
	input \sport1_cfg_TFSgi_d_reg/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[11]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[7]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[8]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[9]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[11]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[12]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[13]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[14]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[15]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[7]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[8]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[9]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[7]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[8]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[9]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[11]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[12]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[13]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[15]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[7]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[0]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[1]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[2]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[3]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[4]/NET0131  ;
	input \sport1_rxctl_ISRa_reg/P0001  ;
	input \sport1_rxctl_LMcnt_reg[0]/NET0131  ;
	input \sport1_rxctl_LMcnt_reg[1]/NET0131  ;
	input \sport1_rxctl_LMcnt_reg[2]/NET0131  ;
	input \sport1_rxctl_LMcnt_reg[3]/NET0131  ;
	input \sport1_rxctl_LMcnt_reg[4]/NET0131  ;
	input \sport1_rxctl_RCS_reg[0]/NET0131  ;
	input \sport1_rxctl_RCS_reg[1]/NET0131  ;
	input \sport1_rxctl_RCS_reg[2]/NET0131  ;
	input \sport1_rxctl_RSreq_reg/NET0131  ;
	input \sport1_rxctl_RXSHT_reg[0]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[10]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[11]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[12]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[13]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[14]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[15]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[1]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[2]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[3]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[4]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[5]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[6]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[7]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[8]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[9]/P0001  ;
	input \sport1_rxctl_RX_reg[0]/P0001  ;
	input \sport1_rxctl_RX_reg[10]/P0001  ;
	input \sport1_rxctl_RX_reg[11]/P0001  ;
	input \sport1_rxctl_RX_reg[12]/P0001  ;
	input \sport1_rxctl_RX_reg[13]/P0001  ;
	input \sport1_rxctl_RX_reg[14]/P0001  ;
	input \sport1_rxctl_RX_reg[15]/P0001  ;
	input \sport1_rxctl_RX_reg[1]/P0001  ;
	input \sport1_rxctl_RX_reg[2]/P0001  ;
	input \sport1_rxctl_RX_reg[3]/P0001  ;
	input \sport1_rxctl_RX_reg[4]/P0001  ;
	input \sport1_rxctl_RX_reg[5]/P0001  ;
	input \sport1_rxctl_RX_reg[6]/P0001  ;
	input \sport1_rxctl_RX_reg[7]/P0001  ;
	input \sport1_rxctl_RX_reg[8]/P0001  ;
	input \sport1_rxctl_RX_reg[9]/P0001  ;
	input \sport1_rxctl_SLOT1_EXT_reg[2]/NET0131  ;
	input \sport1_rxctl_SLOT1_EXT_reg[3]/NET0131  ;
	input \sport1_rxctl_TAG_SLOT_reg/P0001  ;
	input \sport1_rxctl_Wcnt_reg[0]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[1]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[2]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[3]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[4]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[5]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[6]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[7]/NET0131  ;
	input \sport1_rxctl_a_sync1_reg/P0001  ;
	input \sport1_rxctl_a_sync2_reg/P0001  ;
	input \sport1_rxctl_sht2nd_reg/P0001  ;
	input \sport1_txctl_Bcnt_reg[0]/NET0131  ;
	input \sport1_txctl_Bcnt_reg[1]/NET0131  ;
	input \sport1_txctl_Bcnt_reg[2]/NET0131  ;
	input \sport1_txctl_Bcnt_reg[3]/NET0131  ;
	input \sport1_txctl_Bcnt_reg[4]/NET0131  ;
	input \sport1_txctl_SP_EN_D1_reg/P0001  ;
	input \sport1_txctl_TCS_reg[0]/NET0131  ;
	input \sport1_txctl_TCS_reg[1]/NET0131  ;
	input \sport1_txctl_TCS_reg[2]/NET0131  ;
	input \sport1_txctl_TSreq_reg/NET0131  ;
	input \sport1_txctl_TSreqi_reg/NET0131  ;
	input \sport1_txctl_TXSHT_reg[0]/P0001  ;
	input \sport1_txctl_TXSHT_reg[10]/P0001  ;
	input \sport1_txctl_TXSHT_reg[11]/P0001  ;
	input \sport1_txctl_TXSHT_reg[12]/P0001  ;
	input \sport1_txctl_TXSHT_reg[13]/P0001  ;
	input \sport1_txctl_TXSHT_reg[14]/P0001  ;
	input \sport1_txctl_TXSHT_reg[15]/P0001  ;
	input \sport1_txctl_TXSHT_reg[1]/P0001  ;
	input \sport1_txctl_TXSHT_reg[2]/P0001  ;
	input \sport1_txctl_TXSHT_reg[3]/P0001  ;
	input \sport1_txctl_TXSHT_reg[4]/P0001  ;
	input \sport1_txctl_TXSHT_reg[5]/P0001  ;
	input \sport1_txctl_TXSHT_reg[6]/P0001  ;
	input \sport1_txctl_TXSHT_reg[7]/P0001  ;
	input \sport1_txctl_TXSHT_reg[8]/P0001  ;
	input \sport1_txctl_TXSHT_reg[9]/P0001  ;
	input \sport1_txctl_TX_reg[0]/P0001  ;
	input \sport1_txctl_TX_reg[10]/P0001  ;
	input \sport1_txctl_TX_reg[11]/P0001  ;
	input \sport1_txctl_TX_reg[12]/P0001  ;
	input \sport1_txctl_TX_reg[13]/P0001  ;
	input \sport1_txctl_TX_reg[14]/P0001  ;
	input \sport1_txctl_TX_reg[15]/P0001  ;
	input \sport1_txctl_TX_reg[1]/P0001  ;
	input \sport1_txctl_TX_reg[2]/P0001  ;
	input \sport1_txctl_TX_reg[3]/P0001  ;
	input \sport1_txctl_TX_reg[4]/P0001  ;
	input \sport1_txctl_TX_reg[5]/P0001  ;
	input \sport1_txctl_TX_reg[6]/P0001  ;
	input \sport1_txctl_TX_reg[7]/P0001  ;
	input \sport1_txctl_TX_reg[8]/P0001  ;
	input \sport1_txctl_TX_reg[9]/P0001  ;
	input \sport1_txctl_Wcnt_reg[0]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[1]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[2]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[3]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[4]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[5]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[6]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[7]/NET0131  ;
	input \sport1_txctl_c_sync1_reg/P0001  ;
	input \sport1_txctl_c_sync2_reg/P0001  ;
	input \tm_MSTAT5_syn_reg/NET0131  ;
	input \tm_TCR_TMP_reg[0]/NET0131  ;
	input \tm_TCR_TMP_reg[10]/NET0131  ;
	input \tm_TCR_TMP_reg[11]/NET0131  ;
	input \tm_TCR_TMP_reg[12]/NET0131  ;
	input \tm_TCR_TMP_reg[13]/NET0131  ;
	input \tm_TCR_TMP_reg[14]/NET0131  ;
	input \tm_TCR_TMP_reg[15]/NET0131  ;
	input \tm_TCR_TMP_reg[1]/NET0131  ;
	input \tm_TCR_TMP_reg[2]/NET0131  ;
	input \tm_TCR_TMP_reg[3]/NET0131  ;
	input \tm_TCR_TMP_reg[4]/NET0131  ;
	input \tm_TCR_TMP_reg[5]/NET0131  ;
	input \tm_TCR_TMP_reg[6]/NET0131  ;
	input \tm_TCR_TMP_reg[7]/NET0131  ;
	input \tm_TCR_TMP_reg[8]/NET0131  ;
	input \tm_TCR_TMP_reg[9]/NET0131  ;
	input \tm_TINT_GEN1_reg/NET0131  ;
	input \tm_TINT_GEN2_reg/NET0131  ;
	input \tm_TSR_TMP_reg[0]/NET0131  ;
	input \tm_TSR_TMP_reg[1]/NET0131  ;
	input \tm_TSR_TMP_reg[2]/NET0131  ;
	input \tm_TSR_TMP_reg[3]/NET0131  ;
	input \tm_TSR_TMP_reg[4]/NET0131  ;
	input \tm_TSR_TMP_reg[5]/NET0131  ;
	input \tm_TSR_TMP_reg[6]/NET0131  ;
	input \tm_TSR_TMP_reg[7]/NET0131  ;
	input \tm_WR_TCR_KEEP_TO_TMCLK_p_reg/NET0131  ;
	input \tm_WR_TCR_TMP_GEN1_reg/P0001  ;
	input \tm_WR_TCR_TMP_GEN2_reg/P0001  ;
	input \tm_WR_TCR_p_reg/P0001  ;
	input \tm_WR_TSR_KEEP_TO_TMCLK_p_reg/NET0131  ;
	input \tm_WR_TSR_TMP_GEN1_reg/P0001  ;
	input \tm_WR_TSR_TMP_GEN2_reg/P0001  ;
	input \tm_WR_TSR_p_reg/P0001  ;
	input \tm_tcr_reg_DO_reg[0]/NET0131  ;
	input \tm_tcr_reg_DO_reg[10]/NET0131  ;
	input \tm_tcr_reg_DO_reg[11]/NET0131  ;
	input \tm_tcr_reg_DO_reg[12]/NET0131  ;
	input \tm_tcr_reg_DO_reg[13]/NET0131  ;
	input \tm_tcr_reg_DO_reg[14]/NET0131  ;
	input \tm_tcr_reg_DO_reg[15]/NET0131  ;
	input \tm_tcr_reg_DO_reg[1]/NET0131  ;
	input \tm_tcr_reg_DO_reg[2]/NET0131  ;
	input \tm_tcr_reg_DO_reg[3]/NET0131  ;
	input \tm_tcr_reg_DO_reg[4]/NET0131  ;
	input \tm_tcr_reg_DO_reg[5]/NET0131  ;
	input \tm_tcr_reg_DO_reg[6]/NET0131  ;
	input \tm_tcr_reg_DO_reg[7]/NET0131  ;
	input \tm_tcr_reg_DO_reg[8]/NET0131  ;
	input \tm_tcr_reg_DO_reg[9]/NET0131  ;
	input \tm_tpr_reg_DO_reg[0]/NET0131  ;
	input \tm_tpr_reg_DO_reg[10]/NET0131  ;
	input \tm_tpr_reg_DO_reg[11]/NET0131  ;
	input \tm_tpr_reg_DO_reg[12]/NET0131  ;
	input \tm_tpr_reg_DO_reg[13]/NET0131  ;
	input \tm_tpr_reg_DO_reg[14]/NET0131  ;
	input \tm_tpr_reg_DO_reg[15]/NET0131  ;
	input \tm_tpr_reg_DO_reg[1]/NET0131  ;
	input \tm_tpr_reg_DO_reg[2]/NET0131  ;
	input \tm_tpr_reg_DO_reg[3]/NET0131  ;
	input \tm_tpr_reg_DO_reg[4]/NET0131  ;
	input \tm_tpr_reg_DO_reg[5]/NET0131  ;
	input \tm_tpr_reg_DO_reg[6]/NET0131  ;
	input \tm_tpr_reg_DO_reg[7]/NET0131  ;
	input \tm_tpr_reg_DO_reg[8]/NET0131  ;
	input \tm_tpr_reg_DO_reg[9]/NET0131  ;
	input \tm_tsr_reg_DO_reg[0]/NET0131  ;
	input \tm_tsr_reg_DO_reg[1]/NET0131  ;
	input \tm_tsr_reg_DO_reg[2]/NET0131  ;
	input \tm_tsr_reg_DO_reg[3]/NET0131  ;
	input \tm_tsr_reg_DO_reg[4]/NET0131  ;
	input \tm_tsr_reg_DO_reg[5]/NET0131  ;
	input \tm_tsr_reg_DO_reg[6]/NET0131  ;
	input \tm_tsr_reg_DO_reg[7]/NET0131  ;
	input \tm_tsr_reg_DO_reg[8]/NET0131  ;
	output CLKO_pad ;
	output \CMAinx[0]_pad  ;
	output \CMAinx[10]_pad  ;
	output \CMAinx[11]_pad  ;
	output \CMAinx[1]_pad  ;
	output \CMAinx[2]_pad  ;
	output \CMAinx[3]_pad  ;
	output \CMAinx[4]_pad  ;
	output \CMAinx[5]_pad  ;
	output \CMAinx[6]_pad  ;
	output \CMAinx[7]_pad  ;
	output \CMAinx[8]_pad  ;
	output \CMAinx[9]_pad  ;
	output CMSn_pad ;
	output CM_cs_pad ;
	output \CM_wd[0]_pad  ;
	output \CM_wd[10]_pad  ;
	output \CM_wd[11]_pad  ;
	output \CM_wd[12]_pad  ;
	output \CM_wd[13]_pad  ;
	output \CM_wd[14]_pad  ;
	output \CM_wd[15]_pad  ;
	output \CM_wd[16]_pad  ;
	output \CM_wd[17]_pad  ;
	output \CM_wd[18]_pad  ;
	output \CM_wd[19]_pad  ;
	output \CM_wd[1]_pad  ;
	output \CM_wd[20]_pad  ;
	output \CM_wd[21]_pad  ;
	output \CM_wd[22]_pad  ;
	output \CM_wd[23]_pad  ;
	output \CM_wd[2]_pad  ;
	output \CM_wd[3]_pad  ;
	output \CM_wd[4]_pad  ;
	output \CM_wd[5]_pad  ;
	output \CM_wd[6]_pad  ;
	output \CM_wd[7]_pad  ;
	output \CM_wd[8]_pad  ;
	output \CM_wd[9]_pad  ;
	output CM_web_pad ;
	output \CMo_cs0_pad  ;
	output \CMo_cs1_pad  ;
	output \CMo_cs2_pad  ;
	output \CMo_cs3_pad  ;
	output \CMo_cs4_pad  ;
	output \CMo_cs5_pad  ;
	output \CMo_cs6_pad  ;
	output \CMo_cs7_pad  ;
	output \DMAinx[0]_pad  ;
	output \DMAinx[10]_pad  ;
	output \DMAinx[11]_pad  ;
	output \DMAinx[12]_pad  ;
	output \DMAinx[13]_pad  ;
	output \DMAinx[1]_pad  ;
	output \DMAinx[2]_pad  ;
	output \DMAinx[3]_pad  ;
	output \DMAinx[4]_pad  ;
	output \DMAinx[5]_pad  ;
	output \DMAinx[6]_pad  ;
	output \DMAinx[7]_pad  ;
	output \DMAinx[8]_pad  ;
	output \DMAinx[9]_pad  ;
	output DMSn_pad ;
	output DM_cs_pad ;
	output \DM_wd[0]_pad  ;
	output \DM_wd[10]_pad  ;
	output \DM_wd[11]_pad  ;
	output \DM_wd[12]_pad  ;
	output \DM_wd[13]_pad  ;
	output \DM_wd[14]_pad  ;
	output \DM_wd[15]_pad  ;
	output \DM_wd[1]_pad  ;
	output \DM_wd[2]_pad  ;
	output \DM_wd[3]_pad  ;
	output \DM_wd[4]_pad  ;
	output \DM_wd[5]_pad  ;
	output \DM_wd[6]_pad  ;
	output \DM_wd[7]_pad  ;
	output \DM_wd[8]_pad  ;
	output \DM_wd[9]_pad  ;
	output \DMo_cs0_pad  ;
	output \DMo_cs1_pad  ;
	output \DMo_cs2_pad  ;
	output \DMo_cs3_pad  ;
	output \DMo_cs4_pad  ;
	output \DMo_cs5_pad  ;
	output \DMo_cs6_pad  ;
	output \DMo_cs7_pad  ;
	output \DSPCLK_cm1_pad  ;
	output \EA_do[0]_pad  ;
	output \EA_do[10]_pad  ;
	output \EA_do[12]_pad  ;
	output \EA_do[13]_pad  ;
	output \EA_do[14]_pad  ;
	output \EA_do[1]_pad  ;
	output \EA_do[2]_pad  ;
	output \EA_do[3]_pad  ;
	output \EA_do[4]_pad  ;
	output \EA_do[5]_pad  ;
	output \EA_do[6]_pad  ;
	output \EA_do[7]_pad  ;
	output \EA_do[8]_pad  ;
	output \EA_do[9]_pad  ;
	output EA_oe_pad ;
	output \ED_do[0]_pad  ;
	output \ED_do[10]_pad  ;
	output \ED_do[11]_pad  ;
	output \ED_do[12]_pad  ;
	output \ED_do[13]_pad  ;
	output \ED_do[14]_pad  ;
	output \ED_do[15]_pad  ;
	output \ED_do[1]_pad  ;
	output \ED_do[2]_pad  ;
	output \ED_do[3]_pad  ;
	output \ED_do[4]_pad  ;
	output \ED_do[5]_pad  ;
	output \ED_do[6]_pad  ;
	output \ED_do[7]_pad  ;
	output \ED_do[8]_pad  ;
	output \ED_do[9]_pad  ;
	output \ED_oe_14_8_pad  ;
	output \ED_oe_7_0_pad  ;
	output \IAD_do[0]_pad  ;
	output \IAD_do[10]_pad  ;
	output \IAD_do[11]_pad  ;
	output \IAD_do[12]_pad  ;
	output \IAD_do[13]_pad  ;
	output \IAD_do[14]_pad  ;
	output \IAD_do[15]_pad  ;
	output \IAD_do[1]_pad  ;
	output \IAD_do[2]_pad  ;
	output \IAD_do[3]_pad  ;
	output \IAD_do[4]_pad  ;
	output \IAD_do[5]_pad  ;
	output \IAD_do[6]_pad  ;
	output \IAD_do[7]_pad  ;
	output \IAD_do[8]_pad  ;
	output \IAD_do[9]_pad  ;
	output IAD_oe_pad ;
	output IDoe_pad ;
	output IOSn_pad ;
	output \PMAinx[0]_pad  ;
	output \PMAinx[10]_pad  ;
	output \PMAinx[11]_pad  ;
	output \PMAinx[1]_pad  ;
	output \PMAinx[2]_pad  ;
	output \PMAinx[3]_pad  ;
	output \PMAinx[4]_pad  ;
	output \PMAinx[5]_pad  ;
	output \PMAinx[6]_pad  ;
	output \PMAinx[7]_pad  ;
	output \PMAinx[8]_pad  ;
	output \PMAinx[9]_pad  ;
	output \PM_wd[0]_pad  ;
	output \PM_wd[10]_pad  ;
	output \PM_wd[11]_pad  ;
	output \PM_wd[12]_pad  ;
	output \PM_wd[13]_pad  ;
	output \PM_wd[14]_pad  ;
	output \PM_wd[15]_pad  ;
	output \PM_wd[1]_pad  ;
	output \PM_wd[2]_pad  ;
	output \PM_wd[3]_pad  ;
	output \PM_wd[4]_pad  ;
	output \PM_wd[5]_pad  ;
	output \PM_wd[6]_pad  ;
	output \PM_wd[7]_pad  ;
	output \PM_wd[8]_pad  ;
	output \PM_wd[9]_pad  ;
	output \PMo_cs0_pad  ;
	output \PMo_cs1_pad  ;
	output \PMo_cs2_pad  ;
	output \PMo_cs3_pad  ;
	output \PMo_cs4_pad  ;
	output \PMo_cs5_pad  ;
	output \PMo_cs6_pad  ;
	output \PMo_cs7_pad  ;
	output \PMo_oe0_pad  ;
	output \RFS0_pad  ;
	output \RFS1_pad  ;
	output \SCLK0_pad  ;
	output \SCLK1_pad  ;
	output \TD0_pad  ;
	output \TD1_pad  ;
	output \TFS0_pad  ;
	output \TFS1_pad  ;
	output \T_ISn_syn_2  ;
	output WRn_pad ;
	output XTALoffn_pad ;
	output \_al_n0  ;
	output \bdma_BDMA_boot_reg/NET0131_reg_syn_3  ;
	output \bdma_BDMA_boot_reg/n0  ;
	output \bdma_BM_cyc_reg/P0000  ;
	output \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_3  ;
	output \core_c_psq_MGNT_reg/P0001  ;
	output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001_reg_syn_3  ;
	output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001_reg_syn_3  ;
	output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001_reg_syn_3  ;
	output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001_reg_syn_3  ;
	output \core_eu_ec_cun_MVi_pre_C_reg/P0001_reg_syn_3  ;
	output \core_eu_em_mac_em_reg_Sq_E_reg/P0001_reg_syn_3  ;
	output \emc_DMDreg_reg[8]/P0001_reg_syn_3  ;
	output \emc_DMDreg_reg[9]/P0001_reg_syn_3  ;
	output \emc_ECMcs_reg/P0001  ;
	output \emc_PMDreg_reg[8]/P0001_reg_syn_3  ;
	output \emc_PMDreg_reg[9]/P0001_reg_syn_3  ;
	output \g10/_0_  ;
	output \g1000/_0_  ;
	output \g10000/_0_  ;
	output \g10001/_0_  ;
	output \g10002/_0_  ;
	output \g10003/_0_  ;
	output \g10004/_0_  ;
	output \g10005/_0_  ;
	output \g10007/_0_  ;
	output \g10008/_0_  ;
	output \g10009/_0_  ;
	output \g1001/_3_  ;
	output \g10010/_0_  ;
	output \g10011/_0_  ;
	output \g10012/_0_  ;
	output \g10013/_0_  ;
	output \g10014/_0_  ;
	output \g10015/_0_  ;
	output \g10016/_0_  ;
	output \g10017/_0_  ;
	output \g10018/_0_  ;
	output \g10019/_0_  ;
	output \g1002/_3_  ;
	output \g10020/_0_  ;
	output \g10021/_0_  ;
	output \g10022/_0_  ;
	output \g10023/_0_  ;
	output \g10024/_0_  ;
	output \g10025/_0_  ;
	output \g10026/_0_  ;
	output \g10027/_0_  ;
	output \g10028/_0_  ;
	output \g10029/_0_  ;
	output \g1003/_0_  ;
	output \g10030/_0_  ;
	output \g10031/_0_  ;
	output \g10032/_0_  ;
	output \g10033/_0_  ;
	output \g10034/_0_  ;
	output \g10035/_0_  ;
	output \g10036/_0_  ;
	output \g10037/_0_  ;
	output \g10038/_0_  ;
	output \g10039/_0_  ;
	output \g10040/_0_  ;
	output \g10041/_0_  ;
	output \g10042/_0_  ;
	output \g10043/_0_  ;
	output \g10044/_0_  ;
	output \g10045/_0_  ;
	output \g10046/_0_  ;
	output \g10047/_0_  ;
	output \g10048/_0_  ;
	output \g10049/_0_  ;
	output \g10050/_0_  ;
	output \g10051/_0_  ;
	output \g10052/_0_  ;
	output \g10053/_0_  ;
	output \g10054/_0_  ;
	output \g10055/_0_  ;
	output \g10056/_0_  ;
	output \g10057/_0_  ;
	output \g10058/_0_  ;
	output \g10059/_0_  ;
	output \g10060/_0_  ;
	output \g10061/_0_  ;
	output \g10062/_0_  ;
	output \g10063/_0_  ;
	output \g10064/_0_  ;
	output \g10065/_0_  ;
	output \g10066/_0_  ;
	output \g10067/_0_  ;
	output \g10068/_0_  ;
	output \g10069/_0_  ;
	output \g10070/_0_  ;
	output \g10071/_0_  ;
	output \g10072/_0_  ;
	output \g10073/_0_  ;
	output \g10074/_0_  ;
	output \g10075/_0_  ;
	output \g10076/_0_  ;
	output \g10077/_0_  ;
	output \g10078/_0_  ;
	output \g10080/_0_  ;
	output \g10081/_0_  ;
	output \g10083/_0_  ;
	output \g10089/_0_  ;
	output \g1009/_0_  ;
	output \g10090/_0_  ;
	output \g10091/_0_  ;
	output \g10092/_0_  ;
	output \g10093/_0_  ;
	output \g10094/_0_  ;
	output \g1010/_0_  ;
	output \g10108/_3_  ;
	output \g1011/_0_  ;
	output \g10110/_0_  ;
	output \g10111/_0_  ;
	output \g10113/_3_  ;
	output \g10115/_3_  ;
	output \g1013/_0_  ;
	output \g1014/_0_  ;
	output \g10152/_0_  ;
	output \g10153/_0_  ;
	output \g10154/_0_  ;
	output \g10155/_0_  ;
	output \g10156/_0_  ;
	output \g10157/_0_  ;
	output \g10158/_0_  ;
	output \g10159/_0_  ;
	output \g1016/_0_  ;
	output \g10160/_0_  ;
	output \g10161/_0_  ;
	output \g10162/_0_  ;
	output \g10163/_0_  ;
	output \g10164/_0_  ;
	output \g10165/_0_  ;
	output \g1017/_0_  ;
	output \g10170/_3_  ;
	output \g1018/_0_  ;
	output \g10190/_3_  ;
	output \g10194/_3_  ;
	output \g10198/_0_  ;
	output \g10199/_0_  ;
	output \g102/_0_  ;
	output \g103/_0_  ;
	output \g104/_0_  ;
	output \g105/_0_  ;
	output \g10598/_0_  ;
	output \g106/_0_  ;
	output \g10667/_0_  ;
	output \g10683/_0_  ;
	output \g10685/_0_  ;
	output \g107/_0_  ;
	output \g10721/_0_  ;
	output \g10758/_0_  ;
	output \g10765/_0_  ;
	output \g10778/_0_  ;
	output \g10791/_0_  ;
	output \g108/_0_  ;
	output \g10887/_0_  ;
	output \g1089/_0_  ;
	output \g109/_0_  ;
	output \g1090/_0_  ;
	output \g1091/_0_  ;
	output \g1092/_0_  ;
	output \g10923/_0_  ;
	output \g1093/_0_  ;
	output \g10930/_0_  ;
	output \g10931/_0_  ;
	output \g10936/_0_  ;
	output \g1097/_0_  ;
	output \g11/_0_  ;
	output \g110/_0_  ;
	output \g1101/_0_  ;
	output \g11013/_0_  ;
	output \g1102/_0_  ;
	output \g1103/_0_  ;
	output \g11032/_0_  ;
	output \g1104/_0_  ;
	output \g1105/_0_  ;
	output \g1107/_0_  ;
	output \g11074/_0_  ;
	output \g11077/_0_  ;
	output \g1108/_0_  ;
	output \g1109/_0_  ;
	output \g11112/_0_  ;
	output \g11115/_0_  ;
	output \g11116/_0_  ;
	output \g11119/_0_  ;
	output \g11120/_0_  ;
	output \g1113/_0_  ;
	output \g1115/_0_  ;
	output \g1116/_0_  ;
	output \g1117/_0_  ;
	output \g11267/_0_  ;
	output \g11281/_0_  ;
	output \g11287/_0_  ;
	output \g11300/_0_  ;
	output \g11323/_0_  ;
	output \g11325/_2__syn_2  ;
	output \g11345/_2_  ;
	output \g11470/_0_  ;
	output \g11471/_0_  ;
	output \g11472/_0_  ;
	output \g11473/_0_  ;
	output \g11474/_0_  ;
	output \g11476/_0_  ;
	output \g11477/_0_  ;
	output \g11496/_0_  ;
	output \g11497/_0_  ;
	output \g11498/_0_  ;
	output \g11499/_0_  ;
	output \g11500/_0_  ;
	output \g11501/_0_  ;
	output \g11502/_0_  ;
	output \g11503/_0_  ;
	output \g11504/_0_  ;
	output \g11505/_0_  ;
	output \g11506/_0_  ;
	output \g11507/_0_  ;
	output \g11509/_0_  ;
	output \g11510/_0_  ;
	output \g11515/_0_  ;
	output \g11516/_0_  ;
	output \g11520/_0_  ;
	output \g11521/_0_  ;
	output \g11576/_0_  ;
	output \g11577/_0_  ;
	output \g11578/_0_  ;
	output \g11579/_0_  ;
	output \g11580/_0_  ;
	output \g11581/_0_  ;
	output \g11582/_0_  ;
	output \g11583/_0_  ;
	output \g11584/_0_  ;
	output \g11585/_0_  ;
	output \g11586/_0_  ;
	output \g11587/_0_  ;
	output \g11588/_0_  ;
	output \g11589/_0_  ;
	output \g11591/_0_  ;
	output \g11593/_0_  ;
	output \g11595/_0_  ;
	output \g11596/_0_  ;
	output \g11597/_0_  ;
	output \g11605/_0_  ;
	output \g11606/_0_  ;
	output \g11607/_0_  ;
	output \g11608/_0_  ;
	output \g11609/_0_  ;
	output \g11610/_0_  ;
	output \g11611/_0_  ;
	output \g11612/_0_  ;
	output \g11613/_0_  ;
	output \g11615/_0_  ;
	output \g11616/_0_  ;
	output \g11617/_0_  ;
	output \g11651/_3_  ;
	output \g11704/_0_  ;
	output \g11705/_0_  ;
	output \g11709/_0_  ;
	output \g11722/_0_  ;
	output \g11723/_0_  ;
	output \g119/_0_  ;
	output \g1192/_0_  ;
	output \g11994/_0_  ;
	output \g120/_0_  ;
	output \g1200/_0_  ;
	output \g12003/_0_  ;
	output \g1201/_0_  ;
	output \g12019/_0_  ;
	output \g1203/_3_  ;
	output \g1204/_3_  ;
	output \g1207/_0_  ;
	output \g1208/_0_  ;
	output \g12092/_0_  ;
	output \g1210/_0_  ;
	output \g1211/_0_  ;
	output \g1212/_0_  ;
	output \g1213/_0_  ;
	output \g12145/_0_  ;
	output \g12155/_0_  ;
	output \g12186/_0_  ;
	output \g12187/_0_  ;
	output \g12192/_0_  ;
	output \g12201/_0_  ;
	output \g12202/_0_  ;
	output \g12203/_0_  ;
	output \g12204/_0_  ;
	output \g12207/_0_  ;
	output \g12229/_3_  ;
	output \g12267/_0_  ;
	output \g12276/_0_  ;
	output \g12278/_0_  ;
	output \g12279/_0_  ;
	output \g12280/_0_  ;
	output \g12302/_0_  ;
	output \g12316/_0_  ;
	output \g12317/_0_  ;
	output \g12319/_0_  ;
	output \g12328/_3_  ;
	output \g1233/_0_  ;
	output \g12348/_0_  ;
	output \g12351/_0_  ;
	output \g12352/_0_  ;
	output \g12353/_0_  ;
	output \g12354/_0_  ;
	output \g12355/_0_  ;
	output \g1237/_0_  ;
	output \g124/_0_  ;
	output \g12444/_0_  ;
	output \g125/_0_  ;
	output \g12637/_0_  ;
	output \g12639/_0_  ;
	output \g12658/_0_  ;
	output \g12659/_0_  ;
	output \g12660/_0_  ;
	output \g12663/_0_  ;
	output \g12664/_0_  ;
	output \g12665/_0_  ;
	output \g12672/_3_  ;
	output \g12673/_3_  ;
	output \g12674/_3_  ;
	output \g12675/_3_  ;
	output \g12676/_3_  ;
	output \g12677/_3_  ;
	output \g12678/_0_  ;
	output \g12679/_3_  ;
	output \g12697/_3_  ;
	output \g12701/_3_  ;
	output \g12711/_2_  ;
	output \g12713/_2_  ;
	output \g12715/_2_  ;
	output \g12717/_2_  ;
	output \g12718/_2__syn_2  ;
	output \g1272/_0_  ;
	output \g12728/_1__syn_2  ;
	output \g12730/_3_  ;
	output \g12741/_1__syn_2  ;
	output \g12746/_0__syn_2  ;
	output \g12748/_0_  ;
	output \g12749/_0_  ;
	output \g12759/_1__syn_2  ;
	output \g12760/_0_  ;
	output \g12762/_0_  ;
	output \g12763/_0_  ;
	output \g12764/_0_  ;
	output \g12765/_0_  ;
	output \g12766/_0_  ;
	output \g12767/_0_  ;
	output \g12768/_0_  ;
	output \g12769/_0_  ;
	output \g12770/_0_  ;
	output \g12771/_0_  ;
	output \g12772/_0_  ;
	output \g12773/_0_  ;
	output \g12774/_0_  ;
	output \g12775/_0_  ;
	output \g12776/_0_  ;
	output \g12777/_0_  ;
	output \g12778/_0_  ;
	output \g12779/_0_  ;
	output \g1278/_0_  ;
	output \g12780/_0_  ;
	output \g12781/_0_  ;
	output \g12782/_0_  ;
	output \g12783/_0_  ;
	output \g12784/_0_  ;
	output \g12785/_0_  ;
	output \g12786/_0_  ;
	output \g12787/_0_  ;
	output \g12788/_0_  ;
	output \g12789/_0_  ;
	output \g12790/_0_  ;
	output \g12791/_0_  ;
	output \g12792/_0_  ;
	output \g12793/_0_  ;
	output \g12794/_0_  ;
	output \g12795/_0_  ;
	output \g12796/_0_  ;
	output \g12797/_0_  ;
	output \g12798/_0_  ;
	output \g12799/_0_  ;
	output \g12800/_0_  ;
	output \g12801/_0_  ;
	output \g12802/_0_  ;
	output \g12803/_0_  ;
	output \g12804/_0_  ;
	output \g12805/_0_  ;
	output \g12806/_0_  ;
	output \g12807/_0_  ;
	output \g12808/_0_  ;
	output \g12809/_0_  ;
	output \g1281/_0_  ;
	output \g12810/_0_  ;
	output \g12811/_0_  ;
	output \g12812/_0_  ;
	output \g12813/_0_  ;
	output \g12814/_0_  ;
	output \g12815/_0_  ;
	output \g12816/_0_  ;
	output \g12817/_0_  ;
	output \g12818/_0_  ;
	output \g12819/_0_  ;
	output \g1282/_0_  ;
	output \g12820/_0_  ;
	output \g12821/_0_  ;
	output \g12822/_0_  ;
	output \g12823/_0_  ;
	output \g12824/_0_  ;
	output \g12825/_0_  ;
	output \g12826/_0_  ;
	output \g12827/_0_  ;
	output \g12828/_0_  ;
	output \g12829/_0_  ;
	output \g12830/_0_  ;
	output \g12831/_0_  ;
	output \g12832/_0_  ;
	output \g12833/_0_  ;
	output \g12835/_0_  ;
	output \g12836/_0_  ;
	output \g12838/_0_  ;
	output \g12848/_0_  ;
	output \g12849/_0_  ;
	output \g1285/_0_  ;
	output \g12850/_0_  ;
	output \g12857/_0_  ;
	output \g12858/_0_  ;
	output \g12859/_0_  ;
	output \g12861/_0_  ;
	output \g12862/_0_  ;
	output \g12868/_0_  ;
	output \g12869/_0_  ;
	output \g1287/_0_  ;
	output \g12870/_0_  ;
	output \g12871/_0_  ;
	output \g12872/_0_  ;
	output \g12873/_0_  ;
	output \g12874/_0_  ;
	output \g12875/_0_  ;
	output \g12876/_0_  ;
	output \g12877/_0_  ;
	output \g12878/_0_  ;
	output \g12879/_0_  ;
	output \g12880/_0_  ;
	output \g12881/_0_  ;
	output \g12882/_0_  ;
	output \g12883/_0_  ;
	output \g12884/_0_  ;
	output \g12885/_0_  ;
	output \g12886/_0_  ;
	output \g12887/_0_  ;
	output \g12888/_0_  ;
	output \g12889/_0_  ;
	output \g1289/_0_  ;
	output \g12890/_0_  ;
	output \g12891/_0_  ;
	output \g12894/_0_  ;
	output \g12898/_0_  ;
	output \g12899/_0_  ;
	output \g12900/_0_  ;
	output \g12901/_0_  ;
	output \g12902/_0_  ;
	output \g12903/_0_  ;
	output \g12906/_0_  ;
	output \g12907/_0_  ;
	output \g12908/_0_  ;
	output \g12912/_0_  ;
	output \g12913/_0_  ;
	output \g12914/_0_  ;
	output \g12915/_0_  ;
	output \g12916/_0_  ;
	output \g12917/_0_  ;
	output \g12918/_0_  ;
	output \g12919/_0_  ;
	output \g12920/_0_  ;
	output \g12921/_0_  ;
	output \g12922/_0_  ;
	output \g12923/_0_  ;
	output \g12924/_0_  ;
	output \g12925/_0_  ;
	output \g12926/_0_  ;
	output \g12932/_0_  ;
	output \g12933/_0_  ;
	output \g12936/_0_  ;
	output \g12955/_0_  ;
	output \g13015/_0_  ;
	output \g13016/_0_  ;
	output \g13017/_0_  ;
	output \g13018/_0_  ;
	output \g13019/_0_  ;
	output \g13020/_0_  ;
	output \g13021/_0_  ;
	output \g13024/_0_  ;
	output \g13025/_0_  ;
	output \g13027/_0_  ;
	output \g13028/_0_  ;
	output \g13030/_0_  ;
	output \g13031/_0_  ;
	output \g13033/_0_  ;
	output \g13047/_0_  ;
	output \g13060/_0_  ;
	output \g13062/_0_  ;
	output \g13063/_0_  ;
	output \g13064/_0_  ;
	output \g13067/_0_  ;
	output \g13068/_0_  ;
	output \g13069/_0_  ;
	output \g13070/_0_  ;
	output \g13072/_0_  ;
	output \g13094/_0_  ;
	output \g13104/_0_  ;
	output \g13110/_0_  ;
	output \g13114/_0_  ;
	output \g13115/_0_  ;
	output \g13116/_0_  ;
	output \g13117/_0_  ;
	output \g13118/_0_  ;
	output \g13119/_0_  ;
	output \g13120/_0_  ;
	output \g13121/_0_  ;
	output \g13124/_0_  ;
	output \g13125/_0_  ;
	output \g13127/_0_  ;
	output \g13128/_0_  ;
	output \g13129/_0_  ;
	output \g13130/_0_  ;
	output \g13131/_0_  ;
	output \g13132/_0_  ;
	output \g13133/_0_  ;
	output \g13134/_0_  ;
	output \g13138/_0_  ;
	output \g13139/_0_  ;
	output \g13140/_0_  ;
	output \g13141/_0_  ;
	output \g13142/_0_  ;
	output \g13143/_0_  ;
	output \g13144/_0_  ;
	output \g13146/_0_  ;
	output \g13150/_0_  ;
	output \g13152/_0_  ;
	output \g13154/_0_  ;
	output \g13155/_0_  ;
	output \g13156/_0_  ;
	output \g13157/_0_  ;
	output \g13158/_0_  ;
	output \g1320/_3_  ;
	output \g13266/_0_  ;
	output \g13269/_0_  ;
	output \g13274/_0_  ;
	output \g13277/_0_  ;
	output \g13280/_0_  ;
	output \g13283/_0_  ;
	output \g13294/_0_  ;
	output \g13330/_0_  ;
	output \g13333/_0_  ;
	output \g13334/_0_  ;
	output \g13335/_0_  ;
	output \g13336/_0_  ;
	output \g13337/_0_  ;
	output \g13338/_0_  ;
	output \g13345/_0_  ;
	output \g13346/_0_  ;
	output \g13347/_0_  ;
	output \g13348/_0_  ;
	output \g13349/_0_  ;
	output \g13350/_0_  ;
	output \g13351/_0_  ;
	output \g13352/_0_  ;
	output \g13486/_0_  ;
	output \g13488/_0_  ;
	output \g13508/_0_  ;
	output \g13509/_0_  ;
	output \g13510/_0_  ;
	output \g13511/_0_  ;
	output \g13512/_0_  ;
	output \g13513/_0_  ;
	output \g13514/_0_  ;
	output \g13515/_0_  ;
	output \g13516/_0_  ;
	output \g13517/_0_  ;
	output \g13518/_0_  ;
	output \g13519/_0_  ;
	output \g13520/_0_  ;
	output \g13521/_0_  ;
	output \g13540/_0_  ;
	output \g13541/_0_  ;
	output \g13542/_0_  ;
	output \g13543/_0_  ;
	output \g13544/_0_  ;
	output \g13545/_0_  ;
	output \g13546/_0_  ;
	output \g13547/_0_  ;
	output \g13548/_0_  ;
	output \g13549/_0_  ;
	output \g13550/_0_  ;
	output \g13551/_0_  ;
	output \g13552/_0_  ;
	output \g13553/_0_  ;
	output \g13554/_0_  ;
	output \g13555/_0_  ;
	output \g13556/_0_  ;
	output \g13557/_0_  ;
	output \g13558/_0_  ;
	output \g13559/_0_  ;
	output \g13560/_0_  ;
	output \g13561/_0_  ;
	output \g13562/_0_  ;
	output \g13563/_0_  ;
	output \g13564/_0_  ;
	output \g13565/_0_  ;
	output \g13566/_0_  ;
	output \g13567/_0_  ;
	output \g13568/_0_  ;
	output \g13569/_0_  ;
	output \g13570/_0_  ;
	output \g13571/_0_  ;
	output \g13572/_0_  ;
	output \g137/_3_  ;
	output \g1387/_3_  ;
	output \g1388/_3_  ;
	output \g1389/_0_  ;
	output \g139/_0_  ;
	output \g1390/_0_  ;
	output \g1393/_0_  ;
	output \g140/_0_  ;
	output \g141/_0_  ;
	output \g14173/_0_  ;
	output \g14176/_0_  ;
	output \g142/_3_  ;
	output \g14273/_1__syn_2  ;
	output \g14274/_0_  ;
	output \g14280/_0_  ;
	output \g14281/_0_  ;
	output \g143/_3_  ;
	output \g14354/_3__syn_2  ;
	output \g14370/_0_  ;
	output \g14385/_0_  ;
	output \g14386/_0_  ;
	output \g144/_3_  ;
	output \g14407/_0_  ;
	output \g14412/_0_  ;
	output \g14435/_0_  ;
	output \g14439/_0_  ;
	output \g145/_0_  ;
	output \g14522/_0_  ;
	output \g14528/_0_  ;
	output \g14533/_0_  ;
	output \g14581/_1_  ;
	output \g14582/_0_  ;
	output \g146/_3_  ;
	output \g14671/_0_  ;
	output \g14672/_0_  ;
	output \g147/_0_  ;
	output \g1473/_0_  ;
	output \g148/_0_  ;
	output \g14826/_0_  ;
	output \g149/_0_  ;
	output \g14908/_0_  ;
	output \g14911/_0_  ;
	output \g14936/_2_  ;
	output \g1494/_0_  ;
	output \g1495/_0_  ;
	output \g14950/_2_  ;
	output \g14953/_2_  ;
	output \g15003/_0_  ;
	output \g15004/_0_  ;
	output \g15006/_0_  ;
	output \g15007/_0_  ;
	output \g15008/_0_  ;
	output \g15009/_0_  ;
	output \g15010/_0_  ;
	output \g15011/_0_  ;
	output \g15012/_0_  ;
	output \g15013/_0_  ;
	output \g15014/_0_  ;
	output \g15015/_0_  ;
	output \g15016/_0_  ;
	output \g15017/_0_  ;
	output \g15018/_0_  ;
	output \g15019/_0_  ;
	output \g15035/_0_  ;
	output \g15036/_0_  ;
	output \g15038/_0_  ;
	output \g15039/_0_  ;
	output \g15040/_0_  ;
	output \g15041/_0_  ;
	output \g15042/_0_  ;
	output \g15043/_0_  ;
	output \g15044/_0_  ;
	output \g15045/_0_  ;
	output \g15046/_0_  ;
	output \g15056/_00_  ;
	output \g151/_0_  ;
	output \g15193/_0_  ;
	output \g152/_0_  ;
	output \g15256/_0_  ;
	output \g153/_0_  ;
	output \g15393/_0_  ;
	output \g15394/_0_  ;
	output \g15395/_0_  ;
	output \g15396/_0_  ;
	output \g15397/_0_  ;
	output \g15398/_0_  ;
	output \g15399/_0_  ;
	output \g154/_0_  ;
	output \g15400/_0_  ;
	output \g15401/_0_  ;
	output \g15402/_0_  ;
	output \g15403/_0_  ;
	output \g15404/_0_  ;
	output \g15405/_0_  ;
	output \g15406/_0_  ;
	output \g15407/_0_  ;
	output \g15408/_0_  ;
	output \g15473/_0_  ;
	output \g15650/_0_  ;
	output \g15651/_0_  ;
	output \g15652/_0_  ;
	output \g15653/_0_  ;
	output \g15662/_0_  ;
	output \g15663/_0_  ;
	output \g15664/_0_  ;
	output \g15665/_0_  ;
	output \g15666/_0_  ;
	output \g15667/_0_  ;
	output \g15668/_0_  ;
	output \g15669/_0_  ;
	output \g15670/_0_  ;
	output \g15671/_0_  ;
	output \g15672/_0_  ;
	output \g15673/_0_  ;
	output \g15674/_0_  ;
	output \g15675/_0_  ;
	output \g1569/_0_  ;
	output \g1570/_0_  ;
	output \g1575/_0_  ;
	output \g1576/_0_  ;
	output \g15922/_1_  ;
	output \g15970/_0_  ;
	output \g16059/_0_  ;
	output \g1606/_3_  ;
	output \g16124/_0_  ;
	output \g16144/_0_  ;
	output \g16202/_0_  ;
	output \g16214/_0_  ;
	output \g16247/_0_  ;
	output \g16257/_0_  ;
	output \g16274/_1_  ;
	output \g16324/_0_  ;
	output \g16343/_1__syn_2  ;
	output \g16381/_0_  ;
	output \g16383/_0_  ;
	output \g16386/_0_  ;
	output \g16414/_1__syn_2  ;
	output \g16416/_0__syn_2  ;
	output \g16448/_0_  ;
	output \g16460/_1_  ;
	output \g16625/_3_  ;
	output \g16662/_0_  ;
	output \g16668/_1__syn_2  ;
	output \g16692/_0_  ;
	output \g16721/_0_  ;
	output \g16723/_0_  ;
	output \g16725/_0_  ;
	output \g16726/_0_  ;
	output \g16727/_0_  ;
	output \g16728/_0_  ;
	output \g16729/_0_  ;
	output \g16730/_0_  ;
	output \g16731/_0_  ;
	output \g16732/_0_  ;
	output \g16733/_0_  ;
	output \g16734/_0_  ;
	output \g16735/_0_  ;
	output \g16736/_0_  ;
	output \g16737/_0_  ;
	output \g16738/_0_  ;
	output \g16739/_0_  ;
	output \g16740/_0_  ;
	output \g16741/_0_  ;
	output \g16742/_0_  ;
	output \g16743/_0_  ;
	output \g16747/_0_  ;
	output \g16748/_0_  ;
	output \g16749/_0_  ;
	output \g16750/_0_  ;
	output \g16753/_0_  ;
	output \g16754/_0_  ;
	output \g16755/_0_  ;
	output \g16756/_0_  ;
	output \g16757/_0_  ;
	output \g16758/_0_  ;
	output \g16761/_0_  ;
	output \g16765/_0_  ;
	output \g16766/_0_  ;
	output \g16767/_0_  ;
	output \g16768/_0_  ;
	output \g16769/_0_  ;
	output \g16772/_0_  ;
	output \g16785/_0_  ;
	output \g16786/_0_  ;
	output \g16787/_0_  ;
	output \g16788/_0_  ;
	output \g16789/_0_  ;
	output \g16790/_0_  ;
	output \g16791/_0_  ;
	output \g16804/_0_  ;
	output \g16805/_0_  ;
	output \g16806/_0_  ;
	output \g16807/_0_  ;
	output \g16808/_0_  ;
	output \g16809/_0_  ;
	output \g16810/_0_  ;
	output \g16811/_0_  ;
	output \g16812/_0_  ;
	output \g16813/_0_  ;
	output \g16814/_0_  ;
	output \g16815/_0_  ;
	output \g16816/_0_  ;
	output \g16817/_0_  ;
	output \g16819/_0_  ;
	output \g16822/_0_  ;
	output \g16823/_0_  ;
	output \g16824/_0_  ;
	output \g16825/_0_  ;
	output \g16828/_0_  ;
	output \g16829/_0_  ;
	output \g16830/_0_  ;
	output \g16831/_0_  ;
	output \g16832/_0_  ;
	output \g16833/_0_  ;
	output \g16834/_0_  ;
	output \g16835/_0_  ;
	output \g16836/_0_  ;
	output \g16837/_0_  ;
	output \g16840/_0_  ;
	output \g16841/_0_  ;
	output \g16842/_0_  ;
	output \g16843/_0_  ;
	output \g16846/_0_  ;
	output \g16847/_0_  ;
	output \g16848/_0_  ;
	output \g16849/_0_  ;
	output \g16850/_0_  ;
	output \g16851/_0_  ;
	output \g16852/_0_  ;
	output \g16853/_0_  ;
	output \g16854/_0_  ;
	output \g16855/_0_  ;
	output \g16856/_0_  ;
	output \g16857/_0_  ;
	output \g16859/_0_  ;
	output \g16862/_0_  ;
	output \g16865/_0_  ;
	output \g16866/_0_  ;
	output \g16867/_0_  ;
	output \g16868/_0_  ;
	output \g16869/_0_  ;
	output \g16870/_0_  ;
	output \g16871/_0_  ;
	output \g16872/_0_  ;
	output \g16873/_0_  ;
	output \g16874/_0_  ;
	output \g16875/_0_  ;
	output \g16876/_0_  ;
	output \g16877/_0_  ;
	output \g16878/_0_  ;
	output \g16879/_0_  ;
	output \g16880/_0_  ;
	output \g16881/_0_  ;
	output \g16882/_0_  ;
	output \g16884/_0_  ;
	output \g16887/_0_  ;
	output \g16891/_0_  ;
	output \g16892/_0_  ;
	output \g16893/_0_  ;
	output \g16894/_0_  ;
	output \g16895/_0_  ;
	output \g16897/_0_  ;
	output \g16898/_0_  ;
	output \g16899/_0_  ;
	output \g16900/_0_  ;
	output \g16901/_0_  ;
	output \g16902/_0_  ;
	output \g16903/_0_  ;
	output \g16904/_0_  ;
	output \g16905/_0_  ;
	output \g16906/_0_  ;
	output \g16907/_0_  ;
	output \g16908/_0_  ;
	output \g16909/_0_  ;
	output \g16910/_0_  ;
	output \g16912/_0_  ;
	output \g16914/_0_  ;
	output \g16915/_0_  ;
	output \g16950/_0_  ;
	output \g16951/_0_  ;
	output \g16952/_0_  ;
	output \g16953/_0_  ;
	output \g16954/_0_  ;
	output \g16955/_0_  ;
	output \g16956/_0_  ;
	output \g16957/_0_  ;
	output \g16958/_0_  ;
	output \g16959/_0_  ;
	output \g16960/_0_  ;
	output \g16961/_0_  ;
	output \g16962/_0_  ;
	output \g16963/_0_  ;
	output \g16964/_0_  ;
	output \g16965/_0_  ;
	output \g16966/_0_  ;
	output \g16967/_0_  ;
	output \g16968/_0_  ;
	output \g16970/_0_  ;
	output \g17102/_3_  ;
	output \g17106/_0_  ;
	output \g17107/_0_  ;
	output \g17109/_0_  ;
	output \g17110/_0_  ;
	output \g17111/_0_  ;
	output \g17112/_0_  ;
	output \g17115/_0_  ;
	output \g17116/_0_  ;
	output \g17119/_0_  ;
	output \g17120/_0_  ;
	output \g17122/_0_  ;
	output \g17123/_0_  ;
	output \g17124/_0_  ;
	output \g17125/_0_  ;
	output \g17126/_0_  ;
	output \g17127/_0_  ;
	output \g17128/_0_  ;
	output \g17130/_0_  ;
	output \g17131/_0_  ;
	output \g17132/_0_  ;
	output \g17133/_0_  ;
	output \g17134/_0_  ;
	output \g17135/_0_  ;
	output \g17136/_0_  ;
	output \g17137/_0_  ;
	output \g17138/_0_  ;
	output \g17140/_0_  ;
	output \g17141/_0_  ;
	output \g17142/_0_  ;
	output \g17143/_0_  ;
	output \g17144/_0_  ;
	output \g17145/_0_  ;
	output \g17146/_0_  ;
	output \g17147/_0_  ;
	output \g17148/_0_  ;
	output \g17149/_0_  ;
	output \g17150/_0_  ;
	output \g17151/_0_  ;
	output \g17152/_0_  ;
	output \g17153/_0_  ;
	output \g17154/_0_  ;
	output \g17155/_0_  ;
	output \g17157/_0_  ;
	output \g17159/_0_  ;
	output \g17160/_0_  ;
	output \g17161/_0_  ;
	output \g17162/_0_  ;
	output \g17163/_0_  ;
	output \g17164/_0_  ;
	output \g17165/_0_  ;
	output \g17166/_0_  ;
	output \g17168/_0_  ;
	output \g17171/_0_  ;
	output \g17173/_0_  ;
	output \g17177/_0_  ;
	output \g17178/_0_  ;
	output \g17179/_0_  ;
	output \g17180/_0_  ;
	output \g17182/_0_  ;
	output \g17183/_0_  ;
	output \g17184/_0_  ;
	output \g17185/_0_  ;
	output \g17186/_0_  ;
	output \g17188/_0_  ;
	output \g17189/_0_  ;
	output \g17190/_0_  ;
	output \g17191/_0_  ;
	output \g17193/_0_  ;
	output \g17194/_0_  ;
	output \g17195/_0_  ;
	output \g17196/_0_  ;
	output \g17197/_0_  ;
	output \g17198/_0_  ;
	output \g17199/_0_  ;
	output \g17200/_0_  ;
	output \g17201/_0_  ;
	output \g17202/_0_  ;
	output \g17203/_0_  ;
	output \g17204/_0_  ;
	output \g17205/_0_  ;
	output \g17206/_0_  ;
	output \g17207/_0_  ;
	output \g17208/_0_  ;
	output \g17209/_0_  ;
	output \g17210/_0_  ;
	output \g17211/_0_  ;
	output \g17212/_0_  ;
	output \g17213/_0_  ;
	output \g17214/_0_  ;
	output \g17215/_0_  ;
	output \g17216/_0_  ;
	output \g17217/_0_  ;
	output \g17218/_0_  ;
	output \g17219/_0_  ;
	output \g17223/_0_  ;
	output \g17224/_0_  ;
	output \g17225/_0_  ;
	output \g17226/_0_  ;
	output \g17227/_0_  ;
	output \g17228/_0_  ;
	output \g17229/_0_  ;
	output \g17231/_0_  ;
	output \g17232/_0_  ;
	output \g17233/_0_  ;
	output \g17234/_0_  ;
	output \g17237/_0_  ;
	output \g17239/_0_  ;
	output \g17240/_0_  ;
	output \g17243/_0_  ;
	output \g17246/_0_  ;
	output \g17247/_0_  ;
	output \g17248/_0_  ;
	output \g17249/_0_  ;
	output \g17250/_0_  ;
	output \g17251/_0_  ;
	output \g17252/_0_  ;
	output \g17253/_0_  ;
	output \g17254/_0_  ;
	output \g17258/_0_  ;
	output \g17261/_0_  ;
	output \g17262/_0_  ;
	output \g17269/_0_  ;
	output \g17271/_0_  ;
	output \g17274/_0_  ;
	output \g17275/_0_  ;
	output \g17276/_0_  ;
	output \g17277/_0_  ;
	output \g17278/_0_  ;
	output \g17279/_0_  ;
	output \g17280/_0_  ;
	output \g17281/_0_  ;
	output \g17282/_0_  ;
	output \g17283/_0_  ;
	output \g17285/_0_  ;
	output \g17290/_0_  ;
	output \g17292/_0_  ;
	output \g17293/_0_  ;
	output \g17296/_0_  ;
	output \g17297/_0_  ;
	output \g17298/_0_  ;
	output \g173/_0_  ;
	output \g17303/_0_  ;
	output \g17304/_0_  ;
	output \g17305/_0_  ;
	output \g17306/_0_  ;
	output \g17307/_0_  ;
	output \g17308/_0_  ;
	output \g17309/_0_  ;
	output \g17310/_0_  ;
	output \g17311/_0_  ;
	output \g17312/_0_  ;
	output \g17314/_0_  ;
	output \g17315/_0_  ;
	output \g17316/_0_  ;
	output \g17317/_0_  ;
	output \g17318/_0_  ;
	output \g17319/_0_  ;
	output \g17320/_0_  ;
	output \g17321/_0_  ;
	output \g17322/_0_  ;
	output \g17323/_0_  ;
	output \g17324/_0_  ;
	output \g17325/_0_  ;
	output \g17326/_0_  ;
	output \g17327/_0_  ;
	output \g17328/_0_  ;
	output \g17329/_0_  ;
	output \g17330/_0_  ;
	output \g17331/_0_  ;
	output \g17332/_0_  ;
	output \g17333/_0_  ;
	output \g17335/_0_  ;
	output \g17336/_0_  ;
	output \g17337/_0_  ;
	output \g17338/_0_  ;
	output \g17339/_0_  ;
	output \g17340/_0_  ;
	output \g17342/_0_  ;
	output \g17343/_0_  ;
	output \g17347/_0_  ;
	output \g17350/_0_  ;
	output \g17354/_0_  ;
	output \g17356/_0_  ;
	output \g17357/_0_  ;
	output \g17358/_0_  ;
	output \g17359/_0_  ;
	output \g17360/_0_  ;
	output \g17415/_0_  ;
	output \g17441/_0_  ;
	output \g17442/_0_  ;
	output \g17451/_0_  ;
	output \g17457/_0_  ;
	output \g17458/_0_  ;
	output \g17459/_0_  ;
	output \g17460/_0_  ;
	output \g17461/_0_  ;
	output \g17462/_0_  ;
	output \g17463/_0_  ;
	output \g17464/_0_  ;
	output \g17465/_0_  ;
	output \g17466/_0_  ;
	output \g17467/_0_  ;
	output \g17468/_0_  ;
	output \g17469/_0_  ;
	output \g17470/_0_  ;
	output \g17471/_0_  ;
	output \g17472/_0_  ;
	output \g175/_3_  ;
	output \g1750/_0_  ;
	output \g176/_3_  ;
	output \g17619/_0_  ;
	output \g17620/_0_  ;
	output \g1763/_3_  ;
	output \g1764/_3_  ;
	output \g1768/_0_  ;
	output \g1769/_0_  ;
	output \g177/_3_  ;
	output \g17737/_0_  ;
	output \g17747/_0_  ;
	output \g178/_3_  ;
	output \g17814/_1_  ;
	output \g17815/_0_  ;
	output \g17821/_1_  ;
	output \g17821/_1__syn_2  ;
	output \g17872/_0_  ;
	output \g179/_3_  ;
	output \g17902/_0_  ;
	output \g180/_3_  ;
	output \g18020/_1_  ;
	output \g18057/_0_  ;
	output \g18096/_0_  ;
	output \g18099/_0_  ;
	output \g18107/_0_  ;
	output \g18133/_0_  ;
	output \g18140/_1_  ;
	output \g18153/_0_  ;
	output \g182/_0_  ;
	output \g18218/_0_  ;
	output \g18244/_0_  ;
	output \g18262/_0_  ;
	output \g18267/_0_  ;
	output \g18387/_1__syn_2  ;
	output \g184/_0_  ;
	output \g18478/_1_  ;
	output \g18585/_3_  ;
	output \g18608/_0_  ;
	output \g18609/_0_  ;
	output \g18613/_0_  ;
	output \g18618/_0_  ;
	output \g18647/_0_  ;
	output \g18687/_2_  ;
	output \g18707/_0_  ;
	output \g18748/_0_  ;
	output \g18753/_0_  ;
	output \g18758/_0_  ;
	output \g18759/_0_  ;
	output \g18760/_0_  ;
	output \g18761/_0_  ;
	output \g18762/_0_  ;
	output \g18763/_0_  ;
	output \g18764/_0_  ;
	output \g18765/_0_  ;
	output \g18766/_0_  ;
	output \g18767/_0_  ;
	output \g18768/_0_  ;
	output \g18770/_0_  ;
	output \g18771/_0_  ;
	output \g18788/_0_  ;
	output \g18796/_0_  ;
	output \g18800/_0_  ;
	output \g18801/_0_  ;
	output \g18802/_0_  ;
	output \g18803/_0_  ;
	output \g18804/_0_  ;
	output \g18805/_0_  ;
	output \g18807/_0_  ;
	output \g18840/_0_  ;
	output \g18843/_0_  ;
	output \g18844/_0_  ;
	output \g18846/_0_  ;
	output \g18847/_0_  ;
	output \g18848/_0_  ;
	output \g18849/_0_  ;
	output \g18850/_0_  ;
	output \g18851/_0_  ;
	output \g18852/_0_  ;
	output \g18853/_0_  ;
	output \g18854/_0_  ;
	output \g18855/_0_  ;
	output \g18856/_0_  ;
	output \g18858/_0_  ;
	output \g18860/_0_  ;
	output \g18861/_0_  ;
	output \g18863/_0_  ;
	output \g18864/_0_  ;
	output \g18866/_0_  ;
	output \g18867/_0_  ;
	output \g18868/_0_  ;
	output \g18869/_0_  ;
	output \g18870/_0_  ;
	output \g18871/_0_  ;
	output \g18872/_0_  ;
	output \g18873/_0_  ;
	output \g18874/_0_  ;
	output \g18875/_0_  ;
	output \g18876/_0_  ;
	output \g18877/_0_  ;
	output \g18878/_0_  ;
	output \g18879/_0_  ;
	output \g18880/_0_  ;
	output \g18881/_0_  ;
	output \g18882/_0_  ;
	output \g18883/_0_  ;
	output \g18888/_0_  ;
	output \g18892/_0_  ;
	output \g18895/_0_  ;
	output \g18896/_0_  ;
	output \g18897/_0_  ;
	output \g18905/_0_  ;
	output \g18908/_0_  ;
	output \g18909/_0_  ;
	output \g18912/_0_  ;
	output \g18918/_0_  ;
	output \g18919/_0_  ;
	output \g18920/_0_  ;
	output \g18921/_0_  ;
	output \g18922/_0_  ;
	output \g18924/_0_  ;
	output \g18925/_0_  ;
	output \g18927/_0_  ;
	output \g18930/_0_  ;
	output \g18966/_0_  ;
	output \g18968/_0_  ;
	output \g18970/_0_  ;
	output \g18974/_0_  ;
	output \g18975/_0_  ;
	output \g18977/_0_  ;
	output \g18981/_0_  ;
	output \g18983/_0_  ;
	output \g18985/_0_  ;
	output \g18987/_0_  ;
	output \g18989/_0_  ;
	output \g18991/_0_  ;
	output \g18992/_0_  ;
	output \g18993/_0_  ;
	output \g18994/_0_  ;
	output \g18995/_0_  ;
	output \g18996/_0_  ;
	output \g18997/_0_  ;
	output \g18998/_0_  ;
	output \g18999/_0_  ;
	output \g19001/_0_  ;
	output \g19003/_0_  ;
	output \g19005/_0_  ;
	output \g19006/_0_  ;
	output \g19014/_0_  ;
	output \g19016/_0_  ;
	output \g19018/_0_  ;
	output \g19020/_0_  ;
	output \g19022/_0_  ;
	output \g19056/_3_  ;
	output \g19058/_3_  ;
	output \g19060/_3_  ;
	output \g19062/_3_  ;
	output \g1910/_0_  ;
	output \g19186/_0_  ;
	output \g19188/_0_  ;
	output \g19235/_0_  ;
	output \g19239/_0_  ;
	output \g19244/_0_  ;
	output \g19253/_0_  ;
	output \g19254/_0_  ;
	output \g19259/_0_  ;
	output \g19261/_0_  ;
	output \g19267/_0_  ;
	output \g19277/_0_  ;
	output \g19278/_0_  ;
	output \g19280/_0_  ;
	output \g19281/_0_  ;
	output \g19282/_0_  ;
	output \g19283/_0_  ;
	output \g19284/_0_  ;
	output \g19285/_0_  ;
	output \g19286/_0_  ;
	output \g19287/_0_  ;
	output \g19288/_0_  ;
	output \g19289/_0_  ;
	output \g19290/_0_  ;
	output \g19291/_0_  ;
	output \g19292/_0_  ;
	output \g19293/_0_  ;
	output \g19294/_0_  ;
	output \g19295/_0_  ;
	output \g19296/_0_  ;
	output \g19297/_0_  ;
	output \g19298/_0_  ;
	output \g19299/_0_  ;
	output \g19300/_0_  ;
	output \g19301/_0_  ;
	output \g19302/_0_  ;
	output \g19303/_0_  ;
	output \g19304/_0_  ;
	output \g19305/_0_  ;
	output \g19306/_0_  ;
	output \g19307/_0_  ;
	output \g19308/_0_  ;
	output \g19315/_0_  ;
	output \g19316/_0_  ;
	output \g19317/_0_  ;
	output \g19318/_0_  ;
	output \g19319/_0_  ;
	output \g19320/_0_  ;
	output \g19321/_0_  ;
	output \g19322/_0_  ;
	output \g19323/_0_  ;
	output \g19325/_3_  ;
	output \g19326/_3_  ;
	output \g19333/_3_  ;
	output \g19341/_3_  ;
	output \g19347/_3_  ;
	output \g19377/_3_  ;
	output \g19381/_3_  ;
	output \g19393/_0_  ;
	output \g19401/_0_  ;
	output \g19402/_0_  ;
	output \g195/_2_  ;
	output \g19513/_0_  ;
	output \g19514/_0_  ;
	output \g19515/_0_  ;
	output \g19516/_0_  ;
	output \g1952/_3_  ;
	output \g19529/_0_  ;
	output \g19530/_0_  ;
	output \g19531/_0_  ;
	output \g19532/_0_  ;
	output \g19533/_0_  ;
	output \g19534/_0_  ;
	output \g19535/_0_  ;
	output \g19536/_0_  ;
	output \g19537/_0_  ;
	output \g19539/_0_  ;
	output \g19546/_0_  ;
	output \g19552/_0_  ;
	output \g19553/_0_  ;
	output \g19562/_0_  ;
	output \g19563/_0_  ;
	output \g19564/_0_  ;
	output \g19572/_0_  ;
	output \g19575/_0_  ;
	output \g19615/_0_  ;
	output \g19686/_0_  ;
	output \g19688/_0_  ;
	output \g197/_0_  ;
	output \g19729/_0_  ;
	output \g19774/_0_  ;
	output \g19777/_0_  ;
	output \g19791/_0_  ;
	output \g19818/_0_  ;
	output \g19819/_0_  ;
	output \g19828/_0_  ;
	output \g19852/_1_  ;
	output \g19860/_0_  ;
	output \g19861/_0_  ;
	output \g19864/_0_  ;
	output \g19886/_0_  ;
	output \g19887/_0_  ;
	output \g199/_0_  ;
	output \g19908/_0_  ;
	output \g19918/_0_  ;
	output \g19927/_0_  ;
	output \g19933/_0_  ;
	output \g200/_0_  ;
	output \g20019/_0_  ;
	output \g20046/_0_  ;
	output \g20068/_1_  ;
	output \g20080/_1_  ;
	output \g201/_0_  ;
	output \g20137/_0_  ;
	output \g20139/_0_  ;
	output \g20141/_0_  ;
	output \g20152/_1_  ;
	output \g20154/_00_  ;
	output \g202/_0_  ;
	output \g20206/_0_  ;
	output \g20211/_2_  ;
	output \g20217/_2_  ;
	output \g20239/_0_  ;
	output \g20265/_2_  ;
	output \g20266/_0_  ;
	output \g20272/_2_  ;
	output \g20278/_2_  ;
	output \g20283/_0_  ;
	output \g20285/_2_  ;
	output \g20288/_2__syn_2  ;
	output \g20293/_0_  ;
	output \g20295/_2_  ;
	output \g203/_0_  ;
	output \g20302/_2_  ;
	output \g20303/_2_  ;
	output \g20304/_2_  ;
	output \g20311/_2_  ;
	output \g20326/_0_  ;
	output \g20330/_0_  ;
	output \g2034/_0_  ;
	output \g20345/_0_  ;
	output \g20346/_0_  ;
	output \g2035/_0_  ;
	output \g20363/_0_  ;
	output \g20364/_0_  ;
	output \g204/_0_  ;
	output \g2047/_0_  ;
	output \g20483/_0_  ;
	output \g20493/_00_  ;
	output \g205/_0_  ;
	output \g20569/_0_  ;
	output \g20570/_0_  ;
	output \g20571/_0_  ;
	output \g206/_0_  ;
	output \g20613/_0_  ;
	output \g20615/_0_  ;
	output \g20657/_1__syn_2  ;
	output \g20660/_0_  ;
	output \g20685/_0_  ;
	output \g207/_0_  ;
	output \g20713/_1_  ;
	output \g20747/_1_  ;
	output \g20784/_0_  ;
	output \g20820/_1_  ;
	output \g20859/_0_  ;
	output \g20873/_2_  ;
	output \g20886/_0_  ;
	output \g20887/_0_  ;
	output \g20891/_2__syn_2  ;
	output \g20907/_2_  ;
	output \g20936/_2__syn_2  ;
	output \g20937/_1_  ;
	output \g20955/_0_  ;
	output \g20959/_2__syn_2  ;
	output \g20967/_0_  ;
	output \g20971/_2__syn_2  ;
	output \g20974/_1__syn_2  ;
	output \g21015/_1_  ;
	output \g21051/_2_  ;
	output \g21079/_1_  ;
	output \g21081/_1_  ;
	output \g21087/_2__syn_2  ;
	output \g21114/_1_  ;
	output \g21116/_1_  ;
	output \g21120/_2__syn_2  ;
	output \g21147/_0_  ;
	output \g21179/_1_  ;
	output \g21185/_1_  ;
	output \g21223/_0_  ;
	output \g21242/_0_  ;
	output \g21253/_0_  ;
	output \g21257/_0_  ;
	output \g21323/_1_  ;
	output \g21324/_1_  ;
	output \g21366/_0_  ;
	output \g21385/_2_  ;
	output \g21464/_0_  ;
	output \g21475/_3_  ;
	output \g21481/_0_  ;
	output \g21482/_0_  ;
	output \g21494/_3_  ;
	output \g21500/_3_  ;
	output \g21507/_3_  ;
	output \g21511/_3_  ;
	output \g21537/_1_  ;
	output \g21568/_0_  ;
	output \g21591/_0_  ;
	output \g21604/_0_  ;
	output \g21605/_3_  ;
	output \g21606/_0_  ;
	output \g21607/_0_  ;
	output \g21608/_0_  ;
	output \g21609/_0_  ;
	output \g21610/_0_  ;
	output \g21611/_0_  ;
	output \g21612/_0_  ;
	output \g21613/_0_  ;
	output \g21614/_0_  ;
	output \g21615/_0_  ;
	output \g21616/_0_  ;
	output \g21617/_0_  ;
	output \g21618/_0_  ;
	output \g21621/_0_  ;
	output \g21640/_0_  ;
	output \g21678/_0_  ;
	output \g21679/_0_  ;
	output \g21686/_0_  ;
	output \g21692/_3_  ;
	output \g21696/_0_  ;
	output \g21698/_0_  ;
	output \g21702/_3_  ;
	output \g21707/_0_  ;
	output \g21709/_0_  ;
	output \g21728/_0_  ;
	output \g21729/_0_  ;
	output \g21731/_0_  ;
	output \g21732/_0_  ;
	output \g21733/_0_  ;
	output \g21736/_0_  ;
	output \g21744/_3_  ;
	output \g21753/_0_  ;
	output \g21754/_0_  ;
	output \g21755/_0_  ;
	output \g21756/_0_  ;
	output \g21757/_0_  ;
	output \g21759/_0_  ;
	output \g21761/_0_  ;
	output \g21763/_0_  ;
	output \g21764/_0_  ;
	output \g21766/_0_  ;
	output \g2180/_0_  ;
	output \g21853/_3_  ;
	output \g21861/_3_  ;
	output \g21863/_3_  ;
	output \g21869/_3_  ;
	output \g2187/_0_  ;
	output \g21875/_3_  ;
	output \g21877/_3_  ;
	output \g21879/_3_  ;
	output \g2188/_0_  ;
	output \g21900/_0_  ;
	output \g22080/_0_  ;
	output \g22082/_0_  ;
	output \g22135/_0_  ;
	output \g22145/_1_  ;
	output \g22225/_0_  ;
	output \g223/_0_  ;
	output \g22354/_0_  ;
	output \g224/_0_  ;
	output \g22412/_0_  ;
	output \g22415/_1__syn_2  ;
	output \g225/_0_  ;
	output \g2257/_0_  ;
	output \g226/_3_  ;
	output \g22624/_0_  ;
	output \g227/_3_  ;
	output \g22702/_0_  ;
	output \g22919/_1__syn_2  ;
	output \g22933/_0_  ;
	output \g22954/_0_  ;
	output \g22989/_1_  ;
	output \g23529/_0_  ;
	output \g23539/_0_  ;
	output \g2362/_2_  ;
	output \g23766/_0_  ;
	output \g24/_3_  ;
	output \g24018/_0_  ;
	output \g2416/_0_  ;
	output \g2420/_0_  ;
	output \g24213/_0_  ;
	output \g24301/_0_  ;
	output \g2479/_0_  ;
	output \g248/_3_  ;
	output \g2480/_0_  ;
	output \g2481/_0_  ;
	output \g2482/_0_  ;
	output \g2483/_0_  ;
	output \g2484/_0_  ;
	output \g2485/_0_  ;
	output \g2486/_0_  ;
	output \g2487/_0_  ;
	output \g2488/_0_  ;
	output \g249/_3_  ;
	output \g2490/_0_  ;
	output \g2491/_0_  ;
	output \g2492/_0_  ;
	output \g2493/_0_  ;
	output \g2494/_0_  ;
	output \g2495/_0_  ;
	output \g2496/_0_  ;
	output \g2497/_0_  ;
	output \g2507/_0_  ;
	output \g2508/_0_  ;
	output \g2509/_0_  ;
	output \g2510/_0_  ;
	output \g2511/_0_  ;
	output \g2512/_0_  ;
	output \g2513/_0_  ;
	output \g2514/_0_  ;
	output \g2515/_0_  ;
	output \g2516/_0_  ;
	output \g25237/_0_  ;
	output \g2558/_0_  ;
	output \g2562/_0_  ;
	output \g2563/_0_  ;
	output \g2564/_0_  ;
	output \g2565/_0_  ;
	output \g2566/_0_  ;
	output \g2567/_0_  ;
	output \g2699/_0_  ;
	output \g27/_2_  ;
	output \g271/_0_  ;
	output \g272/_3_  ;
	output \g273/_3_  ;
	output \g274/_3_  ;
	output \g275/_3_  ;
	output \g276/_3_  ;
	output \g277/_3_  ;
	output \g2787/_3_  ;
	output \g2788/_3_  ;
	output \g279/_0_  ;
	output \g2795/_0_  ;
	output \g2796/_0_  ;
	output \g280/_0_  ;
	output \g2842/_3_  ;
	output \g29/_1_  ;
	output \g2927/_0_  ;
	output \g2978/_0_  ;
	output \g2979/_0_  ;
	output \g2980/_0_  ;
	output \g2981/_0_  ;
	output \g2982/_0_  ;
	output \g2983/_0_  ;
	output \g2984/_0_  ;
	output \g2985/_0_  ;
	output \g3021/_3_  ;
	output \g3022/_3_  ;
	output \g3023/_3_  ;
	output \g3024/_3_  ;
	output \g3025/_3_  ;
	output \g3026/_3_  ;
	output \g3027/_3_  ;
	output \g3028/_3_  ;
	output \g3029/_3_  ;
	output \g3030/_3_  ;
	output \g3031/_3_  ;
	output \g3032/_3_  ;
	output \g3033/_3_  ;
	output \g3034/_3_  ;
	output \g3035/_3_  ;
	output \g3036/_3_  ;
	output \g3037/_3_  ;
	output \g3038/_3_  ;
	output \g3039/_3_  ;
	output \g3040/_3_  ;
	output \g3041/_3_  ;
	output \g3042/_3_  ;
	output \g3049/_0_  ;
	output \g3050/_0_  ;
	output \g3051/_0_  ;
	output \g3052/_0_  ;
	output \g3053/_0_  ;
	output \g3054/_0_  ;
	output \g3058/_0_  ;
	output \g3059/_0_  ;
	output \g3088/_0_  ;
	output \g3089/_0_  ;
	output \g3090/_0_  ;
	output \g3091/_0_  ;
	output \g3092/_0_  ;
	output \g3093/_0_  ;
	output \g3094/_0_  ;
	output \g3095/_0_  ;
	output \g314/_0_  ;
	output \g3147/_3_  ;
	output \g3148/_3_  ;
	output \g3189/_0_  ;
	output \g3190/_0_  ;
	output \g3191/_0_  ;
	output \g3192/_0_  ;
	output \g3193/_0_  ;
	output \g3194/_0_  ;
	output \g3195/_0_  ;
	output \g3196/_0_  ;
	output \g3197/_0_  ;
	output \g3198/_0_  ;
	output \g3199/_0_  ;
	output \g32/_0_  ;
	output \g320/_3_  ;
	output \g3200/_0_  ;
	output \g3201/_0_  ;
	output \g3202/_0_  ;
	output \g3203/_0_  ;
	output \g3204/_0_  ;
	output \g321/_3_  ;
	output \g325/_3_  ;
	output \g3271/_2_  ;
	output \g33/_0_  ;
	output \g3363/_0_  ;
	output \g3413/_0_  ;
	output \g3414/_0_  ;
	output \g352/_0_  ;
	output \g355/_0_  ;
	output \g356/_3_  ;
	output \g357/_3_  ;
	output \g35_dup/_1_  ;
	output \g36/_3_  ;
	output \g365/_3_  ;
	output \g366/_3_  ;
	output \g367/_3_  ;
	output \g368/_3_  ;
	output \g3687/_0_  ;
	output \g369/_3_  ;
	output \g37/_3_  ;
	output \g370/_3_  ;
	output \g372/_3_  ;
	output \g374/_3_  ;
	output \g3740/_0_  ;
	output \g375/_3_  ;
	output \g376/_3_  ;
	output \g3878/_0_  ;
	output \g3879/_0_  ;
	output \g388/_3_  ;
	output \g3880/_0_  ;
	output \g3881/_0_  ;
	output \g3882/_0_  ;
	output \g389/_3_  ;
	output \g3894/_0_  ;
	output \g3895/_0_  ;
	output \g3896/_0_  ;
	output \g3897/_0_  ;
	output \g3898/_0_  ;
	output \g392/_3_  ;
	output \g393/_3_  ;
	output \g394/_3_  ;
	output \g395/_3_  ;
	output \g396/_3_  ;
	output \g397/_3_  ;
	output \g398/_3_  ;
	output \g399/_3_  ;
	output \g401/_3_  ;
	output \g402/_3_  ;
	output \g404/_3_  ;
	output \g4048/_0_  ;
	output \g405/_3_  ;
	output \g4050/_0_  ;
	output \g406/_3_  ;
	output \g407/_3_  ;
	output \g410/_3_  ;
	output \g411/_3_  ;
	output \g412/_3_  ;
	output \g413/_3_  ;
	output \g415/_3_  ;
	output \g416/_3_  ;
	output \g42/_0_  ;
	output \g4216/_3_  ;
	output \g4217/_3_  ;
	output \g4218/_3_  ;
	output \g4219/_3_  ;
	output \g4296/_0_  ;
	output \g4297/_0_  ;
	output \g4298/_0_  ;
	output \g4299/_0_  ;
	output \g43/_0_  ;
	output \g4300/_0_  ;
	output \g4301/_0_  ;
	output \g4302/_0_  ;
	output \g4303/_0_  ;
	output \g4304/_0_  ;
	output \g4305/_0_  ;
	output \g4306/_0_  ;
	output \g4307/_0_  ;
	output \g4308/_0_  ;
	output \g4309/_0_  ;
	output \g4310/_0_  ;
	output \g4311/_0_  ;
	output \g4312/_0_  ;
	output \g4313/_0_  ;
	output \g4314/_0_  ;
	output \g4315/_0_  ;
	output \g4316/_0_  ;
	output \g4317/_0_  ;
	output \g4318/_0_  ;
	output \g4319/_0_  ;
	output \g4320/_0_  ;
	output \g4321/_0_  ;
	output \g4322/_0_  ;
	output \g4323/_0_  ;
	output \g436/_0_  ;
	output \g44/_0_  ;
	output \g448/_3_  ;
	output \g45/_0_  ;
	output \g4587/_0_  ;
	output \g4588/_0_  ;
	output \g46/_0_  ;
	output \g4601/_0_  ;
	output \g4602/_0_  ;
	output \g4613/_3_  ;
	output \g4614/_3_  ;
	output \g4615/_3_  ;
	output \g463/_0_  ;
	output \g465/_0_  ;
	output \g4653/_0_  ;
	output \g4654/_0_  ;
	output \g4655/_0_  ;
	output \g4656/_0_  ;
	output \g4659/_0_  ;
	output \g466/_0_  ;
	output \g468/_3_  ;
	output \g469/_3_  ;
	output \g4697/_0_  ;
	output \g47/_3_  ;
	output \g470/_0_  ;
	output \g471/_0_  ;
	output \g4755/_0_  ;
	output \g476/_0_  ;
	output \g48/_3_  ;
	output \g480/_00_  ;
	output \g4839/_0_  ;
	output \g4840/_0_  ;
	output \g485/_3_  ;
	output \g4854/_0_  ;
	output \g4855/_0_  ;
	output \g4859/_0_  ;
	output \g486/_3_  ;
	output \g4860/_0_  ;
	output \g4880/_0_  ;
	output \g4881/_0_  ;
	output \g4882/_0_  ;
	output \g4883/_0_  ;
	output \g4884/_0_  ;
	output \g4885/_0_  ;
	output \g4886/_0_  ;
	output \g4887/_0_  ;
	output \g4888/_0_  ;
	output \g49/_0_  ;
	output \g494/_0_  ;
	output \g499/_1_  ;
	output \g50/_0_  ;
	output \g5002/_0_  ;
	output \g5003/_0_  ;
	output \g5009/_0_  ;
	output \g5010/_0_  ;
	output \g5011/_0_  ;
	output \g5014/_0_  ;
	output \g51/_0_  ;
	output \g5105/_0_  ;
	output \g5129/_2_  ;
	output \g5132/_0_  ;
	output \g5135/_0_  ;
	output \g5168/_0_  ;
	output \g5169/_0_  ;
	output \g5173/_0_  ;
	output \g5224/_0_  ;
	output \g5225/_0_  ;
	output \g5226/_0_  ;
	output \g5227/_0_  ;
	output \g5334/_0_  ;
	output \g5335/_0_  ;
	output \g5336/_0_  ;
	output \g5337/_0_  ;
	output \g5338/_0_  ;
	output \g5339/_0_  ;
	output \g5340/_0_  ;
	output \g5341/_0_  ;
	output \g5342/_0_  ;
	output \g5343/_0_  ;
	output \g5344/_0_  ;
	output \g5345/_0_  ;
	output \g5346/_0_  ;
	output \g5347/_0_  ;
	output \g5348/_0_  ;
	output \g5349/_0_  ;
	output \g5395/_0_  ;
	output \g54/_0_  ;
	output \g5434/_0_  ;
	output \g5447/_0_  ;
	output \g5450/_0_  ;
	output \g5451/_0_  ;
	output \g5452/_0_  ;
	output \g5453/_0_  ;
	output \g5454/_0_  ;
	output \g5461/_0_  ;
	output \g5483/_0_  ;
	output \g5484/_0_  ;
	output \g5492/_0_  ;
	output \g5493/_0_  ;
	output \g5496/_3_  ;
	output \g5497/_3_  ;
	output \g55/_0_  ;
	output \g5500/_0_  ;
	output \g5502/_0_  ;
	output \g5503/_0_  ;
	output \g5506/_0_  ;
	output \g5511/_0_  ;
	output \g5518/_0_  ;
	output \g5519/_0_  ;
	output \g5520/_0_  ;
	output \g5522/_0_  ;
	output \g5523/_0_  ;
	output \g5524/_0_  ;
	output \g5525/_0_  ;
	output \g5532/_0_  ;
	output \g5533/_0_  ;
	output \g5534/_0_  ;
	output \g5535/_0_  ;
	output \g5536/_0_  ;
	output \g5537/_0_  ;
	output \g5538/_0_  ;
	output \g5546/_0_  ;
	output \g5555/_00_  ;
	output \g5593/_0_  ;
	output \g5614/_2_  ;
	output \g567/_0_  ;
	output \g5677/_0_  ;
	output \g5678/_0_  ;
	output \g5682/_0_  ;
	output \g5683/_0_  ;
	output \g5684/_0_  ;
	output \g5686/_0_  ;
	output \g5687/_0_  ;
	output \g5689/_0_  ;
	output \g5690/_0_  ;
	output \g5691/_0_  ;
	output \g5692/_0_  ;
	output \g5698/_0_  ;
	output \g5699/_0_  ;
	output \g5700/_0_  ;
	output \g5701/_0_  ;
	output \g5702/_0_  ;
	output \g5703/_0_  ;
	output \g5704/_0_  ;
	output \g5709/_0_  ;
	output \g5711/_0_  ;
	output \g5714/_0_  ;
	output \g572/_0_  ;
	output \g5723/_0_  ;
	output \g5724/_0_  ;
	output \g5725/_0_  ;
	output \g573/_0_  ;
	output \g5739/_0_  ;
	output \g5740/_0_  ;
	output \g575/_0_  ;
	output \g5756/_0_  ;
	output \g5757/_0_  ;
	output \g5758/_0_  ;
	output \g5759/_0_  ;
	output \g576/_0_  ;
	output \g5760/_0_  ;
	output \g5761/_0_  ;
	output \g5762/_0_  ;
	output \g5763/_0_  ;
	output \g577/_0_  ;
	output \g5772/_0_  ;
	output \g5773/_0_  ;
	output \g5774/_0_  ;
	output \g5775/_0_  ;
	output \g5776/_0_  ;
	output \g5777/_0_  ;
	output \g578/_0_  ;
	output \g5781/_0_  ;
	output \g5783/_0_  ;
	output \g5784/_0_  ;
	output \g5785/_0_  ;
	output \g5786/_0_  ;
	output \g5787/_0_  ;
	output \g5788/_0_  ;
	output \g5789/_0_  ;
	output \g579/_0_  ;
	output \g5790/_0_  ;
	output \g5791/_0_  ;
	output \g5792/_0_  ;
	output \g5794/_0_  ;
	output \g5795/_0_  ;
	output \g5796/_0_  ;
	output \g580/_0_  ;
	output \g5801/_0_  ;
	output \g5802/_0_  ;
	output \g5803/_0_  ;
	output \g5804/_0_  ;
	output \g5805/_0_  ;
	output \g581/_0_  ;
	output \g5814/_0_  ;
	output \g582/_0_  ;
	output \g583/_0_  ;
	output \g5849/_3_  ;
	output \g585/_0_  ;
	output \g586/_0_  ;
	output \g587/_0_  ;
	output \g588/_0_  ;
	output \g589/_0_  ;
	output \g590/_0_  ;
	output \g591/_0_  ;
	output \g592/_0_  ;
	output \g593/_0_  ;
	output \g594/_0_  ;
	output \g595/_0_  ;
	output \g596/_0_  ;
	output \g597/_0_  ;
	output \g5971/_0_  ;
	output \g5972/_0_  ;
	output \g5976/_0_  ;
	output \g598/_0_  ;
	output \g5989/_0_  ;
	output \g599/_0_  ;
	output \g600/_0_  ;
	output \g601/_0_  ;
	output \g602/_0_  ;
	output \g603/_0_  ;
	output \g604/_0_  ;
	output \g605/_0_  ;
	output \g6092/_0_  ;
	output \g6093/_2_  ;
	output \g6094/_0_  ;
	output \g6114/_0_  ;
	output \g614/_3_  ;
	output \g6148/_0_  ;
	output \g6149/_0_  ;
	output \g6171/_0_  ;
	output \g6172/_0_  ;
	output \g6173/_0_  ;
	output \g6174/_0_  ;
	output \g6175/_0_  ;
	output \g6176/_0_  ;
	output \g6177/_0_  ;
	output \g6178/_0_  ;
	output \g6179/_0_  ;
	output \g6180/_0_  ;
	output \g6181/_0_  ;
	output \g6182/_0_  ;
	output \g6183/_0_  ;
	output \g6184/_0_  ;
	output \g6185/_0_  ;
	output \g6186/_0_  ;
	output \g6187/_0_  ;
	output \g6193/_0_  ;
	output \g6196/_0_  ;
	output \g6197/_0_  ;
	output \g6198/_3_  ;
	output \g6200/_2_  ;
	output \g6202/_2_  ;
	output \g6203/_3_  ;
	output \g6204/_3_  ;
	output \g6209/_0_  ;
	output \g6211/_0_  ;
	output \g6215/_0_  ;
	output \g6217/_0_  ;
	output \g6219/_0_  ;
	output \g6220/_0_  ;
	output \g6222/_0_  ;
	output \g6224/_0_  ;
	output \g6228/_0_  ;
	output \g6238/_0_  ;
	output \g6239/_0_  ;
	output \g6240/_0_  ;
	output \g6242/_0_  ;
	output \g6243/_0_  ;
	output \g6244/_0_  ;
	output \g6245/_0_  ;
	output \g6246/_0_  ;
	output \g6248/_0_  ;
	output \g6249/_0_  ;
	output \g6259/_0_  ;
	output \g6260/_0_  ;
	output \g6261/_0_  ;
	output \g6262/_0_  ;
	output \g6263/_0_  ;
	output \g6264/_0_  ;
	output \g6265/_0_  ;
	output \g6266/_0_  ;
	output \g6267/_0_  ;
	output \g6268/_0_  ;
	output \g6269/_0_  ;
	output \g6270/_0_  ;
	output \g6271/_0_  ;
	output \g6272/_0_  ;
	output \g6277/_0_  ;
	output \g6318/_0_  ;
	output \g6326/_0_  ;
	output \g6329/_0_  ;
	output \g6330/_0_  ;
	output \g6331/_0_  ;
	output \g6332/_0_  ;
	output \g6333/_0_  ;
	output \g6334/_0_  ;
	output \g6335/_0_  ;
	output \g6336/_0_  ;
	output \g6337/_0_  ;
	output \g6338/_0_  ;
	output \g6339/_0_  ;
	output \g6340/_0_  ;
	output \g6341/_0_  ;
	output \g6342/_0_  ;
	output \g6343/_0_  ;
	output \g6344/_0_  ;
	output \g6345/_0_  ;
	output \g6346/_0_  ;
	output \g6347/_0_  ;
	output \g6348/_0_  ;
	output \g6349/_0_  ;
	output \g6350/_0_  ;
	output \g6351/_0_  ;
	output \g6352/_0_  ;
	output \g6353/_0_  ;
	output \g6354/_0_  ;
	output \g6355/_0_  ;
	output \g6361/_0_  ;
	output \g637/_0_  ;
	output \g638/_0_  ;
	output \g639/_3_  ;
	output \g64/_3_  ;
	output \g640/_3_  ;
	output \g6419/_0_  ;
	output \g6442/_0_  ;
	output \g6442/_1_  ;
	output \g6489/_0_  ;
	output \g6490/_0_  ;
	output \g65/_3_  ;
	output \g6513/_0_  ;
	output \g6515/_0_  ;
	output \g6571/_0_  ;
	output \g6588/_0_  ;
	output \g6589/_0_  ;
	output \g6638/_0_  ;
	output \g6639/_0_  ;
	output \g6653/_0_  ;
	output \g6654/_3_  ;
	output \g6655/_0_  ;
	output \g6656/_0_  ;
	output \g6657/_0_  ;
	output \g6687/_0_  ;
	output \g6688/_0_  ;
	output \g6689/_0_  ;
	output \g6690/_0_  ;
	output \g6691/_0_  ;
	output \g6692/_0_  ;
	output \g6693/_0_  ;
	output \g6694/_0_  ;
	output \g6701/_0_  ;
	output \g6706/_0_  ;
	output \g6711/_0_  ;
	output \g6727/_0_  ;
	output \g6728/_0_  ;
	output \g6736/_0_  ;
	output \g6739/_0_  ;
	output \g6742/_0_  ;
	output \g6746/_0_  ;
	output \g6752/_0_  ;
	output \g6771/_0_  ;
	output \g684/_0_  ;
	output \g685/_0_  ;
	output \g686/_0_  ;
	output \g687/_0_  ;
	output \g688/_0_  ;
	output \g689/_0_  ;
	output \g690/_0_  ;
	output \g691/_0_  ;
	output \g692/_0_  ;
	output \g693/_0_  ;
	output \g696/_3_  ;
	output \g697/_3_  ;
	output \g699/_0_  ;
	output \g7/_0_  ;
	output \g700/_0_  ;
	output \g7005/_0_  ;
	output \g7056/_0_  ;
	output \g7057/_0_  ;
	output \g7058/_0_  ;
	output \g7060/_0_  ;
	output \g7075/_0_  ;
	output \g7086/_0_  ;
	output \g7087/_0_  ;
	output \g7089/_0_  ;
	output \g7108/_0_  ;
	output \g7109/_0_  ;
	output \g7112/_0_  ;
	output \g7172/_2_  ;
	output \g7210/_2_  ;
	output \g7211/_0_  ;
	output \g7212/_0_  ;
	output \g7213/_0_  ;
	output \g7214/_0_  ;
	output \g7215/_0_  ;
	output \g7216/_0_  ;
	output \g7217/_3_  ;
	output \g7218/_0_  ;
	output \g7219/_0_  ;
	output \g7220/_0_  ;
	output \g7222/_0_  ;
	output \g7227/_2_  ;
	output \g723/_3_  ;
	output \g7234/_0_  ;
	output \g7237/_3_  ;
	output \g7238/_3_  ;
	output \g7239/_3_  ;
	output \g724/_3_  ;
	output \g7240/_3_  ;
	output \g7241/_3_  ;
	output \g7242/_3_  ;
	output \g7243/_3_  ;
	output \g7244/_0_  ;
	output \g7245/_0_  ;
	output \g7246/_0_  ;
	output \g7247/_0_  ;
	output \g7248/_0_  ;
	output \g7249/_0_  ;
	output \g7250/_0_  ;
	output \g7251/_0_  ;
	output \g7253/_0_  ;
	output \g7254/_0_  ;
	output \g7255/_0_  ;
	output \g7256/_0_  ;
	output \g7257/_0_  ;
	output \g7258/_0_  ;
	output \g7261/_0_  ;
	output \g7264/_0_  ;
	output \g7265/_0_  ;
	output \g7266/_0_  ;
	output \g7267/_0_  ;
	output \g7268/_0_  ;
	output \g7269/_0_  ;
	output \g7278/_0_  ;
	output \g7279/_0_  ;
	output \g7280/_0_  ;
	output \g7281/_0_  ;
	output \g7282/_0_  ;
	output \g7283/_0_  ;
	output \g7284/_0_  ;
	output \g7285/_0_  ;
	output \g7286/_3_  ;
	output \g7288/_3_  ;
	output \g7291/_0_  ;
	output \g7296/_3_  ;
	output \g73/_0_  ;
	output \g7302/_3_  ;
	output \g7306/_3_  ;
	output \g7310/_3_  ;
	output \g7311/_3_  ;
	output \g7312/_3_  ;
	output \g7313/_3_  ;
	output \g7314/_3_  ;
	output \g7315/_3_  ;
	output \g7316/_3_  ;
	output \g7317/_3_  ;
	output \g7323/_3_  ;
	output \g7324/_3_  ;
	output \g7325/_3_  ;
	output \g7327/_0_  ;
	output \g7362/_0_  ;
	output \g74/_0_  ;
	output \g75/_0_  ;
	output \g7512/_0_  ;
	output \g7513/_0_  ;
	output \g7514/_0_  ;
	output \g7515/_0_  ;
	output \g7516/_0_  ;
	output \g7518/_0_  ;
	output \g7528/_0_  ;
	output \g7529/_0_  ;
	output \g7548/_0_  ;
	output \g7549/_0_  ;
	output \g7550/_0_  ;
	output \g7575/_0_  ;
	output \g7576/_0_  ;
	output \g7577/_0_  ;
	output \g7578/_0_  ;
	output \g7579/_0_  ;
	output \g7580/_0_  ;
	output \g7581/_0_  ;
	output \g7582/_0_  ;
	output \g7583/_0_  ;
	output \g7584/_0_  ;
	output \g7585/_0_  ;
	output \g7586/_0_  ;
	output \g7587/_0_  ;
	output \g7588/_0_  ;
	output \g7589/_0_  ;
	output \g7590/_0_  ;
	output \g7591/_0_  ;
	output \g7592/_0_  ;
	output \g7593/_0_  ;
	output \g7594/_0_  ;
	output \g7595/_0_  ;
	output \g7596/_0_  ;
	output \g7597/_0_  ;
	output \g7598/_0_  ;
	output \g7599/_0_  ;
	output \g76/_0_  ;
	output \g7600/_0_  ;
	output \g7601/_0_  ;
	output \g7602/_0_  ;
	output \g7603/_0_  ;
	output \g7604/_0_  ;
	output \g7614/_0_  ;
	output \g7618/_0_  ;
	output \g762/_0_  ;
	output \g7634/_0_  ;
	output \g766/_0_  ;
	output \g767/_0_  ;
	output \g768/_0_  ;
	output \g769/_0_  ;
	output \g77/_0_  ;
	output \g770/_3_  ;
	output \g771/_3_  ;
	output \g7715/_0_  ;
	output \g774/_0_  ;
	output \g7746/_0_  ;
	output \g7753/_0_  ;
	output \g7754/_0_  ;
	output \g7755/_0_  ;
	output \g7756/_0_  ;
	output \g7757/_0_  ;
	output \g7758/_0_  ;
	output \g7759/_0_  ;
	output \g7760/_0_  ;
	output \g7761/_0_  ;
	output \g7762/_0_  ;
	output \g7763/_0_  ;
	output \g7764/_0_  ;
	output \g7765/_0_  ;
	output \g7766/_0_  ;
	output \g7778/_0_  ;
	output \g7779/_0_  ;
	output \g7780/_0_  ;
	output \g7781/_0_  ;
	output \g7782/_0_  ;
	output \g7784/_0_  ;
	output \g78/_0_  ;
	output \g7800/_0_  ;
	output \g7823/_3_  ;
	output \g7837/_0_  ;
	output \g7841/_0_  ;
	output \g7842/_0_  ;
	output \g7843/_0_  ;
	output \g7844/_0_  ;
	output \g7845/_0_  ;
	output \g7846/_0_  ;
	output \g7847/_0_  ;
	output \g7849/_0_  ;
	output \g7850/_0_  ;
	output \g7852/_0_  ;
	output \g7854/_0_  ;
	output \g7855/_0_  ;
	output \g7857/_0_  ;
	output \g7858/_0_  ;
	output \g7859/_0_  ;
	output \g7860/_0_  ;
	output \g7861/_0_  ;
	output \g7862/_0_  ;
	output \g7863/_0_  ;
	output \g7864/_0_  ;
	output \g7865/_0_  ;
	output \g7866/_0_  ;
	output \g7867/_0_  ;
	output \g7868/_0_  ;
	output \g7869/_0_  ;
	output \g7870/_0_  ;
	output \g7871/_0_  ;
	output \g79211/_3_  ;
	output \g79258/_3_  ;
	output \g79299/_3_  ;
	output \g79316/_2_  ;
	output \g79342/_3_  ;
	output \g79401/_3_  ;
	output \g79452/_3_  ;
	output \g79457/_3_  ;
	output \g7951/_0_  ;
	output \g79541/_3_  ;
	output \g7958/_0_  ;
	output \g79598/_3_  ;
	output \g79654/_3_  ;
	output \g79675/_3_  ;
	output \g7971/_0_  ;
	output \g7972/_0_  ;
	output \g7973/_3_  ;
	output \g79753/_3_  ;
	output \g7976/_3_  ;
	output \g79855/_3_  ;
	output \g79858/_3_  ;
	output \g79997/_3_  ;
	output \g8/_0_  ;
	output \g80008/_3_  ;
	output \g80011/_0_  ;
	output \g80104/_0_  ;
	output \g80172/_1_  ;
	output \g80195/_3_  ;
	output \g80238/_3_  ;
	output \g80290/_2_  ;
	output \g80294/_0_  ;
	output \g80302/_0_  ;
	output \g80327/_0_  ;
	output \g80360/_3_  ;
	output \g80373/_0_  ;
	output \g80401/_0_  ;
	output \g80410/_0_  ;
	output \g80475/_0_  ;
	output \g80476/_0_  ;
	output \g80516/_3_  ;
	output \g80536/_0_  ;
	output \g80537/_0_  ;
	output \g80572/_0_  ;
	output \g80573/_0_  ;
	output \g80609/_2_  ;
	output \g80610/_2_  ;
	output \g80676/_0_  ;
	output \g80798/_0_  ;
	output \g80807/_0_  ;
	output \g80890/_2_  ;
	output \g80904/_0_  ;
	output \g81719/_2_  ;
	output \g81746/_0_  ;
	output \g81775/_0_  ;
	output \g81872/_0_  ;
	output \g81961/_0_  ;
	output \g81968/_0_  ;
	output \g82096/_0_  ;
	output \g82123/_0_  ;
	output \g82147/_0_  ;
	output \g82147/_1_  ;
	output \g82335/_0_  ;
	output \g82338/_2_  ;
	output \g82368/_0_  ;
	output \g82460/_2_  ;
	output \g82469/_0_  ;
	output \g82481/_0_  ;
	output \g82625/_1_  ;
	output \g82711/_0_  ;
	output \g82772/_0_  ;
	output \g82946/_0_  ;
	output \g82947/_0_  ;
	output \g82956/_0_  ;
	output \g83003/_0_  ;
	output \g83006/_1_  ;
	output \g83415/_0_  ;
	output \g83498/_0_  ;
	output \g837/_0_  ;
	output \g838/_0_  ;
	output \g83863/_0_  ;
	output \g839/_0_  ;
	output \g84049/_3_  ;
	output \g84050/_3_  ;
	output \g84077/_2_  ;
	output \g842/_0_  ;
	output \g84245/_0_  ;
	output \g843/_0_  ;
	output \g844/_0_  ;
	output \g84448/_0_  ;
	output \g84478/_3_  ;
	output \g845/_0_  ;
	output \g846/_0_  ;
	output \g847/_0_  ;
	output \g848/_0_  ;
	output \g8487/_0_  ;
	output \g8488/_0_  ;
	output \g8489/_0_  ;
	output \g849/_0_  ;
	output \g8490/_0_  ;
	output \g84904/_0_  ;
	output \g8491/_0_  ;
	output \g8492/_0_  ;
	output \g8493/_0_  ;
	output \g8494/_0_  ;
	output \g8496/_0_  ;
	output \g8517/_0_  ;
	output \g8534/_0_  ;
	output \g8538/_0_  ;
	output \g8540/_0_  ;
	output \g8576/_2_  ;
	output \g8597/_0_  ;
	output \g8598/_0_  ;
	output \g8599/_0_  ;
	output \g8600/_0_  ;
	output \g8601/_0_  ;
	output \g8602/_0_  ;
	output \g8603/_0_  ;
	output \g8605/_0_  ;
	output \g8606/_0_  ;
	output \g8607/_0_  ;
	output \g8608/_0_  ;
	output \g8609/_0_  ;
	output \g8610/_0_  ;
	output \g8611/_0_  ;
	output \g8612/_0_  ;
	output \g8613/_0_  ;
	output \g8614/_0_  ;
	output \g8615/_0_  ;
	output \g8617/_0_  ;
	output \g8643/_0_  ;
	output \g8644/_0_  ;
	output \g8645/_0_  ;
	output \g8646/_0_  ;
	output \g8647/_0_  ;
	output \g8648/_0_  ;
	output \g8650/_0_  ;
	output \g8651/_0_  ;
	output \g8652/_0_  ;
	output \g8653/_0_  ;
	output \g8654/_0_  ;
	output \g8655/_0_  ;
	output \g8656/_0_  ;
	output \g8657/_0_  ;
	output \g8658/_0_  ;
	output \g8659/_0_  ;
	output \g8660/_0_  ;
	output \g8665/_00_  ;
	output \g8666/_00_  ;
	output \g8667/_00_  ;
	output \g8668/_00_  ;
	output \g8669/_00_  ;
	output \g86715/_0_  ;
	output \g86745/_3_  ;
	output \g8691/_0_  ;
	output \g8700/_0_  ;
	output \g8701/_0_  ;
	output \g8702/_0_  ;
	output \g8703/_0_  ;
	output \g8704/_0_  ;
	output \g8705/_0_  ;
	output \g87063/_0_  ;
	output \g87114/_0_  ;
	output \g8712/_0_  ;
	output \g8713/_0_  ;
	output \g8714/_0_  ;
	output \g87171/_1_  ;
	output \g87252/_1_  ;
	output \g87298/_0_  ;
	output \g8730/_0_  ;
	output \g8741/_0_  ;
	output \g8747/_0_  ;
	output \g87480/_0_  ;
	output \g87484/_2_  ;
	output \g87488/_1__syn_2  ;
	output \g8761/_0_  ;
	output \g8762/_0_  ;
	output \g8763/_0_  ;
	output \g8764/_0_  ;
	output \g8765/_0_  ;
	output \g8775/_0_  ;
	output \g8776/_0_  ;
	output \g8777/_0_  ;
	output \g8778/_0_  ;
	output \g8784/_0_  ;
	output \g8804/_0_  ;
	output \g8807/_0_  ;
	output \g8808/_0_  ;
	output \g8809/_0_  ;
	output \g8810/_0_  ;
	output \g8811/_0_  ;
	output \g8812/_0_  ;
	output \g8813/_0_  ;
	output \g8814/_0_  ;
	output \g8815/_0_  ;
	output \g8816/_0_  ;
	output \g8817/_0_  ;
	output \g8818/_0_  ;
	output \g8819/_0_  ;
	output \g8820/_0_  ;
	output \g8821/_0_  ;
	output \g8822/_0_  ;
	output \g8823/_0_  ;
	output \g8824/_0_  ;
	output \g8825/_0_  ;
	output \g8826/_0_  ;
	output \g8827/_0_  ;
	output \g8828/_0_  ;
	output \g8829/_0_  ;
	output \g8830/_0_  ;
	output \g8831/_0_  ;
	output \g8832/_0_  ;
	output \g8833/_0_  ;
	output \g8834/_0_  ;
	output \g8835/_0_  ;
	output \g8836/_0_  ;
	output \g8837/_0_  ;
	output \g8838/_0_  ;
	output \g8839/_0_  ;
	output \g8840/_0_  ;
	output \g8842/_0_  ;
	output \g8843/_0_  ;
	output \g8846/_0_  ;
	output \g8848/_0_  ;
	output \g8857/_0_  ;
	output \g8895/_0_  ;
	output \g8902/_3_  ;
	output \g8903/_3_  ;
	output \g8904/_3_  ;
	output \g8905/_3_  ;
	output \g8906/_3_  ;
	output \g8909/_0_  ;
	output \g8910/_0_  ;
	output \g8911/_0_  ;
	output \g8924/_3_  ;
	output \g8926/_3_  ;
	output \g8927/_3_  ;
	output \g8943/_0_  ;
	output \g8944/_0_  ;
	output \g8958/_3_  ;
	output \g8960/_00_  ;
	output \g8961/_3_  ;
	output \g8965/_0_  ;
	output \g8966/_0_  ;
	output \g8967/_0_  ;
	output \g8968/_0_  ;
	output \g9/_0_  ;
	output \g9123/_0_  ;
	output \g9125/_0_  ;
	output \g9126/_0_  ;
	output \g913/_0_  ;
	output \g915/_0_  ;
	output \g916/_0_  ;
	output \g917/_0_  ;
	output \g918/_0_  ;
	output \g919/_0_  ;
	output \g920/_3_  ;
	output \g921/_3_  ;
	output \g925/_0_  ;
	output \g926/_0_  ;
	output \g927/_0_  ;
	output \g928/_0_  ;
	output \g929/_0_  ;
	output \g930/_0_  ;
	output \g9336/_0_  ;
	output \g9337/_0_  ;
	output \g939/_3_  ;
	output \g9396/_0_  ;
	output \g9397/_0_  ;
	output \g9399/_0_  ;
	output \g9400/_0_  ;
	output \g9401/_0_  ;
	output \g9402/_0_  ;
	output \g9403/_0_  ;
	output \g9404/_0_  ;
	output \g9415/_0_  ;
	output \g9418/_0_  ;
	output \g9419/_0_  ;
	output \g9420/_0_  ;
	output \g9446/_0_  ;
	output \g9465/_0_  ;
	output \g9493/_0_  ;
	output \g9536/_0_  ;
	output \g9537/_0_  ;
	output \g9538/_0_  ;
	output \g9539/_0_  ;
	output \g9540/_0_  ;
	output \g9541/_0_  ;
	output \g9542/_0_  ;
	output \g955/_2_  ;
	output \g9561/_0_  ;
	output \g9562/_0_  ;
	output \g9563/_0_  ;
	output \g9564/_0_  ;
	output \g9565/_0_  ;
	output \g9566/_0_  ;
	output \g9567/_0_  ;
	output \g9568/_0_  ;
	output \g9569/_0_  ;
	output \g9570/_0_  ;
	output \g9571/_0_  ;
	output \g9572/_0_  ;
	output \g9573/_0_  ;
	output \g9574/_0_  ;
	output \g9575/_0_  ;
	output \g9576/_0_  ;
	output \g9577/_0_  ;
	output \g9578/_0_  ;
	output \g9579/_0_  ;
	output \g9580/_0_  ;
	output \g9581/_0_  ;
	output \g9582/_0_  ;
	output \g9583/_0_  ;
	output \g9584/_0_  ;
	output \g9585/_0_  ;
	output \g9586/_0_  ;
	output \g9587/_0_  ;
	output \g9588/_0_  ;
	output \g9589/_0_  ;
	output \g9590/_0_  ;
	output \g9591/_0_  ;
	output \g9592/_0_  ;
	output \g9593/_0_  ;
	output \g9594/_0_  ;
	output \g9595/_0_  ;
	output \g9596/_0_  ;
	output \g9597/_0_  ;
	output \g9598/_0_  ;
	output \g9599/_0_  ;
	output \g9600/_0_  ;
	output \g9601/_0_  ;
	output \g9602/_0_  ;
	output \g9603/_0_  ;
	output \g9604/_0_  ;
	output \g9605/_0_  ;
	output \g9606/_0_  ;
	output \g9607/_0_  ;
	output \g9608/_0_  ;
	output \g9609/_0_  ;
	output \g9610/_0_  ;
	output \g9611/_0_  ;
	output \g9612/_0_  ;
	output \g9613/_0_  ;
	output \g9614/_0_  ;
	output \g9615/_0_  ;
	output \g9616/_0_  ;
	output \g9617/_0_  ;
	output \g9618/_0_  ;
	output \g9619/_0_  ;
	output \g9620/_0_  ;
	output \g9621/_0_  ;
	output \g9622/_0_  ;
	output \g9623/_0_  ;
	output \g9624/_0_  ;
	output \g9625/_0_  ;
	output \g9626/_0_  ;
	output \g9627/_0_  ;
	output \g9628/_0_  ;
	output \g9629/_0_  ;
	output \g9630/_0_  ;
	output \g9631/_0_  ;
	output \g9632/_0_  ;
	output \g9633/_0_  ;
	output \g9634/_0_  ;
	output \g9635/_0_  ;
	output \g9636/_0_  ;
	output \g9637/_0_  ;
	output \g9638/_0_  ;
	output \g9639/_0_  ;
	output \g9640/_0_  ;
	output \g9641/_0_  ;
	output \g9642/_0_  ;
	output \g9643/_0_  ;
	output \g9644/_0_  ;
	output \g9645/_0_  ;
	output \g9646/_0_  ;
	output \g9647/_0_  ;
	output \g9648/_0_  ;
	output \g9649/_0_  ;
	output \g9650/_0_  ;
	output \g9651/_0_  ;
	output \g9652/_0_  ;
	output \g9653/_0_  ;
	output \g9654/_0_  ;
	output \g9655/_0_  ;
	output \g9656/_0_  ;
	output \g9657/_0_  ;
	output \g9658/_0_  ;
	output \g9659/_0_  ;
	output \g9660/_0_  ;
	output \g9661/_0_  ;
	output \g9662/_0_  ;
	output \g9663/_0_  ;
	output \g9664/_0_  ;
	output \g9665/_0_  ;
	output \g9666/_0_  ;
	output \g9667/_0_  ;
	output \g9668/_0_  ;
	output \g9669/_0_  ;
	output \g9670/_0_  ;
	output \g9671/_0_  ;
	output \g9672/_0_  ;
	output \g9673/_0_  ;
	output \g9674/_0_  ;
	output \g9675/_0_  ;
	output \g9676/_0_  ;
	output \g9677/_0_  ;
	output \g9678/_0_  ;
	output \g9681/_0_  ;
	output \g9683/_0_  ;
	output \g9689/_0_  ;
	output \g9692/_0_  ;
	output \g9694/_0_  ;
	output \g9695/_0_  ;
	output \g9701/_0_  ;
	output \g9702/_0_  ;
	output \g9703/_0_  ;
	output \g9704/_0_  ;
	output \g9709/_0_  ;
	output \g9710/_0_  ;
	output \g9711/_0_  ;
	output \g9712/_0_  ;
	output \g9720/_0_  ;
	output \g9721/_0_  ;
	output \g9722/_0_  ;
	output \g9726/_0_  ;
	output \g9733/_0_  ;
	output \g9734/_0_  ;
	output \g9735/_0_  ;
	output \g9736/_0_  ;
	output \g9737/_0_  ;
	output \g9738/_0_  ;
	output \g9739/_0_  ;
	output \g9740/_0_  ;
	output \g9741/_0_  ;
	output \g9742/_0_  ;
	output \g9743/_0_  ;
	output \g9744/_0_  ;
	output \g9745/_0_  ;
	output \g9746/_0_  ;
	output \g9747/_0_  ;
	output \g9748/_0_  ;
	output \g9749/_0_  ;
	output \g9750/_0_  ;
	output \g9751/_0_  ;
	output \g9752/_0_  ;
	output \g9753/_0_  ;
	output \g9754/_0_  ;
	output \g9755/_0_  ;
	output \g9756/_0_  ;
	output \g9757/_0_  ;
	output \g9758/_0_  ;
	output \g9759/_0_  ;
	output \g9760/_0_  ;
	output \g9761/_0_  ;
	output \g9762/_0_  ;
	output \g9763/_0_  ;
	output \g9764/_0_  ;
	output \g9765/_0_  ;
	output \g9766/_0_  ;
	output \g9767/_0_  ;
	output \g9768/_0_  ;
	output \g9769/_0_  ;
	output \g9770/_0_  ;
	output \g9771/_0_  ;
	output \g9772/_0_  ;
	output \g9773/_0_  ;
	output \g9774/_0_  ;
	output \g9775/_0_  ;
	output \g9776/_0_  ;
	output \g9777/_0_  ;
	output \g9778/_0_  ;
	output \g9779/_0_  ;
	output \g9780/_0_  ;
	output \g9781/_0_  ;
	output \g9782/_0_  ;
	output \g9783/_0_  ;
	output \g9784/_0_  ;
	output \g9785/_0_  ;
	output \g9786/_0_  ;
	output \g9787/_0_  ;
	output \g9788/_0_  ;
	output \g9789/_0_  ;
	output \g9790/_0_  ;
	output \g9791/_0_  ;
	output \g9792/_0_  ;
	output \g9793/_0_  ;
	output \g9794/_0_  ;
	output \g9795/_0_  ;
	output \g9796/_0_  ;
	output \g9797/_0_  ;
	output \g9798/_0_  ;
	output \g9799/_0_  ;
	output \g9800/_0_  ;
	output \g9801/_0_  ;
	output \g9802/_0_  ;
	output \g9803/_0_  ;
	output \g9804/_0_  ;
	output \g9805/_0_  ;
	output \g9806/_0_  ;
	output \g9807/_0_  ;
	output \g9808/_0_  ;
	output \g9809/_0_  ;
	output \g9810/_0_  ;
	output \g9811/_0_  ;
	output \g9812/_0_  ;
	output \g9813/_0_  ;
	output \g9814/_0_  ;
	output \g9815/_0_  ;
	output \g9816/_0_  ;
	output \g9817/_0_  ;
	output \g9818/_0_  ;
	output \g9819/_0_  ;
	output \g9820/_0_  ;
	output \g9821/_0_  ;
	output \g9822/_0_  ;
	output \g9823/_0_  ;
	output \g9824/_0_  ;
	output \g9825/_0_  ;
	output \g9826/_0_  ;
	output \g9827/_0_  ;
	output \g9828/_0_  ;
	output \g9829/_0_  ;
	output \g9830/_0_  ;
	output \g9831/_0_  ;
	output \g9832/_0_  ;
	output \g9833/_0_  ;
	output \g9835/_0_  ;
	output \g9836/_0_  ;
	output \g9837/_0_  ;
	output \g9838/_0_  ;
	output \g9839/_0_  ;
	output \g9840/_0_  ;
	output \g9841/_0_  ;
	output \g9842/_0_  ;
	output \g9844/_0_  ;
	output \g9845/_0_  ;
	output \g9846/_0_  ;
	output \g9848/_0_  ;
	output \g9849/_0_  ;
	output \g9850/_0_  ;
	output \g9851/_0_  ;
	output \g9853/_0_  ;
	output \g9854/_0_  ;
	output \g9855/_0_  ;
	output \g9856/_0_  ;
	output \g9857/_0_  ;
	output \g9858/_0_  ;
	output \g9859/_0_  ;
	output \g9860/_0_  ;
	output \g9862/_0_  ;
	output \g9863/_0_  ;
	output \g9864/_0_  ;
	output \g9865/_0_  ;
	output \g9867/_0_  ;
	output \g9868/_0_  ;
	output \g9876/_0_  ;
	output \g9877/_0_  ;
	output \g9878/_0_  ;
	output \g9879/_0_  ;
	output \g9880/_0_  ;
	output \g9881/_0_  ;
	output \g9898/_0_  ;
	output \g9900/_0_  ;
	output \g9901/_0_  ;
	output \g9902/_0_  ;
	output \g9903/_0_  ;
	output \g9904/_0_  ;
	output \g9905/_0_  ;
	output \g9906/_0_  ;
	output \g9907/_0_  ;
	output \g9908/_0_  ;
	output \g9909/_0_  ;
	output \g9910/_0_  ;
	output \g9911/_0_  ;
	output \g9912/_0_  ;
	output \g9913/_0_  ;
	output \g9914/_0_  ;
	output \g9915/_0_  ;
	output \g9916/_0_  ;
	output \g9917/_0_  ;
	output \g9918/_0_  ;
	output \g9919/_0_  ;
	output \g992/_0_  ;
	output \g9920/_0_  ;
	output \g9921/_0_  ;
	output \g9922/_0_  ;
	output \g9923/_0_  ;
	output \g9924/_0_  ;
	output \g9925/_0_  ;
	output \g9926/_0_  ;
	output \g9927/_0_  ;
	output \g9928/_0_  ;
	output \g9929/_0_  ;
	output \g9930/_0_  ;
	output \g9931/_0_  ;
	output \g9932/_0_  ;
	output \g9933/_0_  ;
	output \g9934/_0_  ;
	output \g9935/_0_  ;
	output \g9936/_0_  ;
	output \g9937/_0_  ;
	output \g9938/_0_  ;
	output \g9939/_0_  ;
	output \g9940/_0_  ;
	output \g9941/_0_  ;
	output \g9942/_0_  ;
	output \g9943/_0_  ;
	output \g9944/_0_  ;
	output \g9945/_0_  ;
	output \g9946/_0_  ;
	output \g9947/_0_  ;
	output \g9948/_0_  ;
	output \g9949/_0_  ;
	output \g9950/_0_  ;
	output \g9951/_0_  ;
	output \g9952/_0_  ;
	output \g9953/_0_  ;
	output \g9954/_0_  ;
	output \g9955/_0_  ;
	output \g9956/_0_  ;
	output \g9957/_0_  ;
	output \g9958/_0_  ;
	output \g9959/_0_  ;
	output \g9960/_0_  ;
	output \g9961/_0_  ;
	output \g9962/_0_  ;
	output \g9963/_0_  ;
	output \g9964/_0_  ;
	output \g9965/_0_  ;
	output \g9966/_0_  ;
	output \g9967/_0_  ;
	output \g9968/_0_  ;
	output \g9969/_0_  ;
	output \g9970/_0_  ;
	output \g9971/_0_  ;
	output \g9972/_0_  ;
	output \g9973/_0_  ;
	output \g9974/_0_  ;
	output \g9975/_0_  ;
	output \g9976/_0_  ;
	output \g9977/_0_  ;
	output \g9978/_0_  ;
	output \g9979/_0_  ;
	output \g9980/_0_  ;
	output \g9981/_0_  ;
	output \g9982/_0_  ;
	output \g9983/_0_  ;
	output \g9984/_0_  ;
	output \g9985/_0_  ;
	output \g9987/_0_  ;
	output \g9988/_0_  ;
	output \g9989/_0_  ;
	output \g999/_0_  ;
	output \g9990/_0_  ;
	output \g9991/_0_  ;
	output \g9992/_0_  ;
	output \g9993/_0_  ;
	output \g9994/_0_  ;
	output \g9995/_0_  ;
	output \g9996/_0_  ;
	output \g9997/_0_  ;
	output \g9998/_0_  ;
	output \g9999/_0_  ;
	output \idma_IDMA_boot_reg/NET0131_reg_syn_3  ;
	output \memc_EXTC_Eg_reg/NET0131  ;
	output \memc_EXTC_Eg_reg/NET0131_reg_syn_3  ;
	output \memc_EXTC_Eg_reg/n0  ;
	output \pio_PIO_IN_P_reg[0]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[10]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[11]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[1]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[2]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[3]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[4]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[5]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[6]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[7]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[8]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[9]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[0]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[10]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[2]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[4]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[6]/P0001_reg_syn_3  ;
	output \sice_GO_NXi_reg/NET0131_reg_syn_3  ;
	output \sport0_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  ;
	output \sport0_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  ;
	output \sport1_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  ;
	output \sport1_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  ;
	wire _w23514_ ;
	wire _w23513_ ;
	wire _w23512_ ;
	wire _w23511_ ;
	wire _w23510_ ;
	wire _w23509_ ;
	wire _w23508_ ;
	wire _w23507_ ;
	wire _w23506_ ;
	wire _w23505_ ;
	wire _w23504_ ;
	wire _w23503_ ;
	wire _w23502_ ;
	wire _w23501_ ;
	wire _w23500_ ;
	wire _w23499_ ;
	wire _w23498_ ;
	wire _w23497_ ;
	wire _w23496_ ;
	wire _w23495_ ;
	wire _w23494_ ;
	wire _w23493_ ;
	wire _w23492_ ;
	wire _w23491_ ;
	wire _w23490_ ;
	wire _w23489_ ;
	wire _w23488_ ;
	wire _w23487_ ;
	wire _w23486_ ;
	wire _w23485_ ;
	wire _w23484_ ;
	wire _w23483_ ;
	wire _w23482_ ;
	wire _w23481_ ;
	wire _w23480_ ;
	wire _w23479_ ;
	wire _w23478_ ;
	wire _w23477_ ;
	wire _w23476_ ;
	wire _w23475_ ;
	wire _w23474_ ;
	wire _w23473_ ;
	wire _w23472_ ;
	wire _w23471_ ;
	wire _w23470_ ;
	wire _w23469_ ;
	wire _w23468_ ;
	wire _w23467_ ;
	wire _w23466_ ;
	wire _w23465_ ;
	wire _w23464_ ;
	wire _w23463_ ;
	wire _w23462_ ;
	wire _w23461_ ;
	wire _w23460_ ;
	wire _w23459_ ;
	wire _w23458_ ;
	wire _w23457_ ;
	wire _w23456_ ;
	wire _w23455_ ;
	wire _w23454_ ;
	wire _w23453_ ;
	wire _w23452_ ;
	wire _w23451_ ;
	wire _w23450_ ;
	wire _w23449_ ;
	wire _w23448_ ;
	wire _w23447_ ;
	wire _w23446_ ;
	wire _w23445_ ;
	wire _w23444_ ;
	wire _w23443_ ;
	wire _w23442_ ;
	wire _w23441_ ;
	wire _w23440_ ;
	wire _w23439_ ;
	wire _w23438_ ;
	wire _w23437_ ;
	wire _w23436_ ;
	wire _w23435_ ;
	wire _w23434_ ;
	wire _w23433_ ;
	wire _w23432_ ;
	wire _w23431_ ;
	wire _w23430_ ;
	wire _w23429_ ;
	wire _w23428_ ;
	wire _w23427_ ;
	wire _w23426_ ;
	wire _w23425_ ;
	wire _w23424_ ;
	wire _w23423_ ;
	wire _w23422_ ;
	wire _w23421_ ;
	wire _w23420_ ;
	wire _w23419_ ;
	wire _w23418_ ;
	wire _w23417_ ;
	wire _w23416_ ;
	wire _w23415_ ;
	wire _w23414_ ;
	wire _w23413_ ;
	wire _w23412_ ;
	wire _w23411_ ;
	wire _w23410_ ;
	wire _w23409_ ;
	wire _w23408_ ;
	wire _w23407_ ;
	wire _w23406_ ;
	wire _w23405_ ;
	wire _w23404_ ;
	wire _w23403_ ;
	wire _w23402_ ;
	wire _w23401_ ;
	wire _w23400_ ;
	wire _w23399_ ;
	wire _w23398_ ;
	wire _w23397_ ;
	wire _w23396_ ;
	wire _w23395_ ;
	wire _w23394_ ;
	wire _w23393_ ;
	wire _w23392_ ;
	wire _w23391_ ;
	wire _w23390_ ;
	wire _w23389_ ;
	wire _w23388_ ;
	wire _w23387_ ;
	wire _w23386_ ;
	wire _w23385_ ;
	wire _w23384_ ;
	wire _w23383_ ;
	wire _w23382_ ;
	wire _w23381_ ;
	wire _w23380_ ;
	wire _w23379_ ;
	wire _w23378_ ;
	wire _w23377_ ;
	wire _w23376_ ;
	wire _w23375_ ;
	wire _w23374_ ;
	wire _w23373_ ;
	wire _w23372_ ;
	wire _w23371_ ;
	wire _w23370_ ;
	wire _w23369_ ;
	wire _w23368_ ;
	wire _w23367_ ;
	wire _w23366_ ;
	wire _w23365_ ;
	wire _w23364_ ;
	wire _w23363_ ;
	wire _w23362_ ;
	wire _w23361_ ;
	wire _w23360_ ;
	wire _w23359_ ;
	wire _w23358_ ;
	wire _w23357_ ;
	wire _w23356_ ;
	wire _w23355_ ;
	wire _w23354_ ;
	wire _w23353_ ;
	wire _w23352_ ;
	wire _w23351_ ;
	wire _w23350_ ;
	wire _w23349_ ;
	wire _w23348_ ;
	wire _w23347_ ;
	wire _w23346_ ;
	wire _w23345_ ;
	wire _w23344_ ;
	wire _w23343_ ;
	wire _w23342_ ;
	wire _w23341_ ;
	wire _w23340_ ;
	wire _w23339_ ;
	wire _w23338_ ;
	wire _w23337_ ;
	wire _w23336_ ;
	wire _w23335_ ;
	wire _w23334_ ;
	wire _w23333_ ;
	wire _w23332_ ;
	wire _w23331_ ;
	wire _w23330_ ;
	wire _w23329_ ;
	wire _w23328_ ;
	wire _w23327_ ;
	wire _w23326_ ;
	wire _w23325_ ;
	wire _w23324_ ;
	wire _w23323_ ;
	wire _w23322_ ;
	wire _w23321_ ;
	wire _w23320_ ;
	wire _w23319_ ;
	wire _w23318_ ;
	wire _w23317_ ;
	wire _w23316_ ;
	wire _w23315_ ;
	wire _w23314_ ;
	wire _w23313_ ;
	wire _w23312_ ;
	wire _w23311_ ;
	wire _w23310_ ;
	wire _w23309_ ;
	wire _w23308_ ;
	wire _w23307_ ;
	wire _w23306_ ;
	wire _w23305_ ;
	wire _w23304_ ;
	wire _w23303_ ;
	wire _w23302_ ;
	wire _w23301_ ;
	wire _w23300_ ;
	wire _w23299_ ;
	wire _w23298_ ;
	wire _w23297_ ;
	wire _w23296_ ;
	wire _w23295_ ;
	wire _w23294_ ;
	wire _w23293_ ;
	wire _w23292_ ;
	wire _w23291_ ;
	wire _w23290_ ;
	wire _w23289_ ;
	wire _w23288_ ;
	wire _w23287_ ;
	wire _w23286_ ;
	wire _w23285_ ;
	wire _w23284_ ;
	wire _w23283_ ;
	wire _w23282_ ;
	wire _w23281_ ;
	wire _w23280_ ;
	wire _w23279_ ;
	wire _w23278_ ;
	wire _w23277_ ;
	wire _w23276_ ;
	wire _w23275_ ;
	wire _w23274_ ;
	wire _w23273_ ;
	wire _w23272_ ;
	wire _w23271_ ;
	wire _w23270_ ;
	wire _w23269_ ;
	wire _w23268_ ;
	wire _w23267_ ;
	wire _w23266_ ;
	wire _w23265_ ;
	wire _w23264_ ;
	wire _w23263_ ;
	wire _w23262_ ;
	wire _w23261_ ;
	wire _w23260_ ;
	wire _w23259_ ;
	wire _w23258_ ;
	wire _w23257_ ;
	wire _w23256_ ;
	wire _w23255_ ;
	wire _w23254_ ;
	wire _w23253_ ;
	wire _w23252_ ;
	wire _w23251_ ;
	wire _w23250_ ;
	wire _w23249_ ;
	wire _w23248_ ;
	wire _w23247_ ;
	wire _w23246_ ;
	wire _w23245_ ;
	wire _w23244_ ;
	wire _w23243_ ;
	wire _w23242_ ;
	wire _w23241_ ;
	wire _w23240_ ;
	wire _w23239_ ;
	wire _w23238_ ;
	wire _w23237_ ;
	wire _w23236_ ;
	wire _w23235_ ;
	wire _w23234_ ;
	wire _w23233_ ;
	wire _w23232_ ;
	wire _w23231_ ;
	wire _w23230_ ;
	wire _w23229_ ;
	wire _w23228_ ;
	wire _w23227_ ;
	wire _w23226_ ;
	wire _w23225_ ;
	wire _w23224_ ;
	wire _w23223_ ;
	wire _w23222_ ;
	wire _w23221_ ;
	wire _w23220_ ;
	wire _w23219_ ;
	wire _w23218_ ;
	wire _w23217_ ;
	wire _w23216_ ;
	wire _w23215_ ;
	wire _w23214_ ;
	wire _w23213_ ;
	wire _w23212_ ;
	wire _w23211_ ;
	wire _w23210_ ;
	wire _w23209_ ;
	wire _w23208_ ;
	wire _w23207_ ;
	wire _w23206_ ;
	wire _w23205_ ;
	wire _w23204_ ;
	wire _w23203_ ;
	wire _w23202_ ;
	wire _w23201_ ;
	wire _w23200_ ;
	wire _w23199_ ;
	wire _w23198_ ;
	wire _w23197_ ;
	wire _w23196_ ;
	wire _w23195_ ;
	wire _w23194_ ;
	wire _w23193_ ;
	wire _w23192_ ;
	wire _w23191_ ;
	wire _w23190_ ;
	wire _w23189_ ;
	wire _w23188_ ;
	wire _w23187_ ;
	wire _w23186_ ;
	wire _w23185_ ;
	wire _w23184_ ;
	wire _w23183_ ;
	wire _w23182_ ;
	wire _w23181_ ;
	wire _w23180_ ;
	wire _w23179_ ;
	wire _w23178_ ;
	wire _w23177_ ;
	wire _w23176_ ;
	wire _w23175_ ;
	wire _w23174_ ;
	wire _w23173_ ;
	wire _w23172_ ;
	wire _w23171_ ;
	wire _w23170_ ;
	wire _w23169_ ;
	wire _w23168_ ;
	wire _w23167_ ;
	wire _w23166_ ;
	wire _w23165_ ;
	wire _w23164_ ;
	wire _w23163_ ;
	wire _w23162_ ;
	wire _w23161_ ;
	wire _w23160_ ;
	wire _w23159_ ;
	wire _w23158_ ;
	wire _w23157_ ;
	wire _w23156_ ;
	wire _w23155_ ;
	wire _w23154_ ;
	wire _w23153_ ;
	wire _w23152_ ;
	wire _w23151_ ;
	wire _w23150_ ;
	wire _w23149_ ;
	wire _w23148_ ;
	wire _w23147_ ;
	wire _w23146_ ;
	wire _w23145_ ;
	wire _w23144_ ;
	wire _w23143_ ;
	wire _w23142_ ;
	wire _w23141_ ;
	wire _w23140_ ;
	wire _w23139_ ;
	wire _w23138_ ;
	wire _w23137_ ;
	wire _w23136_ ;
	wire _w23135_ ;
	wire _w23134_ ;
	wire _w23133_ ;
	wire _w23132_ ;
	wire _w23131_ ;
	wire _w23130_ ;
	wire _w23129_ ;
	wire _w23128_ ;
	wire _w23127_ ;
	wire _w23126_ ;
	wire _w23125_ ;
	wire _w23124_ ;
	wire _w23123_ ;
	wire _w23122_ ;
	wire _w23121_ ;
	wire _w23120_ ;
	wire _w23119_ ;
	wire _w23118_ ;
	wire _w23117_ ;
	wire _w23116_ ;
	wire _w23115_ ;
	wire _w23114_ ;
	wire _w23113_ ;
	wire _w23112_ ;
	wire _w23111_ ;
	wire _w23110_ ;
	wire _w23109_ ;
	wire _w23108_ ;
	wire _w23107_ ;
	wire _w23106_ ;
	wire _w23105_ ;
	wire _w23104_ ;
	wire _w23103_ ;
	wire _w23102_ ;
	wire _w23101_ ;
	wire _w23100_ ;
	wire _w23099_ ;
	wire _w23098_ ;
	wire _w23097_ ;
	wire _w23096_ ;
	wire _w23095_ ;
	wire _w23094_ ;
	wire _w23093_ ;
	wire _w23092_ ;
	wire _w23091_ ;
	wire _w23090_ ;
	wire _w23089_ ;
	wire _w23088_ ;
	wire _w23087_ ;
	wire _w23086_ ;
	wire _w23085_ ;
	wire _w23084_ ;
	wire _w23083_ ;
	wire _w23082_ ;
	wire _w23081_ ;
	wire _w23080_ ;
	wire _w23079_ ;
	wire _w23078_ ;
	wire _w23077_ ;
	wire _w23076_ ;
	wire _w23075_ ;
	wire _w23074_ ;
	wire _w23073_ ;
	wire _w23072_ ;
	wire _w23071_ ;
	wire _w23070_ ;
	wire _w23069_ ;
	wire _w23068_ ;
	wire _w23067_ ;
	wire _w23066_ ;
	wire _w23065_ ;
	wire _w23064_ ;
	wire _w23063_ ;
	wire _w23062_ ;
	wire _w23061_ ;
	wire _w23060_ ;
	wire _w23059_ ;
	wire _w23058_ ;
	wire _w23057_ ;
	wire _w23056_ ;
	wire _w23055_ ;
	wire _w23054_ ;
	wire _w23053_ ;
	wire _w23052_ ;
	wire _w23051_ ;
	wire _w23050_ ;
	wire _w23049_ ;
	wire _w23048_ ;
	wire _w23047_ ;
	wire _w23046_ ;
	wire _w23045_ ;
	wire _w23044_ ;
	wire _w23043_ ;
	wire _w23042_ ;
	wire _w23041_ ;
	wire _w23040_ ;
	wire _w23039_ ;
	wire _w23038_ ;
	wire _w23037_ ;
	wire _w23036_ ;
	wire _w23035_ ;
	wire _w23034_ ;
	wire _w23033_ ;
	wire _w23032_ ;
	wire _w23031_ ;
	wire _w23030_ ;
	wire _w23029_ ;
	wire _w23028_ ;
	wire _w23027_ ;
	wire _w23026_ ;
	wire _w23025_ ;
	wire _w23024_ ;
	wire _w23023_ ;
	wire _w23022_ ;
	wire _w23021_ ;
	wire _w23020_ ;
	wire _w23019_ ;
	wire _w23018_ ;
	wire _w23017_ ;
	wire _w23016_ ;
	wire _w23015_ ;
	wire _w23014_ ;
	wire _w23013_ ;
	wire _w23012_ ;
	wire _w23011_ ;
	wire _w23010_ ;
	wire _w23009_ ;
	wire _w23008_ ;
	wire _w23007_ ;
	wire _w23006_ ;
	wire _w23005_ ;
	wire _w23004_ ;
	wire _w23003_ ;
	wire _w23002_ ;
	wire _w23001_ ;
	wire _w23000_ ;
	wire _w22999_ ;
	wire _w22998_ ;
	wire _w22997_ ;
	wire _w22996_ ;
	wire _w22995_ ;
	wire _w22994_ ;
	wire _w22993_ ;
	wire _w22992_ ;
	wire _w22991_ ;
	wire _w22990_ ;
	wire _w22989_ ;
	wire _w22988_ ;
	wire _w22987_ ;
	wire _w22986_ ;
	wire _w22985_ ;
	wire _w22984_ ;
	wire _w22983_ ;
	wire _w22982_ ;
	wire _w22981_ ;
	wire _w22980_ ;
	wire _w22979_ ;
	wire _w22978_ ;
	wire _w22977_ ;
	wire _w22976_ ;
	wire _w22975_ ;
	wire _w22974_ ;
	wire _w22973_ ;
	wire _w22972_ ;
	wire _w22971_ ;
	wire _w22970_ ;
	wire _w22969_ ;
	wire _w22968_ ;
	wire _w22967_ ;
	wire _w22966_ ;
	wire _w22965_ ;
	wire _w22964_ ;
	wire _w22963_ ;
	wire _w22962_ ;
	wire _w22961_ ;
	wire _w22960_ ;
	wire _w22959_ ;
	wire _w22958_ ;
	wire _w22957_ ;
	wire _w22956_ ;
	wire _w22955_ ;
	wire _w22954_ ;
	wire _w22953_ ;
	wire _w22952_ ;
	wire _w22951_ ;
	wire _w22950_ ;
	wire _w22949_ ;
	wire _w22948_ ;
	wire _w22947_ ;
	wire _w22946_ ;
	wire _w22945_ ;
	wire _w22944_ ;
	wire _w22943_ ;
	wire _w22942_ ;
	wire _w22941_ ;
	wire _w22940_ ;
	wire _w22939_ ;
	wire _w22938_ ;
	wire _w22937_ ;
	wire _w22936_ ;
	wire _w22935_ ;
	wire _w22934_ ;
	wire _w22933_ ;
	wire _w22932_ ;
	wire _w22931_ ;
	wire _w22930_ ;
	wire _w22929_ ;
	wire _w22928_ ;
	wire _w22927_ ;
	wire _w22926_ ;
	wire _w22925_ ;
	wire _w22924_ ;
	wire _w22923_ ;
	wire _w22922_ ;
	wire _w22921_ ;
	wire _w22920_ ;
	wire _w22919_ ;
	wire _w22918_ ;
	wire _w22917_ ;
	wire _w22916_ ;
	wire _w22915_ ;
	wire _w22914_ ;
	wire _w22913_ ;
	wire _w22912_ ;
	wire _w22911_ ;
	wire _w22910_ ;
	wire _w22909_ ;
	wire _w22908_ ;
	wire _w22907_ ;
	wire _w22906_ ;
	wire _w22905_ ;
	wire _w22904_ ;
	wire _w22903_ ;
	wire _w22902_ ;
	wire _w22901_ ;
	wire _w22900_ ;
	wire _w22899_ ;
	wire _w22898_ ;
	wire _w22897_ ;
	wire _w22896_ ;
	wire _w22895_ ;
	wire _w22894_ ;
	wire _w22893_ ;
	wire _w22892_ ;
	wire _w22891_ ;
	wire _w22890_ ;
	wire _w22889_ ;
	wire _w22888_ ;
	wire _w22887_ ;
	wire _w22886_ ;
	wire _w22885_ ;
	wire _w22884_ ;
	wire _w22883_ ;
	wire _w22882_ ;
	wire _w22881_ ;
	wire _w22880_ ;
	wire _w22879_ ;
	wire _w22878_ ;
	wire _w22877_ ;
	wire _w22876_ ;
	wire _w22875_ ;
	wire _w22874_ ;
	wire _w22873_ ;
	wire _w22872_ ;
	wire _w22871_ ;
	wire _w22870_ ;
	wire _w22869_ ;
	wire _w22868_ ;
	wire _w22867_ ;
	wire _w22866_ ;
	wire _w22865_ ;
	wire _w22864_ ;
	wire _w22863_ ;
	wire _w22862_ ;
	wire _w22861_ ;
	wire _w22860_ ;
	wire _w22859_ ;
	wire _w22858_ ;
	wire _w22857_ ;
	wire _w22856_ ;
	wire _w22855_ ;
	wire _w22854_ ;
	wire _w22853_ ;
	wire _w22852_ ;
	wire _w22851_ ;
	wire _w22850_ ;
	wire _w22849_ ;
	wire _w22848_ ;
	wire _w22847_ ;
	wire _w22846_ ;
	wire _w22845_ ;
	wire _w22844_ ;
	wire _w22843_ ;
	wire _w22842_ ;
	wire _w22841_ ;
	wire _w22840_ ;
	wire _w22839_ ;
	wire _w22838_ ;
	wire _w22837_ ;
	wire _w22836_ ;
	wire _w22835_ ;
	wire _w22834_ ;
	wire _w22833_ ;
	wire _w22832_ ;
	wire _w22831_ ;
	wire _w22830_ ;
	wire _w22829_ ;
	wire _w22828_ ;
	wire _w22827_ ;
	wire _w22826_ ;
	wire _w22825_ ;
	wire _w22824_ ;
	wire _w22823_ ;
	wire _w22822_ ;
	wire _w22821_ ;
	wire _w22820_ ;
	wire _w22819_ ;
	wire _w22818_ ;
	wire _w22817_ ;
	wire _w22816_ ;
	wire _w22815_ ;
	wire _w22814_ ;
	wire _w22813_ ;
	wire _w22812_ ;
	wire _w22811_ ;
	wire _w22810_ ;
	wire _w22809_ ;
	wire _w22808_ ;
	wire _w22807_ ;
	wire _w22806_ ;
	wire _w22805_ ;
	wire _w22804_ ;
	wire _w22803_ ;
	wire _w22802_ ;
	wire _w22801_ ;
	wire _w22800_ ;
	wire _w22799_ ;
	wire _w22798_ ;
	wire _w22797_ ;
	wire _w22796_ ;
	wire _w22795_ ;
	wire _w22794_ ;
	wire _w22793_ ;
	wire _w22792_ ;
	wire _w22791_ ;
	wire _w22790_ ;
	wire _w22789_ ;
	wire _w22788_ ;
	wire _w22787_ ;
	wire _w22786_ ;
	wire _w22785_ ;
	wire _w22784_ ;
	wire _w22783_ ;
	wire _w22782_ ;
	wire _w22781_ ;
	wire _w22780_ ;
	wire _w22779_ ;
	wire _w22778_ ;
	wire _w22777_ ;
	wire _w22776_ ;
	wire _w22775_ ;
	wire _w22774_ ;
	wire _w22773_ ;
	wire _w22772_ ;
	wire _w22771_ ;
	wire _w22770_ ;
	wire _w22769_ ;
	wire _w22768_ ;
	wire _w22767_ ;
	wire _w22766_ ;
	wire _w22765_ ;
	wire _w22764_ ;
	wire _w22763_ ;
	wire _w22762_ ;
	wire _w22761_ ;
	wire _w22760_ ;
	wire _w22759_ ;
	wire _w22758_ ;
	wire _w22757_ ;
	wire _w22756_ ;
	wire _w22755_ ;
	wire _w22754_ ;
	wire _w22753_ ;
	wire _w22752_ ;
	wire _w22751_ ;
	wire _w22750_ ;
	wire _w22749_ ;
	wire _w22748_ ;
	wire _w22747_ ;
	wire _w22746_ ;
	wire _w22745_ ;
	wire _w22744_ ;
	wire _w22743_ ;
	wire _w22742_ ;
	wire _w22741_ ;
	wire _w22740_ ;
	wire _w22739_ ;
	wire _w22738_ ;
	wire _w22737_ ;
	wire _w22736_ ;
	wire _w22735_ ;
	wire _w22734_ ;
	wire _w22733_ ;
	wire _w22732_ ;
	wire _w22731_ ;
	wire _w22730_ ;
	wire _w22729_ ;
	wire _w22728_ ;
	wire _w22727_ ;
	wire _w22726_ ;
	wire _w22725_ ;
	wire _w22724_ ;
	wire _w22723_ ;
	wire _w22722_ ;
	wire _w22721_ ;
	wire _w22720_ ;
	wire _w22719_ ;
	wire _w22718_ ;
	wire _w22717_ ;
	wire _w22716_ ;
	wire _w22715_ ;
	wire _w22714_ ;
	wire _w22713_ ;
	wire _w22712_ ;
	wire _w22711_ ;
	wire _w22710_ ;
	wire _w22709_ ;
	wire _w22708_ ;
	wire _w22707_ ;
	wire _w22706_ ;
	wire _w22705_ ;
	wire _w22704_ ;
	wire _w22703_ ;
	wire _w22702_ ;
	wire _w22701_ ;
	wire _w22700_ ;
	wire _w22699_ ;
	wire _w22698_ ;
	wire _w22697_ ;
	wire _w22696_ ;
	wire _w22695_ ;
	wire _w22694_ ;
	wire _w22693_ ;
	wire _w22692_ ;
	wire _w22691_ ;
	wire _w22690_ ;
	wire _w22689_ ;
	wire _w22688_ ;
	wire _w22687_ ;
	wire _w22686_ ;
	wire _w22685_ ;
	wire _w22684_ ;
	wire _w22683_ ;
	wire _w22682_ ;
	wire _w22681_ ;
	wire _w22680_ ;
	wire _w22679_ ;
	wire _w22678_ ;
	wire _w22677_ ;
	wire _w22676_ ;
	wire _w22675_ ;
	wire _w22674_ ;
	wire _w22673_ ;
	wire _w22672_ ;
	wire _w22671_ ;
	wire _w22670_ ;
	wire _w22669_ ;
	wire _w22668_ ;
	wire _w22667_ ;
	wire _w22666_ ;
	wire _w22665_ ;
	wire _w22664_ ;
	wire _w22663_ ;
	wire _w22662_ ;
	wire _w22661_ ;
	wire _w22660_ ;
	wire _w22659_ ;
	wire _w22658_ ;
	wire _w22657_ ;
	wire _w22656_ ;
	wire _w22655_ ;
	wire _w22654_ ;
	wire _w22653_ ;
	wire _w22652_ ;
	wire _w22651_ ;
	wire _w22650_ ;
	wire _w22649_ ;
	wire _w22648_ ;
	wire _w22647_ ;
	wire _w22646_ ;
	wire _w22645_ ;
	wire _w22644_ ;
	wire _w22643_ ;
	wire _w22642_ ;
	wire _w22641_ ;
	wire _w22640_ ;
	wire _w22639_ ;
	wire _w22638_ ;
	wire _w22637_ ;
	wire _w22636_ ;
	wire _w22635_ ;
	wire _w22634_ ;
	wire _w22633_ ;
	wire _w22632_ ;
	wire _w22631_ ;
	wire _w22630_ ;
	wire _w22629_ ;
	wire _w22628_ ;
	wire _w22627_ ;
	wire _w22626_ ;
	wire _w22625_ ;
	wire _w22624_ ;
	wire _w22623_ ;
	wire _w22622_ ;
	wire _w22621_ ;
	wire _w22620_ ;
	wire _w22619_ ;
	wire _w22618_ ;
	wire _w22617_ ;
	wire _w22616_ ;
	wire _w22615_ ;
	wire _w22614_ ;
	wire _w22613_ ;
	wire _w22612_ ;
	wire _w22611_ ;
	wire _w22610_ ;
	wire _w22609_ ;
	wire _w22608_ ;
	wire _w22607_ ;
	wire _w22606_ ;
	wire _w22605_ ;
	wire _w22604_ ;
	wire _w22603_ ;
	wire _w22602_ ;
	wire _w22601_ ;
	wire _w22600_ ;
	wire _w22599_ ;
	wire _w22598_ ;
	wire _w22597_ ;
	wire _w22596_ ;
	wire _w22595_ ;
	wire _w22594_ ;
	wire _w22593_ ;
	wire _w22592_ ;
	wire _w22591_ ;
	wire _w22590_ ;
	wire _w22589_ ;
	wire _w22588_ ;
	wire _w22587_ ;
	wire _w22586_ ;
	wire _w22585_ ;
	wire _w22584_ ;
	wire _w22583_ ;
	wire _w22582_ ;
	wire _w22581_ ;
	wire _w22580_ ;
	wire _w22579_ ;
	wire _w22578_ ;
	wire _w22577_ ;
	wire _w22576_ ;
	wire _w22575_ ;
	wire _w22574_ ;
	wire _w22573_ ;
	wire _w22572_ ;
	wire _w22571_ ;
	wire _w22570_ ;
	wire _w22569_ ;
	wire _w22568_ ;
	wire _w22567_ ;
	wire _w22566_ ;
	wire _w22565_ ;
	wire _w22564_ ;
	wire _w22563_ ;
	wire _w22562_ ;
	wire _w22561_ ;
	wire _w22560_ ;
	wire _w22559_ ;
	wire _w22558_ ;
	wire _w22557_ ;
	wire _w22556_ ;
	wire _w22555_ ;
	wire _w22554_ ;
	wire _w22553_ ;
	wire _w22552_ ;
	wire _w22551_ ;
	wire _w22550_ ;
	wire _w22549_ ;
	wire _w22548_ ;
	wire _w22547_ ;
	wire _w22546_ ;
	wire _w22545_ ;
	wire _w22544_ ;
	wire _w22543_ ;
	wire _w22542_ ;
	wire _w22541_ ;
	wire _w22540_ ;
	wire _w22539_ ;
	wire _w22538_ ;
	wire _w22537_ ;
	wire _w22536_ ;
	wire _w22535_ ;
	wire _w22534_ ;
	wire _w22533_ ;
	wire _w22532_ ;
	wire _w22531_ ;
	wire _w22530_ ;
	wire _w22529_ ;
	wire _w22528_ ;
	wire _w22527_ ;
	wire _w22526_ ;
	wire _w22525_ ;
	wire _w22524_ ;
	wire _w22523_ ;
	wire _w22522_ ;
	wire _w22521_ ;
	wire _w22520_ ;
	wire _w22519_ ;
	wire _w22518_ ;
	wire _w22517_ ;
	wire _w22516_ ;
	wire _w22515_ ;
	wire _w22514_ ;
	wire _w22513_ ;
	wire _w22512_ ;
	wire _w22511_ ;
	wire _w22510_ ;
	wire _w22509_ ;
	wire _w22508_ ;
	wire _w22507_ ;
	wire _w22506_ ;
	wire _w22505_ ;
	wire _w22504_ ;
	wire _w22503_ ;
	wire _w22502_ ;
	wire _w22501_ ;
	wire _w22500_ ;
	wire _w22499_ ;
	wire _w22498_ ;
	wire _w22497_ ;
	wire _w22496_ ;
	wire _w22495_ ;
	wire _w22494_ ;
	wire _w22493_ ;
	wire _w22492_ ;
	wire _w22491_ ;
	wire _w22490_ ;
	wire _w22489_ ;
	wire _w22488_ ;
	wire _w22487_ ;
	wire _w22486_ ;
	wire _w22485_ ;
	wire _w22484_ ;
	wire _w22483_ ;
	wire _w22482_ ;
	wire _w22481_ ;
	wire _w22480_ ;
	wire _w22479_ ;
	wire _w22478_ ;
	wire _w22477_ ;
	wire _w22476_ ;
	wire _w22475_ ;
	wire _w22474_ ;
	wire _w22473_ ;
	wire _w22472_ ;
	wire _w22471_ ;
	wire _w22470_ ;
	wire _w22469_ ;
	wire _w22468_ ;
	wire _w22467_ ;
	wire _w22466_ ;
	wire _w22465_ ;
	wire _w22464_ ;
	wire _w22463_ ;
	wire _w22462_ ;
	wire _w22461_ ;
	wire _w22460_ ;
	wire _w22459_ ;
	wire _w22458_ ;
	wire _w22457_ ;
	wire _w22456_ ;
	wire _w22455_ ;
	wire _w22454_ ;
	wire _w22453_ ;
	wire _w22452_ ;
	wire _w22451_ ;
	wire _w22450_ ;
	wire _w22449_ ;
	wire _w22448_ ;
	wire _w22447_ ;
	wire _w22446_ ;
	wire _w22445_ ;
	wire _w22444_ ;
	wire _w22443_ ;
	wire _w22442_ ;
	wire _w22441_ ;
	wire _w22440_ ;
	wire _w22439_ ;
	wire _w22438_ ;
	wire _w22437_ ;
	wire _w22436_ ;
	wire _w22435_ ;
	wire _w22434_ ;
	wire _w22433_ ;
	wire _w22432_ ;
	wire _w22431_ ;
	wire _w22430_ ;
	wire _w22429_ ;
	wire _w22428_ ;
	wire _w22427_ ;
	wire _w22426_ ;
	wire _w22425_ ;
	wire _w22424_ ;
	wire _w22423_ ;
	wire _w22422_ ;
	wire _w22421_ ;
	wire _w22420_ ;
	wire _w22419_ ;
	wire _w22418_ ;
	wire _w22417_ ;
	wire _w22416_ ;
	wire _w22415_ ;
	wire _w22414_ ;
	wire _w22413_ ;
	wire _w22412_ ;
	wire _w22411_ ;
	wire _w22410_ ;
	wire _w22409_ ;
	wire _w22408_ ;
	wire _w22407_ ;
	wire _w22406_ ;
	wire _w22405_ ;
	wire _w22404_ ;
	wire _w22403_ ;
	wire _w22402_ ;
	wire _w22401_ ;
	wire _w22400_ ;
	wire _w22399_ ;
	wire _w22398_ ;
	wire _w22397_ ;
	wire _w22396_ ;
	wire _w22395_ ;
	wire _w22394_ ;
	wire _w22393_ ;
	wire _w22392_ ;
	wire _w22391_ ;
	wire _w22390_ ;
	wire _w22389_ ;
	wire _w22388_ ;
	wire _w22387_ ;
	wire _w22386_ ;
	wire _w22385_ ;
	wire _w22384_ ;
	wire _w22383_ ;
	wire _w22382_ ;
	wire _w22381_ ;
	wire _w22380_ ;
	wire _w22379_ ;
	wire _w22378_ ;
	wire _w22377_ ;
	wire _w22376_ ;
	wire _w22375_ ;
	wire _w22374_ ;
	wire _w22373_ ;
	wire _w22372_ ;
	wire _w22371_ ;
	wire _w22370_ ;
	wire _w22369_ ;
	wire _w22368_ ;
	wire _w22367_ ;
	wire _w22366_ ;
	wire _w22365_ ;
	wire _w22364_ ;
	wire _w22363_ ;
	wire _w22362_ ;
	wire _w22361_ ;
	wire _w22360_ ;
	wire _w22359_ ;
	wire _w22358_ ;
	wire _w22357_ ;
	wire _w22356_ ;
	wire _w22355_ ;
	wire _w22354_ ;
	wire _w22353_ ;
	wire _w22352_ ;
	wire _w22351_ ;
	wire _w22350_ ;
	wire _w22349_ ;
	wire _w22348_ ;
	wire _w22347_ ;
	wire _w22346_ ;
	wire _w22345_ ;
	wire _w22344_ ;
	wire _w22343_ ;
	wire _w22342_ ;
	wire _w22341_ ;
	wire _w22340_ ;
	wire _w22339_ ;
	wire _w22338_ ;
	wire _w22337_ ;
	wire _w22336_ ;
	wire _w22335_ ;
	wire _w22334_ ;
	wire _w22333_ ;
	wire _w22332_ ;
	wire _w22331_ ;
	wire _w22330_ ;
	wire _w22329_ ;
	wire _w22328_ ;
	wire _w22327_ ;
	wire _w22326_ ;
	wire _w22325_ ;
	wire _w22324_ ;
	wire _w22323_ ;
	wire _w22322_ ;
	wire _w22321_ ;
	wire _w22320_ ;
	wire _w22319_ ;
	wire _w22318_ ;
	wire _w22317_ ;
	wire _w22316_ ;
	wire _w22315_ ;
	wire _w22314_ ;
	wire _w22313_ ;
	wire _w22312_ ;
	wire _w22311_ ;
	wire _w22310_ ;
	wire _w22309_ ;
	wire _w22308_ ;
	wire _w22307_ ;
	wire _w22306_ ;
	wire _w22305_ ;
	wire _w22304_ ;
	wire _w22303_ ;
	wire _w22302_ ;
	wire _w22301_ ;
	wire _w22300_ ;
	wire _w22299_ ;
	wire _w22298_ ;
	wire _w22297_ ;
	wire _w22296_ ;
	wire _w22295_ ;
	wire _w22294_ ;
	wire _w22293_ ;
	wire _w22292_ ;
	wire _w22291_ ;
	wire _w22290_ ;
	wire _w22289_ ;
	wire _w22288_ ;
	wire _w22287_ ;
	wire _w22286_ ;
	wire _w22285_ ;
	wire _w22284_ ;
	wire _w22283_ ;
	wire _w22282_ ;
	wire _w22281_ ;
	wire _w22280_ ;
	wire _w22279_ ;
	wire _w22278_ ;
	wire _w22277_ ;
	wire _w22276_ ;
	wire _w22275_ ;
	wire _w22274_ ;
	wire _w22273_ ;
	wire _w22272_ ;
	wire _w22271_ ;
	wire _w22270_ ;
	wire _w22269_ ;
	wire _w22268_ ;
	wire _w22267_ ;
	wire _w22266_ ;
	wire _w22265_ ;
	wire _w22264_ ;
	wire _w22263_ ;
	wire _w22262_ ;
	wire _w22261_ ;
	wire _w22260_ ;
	wire _w22259_ ;
	wire _w22258_ ;
	wire _w22257_ ;
	wire _w22256_ ;
	wire _w22255_ ;
	wire _w22254_ ;
	wire _w22253_ ;
	wire _w22252_ ;
	wire _w22251_ ;
	wire _w22250_ ;
	wire _w22249_ ;
	wire _w22248_ ;
	wire _w22247_ ;
	wire _w22246_ ;
	wire _w22245_ ;
	wire _w22244_ ;
	wire _w22243_ ;
	wire _w22242_ ;
	wire _w22241_ ;
	wire _w22240_ ;
	wire _w22239_ ;
	wire _w22238_ ;
	wire _w22237_ ;
	wire _w22236_ ;
	wire _w22235_ ;
	wire _w22234_ ;
	wire _w22233_ ;
	wire _w22232_ ;
	wire _w22231_ ;
	wire _w22230_ ;
	wire _w22229_ ;
	wire _w22228_ ;
	wire _w22227_ ;
	wire _w22226_ ;
	wire _w22225_ ;
	wire _w22224_ ;
	wire _w22223_ ;
	wire _w22222_ ;
	wire _w22221_ ;
	wire _w22220_ ;
	wire _w22219_ ;
	wire _w22218_ ;
	wire _w22217_ ;
	wire _w22216_ ;
	wire _w22215_ ;
	wire _w22214_ ;
	wire _w22213_ ;
	wire _w22212_ ;
	wire _w22211_ ;
	wire _w22210_ ;
	wire _w22209_ ;
	wire _w22208_ ;
	wire _w22207_ ;
	wire _w22206_ ;
	wire _w22205_ ;
	wire _w22204_ ;
	wire _w22203_ ;
	wire _w22202_ ;
	wire _w22201_ ;
	wire _w22200_ ;
	wire _w22199_ ;
	wire _w22198_ ;
	wire _w22197_ ;
	wire _w22196_ ;
	wire _w22195_ ;
	wire _w22194_ ;
	wire _w22193_ ;
	wire _w22192_ ;
	wire _w22191_ ;
	wire _w22190_ ;
	wire _w22189_ ;
	wire _w22188_ ;
	wire _w22187_ ;
	wire _w22186_ ;
	wire _w22185_ ;
	wire _w22184_ ;
	wire _w22183_ ;
	wire _w22182_ ;
	wire _w22181_ ;
	wire _w22180_ ;
	wire _w22179_ ;
	wire _w22178_ ;
	wire _w22177_ ;
	wire _w22176_ ;
	wire _w22175_ ;
	wire _w22174_ ;
	wire _w22173_ ;
	wire _w22172_ ;
	wire _w22171_ ;
	wire _w22170_ ;
	wire _w22169_ ;
	wire _w22168_ ;
	wire _w22167_ ;
	wire _w22166_ ;
	wire _w22165_ ;
	wire _w22164_ ;
	wire _w22163_ ;
	wire _w22162_ ;
	wire _w22161_ ;
	wire _w22160_ ;
	wire _w22159_ ;
	wire _w22158_ ;
	wire _w22157_ ;
	wire _w22156_ ;
	wire _w22155_ ;
	wire _w22154_ ;
	wire _w22153_ ;
	wire _w22152_ ;
	wire _w22151_ ;
	wire _w22150_ ;
	wire _w22149_ ;
	wire _w22148_ ;
	wire _w22147_ ;
	wire _w22146_ ;
	wire _w22145_ ;
	wire _w22144_ ;
	wire _w22143_ ;
	wire _w22142_ ;
	wire _w22141_ ;
	wire _w22140_ ;
	wire _w22139_ ;
	wire _w22138_ ;
	wire _w22137_ ;
	wire _w22136_ ;
	wire _w22135_ ;
	wire _w22134_ ;
	wire _w22133_ ;
	wire _w22132_ ;
	wire _w22131_ ;
	wire _w22130_ ;
	wire _w22129_ ;
	wire _w22128_ ;
	wire _w22127_ ;
	wire _w22126_ ;
	wire _w22125_ ;
	wire _w22124_ ;
	wire _w22123_ ;
	wire _w22122_ ;
	wire _w22121_ ;
	wire _w22120_ ;
	wire _w22119_ ;
	wire _w22118_ ;
	wire _w22117_ ;
	wire _w22116_ ;
	wire _w22115_ ;
	wire _w22114_ ;
	wire _w22113_ ;
	wire _w22112_ ;
	wire _w22111_ ;
	wire _w22110_ ;
	wire _w22109_ ;
	wire _w22108_ ;
	wire _w22107_ ;
	wire _w22106_ ;
	wire _w22105_ ;
	wire _w22104_ ;
	wire _w22103_ ;
	wire _w22102_ ;
	wire _w22101_ ;
	wire _w22100_ ;
	wire _w22099_ ;
	wire _w22098_ ;
	wire _w22097_ ;
	wire _w22096_ ;
	wire _w22095_ ;
	wire _w22094_ ;
	wire _w22093_ ;
	wire _w22092_ ;
	wire _w22091_ ;
	wire _w22090_ ;
	wire _w22089_ ;
	wire _w22088_ ;
	wire _w22087_ ;
	wire _w22086_ ;
	wire _w22085_ ;
	wire _w22084_ ;
	wire _w22083_ ;
	wire _w22082_ ;
	wire _w22081_ ;
	wire _w22080_ ;
	wire _w22079_ ;
	wire _w22078_ ;
	wire _w22077_ ;
	wire _w22076_ ;
	wire _w22075_ ;
	wire _w22074_ ;
	wire _w22073_ ;
	wire _w22072_ ;
	wire _w22071_ ;
	wire _w22070_ ;
	wire _w22069_ ;
	wire _w22068_ ;
	wire _w22067_ ;
	wire _w22066_ ;
	wire _w22065_ ;
	wire _w22064_ ;
	wire _w22063_ ;
	wire _w22062_ ;
	wire _w22061_ ;
	wire _w22060_ ;
	wire _w22059_ ;
	wire _w22058_ ;
	wire _w22057_ ;
	wire _w22056_ ;
	wire _w22055_ ;
	wire _w22054_ ;
	wire _w22053_ ;
	wire _w22052_ ;
	wire _w22051_ ;
	wire _w22050_ ;
	wire _w22049_ ;
	wire _w22048_ ;
	wire _w22047_ ;
	wire _w22046_ ;
	wire _w22045_ ;
	wire _w22044_ ;
	wire _w22043_ ;
	wire _w22042_ ;
	wire _w22041_ ;
	wire _w22040_ ;
	wire _w22039_ ;
	wire _w22038_ ;
	wire _w22037_ ;
	wire _w22036_ ;
	wire _w22035_ ;
	wire _w22034_ ;
	wire _w22033_ ;
	wire _w22032_ ;
	wire _w22031_ ;
	wire _w22030_ ;
	wire _w22029_ ;
	wire _w22028_ ;
	wire _w22027_ ;
	wire _w22026_ ;
	wire _w22025_ ;
	wire _w22024_ ;
	wire _w22023_ ;
	wire _w22022_ ;
	wire _w22021_ ;
	wire _w22020_ ;
	wire _w22019_ ;
	wire _w22018_ ;
	wire _w22017_ ;
	wire _w22016_ ;
	wire _w22015_ ;
	wire _w22014_ ;
	wire _w22013_ ;
	wire _w22012_ ;
	wire _w22011_ ;
	wire _w22010_ ;
	wire _w22009_ ;
	wire _w22008_ ;
	wire _w22007_ ;
	wire _w22006_ ;
	wire _w22005_ ;
	wire _w22004_ ;
	wire _w22003_ ;
	wire _w22002_ ;
	wire _w22001_ ;
	wire _w22000_ ;
	wire _w21999_ ;
	wire _w21998_ ;
	wire _w21997_ ;
	wire _w21996_ ;
	wire _w21995_ ;
	wire _w21994_ ;
	wire _w21993_ ;
	wire _w21992_ ;
	wire _w21991_ ;
	wire _w21990_ ;
	wire _w21989_ ;
	wire _w21988_ ;
	wire _w21987_ ;
	wire _w21986_ ;
	wire _w21985_ ;
	wire _w21984_ ;
	wire _w21983_ ;
	wire _w21982_ ;
	wire _w21981_ ;
	wire _w21980_ ;
	wire _w21979_ ;
	wire _w21978_ ;
	wire _w21977_ ;
	wire _w21976_ ;
	wire _w21975_ ;
	wire _w21974_ ;
	wire _w21973_ ;
	wire _w21972_ ;
	wire _w21971_ ;
	wire _w21970_ ;
	wire _w21969_ ;
	wire _w21968_ ;
	wire _w21967_ ;
	wire _w21966_ ;
	wire _w21965_ ;
	wire _w21964_ ;
	wire _w21963_ ;
	wire _w21962_ ;
	wire _w21961_ ;
	wire _w21960_ ;
	wire _w21959_ ;
	wire _w21958_ ;
	wire _w21957_ ;
	wire _w21956_ ;
	wire _w21955_ ;
	wire _w21954_ ;
	wire _w21953_ ;
	wire _w21952_ ;
	wire _w21951_ ;
	wire _w21950_ ;
	wire _w21949_ ;
	wire _w21948_ ;
	wire _w21947_ ;
	wire _w21946_ ;
	wire _w21945_ ;
	wire _w21944_ ;
	wire _w21943_ ;
	wire _w21942_ ;
	wire _w21941_ ;
	wire _w21940_ ;
	wire _w21939_ ;
	wire _w21938_ ;
	wire _w21937_ ;
	wire _w21936_ ;
	wire _w21935_ ;
	wire _w21934_ ;
	wire _w21933_ ;
	wire _w21932_ ;
	wire _w21931_ ;
	wire _w21930_ ;
	wire _w21929_ ;
	wire _w21928_ ;
	wire _w21927_ ;
	wire _w21926_ ;
	wire _w21925_ ;
	wire _w21924_ ;
	wire _w21923_ ;
	wire _w21922_ ;
	wire _w21921_ ;
	wire _w21920_ ;
	wire _w21919_ ;
	wire _w21918_ ;
	wire _w21917_ ;
	wire _w21916_ ;
	wire _w21915_ ;
	wire _w21914_ ;
	wire _w21913_ ;
	wire _w21912_ ;
	wire _w21911_ ;
	wire _w21910_ ;
	wire _w21909_ ;
	wire _w21908_ ;
	wire _w21907_ ;
	wire _w21906_ ;
	wire _w21905_ ;
	wire _w21904_ ;
	wire _w21903_ ;
	wire _w21902_ ;
	wire _w21901_ ;
	wire _w21900_ ;
	wire _w21899_ ;
	wire _w21898_ ;
	wire _w21897_ ;
	wire _w21896_ ;
	wire _w21895_ ;
	wire _w21894_ ;
	wire _w21893_ ;
	wire _w21892_ ;
	wire _w21891_ ;
	wire _w21889_ ;
	wire _w21888_ ;
	wire _w21887_ ;
	wire _w21886_ ;
	wire _w21885_ ;
	wire _w21884_ ;
	wire _w21883_ ;
	wire _w21882_ ;
	wire _w21881_ ;
	wire _w21880_ ;
	wire _w21879_ ;
	wire _w21878_ ;
	wire _w21877_ ;
	wire _w21876_ ;
	wire _w21875_ ;
	wire _w21874_ ;
	wire _w21873_ ;
	wire _w21872_ ;
	wire _w21871_ ;
	wire _w21870_ ;
	wire _w21869_ ;
	wire _w21868_ ;
	wire _w21867_ ;
	wire _w21866_ ;
	wire _w21865_ ;
	wire _w21864_ ;
	wire _w21863_ ;
	wire _w21862_ ;
	wire _w21861_ ;
	wire _w21860_ ;
	wire _w21859_ ;
	wire _w21858_ ;
	wire _w21857_ ;
	wire _w21856_ ;
	wire _w21855_ ;
	wire _w21854_ ;
	wire _w21853_ ;
	wire _w21852_ ;
	wire _w21851_ ;
	wire _w21850_ ;
	wire _w21849_ ;
	wire _w21848_ ;
	wire _w21847_ ;
	wire _w21846_ ;
	wire _w21845_ ;
	wire _w21844_ ;
	wire _w21843_ ;
	wire _w21842_ ;
	wire _w21841_ ;
	wire _w21840_ ;
	wire _w21839_ ;
	wire _w21838_ ;
	wire _w21837_ ;
	wire _w21836_ ;
	wire _w21835_ ;
	wire _w21834_ ;
	wire _w21833_ ;
	wire _w21832_ ;
	wire _w21831_ ;
	wire _w21830_ ;
	wire _w21829_ ;
	wire _w21828_ ;
	wire _w21827_ ;
	wire _w21826_ ;
	wire _w21825_ ;
	wire _w21824_ ;
	wire _w21823_ ;
	wire _w21822_ ;
	wire _w21821_ ;
	wire _w21820_ ;
	wire _w21819_ ;
	wire _w21818_ ;
	wire _w21817_ ;
	wire _w21816_ ;
	wire _w21815_ ;
	wire _w21814_ ;
	wire _w21813_ ;
	wire _w21812_ ;
	wire _w21811_ ;
	wire _w21810_ ;
	wire _w21809_ ;
	wire _w21808_ ;
	wire _w21807_ ;
	wire _w21806_ ;
	wire _w21805_ ;
	wire _w21804_ ;
	wire _w21803_ ;
	wire _w21802_ ;
	wire _w21801_ ;
	wire _w21800_ ;
	wire _w21799_ ;
	wire _w21798_ ;
	wire _w21797_ ;
	wire _w21796_ ;
	wire _w21795_ ;
	wire _w21794_ ;
	wire _w21793_ ;
	wire _w21792_ ;
	wire _w21791_ ;
	wire _w21790_ ;
	wire _w21789_ ;
	wire _w21788_ ;
	wire _w21787_ ;
	wire _w21786_ ;
	wire _w21785_ ;
	wire _w21784_ ;
	wire _w21783_ ;
	wire _w21782_ ;
	wire _w21781_ ;
	wire _w21780_ ;
	wire _w21779_ ;
	wire _w21778_ ;
	wire _w21777_ ;
	wire _w21776_ ;
	wire _w21775_ ;
	wire _w21774_ ;
	wire _w21773_ ;
	wire _w21772_ ;
	wire _w21771_ ;
	wire _w21770_ ;
	wire _w21769_ ;
	wire _w21768_ ;
	wire _w21767_ ;
	wire _w21766_ ;
	wire _w21765_ ;
	wire _w21764_ ;
	wire _w21763_ ;
	wire _w21762_ ;
	wire _w21761_ ;
	wire _w21760_ ;
	wire _w21759_ ;
	wire _w21758_ ;
	wire _w21757_ ;
	wire _w21756_ ;
	wire _w21755_ ;
	wire _w21754_ ;
	wire _w21753_ ;
	wire _w21752_ ;
	wire _w21751_ ;
	wire _w21750_ ;
	wire _w21749_ ;
	wire _w21748_ ;
	wire _w21747_ ;
	wire _w21746_ ;
	wire _w21745_ ;
	wire _w21744_ ;
	wire _w21743_ ;
	wire _w21742_ ;
	wire _w21741_ ;
	wire _w21740_ ;
	wire _w21739_ ;
	wire _w21738_ ;
	wire _w21737_ ;
	wire _w21736_ ;
	wire _w21735_ ;
	wire _w21734_ ;
	wire _w21733_ ;
	wire _w21732_ ;
	wire _w21731_ ;
	wire _w21730_ ;
	wire _w21729_ ;
	wire _w21728_ ;
	wire _w21727_ ;
	wire _w21726_ ;
	wire _w21725_ ;
	wire _w21724_ ;
	wire _w21723_ ;
	wire _w21722_ ;
	wire _w21721_ ;
	wire _w21720_ ;
	wire _w21719_ ;
	wire _w21718_ ;
	wire _w21717_ ;
	wire _w21716_ ;
	wire _w21715_ ;
	wire _w21714_ ;
	wire _w21713_ ;
	wire _w21712_ ;
	wire _w21711_ ;
	wire _w21710_ ;
	wire _w21709_ ;
	wire _w21708_ ;
	wire _w21707_ ;
	wire _w21706_ ;
	wire _w21705_ ;
	wire _w21704_ ;
	wire _w21703_ ;
	wire _w21702_ ;
	wire _w21701_ ;
	wire _w21700_ ;
	wire _w21699_ ;
	wire _w21698_ ;
	wire _w21697_ ;
	wire _w21696_ ;
	wire _w21695_ ;
	wire _w21694_ ;
	wire _w21693_ ;
	wire _w21692_ ;
	wire _w21691_ ;
	wire _w21690_ ;
	wire _w21689_ ;
	wire _w21688_ ;
	wire _w21687_ ;
	wire _w21686_ ;
	wire _w21685_ ;
	wire _w21684_ ;
	wire _w21683_ ;
	wire _w21682_ ;
	wire _w21681_ ;
	wire _w21680_ ;
	wire _w21679_ ;
	wire _w21678_ ;
	wire _w21677_ ;
	wire _w21676_ ;
	wire _w21675_ ;
	wire _w21674_ ;
	wire _w21673_ ;
	wire _w21672_ ;
	wire _w21671_ ;
	wire _w21670_ ;
	wire _w21669_ ;
	wire _w21668_ ;
	wire _w21667_ ;
	wire _w21666_ ;
	wire _w21665_ ;
	wire _w21664_ ;
	wire _w21663_ ;
	wire _w21662_ ;
	wire _w21661_ ;
	wire _w21660_ ;
	wire _w21659_ ;
	wire _w21658_ ;
	wire _w21657_ ;
	wire _w21656_ ;
	wire _w21655_ ;
	wire _w21654_ ;
	wire _w21653_ ;
	wire _w21652_ ;
	wire _w21651_ ;
	wire _w21650_ ;
	wire _w21649_ ;
	wire _w21648_ ;
	wire _w21647_ ;
	wire _w21646_ ;
	wire _w21645_ ;
	wire _w21644_ ;
	wire _w21643_ ;
	wire _w21642_ ;
	wire _w21641_ ;
	wire _w21640_ ;
	wire _w21639_ ;
	wire _w21638_ ;
	wire _w21637_ ;
	wire _w21636_ ;
	wire _w21635_ ;
	wire _w21634_ ;
	wire _w21633_ ;
	wire _w21632_ ;
	wire _w21631_ ;
	wire _w21630_ ;
	wire _w21629_ ;
	wire _w21628_ ;
	wire _w21627_ ;
	wire _w21626_ ;
	wire _w21625_ ;
	wire _w21624_ ;
	wire _w21623_ ;
	wire _w21622_ ;
	wire _w21621_ ;
	wire _w21620_ ;
	wire _w21619_ ;
	wire _w21618_ ;
	wire _w21617_ ;
	wire _w21616_ ;
	wire _w21615_ ;
	wire _w21614_ ;
	wire _w21613_ ;
	wire _w21612_ ;
	wire _w21611_ ;
	wire _w21610_ ;
	wire _w21609_ ;
	wire _w21608_ ;
	wire _w21607_ ;
	wire _w21606_ ;
	wire _w21605_ ;
	wire _w21604_ ;
	wire _w21603_ ;
	wire _w21602_ ;
	wire _w21601_ ;
	wire _w21600_ ;
	wire _w21599_ ;
	wire _w21598_ ;
	wire _w21597_ ;
	wire _w21596_ ;
	wire _w21595_ ;
	wire _w21594_ ;
	wire _w21593_ ;
	wire _w21592_ ;
	wire _w21591_ ;
	wire _w21590_ ;
	wire _w21589_ ;
	wire _w21588_ ;
	wire _w21587_ ;
	wire _w21586_ ;
	wire _w21585_ ;
	wire _w21584_ ;
	wire _w21583_ ;
	wire _w21582_ ;
	wire _w21581_ ;
	wire _w21580_ ;
	wire _w21579_ ;
	wire _w21578_ ;
	wire _w21577_ ;
	wire _w21576_ ;
	wire _w21575_ ;
	wire _w21574_ ;
	wire _w21573_ ;
	wire _w21572_ ;
	wire _w21571_ ;
	wire _w21570_ ;
	wire _w21569_ ;
	wire _w21568_ ;
	wire _w21567_ ;
	wire _w21566_ ;
	wire _w21565_ ;
	wire _w21564_ ;
	wire _w21563_ ;
	wire _w21562_ ;
	wire _w21561_ ;
	wire _w21560_ ;
	wire _w21559_ ;
	wire _w21558_ ;
	wire _w21557_ ;
	wire _w21556_ ;
	wire _w21555_ ;
	wire _w21554_ ;
	wire _w21553_ ;
	wire _w21552_ ;
	wire _w21551_ ;
	wire _w21550_ ;
	wire _w21549_ ;
	wire _w21548_ ;
	wire _w21547_ ;
	wire _w21546_ ;
	wire _w21545_ ;
	wire _w21544_ ;
	wire _w21543_ ;
	wire _w21542_ ;
	wire _w21541_ ;
	wire _w21540_ ;
	wire _w21539_ ;
	wire _w21538_ ;
	wire _w21537_ ;
	wire _w21536_ ;
	wire _w21535_ ;
	wire _w21534_ ;
	wire _w21533_ ;
	wire _w21532_ ;
	wire _w21531_ ;
	wire _w21530_ ;
	wire _w21529_ ;
	wire _w21528_ ;
	wire _w21527_ ;
	wire _w21526_ ;
	wire _w21525_ ;
	wire _w21524_ ;
	wire _w21523_ ;
	wire _w21522_ ;
	wire _w21521_ ;
	wire _w21520_ ;
	wire _w21519_ ;
	wire _w21518_ ;
	wire _w21517_ ;
	wire _w21516_ ;
	wire _w21515_ ;
	wire _w21514_ ;
	wire _w21513_ ;
	wire _w21512_ ;
	wire _w21511_ ;
	wire _w21510_ ;
	wire _w21509_ ;
	wire _w21508_ ;
	wire _w21507_ ;
	wire _w21506_ ;
	wire _w21505_ ;
	wire _w21504_ ;
	wire _w21503_ ;
	wire _w21502_ ;
	wire _w21501_ ;
	wire _w21500_ ;
	wire _w21499_ ;
	wire _w21498_ ;
	wire _w21497_ ;
	wire _w21496_ ;
	wire _w21495_ ;
	wire _w21494_ ;
	wire _w21493_ ;
	wire _w21492_ ;
	wire _w21491_ ;
	wire _w21490_ ;
	wire _w21489_ ;
	wire _w21488_ ;
	wire _w21487_ ;
	wire _w21486_ ;
	wire _w21485_ ;
	wire _w21484_ ;
	wire _w21483_ ;
	wire _w21482_ ;
	wire _w21481_ ;
	wire _w21480_ ;
	wire _w21479_ ;
	wire _w21478_ ;
	wire _w21477_ ;
	wire _w21476_ ;
	wire _w21475_ ;
	wire _w21474_ ;
	wire _w21473_ ;
	wire _w21472_ ;
	wire _w21471_ ;
	wire _w21470_ ;
	wire _w21469_ ;
	wire _w21468_ ;
	wire _w21467_ ;
	wire _w21466_ ;
	wire _w21465_ ;
	wire _w21464_ ;
	wire _w21463_ ;
	wire _w21462_ ;
	wire _w21461_ ;
	wire _w21460_ ;
	wire _w21459_ ;
	wire _w21458_ ;
	wire _w21457_ ;
	wire _w21456_ ;
	wire _w21455_ ;
	wire _w21454_ ;
	wire _w21453_ ;
	wire _w21452_ ;
	wire _w21451_ ;
	wire _w21450_ ;
	wire _w21449_ ;
	wire _w21448_ ;
	wire _w21447_ ;
	wire _w21446_ ;
	wire _w21445_ ;
	wire _w21444_ ;
	wire _w21443_ ;
	wire _w21442_ ;
	wire _w21441_ ;
	wire _w21440_ ;
	wire _w21439_ ;
	wire _w21438_ ;
	wire _w21437_ ;
	wire _w21436_ ;
	wire _w21435_ ;
	wire _w21434_ ;
	wire _w21433_ ;
	wire _w21432_ ;
	wire _w21431_ ;
	wire _w21430_ ;
	wire _w21429_ ;
	wire _w21428_ ;
	wire _w21427_ ;
	wire _w21426_ ;
	wire _w21425_ ;
	wire _w21424_ ;
	wire _w21423_ ;
	wire _w21422_ ;
	wire _w21421_ ;
	wire _w21420_ ;
	wire _w21419_ ;
	wire _w21418_ ;
	wire _w21417_ ;
	wire _w21416_ ;
	wire _w21415_ ;
	wire _w21414_ ;
	wire _w21413_ ;
	wire _w21412_ ;
	wire _w21411_ ;
	wire _w21410_ ;
	wire _w21409_ ;
	wire _w21408_ ;
	wire _w21407_ ;
	wire _w21406_ ;
	wire _w21405_ ;
	wire _w21404_ ;
	wire _w21403_ ;
	wire _w21402_ ;
	wire _w21401_ ;
	wire _w21400_ ;
	wire _w21398_ ;
	wire _w21397_ ;
	wire _w21396_ ;
	wire _w21395_ ;
	wire _w21394_ ;
	wire _w21393_ ;
	wire _w21392_ ;
	wire _w21391_ ;
	wire _w21390_ ;
	wire _w21389_ ;
	wire _w21388_ ;
	wire _w21387_ ;
	wire _w21386_ ;
	wire _w21385_ ;
	wire _w21384_ ;
	wire _w21383_ ;
	wire _w21382_ ;
	wire _w21381_ ;
	wire _w21380_ ;
	wire _w21379_ ;
	wire _w21378_ ;
	wire _w21377_ ;
	wire _w21376_ ;
	wire _w21375_ ;
	wire _w21374_ ;
	wire _w21373_ ;
	wire _w21372_ ;
	wire _w21371_ ;
	wire _w21370_ ;
	wire _w21369_ ;
	wire _w21368_ ;
	wire _w21367_ ;
	wire _w21366_ ;
	wire _w21365_ ;
	wire _w21364_ ;
	wire _w21363_ ;
	wire _w21362_ ;
	wire _w21361_ ;
	wire _w21360_ ;
	wire _w21359_ ;
	wire _w21358_ ;
	wire _w21357_ ;
	wire _w21356_ ;
	wire _w21355_ ;
	wire _w21354_ ;
	wire _w21353_ ;
	wire _w21352_ ;
	wire _w21351_ ;
	wire _w21350_ ;
	wire _w21349_ ;
	wire _w21348_ ;
	wire _w21347_ ;
	wire _w21346_ ;
	wire _w21345_ ;
	wire _w21344_ ;
	wire _w21343_ ;
	wire _w21342_ ;
	wire _w21341_ ;
	wire _w21340_ ;
	wire _w21339_ ;
	wire _w21338_ ;
	wire _w21337_ ;
	wire _w21336_ ;
	wire _w21335_ ;
	wire _w21334_ ;
	wire _w21333_ ;
	wire _w21332_ ;
	wire _w21331_ ;
	wire _w21330_ ;
	wire _w21328_ ;
	wire _w21327_ ;
	wire _w21326_ ;
	wire _w21325_ ;
	wire _w21324_ ;
	wire _w21323_ ;
	wire _w21322_ ;
	wire _w21321_ ;
	wire _w21320_ ;
	wire _w21319_ ;
	wire _w21318_ ;
	wire _w21317_ ;
	wire _w21316_ ;
	wire _w21315_ ;
	wire _w21314_ ;
	wire _w21312_ ;
	wire _w21310_ ;
	wire _w21308_ ;
	wire _w21306_ ;
	wire _w21304_ ;
	wire _w21302_ ;
	wire _w21300_ ;
	wire _w21299_ ;
	wire _w21298_ ;
	wire _w21297_ ;
	wire _w21296_ ;
	wire _w21295_ ;
	wire _w21294_ ;
	wire _w21293_ ;
	wire _w21292_ ;
	wire _w21291_ ;
	wire _w21290_ ;
	wire _w21289_ ;
	wire _w21288_ ;
	wire _w21287_ ;
	wire _w21286_ ;
	wire _w21285_ ;
	wire _w21284_ ;
	wire _w21283_ ;
	wire _w21282_ ;
	wire _w21281_ ;
	wire _w21280_ ;
	wire _w21279_ ;
	wire _w21278_ ;
	wire _w21277_ ;
	wire _w21276_ ;
	wire _w21275_ ;
	wire _w21274_ ;
	wire _w21273_ ;
	wire _w21272_ ;
	wire _w21271_ ;
	wire _w21270_ ;
	wire _w21269_ ;
	wire _w21268_ ;
	wire _w21267_ ;
	wire _w21266_ ;
	wire _w21265_ ;
	wire _w21264_ ;
	wire _w21263_ ;
	wire _w21262_ ;
	wire _w21261_ ;
	wire _w21260_ ;
	wire _w21259_ ;
	wire _w21258_ ;
	wire _w21257_ ;
	wire _w21256_ ;
	wire _w21255_ ;
	wire _w21254_ ;
	wire _w21253_ ;
	wire _w21252_ ;
	wire _w21251_ ;
	wire _w21250_ ;
	wire _w21249_ ;
	wire _w21248_ ;
	wire _w21247_ ;
	wire _w21246_ ;
	wire _w21245_ ;
	wire _w21244_ ;
	wire _w21243_ ;
	wire _w21242_ ;
	wire _w21241_ ;
	wire _w21240_ ;
	wire _w21239_ ;
	wire _w21238_ ;
	wire _w21237_ ;
	wire _w21236_ ;
	wire _w21235_ ;
	wire _w21234_ ;
	wire _w21233_ ;
	wire _w21232_ ;
	wire _w21231_ ;
	wire _w21230_ ;
	wire _w21229_ ;
	wire _w21228_ ;
	wire _w21227_ ;
	wire _w21226_ ;
	wire _w21225_ ;
	wire _w21224_ ;
	wire _w21223_ ;
	wire _w21222_ ;
	wire _w21221_ ;
	wire _w21220_ ;
	wire _w21219_ ;
	wire _w21218_ ;
	wire _w21217_ ;
	wire _w21216_ ;
	wire _w21215_ ;
	wire _w21214_ ;
	wire _w21213_ ;
	wire _w21212_ ;
	wire _w21211_ ;
	wire _w21210_ ;
	wire _w21209_ ;
	wire _w21208_ ;
	wire _w21207_ ;
	wire _w21206_ ;
	wire _w21205_ ;
	wire _w21204_ ;
	wire _w21203_ ;
	wire _w21202_ ;
	wire _w21201_ ;
	wire _w21200_ ;
	wire _w21199_ ;
	wire _w21198_ ;
	wire _w21197_ ;
	wire _w21196_ ;
	wire _w21195_ ;
	wire _w21194_ ;
	wire _w21193_ ;
	wire _w21192_ ;
	wire _w21191_ ;
	wire _w21190_ ;
	wire _w21189_ ;
	wire _w21188_ ;
	wire _w21187_ ;
	wire _w21186_ ;
	wire _w21185_ ;
	wire _w21184_ ;
	wire _w21183_ ;
	wire _w21182_ ;
	wire _w21181_ ;
	wire _w21180_ ;
	wire _w21179_ ;
	wire _w21178_ ;
	wire _w21177_ ;
	wire _w21176_ ;
	wire _w21175_ ;
	wire _w21174_ ;
	wire _w21173_ ;
	wire _w21172_ ;
	wire _w21171_ ;
	wire _w21170_ ;
	wire _w21169_ ;
	wire _w21168_ ;
	wire _w21167_ ;
	wire _w21166_ ;
	wire _w21165_ ;
	wire _w21164_ ;
	wire _w21163_ ;
	wire _w21162_ ;
	wire _w21161_ ;
	wire _w21160_ ;
	wire _w21159_ ;
	wire _w21158_ ;
	wire _w21157_ ;
	wire _w21156_ ;
	wire _w21155_ ;
	wire _w21154_ ;
	wire _w21153_ ;
	wire _w21152_ ;
	wire _w21151_ ;
	wire _w21150_ ;
	wire _w21149_ ;
	wire _w21148_ ;
	wire _w21147_ ;
	wire _w21146_ ;
	wire _w21145_ ;
	wire _w21144_ ;
	wire _w21143_ ;
	wire _w21142_ ;
	wire _w21141_ ;
	wire _w21140_ ;
	wire _w21139_ ;
	wire _w21138_ ;
	wire _w21137_ ;
	wire _w21136_ ;
	wire _w21135_ ;
	wire _w21134_ ;
	wire _w21133_ ;
	wire _w21132_ ;
	wire _w21131_ ;
	wire _w21130_ ;
	wire _w21129_ ;
	wire _w21128_ ;
	wire _w21127_ ;
	wire _w21126_ ;
	wire _w21125_ ;
	wire _w21124_ ;
	wire _w21123_ ;
	wire _w21122_ ;
	wire _w21121_ ;
	wire _w21120_ ;
	wire _w21119_ ;
	wire _w21118_ ;
	wire _w21117_ ;
	wire _w21116_ ;
	wire _w21115_ ;
	wire _w21114_ ;
	wire _w21113_ ;
	wire _w21112_ ;
	wire _w21111_ ;
	wire _w21110_ ;
	wire _w21109_ ;
	wire _w21108_ ;
	wire _w21107_ ;
	wire _w21106_ ;
	wire _w21105_ ;
	wire _w21104_ ;
	wire _w21103_ ;
	wire _w21102_ ;
	wire _w21101_ ;
	wire _w21100_ ;
	wire _w21099_ ;
	wire _w21098_ ;
	wire _w21097_ ;
	wire _w21096_ ;
	wire _w21095_ ;
	wire _w21094_ ;
	wire _w21093_ ;
	wire _w21092_ ;
	wire _w21091_ ;
	wire _w21090_ ;
	wire _w21089_ ;
	wire _w21088_ ;
	wire _w21087_ ;
	wire _w21086_ ;
	wire _w21085_ ;
	wire _w21084_ ;
	wire _w21083_ ;
	wire _w21082_ ;
	wire _w21081_ ;
	wire _w21080_ ;
	wire _w21079_ ;
	wire _w21078_ ;
	wire _w21077_ ;
	wire _w21076_ ;
	wire _w21075_ ;
	wire _w21074_ ;
	wire _w21073_ ;
	wire _w21072_ ;
	wire _w21071_ ;
	wire _w21070_ ;
	wire _w21069_ ;
	wire _w21068_ ;
	wire _w21067_ ;
	wire _w21066_ ;
	wire _w21065_ ;
	wire _w21064_ ;
	wire _w21063_ ;
	wire _w21062_ ;
	wire _w21061_ ;
	wire _w21060_ ;
	wire _w21059_ ;
	wire _w21058_ ;
	wire _w21057_ ;
	wire _w21056_ ;
	wire _w21055_ ;
	wire _w21054_ ;
	wire _w21053_ ;
	wire _w21052_ ;
	wire _w21051_ ;
	wire _w21050_ ;
	wire _w21049_ ;
	wire _w21048_ ;
	wire _w21047_ ;
	wire _w21046_ ;
	wire _w21045_ ;
	wire _w21044_ ;
	wire _w21043_ ;
	wire _w21042_ ;
	wire _w21041_ ;
	wire _w21040_ ;
	wire _w21039_ ;
	wire _w21038_ ;
	wire _w21037_ ;
	wire _w21036_ ;
	wire _w21035_ ;
	wire _w21034_ ;
	wire _w21033_ ;
	wire _w21032_ ;
	wire _w21031_ ;
	wire _w21030_ ;
	wire _w21029_ ;
	wire _w21028_ ;
	wire _w21027_ ;
	wire _w21026_ ;
	wire _w21025_ ;
	wire _w21024_ ;
	wire _w21023_ ;
	wire _w21022_ ;
	wire _w21021_ ;
	wire _w21020_ ;
	wire _w21019_ ;
	wire _w21018_ ;
	wire _w21017_ ;
	wire _w21016_ ;
	wire _w21015_ ;
	wire _w21014_ ;
	wire _w21013_ ;
	wire _w21012_ ;
	wire _w21011_ ;
	wire _w21010_ ;
	wire _w21009_ ;
	wire _w21008_ ;
	wire _w21007_ ;
	wire _w21006_ ;
	wire _w21005_ ;
	wire _w21004_ ;
	wire _w21003_ ;
	wire _w21002_ ;
	wire _w21001_ ;
	wire _w21000_ ;
	wire _w20999_ ;
	wire _w20998_ ;
	wire _w20997_ ;
	wire _w20996_ ;
	wire _w20995_ ;
	wire _w20994_ ;
	wire _w20993_ ;
	wire _w20992_ ;
	wire _w20991_ ;
	wire _w20990_ ;
	wire _w20989_ ;
	wire _w20988_ ;
	wire _w20987_ ;
	wire _w20986_ ;
	wire _w20985_ ;
	wire _w20984_ ;
	wire _w20983_ ;
	wire _w20982_ ;
	wire _w20981_ ;
	wire _w20980_ ;
	wire _w20979_ ;
	wire _w20978_ ;
	wire _w20977_ ;
	wire _w20976_ ;
	wire _w20975_ ;
	wire _w20974_ ;
	wire _w20973_ ;
	wire _w20972_ ;
	wire _w20971_ ;
	wire _w20970_ ;
	wire _w20969_ ;
	wire _w20968_ ;
	wire _w20967_ ;
	wire _w20966_ ;
	wire _w20965_ ;
	wire _w20964_ ;
	wire _w20963_ ;
	wire _w20962_ ;
	wire _w20961_ ;
	wire _w20960_ ;
	wire _w20959_ ;
	wire _w20958_ ;
	wire _w20957_ ;
	wire _w20956_ ;
	wire _w20955_ ;
	wire _w20954_ ;
	wire _w20953_ ;
	wire _w20952_ ;
	wire _w20951_ ;
	wire _w20950_ ;
	wire _w20949_ ;
	wire _w20948_ ;
	wire _w20947_ ;
	wire _w20946_ ;
	wire _w20945_ ;
	wire _w20944_ ;
	wire _w20943_ ;
	wire _w20942_ ;
	wire _w20941_ ;
	wire _w20940_ ;
	wire _w20939_ ;
	wire _w20938_ ;
	wire _w20937_ ;
	wire _w20936_ ;
	wire _w20935_ ;
	wire _w20934_ ;
	wire _w20933_ ;
	wire _w20932_ ;
	wire _w20931_ ;
	wire _w20930_ ;
	wire _w20929_ ;
	wire _w20928_ ;
	wire _w20927_ ;
	wire _w20926_ ;
	wire _w20925_ ;
	wire _w20924_ ;
	wire _w20923_ ;
	wire _w20922_ ;
	wire _w20921_ ;
	wire _w20920_ ;
	wire _w20919_ ;
	wire _w20918_ ;
	wire _w20917_ ;
	wire _w20916_ ;
	wire _w20915_ ;
	wire _w20914_ ;
	wire _w20913_ ;
	wire _w20912_ ;
	wire _w20911_ ;
	wire _w20910_ ;
	wire _w20909_ ;
	wire _w20908_ ;
	wire _w20907_ ;
	wire _w20906_ ;
	wire _w20905_ ;
	wire _w20904_ ;
	wire _w20903_ ;
	wire _w20902_ ;
	wire _w20901_ ;
	wire _w20900_ ;
	wire _w20899_ ;
	wire _w20898_ ;
	wire _w20897_ ;
	wire _w20896_ ;
	wire _w20895_ ;
	wire _w20894_ ;
	wire _w20893_ ;
	wire _w20892_ ;
	wire _w20891_ ;
	wire _w20890_ ;
	wire _w20889_ ;
	wire _w20888_ ;
	wire _w20887_ ;
	wire _w20886_ ;
	wire _w20885_ ;
	wire _w20884_ ;
	wire _w20883_ ;
	wire _w20882_ ;
	wire _w20881_ ;
	wire _w20880_ ;
	wire _w20879_ ;
	wire _w20878_ ;
	wire _w20877_ ;
	wire _w20876_ ;
	wire _w20875_ ;
	wire _w20874_ ;
	wire _w20873_ ;
	wire _w20872_ ;
	wire _w20871_ ;
	wire _w20870_ ;
	wire _w20869_ ;
	wire _w20868_ ;
	wire _w20867_ ;
	wire _w20866_ ;
	wire _w20865_ ;
	wire _w20864_ ;
	wire _w20863_ ;
	wire _w20862_ ;
	wire _w20861_ ;
	wire _w20860_ ;
	wire _w20859_ ;
	wire _w20858_ ;
	wire _w20857_ ;
	wire _w20856_ ;
	wire _w20855_ ;
	wire _w20854_ ;
	wire _w20853_ ;
	wire _w20852_ ;
	wire _w20851_ ;
	wire _w20850_ ;
	wire _w20849_ ;
	wire _w20848_ ;
	wire _w20847_ ;
	wire _w20846_ ;
	wire _w20845_ ;
	wire _w20844_ ;
	wire _w20843_ ;
	wire _w20842_ ;
	wire _w20841_ ;
	wire _w20840_ ;
	wire _w20839_ ;
	wire _w20838_ ;
	wire _w20837_ ;
	wire _w20836_ ;
	wire _w20835_ ;
	wire _w20834_ ;
	wire _w20833_ ;
	wire _w20832_ ;
	wire _w20831_ ;
	wire _w20830_ ;
	wire _w20829_ ;
	wire _w20828_ ;
	wire _w20827_ ;
	wire _w20826_ ;
	wire _w20825_ ;
	wire _w20824_ ;
	wire _w20823_ ;
	wire _w20822_ ;
	wire _w20821_ ;
	wire _w20820_ ;
	wire _w20819_ ;
	wire _w20818_ ;
	wire _w20817_ ;
	wire _w20816_ ;
	wire _w20815_ ;
	wire _w20814_ ;
	wire _w20813_ ;
	wire _w20812_ ;
	wire _w20811_ ;
	wire _w20810_ ;
	wire _w20809_ ;
	wire _w20808_ ;
	wire _w20807_ ;
	wire _w20806_ ;
	wire _w20805_ ;
	wire _w20804_ ;
	wire _w20803_ ;
	wire _w20802_ ;
	wire _w20801_ ;
	wire _w20800_ ;
	wire _w20799_ ;
	wire _w20798_ ;
	wire _w20797_ ;
	wire _w20796_ ;
	wire _w20795_ ;
	wire _w20794_ ;
	wire _w20793_ ;
	wire _w20792_ ;
	wire _w20791_ ;
	wire _w20790_ ;
	wire _w20789_ ;
	wire _w20788_ ;
	wire _w20787_ ;
	wire _w20786_ ;
	wire _w20785_ ;
	wire _w20784_ ;
	wire _w20783_ ;
	wire _w20782_ ;
	wire _w20781_ ;
	wire _w20780_ ;
	wire _w20779_ ;
	wire _w20778_ ;
	wire _w20777_ ;
	wire _w20776_ ;
	wire _w20775_ ;
	wire _w20774_ ;
	wire _w20773_ ;
	wire _w20772_ ;
	wire _w20771_ ;
	wire _w20770_ ;
	wire _w20769_ ;
	wire _w20768_ ;
	wire _w20767_ ;
	wire _w20766_ ;
	wire _w20765_ ;
	wire _w20764_ ;
	wire _w20763_ ;
	wire _w20762_ ;
	wire _w20761_ ;
	wire _w20760_ ;
	wire _w20759_ ;
	wire _w20758_ ;
	wire _w20757_ ;
	wire _w20756_ ;
	wire _w20755_ ;
	wire _w20754_ ;
	wire _w20753_ ;
	wire _w20752_ ;
	wire _w20751_ ;
	wire _w20750_ ;
	wire _w20749_ ;
	wire _w20748_ ;
	wire _w20747_ ;
	wire _w20746_ ;
	wire _w20745_ ;
	wire _w20744_ ;
	wire _w20743_ ;
	wire _w20742_ ;
	wire _w20741_ ;
	wire _w20740_ ;
	wire _w20739_ ;
	wire _w20738_ ;
	wire _w20737_ ;
	wire _w20736_ ;
	wire _w20735_ ;
	wire _w20734_ ;
	wire _w20733_ ;
	wire _w20732_ ;
	wire _w20731_ ;
	wire _w20730_ ;
	wire _w20729_ ;
	wire _w20728_ ;
	wire _w20727_ ;
	wire _w20726_ ;
	wire _w20725_ ;
	wire _w20724_ ;
	wire _w20723_ ;
	wire _w20722_ ;
	wire _w20721_ ;
	wire _w20720_ ;
	wire _w20719_ ;
	wire _w20718_ ;
	wire _w20717_ ;
	wire _w20716_ ;
	wire _w20715_ ;
	wire _w20714_ ;
	wire _w20713_ ;
	wire _w20712_ ;
	wire _w20711_ ;
	wire _w20710_ ;
	wire _w20709_ ;
	wire _w20708_ ;
	wire _w20707_ ;
	wire _w20706_ ;
	wire _w20705_ ;
	wire _w20704_ ;
	wire _w20703_ ;
	wire _w20702_ ;
	wire _w20701_ ;
	wire _w20700_ ;
	wire _w20699_ ;
	wire _w20698_ ;
	wire _w20697_ ;
	wire _w20696_ ;
	wire _w20695_ ;
	wire _w20694_ ;
	wire _w20693_ ;
	wire _w20692_ ;
	wire _w20691_ ;
	wire _w20690_ ;
	wire _w20689_ ;
	wire _w20688_ ;
	wire _w20687_ ;
	wire _w20686_ ;
	wire _w20685_ ;
	wire _w20684_ ;
	wire _w20683_ ;
	wire _w20682_ ;
	wire _w20681_ ;
	wire _w20680_ ;
	wire _w20679_ ;
	wire _w20678_ ;
	wire _w20677_ ;
	wire _w20676_ ;
	wire _w20675_ ;
	wire _w20674_ ;
	wire _w20673_ ;
	wire _w20672_ ;
	wire _w20671_ ;
	wire _w20670_ ;
	wire _w20669_ ;
	wire _w20668_ ;
	wire _w20667_ ;
	wire _w20666_ ;
	wire _w20665_ ;
	wire _w20664_ ;
	wire _w20663_ ;
	wire _w20662_ ;
	wire _w20661_ ;
	wire _w20660_ ;
	wire _w20659_ ;
	wire _w20658_ ;
	wire _w20657_ ;
	wire _w20656_ ;
	wire _w20655_ ;
	wire _w20654_ ;
	wire _w20653_ ;
	wire _w20652_ ;
	wire _w20651_ ;
	wire _w20650_ ;
	wire _w20649_ ;
	wire _w20648_ ;
	wire _w20647_ ;
	wire _w20646_ ;
	wire _w20645_ ;
	wire _w20644_ ;
	wire _w20643_ ;
	wire _w20642_ ;
	wire _w20641_ ;
	wire _w20640_ ;
	wire _w20639_ ;
	wire _w20638_ ;
	wire _w20637_ ;
	wire _w20636_ ;
	wire _w20635_ ;
	wire _w20634_ ;
	wire _w20633_ ;
	wire _w20632_ ;
	wire _w20631_ ;
	wire _w20630_ ;
	wire _w20629_ ;
	wire _w20628_ ;
	wire _w20627_ ;
	wire _w20626_ ;
	wire _w20625_ ;
	wire _w20624_ ;
	wire _w20623_ ;
	wire _w20622_ ;
	wire _w20621_ ;
	wire _w20620_ ;
	wire _w20619_ ;
	wire _w20618_ ;
	wire _w20617_ ;
	wire _w20616_ ;
	wire _w20615_ ;
	wire _w20614_ ;
	wire _w20613_ ;
	wire _w20612_ ;
	wire _w20611_ ;
	wire _w20610_ ;
	wire _w20609_ ;
	wire _w20608_ ;
	wire _w20607_ ;
	wire _w20606_ ;
	wire _w20605_ ;
	wire _w20604_ ;
	wire _w20603_ ;
	wire _w20602_ ;
	wire _w20601_ ;
	wire _w20600_ ;
	wire _w20599_ ;
	wire _w20598_ ;
	wire _w20597_ ;
	wire _w20596_ ;
	wire _w20595_ ;
	wire _w20594_ ;
	wire _w20593_ ;
	wire _w20592_ ;
	wire _w20591_ ;
	wire _w20590_ ;
	wire _w20589_ ;
	wire _w20588_ ;
	wire _w20587_ ;
	wire _w20586_ ;
	wire _w20585_ ;
	wire _w20584_ ;
	wire _w20583_ ;
	wire _w20582_ ;
	wire _w20581_ ;
	wire _w20580_ ;
	wire _w20579_ ;
	wire _w20578_ ;
	wire _w20577_ ;
	wire _w20576_ ;
	wire _w20575_ ;
	wire _w20574_ ;
	wire _w20573_ ;
	wire _w20572_ ;
	wire _w20571_ ;
	wire _w20570_ ;
	wire _w20569_ ;
	wire _w20568_ ;
	wire _w20567_ ;
	wire _w20566_ ;
	wire _w20565_ ;
	wire _w20564_ ;
	wire _w20563_ ;
	wire _w20562_ ;
	wire _w20561_ ;
	wire _w20560_ ;
	wire _w20559_ ;
	wire _w20558_ ;
	wire _w20557_ ;
	wire _w20556_ ;
	wire _w20555_ ;
	wire _w20554_ ;
	wire _w20553_ ;
	wire _w20552_ ;
	wire _w20551_ ;
	wire _w20550_ ;
	wire _w20549_ ;
	wire _w20548_ ;
	wire _w20547_ ;
	wire _w20546_ ;
	wire _w20545_ ;
	wire _w20544_ ;
	wire _w20543_ ;
	wire _w20542_ ;
	wire _w20541_ ;
	wire _w20540_ ;
	wire _w20539_ ;
	wire _w20538_ ;
	wire _w20537_ ;
	wire _w20536_ ;
	wire _w20535_ ;
	wire _w20534_ ;
	wire _w20533_ ;
	wire _w20532_ ;
	wire _w20531_ ;
	wire _w20530_ ;
	wire _w20529_ ;
	wire _w20528_ ;
	wire _w20527_ ;
	wire _w20526_ ;
	wire _w20525_ ;
	wire _w20524_ ;
	wire _w20523_ ;
	wire _w20522_ ;
	wire _w20521_ ;
	wire _w20520_ ;
	wire _w20519_ ;
	wire _w20518_ ;
	wire _w20517_ ;
	wire _w20516_ ;
	wire _w20515_ ;
	wire _w20514_ ;
	wire _w20513_ ;
	wire _w20512_ ;
	wire _w20511_ ;
	wire _w20510_ ;
	wire _w20509_ ;
	wire _w20508_ ;
	wire _w20507_ ;
	wire _w20506_ ;
	wire _w20505_ ;
	wire _w20504_ ;
	wire _w20503_ ;
	wire _w20502_ ;
	wire _w20501_ ;
	wire _w20500_ ;
	wire _w20499_ ;
	wire _w20498_ ;
	wire _w20497_ ;
	wire _w20496_ ;
	wire _w20495_ ;
	wire _w20494_ ;
	wire _w20493_ ;
	wire _w20492_ ;
	wire _w20491_ ;
	wire _w20490_ ;
	wire _w20489_ ;
	wire _w20488_ ;
	wire _w20487_ ;
	wire _w20486_ ;
	wire _w20485_ ;
	wire _w20484_ ;
	wire _w20483_ ;
	wire _w20482_ ;
	wire _w20481_ ;
	wire _w20480_ ;
	wire _w20479_ ;
	wire _w20478_ ;
	wire _w20477_ ;
	wire _w20476_ ;
	wire _w20475_ ;
	wire _w20474_ ;
	wire _w20473_ ;
	wire _w20472_ ;
	wire _w20471_ ;
	wire _w20470_ ;
	wire _w20469_ ;
	wire _w20468_ ;
	wire _w20467_ ;
	wire _w20466_ ;
	wire _w20465_ ;
	wire _w20464_ ;
	wire _w20463_ ;
	wire _w20462_ ;
	wire _w20461_ ;
	wire _w20460_ ;
	wire _w20459_ ;
	wire _w20458_ ;
	wire _w20457_ ;
	wire _w20456_ ;
	wire _w20455_ ;
	wire _w20454_ ;
	wire _w20453_ ;
	wire _w20452_ ;
	wire _w20451_ ;
	wire _w20450_ ;
	wire _w20449_ ;
	wire _w20448_ ;
	wire _w20447_ ;
	wire _w20446_ ;
	wire _w20445_ ;
	wire _w20444_ ;
	wire _w20443_ ;
	wire _w20442_ ;
	wire _w20441_ ;
	wire _w20440_ ;
	wire _w20439_ ;
	wire _w20438_ ;
	wire _w20437_ ;
	wire _w20436_ ;
	wire _w20435_ ;
	wire _w20434_ ;
	wire _w20433_ ;
	wire _w20432_ ;
	wire _w20431_ ;
	wire _w20430_ ;
	wire _w20429_ ;
	wire _w20428_ ;
	wire _w20427_ ;
	wire _w20426_ ;
	wire _w20425_ ;
	wire _w20424_ ;
	wire _w20423_ ;
	wire _w20422_ ;
	wire _w20421_ ;
	wire _w20420_ ;
	wire _w20419_ ;
	wire _w20418_ ;
	wire _w20417_ ;
	wire _w20416_ ;
	wire _w20415_ ;
	wire _w20414_ ;
	wire _w20413_ ;
	wire _w20412_ ;
	wire _w20411_ ;
	wire _w20410_ ;
	wire _w20409_ ;
	wire _w20408_ ;
	wire _w20407_ ;
	wire _w20406_ ;
	wire _w20405_ ;
	wire _w20404_ ;
	wire _w20403_ ;
	wire _w20402_ ;
	wire _w20401_ ;
	wire _w20400_ ;
	wire _w20399_ ;
	wire _w20398_ ;
	wire _w20397_ ;
	wire _w20396_ ;
	wire _w20395_ ;
	wire _w20394_ ;
	wire _w20393_ ;
	wire _w20392_ ;
	wire _w20391_ ;
	wire _w20390_ ;
	wire _w20389_ ;
	wire _w20388_ ;
	wire _w20387_ ;
	wire _w20386_ ;
	wire _w20385_ ;
	wire _w20384_ ;
	wire _w20383_ ;
	wire _w20382_ ;
	wire _w20381_ ;
	wire _w20380_ ;
	wire _w20379_ ;
	wire _w20378_ ;
	wire _w20377_ ;
	wire _w20376_ ;
	wire _w20375_ ;
	wire _w20374_ ;
	wire _w20373_ ;
	wire _w20372_ ;
	wire _w20371_ ;
	wire _w20370_ ;
	wire _w20369_ ;
	wire _w20368_ ;
	wire _w20367_ ;
	wire _w20366_ ;
	wire _w20365_ ;
	wire _w20364_ ;
	wire _w20363_ ;
	wire _w20362_ ;
	wire _w20361_ ;
	wire _w20360_ ;
	wire _w20359_ ;
	wire _w20358_ ;
	wire _w20357_ ;
	wire _w20356_ ;
	wire _w20355_ ;
	wire _w20354_ ;
	wire _w20353_ ;
	wire _w20352_ ;
	wire _w20351_ ;
	wire _w20350_ ;
	wire _w20349_ ;
	wire _w20348_ ;
	wire _w20347_ ;
	wire _w20346_ ;
	wire _w20345_ ;
	wire _w20344_ ;
	wire _w20343_ ;
	wire _w20342_ ;
	wire _w20341_ ;
	wire _w20340_ ;
	wire _w20339_ ;
	wire _w20338_ ;
	wire _w20337_ ;
	wire _w20336_ ;
	wire _w20335_ ;
	wire _w20334_ ;
	wire _w20333_ ;
	wire _w20332_ ;
	wire _w20331_ ;
	wire _w20330_ ;
	wire _w20329_ ;
	wire _w20328_ ;
	wire _w20327_ ;
	wire _w20326_ ;
	wire _w20325_ ;
	wire _w20324_ ;
	wire _w20323_ ;
	wire _w20322_ ;
	wire _w20321_ ;
	wire _w20320_ ;
	wire _w20319_ ;
	wire _w20318_ ;
	wire _w20317_ ;
	wire _w20316_ ;
	wire _w20315_ ;
	wire _w20314_ ;
	wire _w20313_ ;
	wire _w20312_ ;
	wire _w20311_ ;
	wire _w20310_ ;
	wire _w20309_ ;
	wire _w20308_ ;
	wire _w20307_ ;
	wire _w20306_ ;
	wire _w20305_ ;
	wire _w20304_ ;
	wire _w20303_ ;
	wire _w20302_ ;
	wire _w20301_ ;
	wire _w20300_ ;
	wire _w20299_ ;
	wire _w20298_ ;
	wire _w20297_ ;
	wire _w20296_ ;
	wire _w20295_ ;
	wire _w20294_ ;
	wire _w20293_ ;
	wire _w20292_ ;
	wire _w20291_ ;
	wire _w20290_ ;
	wire _w20289_ ;
	wire _w20288_ ;
	wire _w20287_ ;
	wire _w20286_ ;
	wire _w20285_ ;
	wire _w20284_ ;
	wire _w20283_ ;
	wire _w20282_ ;
	wire _w20281_ ;
	wire _w20280_ ;
	wire _w20279_ ;
	wire _w20278_ ;
	wire _w20277_ ;
	wire _w20276_ ;
	wire _w20275_ ;
	wire _w20274_ ;
	wire _w20273_ ;
	wire _w20272_ ;
	wire _w20271_ ;
	wire _w20270_ ;
	wire _w20269_ ;
	wire _w20268_ ;
	wire _w20267_ ;
	wire _w20266_ ;
	wire _w20265_ ;
	wire _w20264_ ;
	wire _w20263_ ;
	wire _w20262_ ;
	wire _w20261_ ;
	wire _w20260_ ;
	wire _w20259_ ;
	wire _w20258_ ;
	wire _w20257_ ;
	wire _w20256_ ;
	wire _w20255_ ;
	wire _w20254_ ;
	wire _w20253_ ;
	wire _w20252_ ;
	wire _w20251_ ;
	wire _w20250_ ;
	wire _w20249_ ;
	wire _w20248_ ;
	wire _w20247_ ;
	wire _w20246_ ;
	wire _w20245_ ;
	wire _w20244_ ;
	wire _w20243_ ;
	wire _w20242_ ;
	wire _w20241_ ;
	wire _w20240_ ;
	wire _w20239_ ;
	wire _w20238_ ;
	wire _w20237_ ;
	wire _w20236_ ;
	wire _w20235_ ;
	wire _w20234_ ;
	wire _w20233_ ;
	wire _w20232_ ;
	wire _w20231_ ;
	wire _w20230_ ;
	wire _w20229_ ;
	wire _w20228_ ;
	wire _w20227_ ;
	wire _w20226_ ;
	wire _w20225_ ;
	wire _w20224_ ;
	wire _w20223_ ;
	wire _w20222_ ;
	wire _w20221_ ;
	wire _w20220_ ;
	wire _w20219_ ;
	wire _w20218_ ;
	wire _w20217_ ;
	wire _w20216_ ;
	wire _w20215_ ;
	wire _w20214_ ;
	wire _w20213_ ;
	wire _w20212_ ;
	wire _w20211_ ;
	wire _w20210_ ;
	wire _w20209_ ;
	wire _w20208_ ;
	wire _w20207_ ;
	wire _w20206_ ;
	wire _w20205_ ;
	wire _w20204_ ;
	wire _w20203_ ;
	wire _w20202_ ;
	wire _w20201_ ;
	wire _w20200_ ;
	wire _w20199_ ;
	wire _w20198_ ;
	wire _w20197_ ;
	wire _w20196_ ;
	wire _w20195_ ;
	wire _w20194_ ;
	wire _w20193_ ;
	wire _w20192_ ;
	wire _w20191_ ;
	wire _w20190_ ;
	wire _w20189_ ;
	wire _w20188_ ;
	wire _w20187_ ;
	wire _w20186_ ;
	wire _w20185_ ;
	wire _w20184_ ;
	wire _w20183_ ;
	wire _w20182_ ;
	wire _w20181_ ;
	wire _w20180_ ;
	wire _w20179_ ;
	wire _w20178_ ;
	wire _w20177_ ;
	wire _w20176_ ;
	wire _w20175_ ;
	wire _w20174_ ;
	wire _w20173_ ;
	wire _w20172_ ;
	wire _w20171_ ;
	wire _w20170_ ;
	wire _w20169_ ;
	wire _w20168_ ;
	wire _w20167_ ;
	wire _w20166_ ;
	wire _w20165_ ;
	wire _w20164_ ;
	wire _w20163_ ;
	wire _w20162_ ;
	wire _w20161_ ;
	wire _w20160_ ;
	wire _w20159_ ;
	wire _w20158_ ;
	wire _w20157_ ;
	wire _w20156_ ;
	wire _w20155_ ;
	wire _w20154_ ;
	wire _w20153_ ;
	wire _w20152_ ;
	wire _w20151_ ;
	wire _w20150_ ;
	wire _w20149_ ;
	wire _w20148_ ;
	wire _w20147_ ;
	wire _w20146_ ;
	wire _w20145_ ;
	wire _w20144_ ;
	wire _w20143_ ;
	wire _w20142_ ;
	wire _w20141_ ;
	wire _w20140_ ;
	wire _w20139_ ;
	wire _w20138_ ;
	wire _w20137_ ;
	wire _w20136_ ;
	wire _w20135_ ;
	wire _w20134_ ;
	wire _w20133_ ;
	wire _w20132_ ;
	wire _w20131_ ;
	wire _w20130_ ;
	wire _w20129_ ;
	wire _w20128_ ;
	wire _w20127_ ;
	wire _w20126_ ;
	wire _w20125_ ;
	wire _w20124_ ;
	wire _w20123_ ;
	wire _w20122_ ;
	wire _w20121_ ;
	wire _w20120_ ;
	wire _w20119_ ;
	wire _w20118_ ;
	wire _w20117_ ;
	wire _w20116_ ;
	wire _w20115_ ;
	wire _w20114_ ;
	wire _w20113_ ;
	wire _w20112_ ;
	wire _w20111_ ;
	wire _w20110_ ;
	wire _w20109_ ;
	wire _w20108_ ;
	wire _w20107_ ;
	wire _w20106_ ;
	wire _w20105_ ;
	wire _w20104_ ;
	wire _w20103_ ;
	wire _w20102_ ;
	wire _w20101_ ;
	wire _w20100_ ;
	wire _w20099_ ;
	wire _w20098_ ;
	wire _w20097_ ;
	wire _w20096_ ;
	wire _w20095_ ;
	wire _w20094_ ;
	wire _w20093_ ;
	wire _w20092_ ;
	wire _w20091_ ;
	wire _w20090_ ;
	wire _w20089_ ;
	wire _w20088_ ;
	wire _w20087_ ;
	wire _w20086_ ;
	wire _w20085_ ;
	wire _w20084_ ;
	wire _w20083_ ;
	wire _w20082_ ;
	wire _w20081_ ;
	wire _w20080_ ;
	wire _w20079_ ;
	wire _w20078_ ;
	wire _w20077_ ;
	wire _w20076_ ;
	wire _w20075_ ;
	wire _w20074_ ;
	wire _w20073_ ;
	wire _w20072_ ;
	wire _w20071_ ;
	wire _w20070_ ;
	wire _w20069_ ;
	wire _w20068_ ;
	wire _w20067_ ;
	wire _w20066_ ;
	wire _w20065_ ;
	wire _w20064_ ;
	wire _w20063_ ;
	wire _w20062_ ;
	wire _w20061_ ;
	wire _w20060_ ;
	wire _w20059_ ;
	wire _w20058_ ;
	wire _w20057_ ;
	wire _w20056_ ;
	wire _w20055_ ;
	wire _w20054_ ;
	wire _w20053_ ;
	wire _w20052_ ;
	wire _w20051_ ;
	wire _w20050_ ;
	wire _w20049_ ;
	wire _w20048_ ;
	wire _w20047_ ;
	wire _w20046_ ;
	wire _w20045_ ;
	wire _w20044_ ;
	wire _w20043_ ;
	wire _w20042_ ;
	wire _w20041_ ;
	wire _w20040_ ;
	wire _w20039_ ;
	wire _w20038_ ;
	wire _w20037_ ;
	wire _w20036_ ;
	wire _w20035_ ;
	wire _w20034_ ;
	wire _w20033_ ;
	wire _w20032_ ;
	wire _w20031_ ;
	wire _w20030_ ;
	wire _w20029_ ;
	wire _w20028_ ;
	wire _w20027_ ;
	wire _w20026_ ;
	wire _w20025_ ;
	wire _w20024_ ;
	wire _w20023_ ;
	wire _w20022_ ;
	wire _w20021_ ;
	wire _w20020_ ;
	wire _w20019_ ;
	wire _w20018_ ;
	wire _w20017_ ;
	wire _w20016_ ;
	wire _w20015_ ;
	wire _w20014_ ;
	wire _w20013_ ;
	wire _w20012_ ;
	wire _w20011_ ;
	wire _w20010_ ;
	wire _w20009_ ;
	wire _w20008_ ;
	wire _w20007_ ;
	wire _w20006_ ;
	wire _w20005_ ;
	wire _w20004_ ;
	wire _w20003_ ;
	wire _w20002_ ;
	wire _w20001_ ;
	wire _w20000_ ;
	wire _w19999_ ;
	wire _w19998_ ;
	wire _w19997_ ;
	wire _w19996_ ;
	wire _w19995_ ;
	wire _w19994_ ;
	wire _w19993_ ;
	wire _w19992_ ;
	wire _w19991_ ;
	wire _w19990_ ;
	wire _w19989_ ;
	wire _w19988_ ;
	wire _w19987_ ;
	wire _w19986_ ;
	wire _w19985_ ;
	wire _w19984_ ;
	wire _w19983_ ;
	wire _w19982_ ;
	wire _w19981_ ;
	wire _w19980_ ;
	wire _w19979_ ;
	wire _w19978_ ;
	wire _w19977_ ;
	wire _w19976_ ;
	wire _w19975_ ;
	wire _w19974_ ;
	wire _w19973_ ;
	wire _w19972_ ;
	wire _w19971_ ;
	wire _w19970_ ;
	wire _w19969_ ;
	wire _w19968_ ;
	wire _w19967_ ;
	wire _w19966_ ;
	wire _w19965_ ;
	wire _w19964_ ;
	wire _w19963_ ;
	wire _w19962_ ;
	wire _w19961_ ;
	wire _w19960_ ;
	wire _w19959_ ;
	wire _w19958_ ;
	wire _w19957_ ;
	wire _w19956_ ;
	wire _w19955_ ;
	wire _w19954_ ;
	wire _w19953_ ;
	wire _w19952_ ;
	wire _w19951_ ;
	wire _w19950_ ;
	wire _w19949_ ;
	wire _w19948_ ;
	wire _w19947_ ;
	wire _w19946_ ;
	wire _w19945_ ;
	wire _w19944_ ;
	wire _w19943_ ;
	wire _w19942_ ;
	wire _w19941_ ;
	wire _w19940_ ;
	wire _w19939_ ;
	wire _w19938_ ;
	wire _w19937_ ;
	wire _w19936_ ;
	wire _w19935_ ;
	wire _w19934_ ;
	wire _w19933_ ;
	wire _w19932_ ;
	wire _w19931_ ;
	wire _w19930_ ;
	wire _w19929_ ;
	wire _w19928_ ;
	wire _w19927_ ;
	wire _w19926_ ;
	wire _w19925_ ;
	wire _w19924_ ;
	wire _w19923_ ;
	wire _w19922_ ;
	wire _w19921_ ;
	wire _w19920_ ;
	wire _w19919_ ;
	wire _w19918_ ;
	wire _w19917_ ;
	wire _w19916_ ;
	wire _w19915_ ;
	wire _w19914_ ;
	wire _w19913_ ;
	wire _w19912_ ;
	wire _w19911_ ;
	wire _w19910_ ;
	wire _w19909_ ;
	wire _w19908_ ;
	wire _w19907_ ;
	wire _w19906_ ;
	wire _w19905_ ;
	wire _w19904_ ;
	wire _w19903_ ;
	wire _w19902_ ;
	wire _w19901_ ;
	wire _w19900_ ;
	wire _w19899_ ;
	wire _w19898_ ;
	wire _w19897_ ;
	wire _w19896_ ;
	wire _w19895_ ;
	wire _w19894_ ;
	wire _w19893_ ;
	wire _w19892_ ;
	wire _w19891_ ;
	wire _w19890_ ;
	wire _w19889_ ;
	wire _w19888_ ;
	wire _w19887_ ;
	wire _w19886_ ;
	wire _w19885_ ;
	wire _w19884_ ;
	wire _w19883_ ;
	wire _w19882_ ;
	wire _w19881_ ;
	wire _w19880_ ;
	wire _w19879_ ;
	wire _w19878_ ;
	wire _w19877_ ;
	wire _w19876_ ;
	wire _w19875_ ;
	wire _w19874_ ;
	wire _w19873_ ;
	wire _w19872_ ;
	wire _w19871_ ;
	wire _w19870_ ;
	wire _w19869_ ;
	wire _w19868_ ;
	wire _w19867_ ;
	wire _w19866_ ;
	wire _w19865_ ;
	wire _w19864_ ;
	wire _w19863_ ;
	wire _w19862_ ;
	wire _w19861_ ;
	wire _w19860_ ;
	wire _w19859_ ;
	wire _w19858_ ;
	wire _w19857_ ;
	wire _w19856_ ;
	wire _w19855_ ;
	wire _w19854_ ;
	wire _w19853_ ;
	wire _w19852_ ;
	wire _w19851_ ;
	wire _w19850_ ;
	wire _w19849_ ;
	wire _w19848_ ;
	wire _w19847_ ;
	wire _w19846_ ;
	wire _w19845_ ;
	wire _w19844_ ;
	wire _w19843_ ;
	wire _w19842_ ;
	wire _w19841_ ;
	wire _w19840_ ;
	wire _w19839_ ;
	wire _w19838_ ;
	wire _w19837_ ;
	wire _w19836_ ;
	wire _w19835_ ;
	wire _w19834_ ;
	wire _w19833_ ;
	wire _w19832_ ;
	wire _w19831_ ;
	wire _w19830_ ;
	wire _w19829_ ;
	wire _w19828_ ;
	wire _w19827_ ;
	wire _w19826_ ;
	wire _w19825_ ;
	wire _w19824_ ;
	wire _w19823_ ;
	wire _w19822_ ;
	wire _w19821_ ;
	wire _w19820_ ;
	wire _w19819_ ;
	wire _w19818_ ;
	wire _w19817_ ;
	wire _w19816_ ;
	wire _w19815_ ;
	wire _w19814_ ;
	wire _w19813_ ;
	wire _w19812_ ;
	wire _w19811_ ;
	wire _w19810_ ;
	wire _w19809_ ;
	wire _w19808_ ;
	wire _w19807_ ;
	wire _w19806_ ;
	wire _w19805_ ;
	wire _w19804_ ;
	wire _w19803_ ;
	wire _w19802_ ;
	wire _w19801_ ;
	wire _w19800_ ;
	wire _w19799_ ;
	wire _w19798_ ;
	wire _w19797_ ;
	wire _w19796_ ;
	wire _w19795_ ;
	wire _w19794_ ;
	wire _w19793_ ;
	wire _w19792_ ;
	wire _w19791_ ;
	wire _w19790_ ;
	wire _w19789_ ;
	wire _w19788_ ;
	wire _w19787_ ;
	wire _w19786_ ;
	wire _w19785_ ;
	wire _w19784_ ;
	wire _w19783_ ;
	wire _w19782_ ;
	wire _w19781_ ;
	wire _w19780_ ;
	wire _w19779_ ;
	wire _w19778_ ;
	wire _w19777_ ;
	wire _w19776_ ;
	wire _w19775_ ;
	wire _w19774_ ;
	wire _w19773_ ;
	wire _w19772_ ;
	wire _w19771_ ;
	wire _w19770_ ;
	wire _w19769_ ;
	wire _w19768_ ;
	wire _w19767_ ;
	wire _w19766_ ;
	wire _w19765_ ;
	wire _w19764_ ;
	wire _w19763_ ;
	wire _w19762_ ;
	wire _w19761_ ;
	wire _w19760_ ;
	wire _w19759_ ;
	wire _w19758_ ;
	wire _w19757_ ;
	wire _w19756_ ;
	wire _w19755_ ;
	wire _w19754_ ;
	wire _w19753_ ;
	wire _w19752_ ;
	wire _w19751_ ;
	wire _w19750_ ;
	wire _w19749_ ;
	wire _w19748_ ;
	wire _w19747_ ;
	wire _w19746_ ;
	wire _w19745_ ;
	wire _w19744_ ;
	wire _w19743_ ;
	wire _w19742_ ;
	wire _w19741_ ;
	wire _w19740_ ;
	wire _w19739_ ;
	wire _w19738_ ;
	wire _w19737_ ;
	wire _w19736_ ;
	wire _w19735_ ;
	wire _w19734_ ;
	wire _w19733_ ;
	wire _w19732_ ;
	wire _w19731_ ;
	wire _w19730_ ;
	wire _w19729_ ;
	wire _w19728_ ;
	wire _w19727_ ;
	wire _w19726_ ;
	wire _w19725_ ;
	wire _w19724_ ;
	wire _w19723_ ;
	wire _w19722_ ;
	wire _w19721_ ;
	wire _w19720_ ;
	wire _w19719_ ;
	wire _w19718_ ;
	wire _w19717_ ;
	wire _w19716_ ;
	wire _w19715_ ;
	wire _w19714_ ;
	wire _w19713_ ;
	wire _w19712_ ;
	wire _w19711_ ;
	wire _w19710_ ;
	wire _w19709_ ;
	wire _w19708_ ;
	wire _w19707_ ;
	wire _w19706_ ;
	wire _w19705_ ;
	wire _w19704_ ;
	wire _w19703_ ;
	wire _w19702_ ;
	wire _w19701_ ;
	wire _w19700_ ;
	wire _w19699_ ;
	wire _w19698_ ;
	wire _w19697_ ;
	wire _w19696_ ;
	wire _w19695_ ;
	wire _w19694_ ;
	wire _w19693_ ;
	wire _w19692_ ;
	wire _w19691_ ;
	wire _w19690_ ;
	wire _w19689_ ;
	wire _w19688_ ;
	wire _w19687_ ;
	wire _w19686_ ;
	wire _w19685_ ;
	wire _w19684_ ;
	wire _w19683_ ;
	wire _w19682_ ;
	wire _w19681_ ;
	wire _w19680_ ;
	wire _w19679_ ;
	wire _w19678_ ;
	wire _w19677_ ;
	wire _w19676_ ;
	wire _w19675_ ;
	wire _w19674_ ;
	wire _w19673_ ;
	wire _w19672_ ;
	wire _w19671_ ;
	wire _w19670_ ;
	wire _w19669_ ;
	wire _w19668_ ;
	wire _w19667_ ;
	wire _w19666_ ;
	wire _w19665_ ;
	wire _w19664_ ;
	wire _w19663_ ;
	wire _w19662_ ;
	wire _w19661_ ;
	wire _w19660_ ;
	wire _w19659_ ;
	wire _w19658_ ;
	wire _w19657_ ;
	wire _w19656_ ;
	wire _w19655_ ;
	wire _w19654_ ;
	wire _w19653_ ;
	wire _w19652_ ;
	wire _w19651_ ;
	wire _w19650_ ;
	wire _w19649_ ;
	wire _w19648_ ;
	wire _w19647_ ;
	wire _w19646_ ;
	wire _w19645_ ;
	wire _w19644_ ;
	wire _w19643_ ;
	wire _w19642_ ;
	wire _w19641_ ;
	wire _w19640_ ;
	wire _w19639_ ;
	wire _w19638_ ;
	wire _w19637_ ;
	wire _w19636_ ;
	wire _w19635_ ;
	wire _w19634_ ;
	wire _w19633_ ;
	wire _w19632_ ;
	wire _w19631_ ;
	wire _w19630_ ;
	wire _w19629_ ;
	wire _w19628_ ;
	wire _w19627_ ;
	wire _w19626_ ;
	wire _w19625_ ;
	wire _w19624_ ;
	wire _w19623_ ;
	wire _w19622_ ;
	wire _w19621_ ;
	wire _w19620_ ;
	wire _w19619_ ;
	wire _w19618_ ;
	wire _w19617_ ;
	wire _w19616_ ;
	wire _w19615_ ;
	wire _w19614_ ;
	wire _w19613_ ;
	wire _w19612_ ;
	wire _w19611_ ;
	wire _w19610_ ;
	wire _w19609_ ;
	wire _w19608_ ;
	wire _w19607_ ;
	wire _w19606_ ;
	wire _w19605_ ;
	wire _w19604_ ;
	wire _w19603_ ;
	wire _w19602_ ;
	wire _w19601_ ;
	wire _w19600_ ;
	wire _w19599_ ;
	wire _w19598_ ;
	wire _w19597_ ;
	wire _w19596_ ;
	wire _w19595_ ;
	wire _w19594_ ;
	wire _w19593_ ;
	wire _w19592_ ;
	wire _w19591_ ;
	wire _w19590_ ;
	wire _w19589_ ;
	wire _w19588_ ;
	wire _w19587_ ;
	wire _w19586_ ;
	wire _w19585_ ;
	wire _w19584_ ;
	wire _w19583_ ;
	wire _w19582_ ;
	wire _w19581_ ;
	wire _w19580_ ;
	wire _w19579_ ;
	wire _w19578_ ;
	wire _w19577_ ;
	wire _w19576_ ;
	wire _w19575_ ;
	wire _w19574_ ;
	wire _w19573_ ;
	wire _w19572_ ;
	wire _w19571_ ;
	wire _w19570_ ;
	wire _w19569_ ;
	wire _w19568_ ;
	wire _w19567_ ;
	wire _w19566_ ;
	wire _w19565_ ;
	wire _w19564_ ;
	wire _w19563_ ;
	wire _w19562_ ;
	wire _w19561_ ;
	wire _w19560_ ;
	wire _w19559_ ;
	wire _w19558_ ;
	wire _w19557_ ;
	wire _w19556_ ;
	wire _w19555_ ;
	wire _w19554_ ;
	wire _w19553_ ;
	wire _w19552_ ;
	wire _w19551_ ;
	wire _w19550_ ;
	wire _w19549_ ;
	wire _w19548_ ;
	wire _w19547_ ;
	wire _w19546_ ;
	wire _w19545_ ;
	wire _w19544_ ;
	wire _w19543_ ;
	wire _w19542_ ;
	wire _w19541_ ;
	wire _w19540_ ;
	wire _w19539_ ;
	wire _w19538_ ;
	wire _w19537_ ;
	wire _w19536_ ;
	wire _w19535_ ;
	wire _w19534_ ;
	wire _w19533_ ;
	wire _w19532_ ;
	wire _w19531_ ;
	wire _w19530_ ;
	wire _w19529_ ;
	wire _w19528_ ;
	wire _w19527_ ;
	wire _w19526_ ;
	wire _w19525_ ;
	wire _w19524_ ;
	wire _w19523_ ;
	wire _w19522_ ;
	wire _w19521_ ;
	wire _w19520_ ;
	wire _w19519_ ;
	wire _w19518_ ;
	wire _w19517_ ;
	wire _w19516_ ;
	wire _w19515_ ;
	wire _w19514_ ;
	wire _w19513_ ;
	wire _w19512_ ;
	wire _w19511_ ;
	wire _w19510_ ;
	wire _w19509_ ;
	wire _w19508_ ;
	wire _w19507_ ;
	wire _w19506_ ;
	wire _w19505_ ;
	wire _w19504_ ;
	wire _w19503_ ;
	wire _w19502_ ;
	wire _w19501_ ;
	wire _w19500_ ;
	wire _w19499_ ;
	wire _w19498_ ;
	wire _w19497_ ;
	wire _w19496_ ;
	wire _w19495_ ;
	wire _w19494_ ;
	wire _w19493_ ;
	wire _w19492_ ;
	wire _w19491_ ;
	wire _w19490_ ;
	wire _w19489_ ;
	wire _w19488_ ;
	wire _w19487_ ;
	wire _w19486_ ;
	wire _w19485_ ;
	wire _w19484_ ;
	wire _w19483_ ;
	wire _w19482_ ;
	wire _w19481_ ;
	wire _w19480_ ;
	wire _w19479_ ;
	wire _w19478_ ;
	wire _w19477_ ;
	wire _w19476_ ;
	wire _w19475_ ;
	wire _w19474_ ;
	wire _w19473_ ;
	wire _w19472_ ;
	wire _w19471_ ;
	wire _w19470_ ;
	wire _w19469_ ;
	wire _w19468_ ;
	wire _w19467_ ;
	wire _w19466_ ;
	wire _w19465_ ;
	wire _w19464_ ;
	wire _w19463_ ;
	wire _w19462_ ;
	wire _w19461_ ;
	wire _w19460_ ;
	wire _w19459_ ;
	wire _w19458_ ;
	wire _w19457_ ;
	wire _w19456_ ;
	wire _w19455_ ;
	wire _w19454_ ;
	wire _w19453_ ;
	wire _w19452_ ;
	wire _w19451_ ;
	wire _w19450_ ;
	wire _w19449_ ;
	wire _w19448_ ;
	wire _w19447_ ;
	wire _w19446_ ;
	wire _w19445_ ;
	wire _w19444_ ;
	wire _w19443_ ;
	wire _w19442_ ;
	wire _w19441_ ;
	wire _w19440_ ;
	wire _w19439_ ;
	wire _w19438_ ;
	wire _w19437_ ;
	wire _w19436_ ;
	wire _w19435_ ;
	wire _w19434_ ;
	wire _w19433_ ;
	wire _w19432_ ;
	wire _w19431_ ;
	wire _w19430_ ;
	wire _w19429_ ;
	wire _w19428_ ;
	wire _w19427_ ;
	wire _w19426_ ;
	wire _w19425_ ;
	wire _w19424_ ;
	wire _w19423_ ;
	wire _w19422_ ;
	wire _w19421_ ;
	wire _w19420_ ;
	wire _w19419_ ;
	wire _w19418_ ;
	wire _w19417_ ;
	wire _w19416_ ;
	wire _w19415_ ;
	wire _w19414_ ;
	wire _w19413_ ;
	wire _w19412_ ;
	wire _w19411_ ;
	wire _w19410_ ;
	wire _w19409_ ;
	wire _w19408_ ;
	wire _w19407_ ;
	wire _w19406_ ;
	wire _w19405_ ;
	wire _w19404_ ;
	wire _w19403_ ;
	wire _w19402_ ;
	wire _w19401_ ;
	wire _w19400_ ;
	wire _w19399_ ;
	wire _w19398_ ;
	wire _w19397_ ;
	wire _w19396_ ;
	wire _w19395_ ;
	wire _w19394_ ;
	wire _w19393_ ;
	wire _w19392_ ;
	wire _w19391_ ;
	wire _w19390_ ;
	wire _w19389_ ;
	wire _w19388_ ;
	wire _w19387_ ;
	wire _w19386_ ;
	wire _w19385_ ;
	wire _w19384_ ;
	wire _w19383_ ;
	wire _w19382_ ;
	wire _w19381_ ;
	wire _w19380_ ;
	wire _w19379_ ;
	wire _w19378_ ;
	wire _w19377_ ;
	wire _w19376_ ;
	wire _w19375_ ;
	wire _w19374_ ;
	wire _w19373_ ;
	wire _w19372_ ;
	wire _w19371_ ;
	wire _w19370_ ;
	wire _w19369_ ;
	wire _w19368_ ;
	wire _w19367_ ;
	wire _w19366_ ;
	wire _w19365_ ;
	wire _w19364_ ;
	wire _w19363_ ;
	wire _w19362_ ;
	wire _w19361_ ;
	wire _w19360_ ;
	wire _w19359_ ;
	wire _w19358_ ;
	wire _w19357_ ;
	wire _w19356_ ;
	wire _w19355_ ;
	wire _w19354_ ;
	wire _w19353_ ;
	wire _w19352_ ;
	wire _w19351_ ;
	wire _w19350_ ;
	wire _w19349_ ;
	wire _w19348_ ;
	wire _w19347_ ;
	wire _w19346_ ;
	wire _w19345_ ;
	wire _w19344_ ;
	wire _w19343_ ;
	wire _w19342_ ;
	wire _w19341_ ;
	wire _w19340_ ;
	wire _w19339_ ;
	wire _w19338_ ;
	wire _w19337_ ;
	wire _w19336_ ;
	wire _w19335_ ;
	wire _w19334_ ;
	wire _w19333_ ;
	wire _w19332_ ;
	wire _w19331_ ;
	wire _w19330_ ;
	wire _w19329_ ;
	wire _w19328_ ;
	wire _w19327_ ;
	wire _w19326_ ;
	wire _w19325_ ;
	wire _w19324_ ;
	wire _w19323_ ;
	wire _w19322_ ;
	wire _w19321_ ;
	wire _w19320_ ;
	wire _w19319_ ;
	wire _w19318_ ;
	wire _w19317_ ;
	wire _w19316_ ;
	wire _w19315_ ;
	wire _w19314_ ;
	wire _w19313_ ;
	wire _w19312_ ;
	wire _w19311_ ;
	wire _w19310_ ;
	wire _w19309_ ;
	wire _w19308_ ;
	wire _w19307_ ;
	wire _w19306_ ;
	wire _w19305_ ;
	wire _w19304_ ;
	wire _w19303_ ;
	wire _w19302_ ;
	wire _w19301_ ;
	wire _w19300_ ;
	wire _w19299_ ;
	wire _w19298_ ;
	wire _w19297_ ;
	wire _w19296_ ;
	wire _w19295_ ;
	wire _w19294_ ;
	wire _w19293_ ;
	wire _w19292_ ;
	wire _w19291_ ;
	wire _w19290_ ;
	wire _w19289_ ;
	wire _w19288_ ;
	wire _w19287_ ;
	wire _w19286_ ;
	wire _w19285_ ;
	wire _w19284_ ;
	wire _w19283_ ;
	wire _w19282_ ;
	wire _w19281_ ;
	wire _w19280_ ;
	wire _w19279_ ;
	wire _w19278_ ;
	wire _w19277_ ;
	wire _w19276_ ;
	wire _w19275_ ;
	wire _w19274_ ;
	wire _w19273_ ;
	wire _w19272_ ;
	wire _w19271_ ;
	wire _w19270_ ;
	wire _w19269_ ;
	wire _w19268_ ;
	wire _w19267_ ;
	wire _w19266_ ;
	wire _w19265_ ;
	wire _w19264_ ;
	wire _w19263_ ;
	wire _w19262_ ;
	wire _w19261_ ;
	wire _w19260_ ;
	wire _w19259_ ;
	wire _w19258_ ;
	wire _w19257_ ;
	wire _w19256_ ;
	wire _w19255_ ;
	wire _w19254_ ;
	wire _w19253_ ;
	wire _w19252_ ;
	wire _w19251_ ;
	wire _w19250_ ;
	wire _w19249_ ;
	wire _w19248_ ;
	wire _w19247_ ;
	wire _w19246_ ;
	wire _w19245_ ;
	wire _w19244_ ;
	wire _w19243_ ;
	wire _w19242_ ;
	wire _w19241_ ;
	wire _w19240_ ;
	wire _w19239_ ;
	wire _w19238_ ;
	wire _w19237_ ;
	wire _w19236_ ;
	wire _w19235_ ;
	wire _w19234_ ;
	wire _w19233_ ;
	wire _w19232_ ;
	wire _w19231_ ;
	wire _w19230_ ;
	wire _w19229_ ;
	wire _w19228_ ;
	wire _w19227_ ;
	wire _w19226_ ;
	wire _w19225_ ;
	wire _w19224_ ;
	wire _w19223_ ;
	wire _w19222_ ;
	wire _w19221_ ;
	wire _w19220_ ;
	wire _w19219_ ;
	wire _w19218_ ;
	wire _w19217_ ;
	wire _w19216_ ;
	wire _w19215_ ;
	wire _w19214_ ;
	wire _w19213_ ;
	wire _w19212_ ;
	wire _w19211_ ;
	wire _w19210_ ;
	wire _w19209_ ;
	wire _w19208_ ;
	wire _w19207_ ;
	wire _w19206_ ;
	wire _w19205_ ;
	wire _w19204_ ;
	wire _w19203_ ;
	wire _w19202_ ;
	wire _w19201_ ;
	wire _w19200_ ;
	wire _w19199_ ;
	wire _w19198_ ;
	wire _w19197_ ;
	wire _w19196_ ;
	wire _w19195_ ;
	wire _w19194_ ;
	wire _w19193_ ;
	wire _w19192_ ;
	wire _w19191_ ;
	wire _w19190_ ;
	wire _w19189_ ;
	wire _w19188_ ;
	wire _w19187_ ;
	wire _w19186_ ;
	wire _w19185_ ;
	wire _w19184_ ;
	wire _w19183_ ;
	wire _w19182_ ;
	wire _w19181_ ;
	wire _w19180_ ;
	wire _w19179_ ;
	wire _w19178_ ;
	wire _w19177_ ;
	wire _w19176_ ;
	wire _w19175_ ;
	wire _w19174_ ;
	wire _w19173_ ;
	wire _w19172_ ;
	wire _w19171_ ;
	wire _w19170_ ;
	wire _w19169_ ;
	wire _w19168_ ;
	wire _w19167_ ;
	wire _w19166_ ;
	wire _w19165_ ;
	wire _w19164_ ;
	wire _w19163_ ;
	wire _w19162_ ;
	wire _w19161_ ;
	wire _w19160_ ;
	wire _w19159_ ;
	wire _w19158_ ;
	wire _w19157_ ;
	wire _w19156_ ;
	wire _w19155_ ;
	wire _w19154_ ;
	wire _w19153_ ;
	wire _w19152_ ;
	wire _w19151_ ;
	wire _w19150_ ;
	wire _w19149_ ;
	wire _w19148_ ;
	wire _w19147_ ;
	wire _w19146_ ;
	wire _w19145_ ;
	wire _w19144_ ;
	wire _w19143_ ;
	wire _w19142_ ;
	wire _w19141_ ;
	wire _w19140_ ;
	wire _w19139_ ;
	wire _w19138_ ;
	wire _w19137_ ;
	wire _w19136_ ;
	wire _w19135_ ;
	wire _w19134_ ;
	wire _w19133_ ;
	wire _w19132_ ;
	wire _w19131_ ;
	wire _w19130_ ;
	wire _w19129_ ;
	wire _w19128_ ;
	wire _w19127_ ;
	wire _w19126_ ;
	wire _w19125_ ;
	wire _w19124_ ;
	wire _w19123_ ;
	wire _w19122_ ;
	wire _w19121_ ;
	wire _w19120_ ;
	wire _w19119_ ;
	wire _w19118_ ;
	wire _w19117_ ;
	wire _w19116_ ;
	wire _w19115_ ;
	wire _w19114_ ;
	wire _w19113_ ;
	wire _w19112_ ;
	wire _w19111_ ;
	wire _w19110_ ;
	wire _w19109_ ;
	wire _w19108_ ;
	wire _w19107_ ;
	wire _w19106_ ;
	wire _w19105_ ;
	wire _w19104_ ;
	wire _w19103_ ;
	wire _w19102_ ;
	wire _w19101_ ;
	wire _w19100_ ;
	wire _w19099_ ;
	wire _w19098_ ;
	wire _w19097_ ;
	wire _w19096_ ;
	wire _w19095_ ;
	wire _w19094_ ;
	wire _w19093_ ;
	wire _w19092_ ;
	wire _w19091_ ;
	wire _w19090_ ;
	wire _w19089_ ;
	wire _w19088_ ;
	wire _w19087_ ;
	wire _w19086_ ;
	wire _w19085_ ;
	wire _w19084_ ;
	wire _w19083_ ;
	wire _w19082_ ;
	wire _w19081_ ;
	wire _w19080_ ;
	wire _w19079_ ;
	wire _w19078_ ;
	wire _w19077_ ;
	wire _w19076_ ;
	wire _w19075_ ;
	wire _w19074_ ;
	wire _w19073_ ;
	wire _w19072_ ;
	wire _w19071_ ;
	wire _w19070_ ;
	wire _w19069_ ;
	wire _w19068_ ;
	wire _w19067_ ;
	wire _w19066_ ;
	wire _w19065_ ;
	wire _w19064_ ;
	wire _w19063_ ;
	wire _w19062_ ;
	wire _w19061_ ;
	wire _w19060_ ;
	wire _w19059_ ;
	wire _w19058_ ;
	wire _w19057_ ;
	wire _w19056_ ;
	wire _w19055_ ;
	wire _w19054_ ;
	wire _w19053_ ;
	wire _w19052_ ;
	wire _w19051_ ;
	wire _w19050_ ;
	wire _w19049_ ;
	wire _w19048_ ;
	wire _w19047_ ;
	wire _w19046_ ;
	wire _w19045_ ;
	wire _w19044_ ;
	wire _w19043_ ;
	wire _w19042_ ;
	wire _w19041_ ;
	wire _w19040_ ;
	wire _w19039_ ;
	wire _w19038_ ;
	wire _w19037_ ;
	wire _w19036_ ;
	wire _w19035_ ;
	wire _w19034_ ;
	wire _w19033_ ;
	wire _w19032_ ;
	wire _w19031_ ;
	wire _w19030_ ;
	wire _w19029_ ;
	wire _w19028_ ;
	wire _w19027_ ;
	wire _w19026_ ;
	wire _w19025_ ;
	wire _w19024_ ;
	wire _w19023_ ;
	wire _w19022_ ;
	wire _w19021_ ;
	wire _w19020_ ;
	wire _w19019_ ;
	wire _w19018_ ;
	wire _w19017_ ;
	wire _w19016_ ;
	wire _w19015_ ;
	wire _w19014_ ;
	wire _w19013_ ;
	wire _w19012_ ;
	wire _w19011_ ;
	wire _w19010_ ;
	wire _w19009_ ;
	wire _w19008_ ;
	wire _w19007_ ;
	wire _w19006_ ;
	wire _w19005_ ;
	wire _w19004_ ;
	wire _w19003_ ;
	wire _w19002_ ;
	wire _w19001_ ;
	wire _w19000_ ;
	wire _w18999_ ;
	wire _w18998_ ;
	wire _w18997_ ;
	wire _w18996_ ;
	wire _w18995_ ;
	wire _w18994_ ;
	wire _w18993_ ;
	wire _w18992_ ;
	wire _w18991_ ;
	wire _w18990_ ;
	wire _w18989_ ;
	wire _w18988_ ;
	wire _w18987_ ;
	wire _w18986_ ;
	wire _w18985_ ;
	wire _w18984_ ;
	wire _w18983_ ;
	wire _w18982_ ;
	wire _w18981_ ;
	wire _w18980_ ;
	wire _w18979_ ;
	wire _w18978_ ;
	wire _w18977_ ;
	wire _w18976_ ;
	wire _w18975_ ;
	wire _w18974_ ;
	wire _w18973_ ;
	wire _w18972_ ;
	wire _w18971_ ;
	wire _w18970_ ;
	wire _w18969_ ;
	wire _w18968_ ;
	wire _w18967_ ;
	wire _w18966_ ;
	wire _w18965_ ;
	wire _w18964_ ;
	wire _w18963_ ;
	wire _w18962_ ;
	wire _w18961_ ;
	wire _w18960_ ;
	wire _w18959_ ;
	wire _w18958_ ;
	wire _w18957_ ;
	wire _w18956_ ;
	wire _w18955_ ;
	wire _w18954_ ;
	wire _w18953_ ;
	wire _w18952_ ;
	wire _w18951_ ;
	wire _w18950_ ;
	wire _w18949_ ;
	wire _w18948_ ;
	wire _w18947_ ;
	wire _w18946_ ;
	wire _w18945_ ;
	wire _w18944_ ;
	wire _w18943_ ;
	wire _w18942_ ;
	wire _w18941_ ;
	wire _w18940_ ;
	wire _w18939_ ;
	wire _w18938_ ;
	wire _w18937_ ;
	wire _w18936_ ;
	wire _w18935_ ;
	wire _w18934_ ;
	wire _w18933_ ;
	wire _w18932_ ;
	wire _w18931_ ;
	wire _w18930_ ;
	wire _w18929_ ;
	wire _w18928_ ;
	wire _w18927_ ;
	wire _w18926_ ;
	wire _w18925_ ;
	wire _w18924_ ;
	wire _w18923_ ;
	wire _w18922_ ;
	wire _w18921_ ;
	wire _w18920_ ;
	wire _w18919_ ;
	wire _w18918_ ;
	wire _w18917_ ;
	wire _w18916_ ;
	wire _w18915_ ;
	wire _w18914_ ;
	wire _w18913_ ;
	wire _w18912_ ;
	wire _w18911_ ;
	wire _w18910_ ;
	wire _w18909_ ;
	wire _w18908_ ;
	wire _w18907_ ;
	wire _w18906_ ;
	wire _w18905_ ;
	wire _w18904_ ;
	wire _w18903_ ;
	wire _w18902_ ;
	wire _w18901_ ;
	wire _w18900_ ;
	wire _w18899_ ;
	wire _w18898_ ;
	wire _w18897_ ;
	wire _w18896_ ;
	wire _w18895_ ;
	wire _w18894_ ;
	wire _w18893_ ;
	wire _w18892_ ;
	wire _w18891_ ;
	wire _w18890_ ;
	wire _w18889_ ;
	wire _w18888_ ;
	wire _w18887_ ;
	wire _w18886_ ;
	wire _w18885_ ;
	wire _w18884_ ;
	wire _w18883_ ;
	wire _w18882_ ;
	wire _w18881_ ;
	wire _w18880_ ;
	wire _w18879_ ;
	wire _w18878_ ;
	wire _w18877_ ;
	wire _w18876_ ;
	wire _w18875_ ;
	wire _w18874_ ;
	wire _w18873_ ;
	wire _w18872_ ;
	wire _w18871_ ;
	wire _w18870_ ;
	wire _w18869_ ;
	wire _w18868_ ;
	wire _w18867_ ;
	wire _w18866_ ;
	wire _w18865_ ;
	wire _w18864_ ;
	wire _w18863_ ;
	wire _w18862_ ;
	wire _w18861_ ;
	wire _w18860_ ;
	wire _w18859_ ;
	wire _w18858_ ;
	wire _w18857_ ;
	wire _w18856_ ;
	wire _w18855_ ;
	wire _w18854_ ;
	wire _w18853_ ;
	wire _w18852_ ;
	wire _w18851_ ;
	wire _w18850_ ;
	wire _w18849_ ;
	wire _w18848_ ;
	wire _w18847_ ;
	wire _w18846_ ;
	wire _w18845_ ;
	wire _w18844_ ;
	wire _w18843_ ;
	wire _w18842_ ;
	wire _w18841_ ;
	wire _w18840_ ;
	wire _w18839_ ;
	wire _w18838_ ;
	wire _w18837_ ;
	wire _w18836_ ;
	wire _w18835_ ;
	wire _w18834_ ;
	wire _w18833_ ;
	wire _w18832_ ;
	wire _w18831_ ;
	wire _w18830_ ;
	wire _w18829_ ;
	wire _w18828_ ;
	wire _w18827_ ;
	wire _w18826_ ;
	wire _w18825_ ;
	wire _w18824_ ;
	wire _w18823_ ;
	wire _w18822_ ;
	wire _w18821_ ;
	wire _w18820_ ;
	wire _w18819_ ;
	wire _w18818_ ;
	wire _w18817_ ;
	wire _w18816_ ;
	wire _w18815_ ;
	wire _w18814_ ;
	wire _w18813_ ;
	wire _w18812_ ;
	wire _w18811_ ;
	wire _w18810_ ;
	wire _w18809_ ;
	wire _w18808_ ;
	wire _w18807_ ;
	wire _w18806_ ;
	wire _w18805_ ;
	wire _w18804_ ;
	wire _w18803_ ;
	wire _w18802_ ;
	wire _w18801_ ;
	wire _w18800_ ;
	wire _w18799_ ;
	wire _w18798_ ;
	wire _w18797_ ;
	wire _w18796_ ;
	wire _w18795_ ;
	wire _w18794_ ;
	wire _w18793_ ;
	wire _w18792_ ;
	wire _w18791_ ;
	wire _w18790_ ;
	wire _w18789_ ;
	wire _w18788_ ;
	wire _w18787_ ;
	wire _w18786_ ;
	wire _w18785_ ;
	wire _w18784_ ;
	wire _w18783_ ;
	wire _w18782_ ;
	wire _w18781_ ;
	wire _w18780_ ;
	wire _w18779_ ;
	wire _w18778_ ;
	wire _w18777_ ;
	wire _w18776_ ;
	wire _w18775_ ;
	wire _w18774_ ;
	wire _w18773_ ;
	wire _w18772_ ;
	wire _w18771_ ;
	wire _w18770_ ;
	wire _w18769_ ;
	wire _w18768_ ;
	wire _w18767_ ;
	wire _w18766_ ;
	wire _w18765_ ;
	wire _w18764_ ;
	wire _w18763_ ;
	wire _w18762_ ;
	wire _w18761_ ;
	wire _w18760_ ;
	wire _w18759_ ;
	wire _w18758_ ;
	wire _w18757_ ;
	wire _w18756_ ;
	wire _w18755_ ;
	wire _w18754_ ;
	wire _w18753_ ;
	wire _w18752_ ;
	wire _w18751_ ;
	wire _w18750_ ;
	wire _w18749_ ;
	wire _w18748_ ;
	wire _w18747_ ;
	wire _w18746_ ;
	wire _w18745_ ;
	wire _w18744_ ;
	wire _w18743_ ;
	wire _w18742_ ;
	wire _w18741_ ;
	wire _w18740_ ;
	wire _w18739_ ;
	wire _w18738_ ;
	wire _w18737_ ;
	wire _w18736_ ;
	wire _w18735_ ;
	wire _w18734_ ;
	wire _w18733_ ;
	wire _w18732_ ;
	wire _w18731_ ;
	wire _w18730_ ;
	wire _w18729_ ;
	wire _w18728_ ;
	wire _w18727_ ;
	wire _w18726_ ;
	wire _w18725_ ;
	wire _w18724_ ;
	wire _w18723_ ;
	wire _w18722_ ;
	wire _w18721_ ;
	wire _w18720_ ;
	wire _w18719_ ;
	wire _w18718_ ;
	wire _w18717_ ;
	wire _w18716_ ;
	wire _w18715_ ;
	wire _w18714_ ;
	wire _w18713_ ;
	wire _w18712_ ;
	wire _w18711_ ;
	wire _w18710_ ;
	wire _w18709_ ;
	wire _w18708_ ;
	wire _w18707_ ;
	wire _w18706_ ;
	wire _w18705_ ;
	wire _w18704_ ;
	wire _w18703_ ;
	wire _w18702_ ;
	wire _w18701_ ;
	wire _w18700_ ;
	wire _w18699_ ;
	wire _w18698_ ;
	wire _w18697_ ;
	wire _w18696_ ;
	wire _w18695_ ;
	wire _w18694_ ;
	wire _w18693_ ;
	wire _w18692_ ;
	wire _w18691_ ;
	wire _w18690_ ;
	wire _w18689_ ;
	wire _w18688_ ;
	wire _w18687_ ;
	wire _w18686_ ;
	wire _w18685_ ;
	wire _w18684_ ;
	wire _w18683_ ;
	wire _w18682_ ;
	wire _w18681_ ;
	wire _w18680_ ;
	wire _w18679_ ;
	wire _w18678_ ;
	wire _w18677_ ;
	wire _w18676_ ;
	wire _w18675_ ;
	wire _w18674_ ;
	wire _w18673_ ;
	wire _w18672_ ;
	wire _w18671_ ;
	wire _w18670_ ;
	wire _w18669_ ;
	wire _w18668_ ;
	wire _w18667_ ;
	wire _w18666_ ;
	wire _w18665_ ;
	wire _w18664_ ;
	wire _w18663_ ;
	wire _w18662_ ;
	wire _w18661_ ;
	wire _w18660_ ;
	wire _w18659_ ;
	wire _w18658_ ;
	wire _w18657_ ;
	wire _w18656_ ;
	wire _w18655_ ;
	wire _w18654_ ;
	wire _w18653_ ;
	wire _w18652_ ;
	wire _w18651_ ;
	wire _w18650_ ;
	wire _w18649_ ;
	wire _w18648_ ;
	wire _w18647_ ;
	wire _w18646_ ;
	wire _w18645_ ;
	wire _w18644_ ;
	wire _w18643_ ;
	wire _w18642_ ;
	wire _w18641_ ;
	wire _w18640_ ;
	wire _w18639_ ;
	wire _w18638_ ;
	wire _w18637_ ;
	wire _w18636_ ;
	wire _w18635_ ;
	wire _w18634_ ;
	wire _w18633_ ;
	wire _w18632_ ;
	wire _w18631_ ;
	wire _w18630_ ;
	wire _w18629_ ;
	wire _w18628_ ;
	wire _w18627_ ;
	wire _w18626_ ;
	wire _w18625_ ;
	wire _w18624_ ;
	wire _w18623_ ;
	wire _w18622_ ;
	wire _w18621_ ;
	wire _w18620_ ;
	wire _w18619_ ;
	wire _w18618_ ;
	wire _w18617_ ;
	wire _w18616_ ;
	wire _w18615_ ;
	wire _w18614_ ;
	wire _w18613_ ;
	wire _w18612_ ;
	wire _w18611_ ;
	wire _w18610_ ;
	wire _w18609_ ;
	wire _w18608_ ;
	wire _w18607_ ;
	wire _w18606_ ;
	wire _w18605_ ;
	wire _w18604_ ;
	wire _w18603_ ;
	wire _w18602_ ;
	wire _w18601_ ;
	wire _w18600_ ;
	wire _w18599_ ;
	wire _w18598_ ;
	wire _w18597_ ;
	wire _w18596_ ;
	wire _w18595_ ;
	wire _w18594_ ;
	wire _w18593_ ;
	wire _w18592_ ;
	wire _w18591_ ;
	wire _w18590_ ;
	wire _w18589_ ;
	wire _w18588_ ;
	wire _w18587_ ;
	wire _w18586_ ;
	wire _w18585_ ;
	wire _w18584_ ;
	wire _w18583_ ;
	wire _w18582_ ;
	wire _w18581_ ;
	wire _w18580_ ;
	wire _w18579_ ;
	wire _w18578_ ;
	wire _w18577_ ;
	wire _w18576_ ;
	wire _w18575_ ;
	wire _w18574_ ;
	wire _w18573_ ;
	wire _w18572_ ;
	wire _w18571_ ;
	wire _w18570_ ;
	wire _w18569_ ;
	wire _w18568_ ;
	wire _w18567_ ;
	wire _w18566_ ;
	wire _w18565_ ;
	wire _w18564_ ;
	wire _w18563_ ;
	wire _w18562_ ;
	wire _w18561_ ;
	wire _w18560_ ;
	wire _w18559_ ;
	wire _w18558_ ;
	wire _w18557_ ;
	wire _w18556_ ;
	wire _w18555_ ;
	wire _w18554_ ;
	wire _w18553_ ;
	wire _w18552_ ;
	wire _w18551_ ;
	wire _w18550_ ;
	wire _w18549_ ;
	wire _w18548_ ;
	wire _w18547_ ;
	wire _w18546_ ;
	wire _w18545_ ;
	wire _w18544_ ;
	wire _w18543_ ;
	wire _w18542_ ;
	wire _w18541_ ;
	wire _w18540_ ;
	wire _w18539_ ;
	wire _w18538_ ;
	wire _w18537_ ;
	wire _w18536_ ;
	wire _w18535_ ;
	wire _w18534_ ;
	wire _w18533_ ;
	wire _w18532_ ;
	wire _w18531_ ;
	wire _w18530_ ;
	wire _w18529_ ;
	wire _w18528_ ;
	wire _w18527_ ;
	wire _w18526_ ;
	wire _w18525_ ;
	wire _w18524_ ;
	wire _w18523_ ;
	wire _w18522_ ;
	wire _w18521_ ;
	wire _w18520_ ;
	wire _w18519_ ;
	wire _w18518_ ;
	wire _w18517_ ;
	wire _w18516_ ;
	wire _w18515_ ;
	wire _w18514_ ;
	wire _w18513_ ;
	wire _w18512_ ;
	wire _w18511_ ;
	wire _w18510_ ;
	wire _w18509_ ;
	wire _w18508_ ;
	wire _w18507_ ;
	wire _w18506_ ;
	wire _w18505_ ;
	wire _w18504_ ;
	wire _w18503_ ;
	wire _w18502_ ;
	wire _w18501_ ;
	wire _w18500_ ;
	wire _w18499_ ;
	wire _w18498_ ;
	wire _w18497_ ;
	wire _w18496_ ;
	wire _w18495_ ;
	wire _w18494_ ;
	wire _w18493_ ;
	wire _w18492_ ;
	wire _w18491_ ;
	wire _w18490_ ;
	wire _w18489_ ;
	wire _w18488_ ;
	wire _w18487_ ;
	wire _w18486_ ;
	wire _w18485_ ;
	wire _w18484_ ;
	wire _w18483_ ;
	wire _w18482_ ;
	wire _w18481_ ;
	wire _w18480_ ;
	wire _w18479_ ;
	wire _w18478_ ;
	wire _w18477_ ;
	wire _w18476_ ;
	wire _w18475_ ;
	wire _w18474_ ;
	wire _w18473_ ;
	wire _w18472_ ;
	wire _w18471_ ;
	wire _w18470_ ;
	wire _w18469_ ;
	wire _w18468_ ;
	wire _w18467_ ;
	wire _w18466_ ;
	wire _w18465_ ;
	wire _w18464_ ;
	wire _w18463_ ;
	wire _w18462_ ;
	wire _w18461_ ;
	wire _w18460_ ;
	wire _w18459_ ;
	wire _w18458_ ;
	wire _w18457_ ;
	wire _w18456_ ;
	wire _w18455_ ;
	wire _w18454_ ;
	wire _w18453_ ;
	wire _w18452_ ;
	wire _w18451_ ;
	wire _w18450_ ;
	wire _w18449_ ;
	wire _w18448_ ;
	wire _w18447_ ;
	wire _w18446_ ;
	wire _w18445_ ;
	wire _w18444_ ;
	wire _w18443_ ;
	wire _w18442_ ;
	wire _w18441_ ;
	wire _w18440_ ;
	wire _w18439_ ;
	wire _w18438_ ;
	wire _w18437_ ;
	wire _w18436_ ;
	wire _w18435_ ;
	wire _w18434_ ;
	wire _w18433_ ;
	wire _w18432_ ;
	wire _w18431_ ;
	wire _w18430_ ;
	wire _w18429_ ;
	wire _w18428_ ;
	wire _w18427_ ;
	wire _w18426_ ;
	wire _w18425_ ;
	wire _w18424_ ;
	wire _w18423_ ;
	wire _w18422_ ;
	wire _w18421_ ;
	wire _w18420_ ;
	wire _w18419_ ;
	wire _w18418_ ;
	wire _w18417_ ;
	wire _w18416_ ;
	wire _w18415_ ;
	wire _w18414_ ;
	wire _w18413_ ;
	wire _w18412_ ;
	wire _w18411_ ;
	wire _w18410_ ;
	wire _w18409_ ;
	wire _w18408_ ;
	wire _w18407_ ;
	wire _w18406_ ;
	wire _w18405_ ;
	wire _w18404_ ;
	wire _w18403_ ;
	wire _w18402_ ;
	wire _w18401_ ;
	wire _w18400_ ;
	wire _w18399_ ;
	wire _w18398_ ;
	wire _w18397_ ;
	wire _w18396_ ;
	wire _w18395_ ;
	wire _w18394_ ;
	wire _w18393_ ;
	wire _w18392_ ;
	wire _w18391_ ;
	wire _w18390_ ;
	wire _w18389_ ;
	wire _w18388_ ;
	wire _w18387_ ;
	wire _w18386_ ;
	wire _w18385_ ;
	wire _w18384_ ;
	wire _w18383_ ;
	wire _w18382_ ;
	wire _w18381_ ;
	wire _w18380_ ;
	wire _w18379_ ;
	wire _w18378_ ;
	wire _w18377_ ;
	wire _w18376_ ;
	wire _w18375_ ;
	wire _w18374_ ;
	wire _w18373_ ;
	wire _w18372_ ;
	wire _w18371_ ;
	wire _w18370_ ;
	wire _w18369_ ;
	wire _w18368_ ;
	wire _w18367_ ;
	wire _w18366_ ;
	wire _w18365_ ;
	wire _w18364_ ;
	wire _w18363_ ;
	wire _w18362_ ;
	wire _w18361_ ;
	wire _w18360_ ;
	wire _w18359_ ;
	wire _w18358_ ;
	wire _w18357_ ;
	wire _w18356_ ;
	wire _w18355_ ;
	wire _w18354_ ;
	wire _w18353_ ;
	wire _w18352_ ;
	wire _w18351_ ;
	wire _w18350_ ;
	wire _w18349_ ;
	wire _w18348_ ;
	wire _w18347_ ;
	wire _w18346_ ;
	wire _w18345_ ;
	wire _w18344_ ;
	wire _w18343_ ;
	wire _w18342_ ;
	wire _w18341_ ;
	wire _w18340_ ;
	wire _w18339_ ;
	wire _w18338_ ;
	wire _w18337_ ;
	wire _w18336_ ;
	wire _w18335_ ;
	wire _w18334_ ;
	wire _w18333_ ;
	wire _w18332_ ;
	wire _w18331_ ;
	wire _w18330_ ;
	wire _w18329_ ;
	wire _w18328_ ;
	wire _w18327_ ;
	wire _w18326_ ;
	wire _w18325_ ;
	wire _w18324_ ;
	wire _w18323_ ;
	wire _w18322_ ;
	wire _w18321_ ;
	wire _w18320_ ;
	wire _w18319_ ;
	wire _w18318_ ;
	wire _w18317_ ;
	wire _w18316_ ;
	wire _w18315_ ;
	wire _w18314_ ;
	wire _w18313_ ;
	wire _w18312_ ;
	wire _w18311_ ;
	wire _w18310_ ;
	wire _w18309_ ;
	wire _w18308_ ;
	wire _w18307_ ;
	wire _w18306_ ;
	wire _w18305_ ;
	wire _w18304_ ;
	wire _w18303_ ;
	wire _w18302_ ;
	wire _w18301_ ;
	wire _w18300_ ;
	wire _w18299_ ;
	wire _w18298_ ;
	wire _w18297_ ;
	wire _w18296_ ;
	wire _w18295_ ;
	wire _w18294_ ;
	wire _w18293_ ;
	wire _w18292_ ;
	wire _w18291_ ;
	wire _w18290_ ;
	wire _w18289_ ;
	wire _w18288_ ;
	wire _w18287_ ;
	wire _w18286_ ;
	wire _w18285_ ;
	wire _w18284_ ;
	wire _w18283_ ;
	wire _w18282_ ;
	wire _w18281_ ;
	wire _w18280_ ;
	wire _w18279_ ;
	wire _w18278_ ;
	wire _w18277_ ;
	wire _w18276_ ;
	wire _w18275_ ;
	wire _w18274_ ;
	wire _w18273_ ;
	wire _w18272_ ;
	wire _w18271_ ;
	wire _w18270_ ;
	wire _w18269_ ;
	wire _w18268_ ;
	wire _w18267_ ;
	wire _w18266_ ;
	wire _w18265_ ;
	wire _w18264_ ;
	wire _w18263_ ;
	wire _w18262_ ;
	wire _w18261_ ;
	wire _w18260_ ;
	wire _w18259_ ;
	wire _w18258_ ;
	wire _w18257_ ;
	wire _w18256_ ;
	wire _w18255_ ;
	wire _w18254_ ;
	wire _w18253_ ;
	wire _w18252_ ;
	wire _w18251_ ;
	wire _w18250_ ;
	wire _w18249_ ;
	wire _w18248_ ;
	wire _w18247_ ;
	wire _w18246_ ;
	wire _w18245_ ;
	wire _w18244_ ;
	wire _w18243_ ;
	wire _w18242_ ;
	wire _w18241_ ;
	wire _w18240_ ;
	wire _w18239_ ;
	wire _w18238_ ;
	wire _w18237_ ;
	wire _w18236_ ;
	wire _w18235_ ;
	wire _w18234_ ;
	wire _w18233_ ;
	wire _w18232_ ;
	wire _w18231_ ;
	wire _w18230_ ;
	wire _w18229_ ;
	wire _w18228_ ;
	wire _w18227_ ;
	wire _w18226_ ;
	wire _w18225_ ;
	wire _w18224_ ;
	wire _w18223_ ;
	wire _w18222_ ;
	wire _w18221_ ;
	wire _w18220_ ;
	wire _w18219_ ;
	wire _w18218_ ;
	wire _w18217_ ;
	wire _w18216_ ;
	wire _w18215_ ;
	wire _w18214_ ;
	wire _w18213_ ;
	wire _w18212_ ;
	wire _w18211_ ;
	wire _w18210_ ;
	wire _w18209_ ;
	wire _w18208_ ;
	wire _w18207_ ;
	wire _w18206_ ;
	wire _w18205_ ;
	wire _w18204_ ;
	wire _w18203_ ;
	wire _w18202_ ;
	wire _w18201_ ;
	wire _w18200_ ;
	wire _w18199_ ;
	wire _w18198_ ;
	wire _w18197_ ;
	wire _w18196_ ;
	wire _w18195_ ;
	wire _w18194_ ;
	wire _w18193_ ;
	wire _w18192_ ;
	wire _w18191_ ;
	wire _w18190_ ;
	wire _w18189_ ;
	wire _w18188_ ;
	wire _w18187_ ;
	wire _w18186_ ;
	wire _w18185_ ;
	wire _w18184_ ;
	wire _w18183_ ;
	wire _w18182_ ;
	wire _w18181_ ;
	wire _w18180_ ;
	wire _w18179_ ;
	wire _w18178_ ;
	wire _w18177_ ;
	wire _w18176_ ;
	wire _w18175_ ;
	wire _w18174_ ;
	wire _w18173_ ;
	wire _w18172_ ;
	wire _w18171_ ;
	wire _w18170_ ;
	wire _w18169_ ;
	wire _w18168_ ;
	wire _w18167_ ;
	wire _w18166_ ;
	wire _w18165_ ;
	wire _w18164_ ;
	wire _w18163_ ;
	wire _w18162_ ;
	wire _w18161_ ;
	wire _w18160_ ;
	wire _w18159_ ;
	wire _w18158_ ;
	wire _w18157_ ;
	wire _w18156_ ;
	wire _w18155_ ;
	wire _w18154_ ;
	wire _w18153_ ;
	wire _w18152_ ;
	wire _w18151_ ;
	wire _w18150_ ;
	wire _w18149_ ;
	wire _w18148_ ;
	wire _w18147_ ;
	wire _w18146_ ;
	wire _w18145_ ;
	wire _w18144_ ;
	wire _w18143_ ;
	wire _w18142_ ;
	wire _w18141_ ;
	wire _w18140_ ;
	wire _w18139_ ;
	wire _w18138_ ;
	wire _w18137_ ;
	wire _w18136_ ;
	wire _w18135_ ;
	wire _w18134_ ;
	wire _w18133_ ;
	wire _w18132_ ;
	wire _w18131_ ;
	wire _w18130_ ;
	wire _w18129_ ;
	wire _w18128_ ;
	wire _w18127_ ;
	wire _w18126_ ;
	wire _w18125_ ;
	wire _w18124_ ;
	wire _w18123_ ;
	wire _w18122_ ;
	wire _w18121_ ;
	wire _w18120_ ;
	wire _w18119_ ;
	wire _w18118_ ;
	wire _w18117_ ;
	wire _w18116_ ;
	wire _w18115_ ;
	wire _w18114_ ;
	wire _w18113_ ;
	wire _w18112_ ;
	wire _w18111_ ;
	wire _w18110_ ;
	wire _w18109_ ;
	wire _w18108_ ;
	wire _w18107_ ;
	wire _w18106_ ;
	wire _w18105_ ;
	wire _w18104_ ;
	wire _w18103_ ;
	wire _w18102_ ;
	wire _w18101_ ;
	wire _w18100_ ;
	wire _w18099_ ;
	wire _w18098_ ;
	wire _w18097_ ;
	wire _w18096_ ;
	wire _w18095_ ;
	wire _w18094_ ;
	wire _w18093_ ;
	wire _w18092_ ;
	wire _w18091_ ;
	wire _w18090_ ;
	wire _w18089_ ;
	wire _w18088_ ;
	wire _w18087_ ;
	wire _w18086_ ;
	wire _w18085_ ;
	wire _w18084_ ;
	wire _w18083_ ;
	wire _w18082_ ;
	wire _w18081_ ;
	wire _w18080_ ;
	wire _w18079_ ;
	wire _w18078_ ;
	wire _w18077_ ;
	wire _w18076_ ;
	wire _w18075_ ;
	wire _w18074_ ;
	wire _w18073_ ;
	wire _w18072_ ;
	wire _w18071_ ;
	wire _w18070_ ;
	wire _w18069_ ;
	wire _w18068_ ;
	wire _w18067_ ;
	wire _w18066_ ;
	wire _w18065_ ;
	wire _w18064_ ;
	wire _w18063_ ;
	wire _w18062_ ;
	wire _w18061_ ;
	wire _w18060_ ;
	wire _w18059_ ;
	wire _w18058_ ;
	wire _w18057_ ;
	wire _w18056_ ;
	wire _w18055_ ;
	wire _w18054_ ;
	wire _w18053_ ;
	wire _w18052_ ;
	wire _w18051_ ;
	wire _w18050_ ;
	wire _w18049_ ;
	wire _w18048_ ;
	wire _w18047_ ;
	wire _w18046_ ;
	wire _w18045_ ;
	wire _w18044_ ;
	wire _w18043_ ;
	wire _w18042_ ;
	wire _w18041_ ;
	wire _w18040_ ;
	wire _w18039_ ;
	wire _w18038_ ;
	wire _w18037_ ;
	wire _w18036_ ;
	wire _w18035_ ;
	wire _w18034_ ;
	wire _w18033_ ;
	wire _w18032_ ;
	wire _w18031_ ;
	wire _w18030_ ;
	wire _w18029_ ;
	wire _w18028_ ;
	wire _w18027_ ;
	wire _w18026_ ;
	wire _w18025_ ;
	wire _w18024_ ;
	wire _w18023_ ;
	wire _w18022_ ;
	wire _w18021_ ;
	wire _w18020_ ;
	wire _w18019_ ;
	wire _w18018_ ;
	wire _w18017_ ;
	wire _w18016_ ;
	wire _w18015_ ;
	wire _w18014_ ;
	wire _w18013_ ;
	wire _w18012_ ;
	wire _w18011_ ;
	wire _w18010_ ;
	wire _w18009_ ;
	wire _w18008_ ;
	wire _w18007_ ;
	wire _w18006_ ;
	wire _w18005_ ;
	wire _w18004_ ;
	wire _w18003_ ;
	wire _w18002_ ;
	wire _w18001_ ;
	wire _w18000_ ;
	wire _w17999_ ;
	wire _w17998_ ;
	wire _w17997_ ;
	wire _w17996_ ;
	wire _w17995_ ;
	wire _w17994_ ;
	wire _w17993_ ;
	wire _w17992_ ;
	wire _w17991_ ;
	wire _w17990_ ;
	wire _w17989_ ;
	wire _w17988_ ;
	wire _w17987_ ;
	wire _w17986_ ;
	wire _w17985_ ;
	wire _w17984_ ;
	wire _w17983_ ;
	wire _w17982_ ;
	wire _w17981_ ;
	wire _w17980_ ;
	wire _w17979_ ;
	wire _w17978_ ;
	wire _w17977_ ;
	wire _w17976_ ;
	wire _w17975_ ;
	wire _w17974_ ;
	wire _w17973_ ;
	wire _w17972_ ;
	wire _w17971_ ;
	wire _w17970_ ;
	wire _w17969_ ;
	wire _w17968_ ;
	wire _w17967_ ;
	wire _w17966_ ;
	wire _w17965_ ;
	wire _w17964_ ;
	wire _w17963_ ;
	wire _w17962_ ;
	wire _w17961_ ;
	wire _w17960_ ;
	wire _w17959_ ;
	wire _w17958_ ;
	wire _w17957_ ;
	wire _w17956_ ;
	wire _w17955_ ;
	wire _w17954_ ;
	wire _w17953_ ;
	wire _w17952_ ;
	wire _w17951_ ;
	wire _w17950_ ;
	wire _w17949_ ;
	wire _w17948_ ;
	wire _w17947_ ;
	wire _w17946_ ;
	wire _w17945_ ;
	wire _w17944_ ;
	wire _w17943_ ;
	wire _w17942_ ;
	wire _w17941_ ;
	wire _w17940_ ;
	wire _w17939_ ;
	wire _w17938_ ;
	wire _w17937_ ;
	wire _w17936_ ;
	wire _w17935_ ;
	wire _w17934_ ;
	wire _w17933_ ;
	wire _w17932_ ;
	wire _w17931_ ;
	wire _w17930_ ;
	wire _w17929_ ;
	wire _w17928_ ;
	wire _w17927_ ;
	wire _w17926_ ;
	wire _w17925_ ;
	wire _w17924_ ;
	wire _w17923_ ;
	wire _w17922_ ;
	wire _w17921_ ;
	wire _w17920_ ;
	wire _w17919_ ;
	wire _w17918_ ;
	wire _w17917_ ;
	wire _w17916_ ;
	wire _w17915_ ;
	wire _w17914_ ;
	wire _w17913_ ;
	wire _w17912_ ;
	wire _w17911_ ;
	wire _w17910_ ;
	wire _w17909_ ;
	wire _w17908_ ;
	wire _w17907_ ;
	wire _w17906_ ;
	wire _w17905_ ;
	wire _w17904_ ;
	wire _w17903_ ;
	wire _w17902_ ;
	wire _w17901_ ;
	wire _w17900_ ;
	wire _w17899_ ;
	wire _w17898_ ;
	wire _w17897_ ;
	wire _w17896_ ;
	wire _w17895_ ;
	wire _w17894_ ;
	wire _w17893_ ;
	wire _w17892_ ;
	wire _w17891_ ;
	wire _w17890_ ;
	wire _w17889_ ;
	wire _w17888_ ;
	wire _w17887_ ;
	wire _w17886_ ;
	wire _w17885_ ;
	wire _w17884_ ;
	wire _w17883_ ;
	wire _w17882_ ;
	wire _w17881_ ;
	wire _w17880_ ;
	wire _w17879_ ;
	wire _w17878_ ;
	wire _w17877_ ;
	wire _w17876_ ;
	wire _w17875_ ;
	wire _w17874_ ;
	wire _w17873_ ;
	wire _w17872_ ;
	wire _w17871_ ;
	wire _w17870_ ;
	wire _w17869_ ;
	wire _w17868_ ;
	wire _w17867_ ;
	wire _w17866_ ;
	wire _w17865_ ;
	wire _w17864_ ;
	wire _w17863_ ;
	wire _w17862_ ;
	wire _w17861_ ;
	wire _w17860_ ;
	wire _w17859_ ;
	wire _w17858_ ;
	wire _w17857_ ;
	wire _w17856_ ;
	wire _w17855_ ;
	wire _w17854_ ;
	wire _w17853_ ;
	wire _w17852_ ;
	wire _w17851_ ;
	wire _w17850_ ;
	wire _w17849_ ;
	wire _w17848_ ;
	wire _w17847_ ;
	wire _w17846_ ;
	wire _w17845_ ;
	wire _w17844_ ;
	wire _w17843_ ;
	wire _w17842_ ;
	wire _w17841_ ;
	wire _w17840_ ;
	wire _w17839_ ;
	wire _w17838_ ;
	wire _w17837_ ;
	wire _w17836_ ;
	wire _w17835_ ;
	wire _w17834_ ;
	wire _w17833_ ;
	wire _w17832_ ;
	wire _w17831_ ;
	wire _w17830_ ;
	wire _w17829_ ;
	wire _w17828_ ;
	wire _w17827_ ;
	wire _w17826_ ;
	wire _w17825_ ;
	wire _w17824_ ;
	wire _w17823_ ;
	wire _w17822_ ;
	wire _w17821_ ;
	wire _w17820_ ;
	wire _w17819_ ;
	wire _w17818_ ;
	wire _w17817_ ;
	wire _w17816_ ;
	wire _w17815_ ;
	wire _w17814_ ;
	wire _w17813_ ;
	wire _w17812_ ;
	wire _w17811_ ;
	wire _w17810_ ;
	wire _w17809_ ;
	wire _w17808_ ;
	wire _w17807_ ;
	wire _w17806_ ;
	wire _w17805_ ;
	wire _w17804_ ;
	wire _w17803_ ;
	wire _w17802_ ;
	wire _w17801_ ;
	wire _w17800_ ;
	wire _w17799_ ;
	wire _w17798_ ;
	wire _w17797_ ;
	wire _w17796_ ;
	wire _w17795_ ;
	wire _w17794_ ;
	wire _w17793_ ;
	wire _w17792_ ;
	wire _w17791_ ;
	wire _w17790_ ;
	wire _w17789_ ;
	wire _w17788_ ;
	wire _w17787_ ;
	wire _w17786_ ;
	wire _w17785_ ;
	wire _w17784_ ;
	wire _w17783_ ;
	wire _w17782_ ;
	wire _w17781_ ;
	wire _w17780_ ;
	wire _w17779_ ;
	wire _w17778_ ;
	wire _w17777_ ;
	wire _w17776_ ;
	wire _w17775_ ;
	wire _w17774_ ;
	wire _w17773_ ;
	wire _w17772_ ;
	wire _w17771_ ;
	wire _w17770_ ;
	wire _w17769_ ;
	wire _w17768_ ;
	wire _w17767_ ;
	wire _w17766_ ;
	wire _w17765_ ;
	wire _w17764_ ;
	wire _w17763_ ;
	wire _w17762_ ;
	wire _w17761_ ;
	wire _w17760_ ;
	wire _w17759_ ;
	wire _w17758_ ;
	wire _w17757_ ;
	wire _w17756_ ;
	wire _w17755_ ;
	wire _w17754_ ;
	wire _w17753_ ;
	wire _w17752_ ;
	wire _w17751_ ;
	wire _w17750_ ;
	wire _w17749_ ;
	wire _w17748_ ;
	wire _w17747_ ;
	wire _w17746_ ;
	wire _w17745_ ;
	wire _w17744_ ;
	wire _w17743_ ;
	wire _w17742_ ;
	wire _w17741_ ;
	wire _w17740_ ;
	wire _w17739_ ;
	wire _w17738_ ;
	wire _w17737_ ;
	wire _w17736_ ;
	wire _w17735_ ;
	wire _w17734_ ;
	wire _w17733_ ;
	wire _w17732_ ;
	wire _w17731_ ;
	wire _w17730_ ;
	wire _w17729_ ;
	wire _w17728_ ;
	wire _w17727_ ;
	wire _w17726_ ;
	wire _w17725_ ;
	wire _w17724_ ;
	wire _w17723_ ;
	wire _w17722_ ;
	wire _w17721_ ;
	wire _w17720_ ;
	wire _w17719_ ;
	wire _w17718_ ;
	wire _w17717_ ;
	wire _w17716_ ;
	wire _w17715_ ;
	wire _w17714_ ;
	wire _w17713_ ;
	wire _w17712_ ;
	wire _w17711_ ;
	wire _w17710_ ;
	wire _w17709_ ;
	wire _w17708_ ;
	wire _w17707_ ;
	wire _w17706_ ;
	wire _w17705_ ;
	wire _w17704_ ;
	wire _w17703_ ;
	wire _w17702_ ;
	wire _w17701_ ;
	wire _w17700_ ;
	wire _w17699_ ;
	wire _w17698_ ;
	wire _w17697_ ;
	wire _w17696_ ;
	wire _w17695_ ;
	wire _w17694_ ;
	wire _w17693_ ;
	wire _w17692_ ;
	wire _w17691_ ;
	wire _w17690_ ;
	wire _w17689_ ;
	wire _w17688_ ;
	wire _w17687_ ;
	wire _w17686_ ;
	wire _w17685_ ;
	wire _w17684_ ;
	wire _w17683_ ;
	wire _w17682_ ;
	wire _w17681_ ;
	wire _w17680_ ;
	wire _w17679_ ;
	wire _w17678_ ;
	wire _w17677_ ;
	wire _w17676_ ;
	wire _w17675_ ;
	wire _w17674_ ;
	wire _w17673_ ;
	wire _w17672_ ;
	wire _w17671_ ;
	wire _w17670_ ;
	wire _w17669_ ;
	wire _w17668_ ;
	wire _w17667_ ;
	wire _w17666_ ;
	wire _w17665_ ;
	wire _w17664_ ;
	wire _w17663_ ;
	wire _w17662_ ;
	wire _w17661_ ;
	wire _w17660_ ;
	wire _w17659_ ;
	wire _w17658_ ;
	wire _w17657_ ;
	wire _w17656_ ;
	wire _w17655_ ;
	wire _w17654_ ;
	wire _w17653_ ;
	wire _w17652_ ;
	wire _w17651_ ;
	wire _w17650_ ;
	wire _w17649_ ;
	wire _w17648_ ;
	wire _w17647_ ;
	wire _w17646_ ;
	wire _w17645_ ;
	wire _w17644_ ;
	wire _w17643_ ;
	wire _w17642_ ;
	wire _w17641_ ;
	wire _w17640_ ;
	wire _w17639_ ;
	wire _w17638_ ;
	wire _w17637_ ;
	wire _w17636_ ;
	wire _w17635_ ;
	wire _w17634_ ;
	wire _w17633_ ;
	wire _w17632_ ;
	wire _w17631_ ;
	wire _w17630_ ;
	wire _w17629_ ;
	wire _w17628_ ;
	wire _w17627_ ;
	wire _w17626_ ;
	wire _w17625_ ;
	wire _w17624_ ;
	wire _w17623_ ;
	wire _w17622_ ;
	wire _w17621_ ;
	wire _w17620_ ;
	wire _w17619_ ;
	wire _w17618_ ;
	wire _w17617_ ;
	wire _w17616_ ;
	wire _w17615_ ;
	wire _w17614_ ;
	wire _w17613_ ;
	wire _w17612_ ;
	wire _w17611_ ;
	wire _w17610_ ;
	wire _w17609_ ;
	wire _w17608_ ;
	wire _w17607_ ;
	wire _w17606_ ;
	wire _w17605_ ;
	wire _w17604_ ;
	wire _w17603_ ;
	wire _w17602_ ;
	wire _w17601_ ;
	wire _w17600_ ;
	wire _w17599_ ;
	wire _w17598_ ;
	wire _w17597_ ;
	wire _w17596_ ;
	wire _w17595_ ;
	wire _w17594_ ;
	wire _w17593_ ;
	wire _w17592_ ;
	wire _w17591_ ;
	wire _w17590_ ;
	wire _w17589_ ;
	wire _w17588_ ;
	wire _w17587_ ;
	wire _w17586_ ;
	wire _w17585_ ;
	wire _w17584_ ;
	wire _w17583_ ;
	wire _w17582_ ;
	wire _w17581_ ;
	wire _w17580_ ;
	wire _w17579_ ;
	wire _w17578_ ;
	wire _w17577_ ;
	wire _w17576_ ;
	wire _w17575_ ;
	wire _w17574_ ;
	wire _w17573_ ;
	wire _w17572_ ;
	wire _w17571_ ;
	wire _w17570_ ;
	wire _w17569_ ;
	wire _w17568_ ;
	wire _w17567_ ;
	wire _w17566_ ;
	wire _w17565_ ;
	wire _w17564_ ;
	wire _w17563_ ;
	wire _w17562_ ;
	wire _w17561_ ;
	wire _w17560_ ;
	wire _w17559_ ;
	wire _w17558_ ;
	wire _w17557_ ;
	wire _w17556_ ;
	wire _w17555_ ;
	wire _w17554_ ;
	wire _w17553_ ;
	wire _w17552_ ;
	wire _w17551_ ;
	wire _w17550_ ;
	wire _w17549_ ;
	wire _w17548_ ;
	wire _w17547_ ;
	wire _w17546_ ;
	wire _w17545_ ;
	wire _w17544_ ;
	wire _w17543_ ;
	wire _w17542_ ;
	wire _w17541_ ;
	wire _w17540_ ;
	wire _w17539_ ;
	wire _w17538_ ;
	wire _w17537_ ;
	wire _w17536_ ;
	wire _w17535_ ;
	wire _w17534_ ;
	wire _w17533_ ;
	wire _w17532_ ;
	wire _w17531_ ;
	wire _w17530_ ;
	wire _w17529_ ;
	wire _w17528_ ;
	wire _w17527_ ;
	wire _w17526_ ;
	wire _w17525_ ;
	wire _w17524_ ;
	wire _w17523_ ;
	wire _w17522_ ;
	wire _w17521_ ;
	wire _w17520_ ;
	wire _w17519_ ;
	wire _w17518_ ;
	wire _w17517_ ;
	wire _w17516_ ;
	wire _w17515_ ;
	wire _w17514_ ;
	wire _w17513_ ;
	wire _w17512_ ;
	wire _w17511_ ;
	wire _w17510_ ;
	wire _w17509_ ;
	wire _w17508_ ;
	wire _w17507_ ;
	wire _w17506_ ;
	wire _w17505_ ;
	wire _w17504_ ;
	wire _w17503_ ;
	wire _w17502_ ;
	wire _w17501_ ;
	wire _w17500_ ;
	wire _w17499_ ;
	wire _w17498_ ;
	wire _w17497_ ;
	wire _w17496_ ;
	wire _w17495_ ;
	wire _w17494_ ;
	wire _w17493_ ;
	wire _w17492_ ;
	wire _w17491_ ;
	wire _w17490_ ;
	wire _w17489_ ;
	wire _w17488_ ;
	wire _w17487_ ;
	wire _w17486_ ;
	wire _w17485_ ;
	wire _w17484_ ;
	wire _w17483_ ;
	wire _w17482_ ;
	wire _w17481_ ;
	wire _w17480_ ;
	wire _w17479_ ;
	wire _w17478_ ;
	wire _w17477_ ;
	wire _w17476_ ;
	wire _w17475_ ;
	wire _w17474_ ;
	wire _w17473_ ;
	wire _w17472_ ;
	wire _w17471_ ;
	wire _w17470_ ;
	wire _w17469_ ;
	wire _w17468_ ;
	wire _w17467_ ;
	wire _w17466_ ;
	wire _w17465_ ;
	wire _w17464_ ;
	wire _w17463_ ;
	wire _w17462_ ;
	wire _w17461_ ;
	wire _w17460_ ;
	wire _w17459_ ;
	wire _w17458_ ;
	wire _w17457_ ;
	wire _w17456_ ;
	wire _w17455_ ;
	wire _w17454_ ;
	wire _w17453_ ;
	wire _w17452_ ;
	wire _w17451_ ;
	wire _w17450_ ;
	wire _w17449_ ;
	wire _w17448_ ;
	wire _w17447_ ;
	wire _w17446_ ;
	wire _w17445_ ;
	wire _w17444_ ;
	wire _w17443_ ;
	wire _w17442_ ;
	wire _w17441_ ;
	wire _w17440_ ;
	wire _w17439_ ;
	wire _w17438_ ;
	wire _w17437_ ;
	wire _w17436_ ;
	wire _w17435_ ;
	wire _w17434_ ;
	wire _w17433_ ;
	wire _w17432_ ;
	wire _w17431_ ;
	wire _w17430_ ;
	wire _w17429_ ;
	wire _w17428_ ;
	wire _w17427_ ;
	wire _w17426_ ;
	wire _w17425_ ;
	wire _w17424_ ;
	wire _w17423_ ;
	wire _w17422_ ;
	wire _w17421_ ;
	wire _w17420_ ;
	wire _w17419_ ;
	wire _w17418_ ;
	wire _w17417_ ;
	wire _w17416_ ;
	wire _w17415_ ;
	wire _w17414_ ;
	wire _w17413_ ;
	wire _w17412_ ;
	wire _w17411_ ;
	wire _w17410_ ;
	wire _w17409_ ;
	wire _w17408_ ;
	wire _w17407_ ;
	wire _w17406_ ;
	wire _w17405_ ;
	wire _w17404_ ;
	wire _w17403_ ;
	wire _w17402_ ;
	wire _w17401_ ;
	wire _w17400_ ;
	wire _w17399_ ;
	wire _w17398_ ;
	wire _w17397_ ;
	wire _w17396_ ;
	wire _w17395_ ;
	wire _w17394_ ;
	wire _w17393_ ;
	wire _w17392_ ;
	wire _w17391_ ;
	wire _w17390_ ;
	wire _w17389_ ;
	wire _w17388_ ;
	wire _w17387_ ;
	wire _w17386_ ;
	wire _w17385_ ;
	wire _w17384_ ;
	wire _w17383_ ;
	wire _w17382_ ;
	wire _w17381_ ;
	wire _w17380_ ;
	wire _w17379_ ;
	wire _w17378_ ;
	wire _w17377_ ;
	wire _w17376_ ;
	wire _w17375_ ;
	wire _w17374_ ;
	wire _w17373_ ;
	wire _w17372_ ;
	wire _w17371_ ;
	wire _w17370_ ;
	wire _w17369_ ;
	wire _w17368_ ;
	wire _w17367_ ;
	wire _w17366_ ;
	wire _w17365_ ;
	wire _w17364_ ;
	wire _w17363_ ;
	wire _w17362_ ;
	wire _w17361_ ;
	wire _w17360_ ;
	wire _w17359_ ;
	wire _w17358_ ;
	wire _w17357_ ;
	wire _w17356_ ;
	wire _w17355_ ;
	wire _w17354_ ;
	wire _w17353_ ;
	wire _w17352_ ;
	wire _w17351_ ;
	wire _w17350_ ;
	wire _w17349_ ;
	wire _w17348_ ;
	wire _w17347_ ;
	wire _w17346_ ;
	wire _w17345_ ;
	wire _w17344_ ;
	wire _w17343_ ;
	wire _w17342_ ;
	wire _w17341_ ;
	wire _w17340_ ;
	wire _w17339_ ;
	wire _w17338_ ;
	wire _w17337_ ;
	wire _w17336_ ;
	wire _w17335_ ;
	wire _w17334_ ;
	wire _w17333_ ;
	wire _w17332_ ;
	wire _w17331_ ;
	wire _w17330_ ;
	wire _w17329_ ;
	wire _w17328_ ;
	wire _w17327_ ;
	wire _w17326_ ;
	wire _w17325_ ;
	wire _w17324_ ;
	wire _w17323_ ;
	wire _w17322_ ;
	wire _w17321_ ;
	wire _w17320_ ;
	wire _w17319_ ;
	wire _w17318_ ;
	wire _w17317_ ;
	wire _w17316_ ;
	wire _w17315_ ;
	wire _w17314_ ;
	wire _w17313_ ;
	wire _w17312_ ;
	wire _w17311_ ;
	wire _w17310_ ;
	wire _w17309_ ;
	wire _w17308_ ;
	wire _w17307_ ;
	wire _w17306_ ;
	wire _w17305_ ;
	wire _w17304_ ;
	wire _w17303_ ;
	wire _w17302_ ;
	wire _w17301_ ;
	wire _w17300_ ;
	wire _w17299_ ;
	wire _w17298_ ;
	wire _w17297_ ;
	wire _w17296_ ;
	wire _w17295_ ;
	wire _w17294_ ;
	wire _w17293_ ;
	wire _w17292_ ;
	wire _w17291_ ;
	wire _w17290_ ;
	wire _w17289_ ;
	wire _w17288_ ;
	wire _w17287_ ;
	wire _w17286_ ;
	wire _w17285_ ;
	wire _w17284_ ;
	wire _w17283_ ;
	wire _w17282_ ;
	wire _w17281_ ;
	wire _w17280_ ;
	wire _w17279_ ;
	wire _w17278_ ;
	wire _w17277_ ;
	wire _w17276_ ;
	wire _w17275_ ;
	wire _w17274_ ;
	wire _w17273_ ;
	wire _w17272_ ;
	wire _w17271_ ;
	wire _w17270_ ;
	wire _w17269_ ;
	wire _w17268_ ;
	wire _w17267_ ;
	wire _w17266_ ;
	wire _w17265_ ;
	wire _w17264_ ;
	wire _w17263_ ;
	wire _w17262_ ;
	wire _w17261_ ;
	wire _w17260_ ;
	wire _w17259_ ;
	wire _w17258_ ;
	wire _w17257_ ;
	wire _w17256_ ;
	wire _w17255_ ;
	wire _w17254_ ;
	wire _w17253_ ;
	wire _w17252_ ;
	wire _w17251_ ;
	wire _w17250_ ;
	wire _w17249_ ;
	wire _w17248_ ;
	wire _w17247_ ;
	wire _w17246_ ;
	wire _w17245_ ;
	wire _w17244_ ;
	wire _w17243_ ;
	wire _w17242_ ;
	wire _w17241_ ;
	wire _w17240_ ;
	wire _w17239_ ;
	wire _w17238_ ;
	wire _w17237_ ;
	wire _w17236_ ;
	wire _w17235_ ;
	wire _w17234_ ;
	wire _w17233_ ;
	wire _w17232_ ;
	wire _w17231_ ;
	wire _w17230_ ;
	wire _w17229_ ;
	wire _w17228_ ;
	wire _w17227_ ;
	wire _w17226_ ;
	wire _w17225_ ;
	wire _w17224_ ;
	wire _w17223_ ;
	wire _w17222_ ;
	wire _w17221_ ;
	wire _w17220_ ;
	wire _w17219_ ;
	wire _w17218_ ;
	wire _w17217_ ;
	wire _w17216_ ;
	wire _w17215_ ;
	wire _w17214_ ;
	wire _w17213_ ;
	wire _w17212_ ;
	wire _w17211_ ;
	wire _w17210_ ;
	wire _w17209_ ;
	wire _w17208_ ;
	wire _w17207_ ;
	wire _w17206_ ;
	wire _w17205_ ;
	wire _w17204_ ;
	wire _w17203_ ;
	wire _w17202_ ;
	wire _w17201_ ;
	wire _w17200_ ;
	wire _w17199_ ;
	wire _w17198_ ;
	wire _w17197_ ;
	wire _w17196_ ;
	wire _w17195_ ;
	wire _w17194_ ;
	wire _w17193_ ;
	wire _w17192_ ;
	wire _w17191_ ;
	wire _w17190_ ;
	wire _w17189_ ;
	wire _w17188_ ;
	wire _w17187_ ;
	wire _w17186_ ;
	wire _w17185_ ;
	wire _w17184_ ;
	wire _w17183_ ;
	wire _w17182_ ;
	wire _w17181_ ;
	wire _w17180_ ;
	wire _w17179_ ;
	wire _w17178_ ;
	wire _w17177_ ;
	wire _w17176_ ;
	wire _w17175_ ;
	wire _w17174_ ;
	wire _w17173_ ;
	wire _w17172_ ;
	wire _w17171_ ;
	wire _w17170_ ;
	wire _w17169_ ;
	wire _w17168_ ;
	wire _w17167_ ;
	wire _w17166_ ;
	wire _w17165_ ;
	wire _w17164_ ;
	wire _w17163_ ;
	wire _w17162_ ;
	wire _w17161_ ;
	wire _w17160_ ;
	wire _w17159_ ;
	wire _w17158_ ;
	wire _w17157_ ;
	wire _w17156_ ;
	wire _w17155_ ;
	wire _w17154_ ;
	wire _w17153_ ;
	wire _w17152_ ;
	wire _w17151_ ;
	wire _w17150_ ;
	wire _w17149_ ;
	wire _w17148_ ;
	wire _w17147_ ;
	wire _w17146_ ;
	wire _w17145_ ;
	wire _w17144_ ;
	wire _w17143_ ;
	wire _w17142_ ;
	wire _w17141_ ;
	wire _w17140_ ;
	wire _w17139_ ;
	wire _w17138_ ;
	wire _w17137_ ;
	wire _w17136_ ;
	wire _w17135_ ;
	wire _w17134_ ;
	wire _w17133_ ;
	wire _w17132_ ;
	wire _w17131_ ;
	wire _w17130_ ;
	wire _w17129_ ;
	wire _w17128_ ;
	wire _w17127_ ;
	wire _w17126_ ;
	wire _w17125_ ;
	wire _w17124_ ;
	wire _w17123_ ;
	wire _w17122_ ;
	wire _w17121_ ;
	wire _w17120_ ;
	wire _w17119_ ;
	wire _w17118_ ;
	wire _w17117_ ;
	wire _w17116_ ;
	wire _w17115_ ;
	wire _w17114_ ;
	wire _w17113_ ;
	wire _w17112_ ;
	wire _w17111_ ;
	wire _w17110_ ;
	wire _w17109_ ;
	wire _w17108_ ;
	wire _w17107_ ;
	wire _w17106_ ;
	wire _w17105_ ;
	wire _w17104_ ;
	wire _w17103_ ;
	wire _w17102_ ;
	wire _w17101_ ;
	wire _w17100_ ;
	wire _w17099_ ;
	wire _w17098_ ;
	wire _w17097_ ;
	wire _w17096_ ;
	wire _w17095_ ;
	wire _w17094_ ;
	wire _w17093_ ;
	wire _w17092_ ;
	wire _w17091_ ;
	wire _w17090_ ;
	wire _w17089_ ;
	wire _w17088_ ;
	wire _w17087_ ;
	wire _w17086_ ;
	wire _w17085_ ;
	wire _w17084_ ;
	wire _w17083_ ;
	wire _w17082_ ;
	wire _w17081_ ;
	wire _w17080_ ;
	wire _w17079_ ;
	wire _w17078_ ;
	wire _w17077_ ;
	wire _w17076_ ;
	wire _w17075_ ;
	wire _w17074_ ;
	wire _w17073_ ;
	wire _w17072_ ;
	wire _w17071_ ;
	wire _w17070_ ;
	wire _w17069_ ;
	wire _w17068_ ;
	wire _w17067_ ;
	wire _w17066_ ;
	wire _w17065_ ;
	wire _w17064_ ;
	wire _w17063_ ;
	wire _w17062_ ;
	wire _w17061_ ;
	wire _w17060_ ;
	wire _w17059_ ;
	wire _w17058_ ;
	wire _w17057_ ;
	wire _w17056_ ;
	wire _w17055_ ;
	wire _w17054_ ;
	wire _w17053_ ;
	wire _w17052_ ;
	wire _w17051_ ;
	wire _w17050_ ;
	wire _w17049_ ;
	wire _w17048_ ;
	wire _w17047_ ;
	wire _w17046_ ;
	wire _w17045_ ;
	wire _w17044_ ;
	wire _w17043_ ;
	wire _w17042_ ;
	wire _w17041_ ;
	wire _w17040_ ;
	wire _w17039_ ;
	wire _w17038_ ;
	wire _w17037_ ;
	wire _w17036_ ;
	wire _w17035_ ;
	wire _w17034_ ;
	wire _w17033_ ;
	wire _w17032_ ;
	wire _w17031_ ;
	wire _w17030_ ;
	wire _w17029_ ;
	wire _w17028_ ;
	wire _w17027_ ;
	wire _w17026_ ;
	wire _w17025_ ;
	wire _w17024_ ;
	wire _w17023_ ;
	wire _w17022_ ;
	wire _w17021_ ;
	wire _w17020_ ;
	wire _w17019_ ;
	wire _w17018_ ;
	wire _w17017_ ;
	wire _w17016_ ;
	wire _w17015_ ;
	wire _w17014_ ;
	wire _w17013_ ;
	wire _w17012_ ;
	wire _w17011_ ;
	wire _w17010_ ;
	wire _w17009_ ;
	wire _w17008_ ;
	wire _w17007_ ;
	wire _w17006_ ;
	wire _w17005_ ;
	wire _w17004_ ;
	wire _w17003_ ;
	wire _w17002_ ;
	wire _w17001_ ;
	wire _w17000_ ;
	wire _w16999_ ;
	wire _w16998_ ;
	wire _w16997_ ;
	wire _w16996_ ;
	wire _w16995_ ;
	wire _w16994_ ;
	wire _w16993_ ;
	wire _w16992_ ;
	wire _w16991_ ;
	wire _w16990_ ;
	wire _w16989_ ;
	wire _w16988_ ;
	wire _w16987_ ;
	wire _w16986_ ;
	wire _w16985_ ;
	wire _w16984_ ;
	wire _w16983_ ;
	wire _w16982_ ;
	wire _w16981_ ;
	wire _w16980_ ;
	wire _w16979_ ;
	wire _w16978_ ;
	wire _w16977_ ;
	wire _w16976_ ;
	wire _w16975_ ;
	wire _w16974_ ;
	wire _w16973_ ;
	wire _w16972_ ;
	wire _w16971_ ;
	wire _w16970_ ;
	wire _w16969_ ;
	wire _w16968_ ;
	wire _w16967_ ;
	wire _w16966_ ;
	wire _w16965_ ;
	wire _w16964_ ;
	wire _w16963_ ;
	wire _w16962_ ;
	wire _w16961_ ;
	wire _w16960_ ;
	wire _w16959_ ;
	wire _w16958_ ;
	wire _w16957_ ;
	wire _w16956_ ;
	wire _w16955_ ;
	wire _w16954_ ;
	wire _w16953_ ;
	wire _w16952_ ;
	wire _w16951_ ;
	wire _w16950_ ;
	wire _w16949_ ;
	wire _w16948_ ;
	wire _w16947_ ;
	wire _w16946_ ;
	wire _w16945_ ;
	wire _w16944_ ;
	wire _w16943_ ;
	wire _w16942_ ;
	wire _w16941_ ;
	wire _w16940_ ;
	wire _w16939_ ;
	wire _w16938_ ;
	wire _w16937_ ;
	wire _w16936_ ;
	wire _w16935_ ;
	wire _w16934_ ;
	wire _w16933_ ;
	wire _w16932_ ;
	wire _w16931_ ;
	wire _w16930_ ;
	wire _w16929_ ;
	wire _w16928_ ;
	wire _w16927_ ;
	wire _w16926_ ;
	wire _w16925_ ;
	wire _w16924_ ;
	wire _w16923_ ;
	wire _w16922_ ;
	wire _w16921_ ;
	wire _w16920_ ;
	wire _w16919_ ;
	wire _w16918_ ;
	wire _w16917_ ;
	wire _w16916_ ;
	wire _w16915_ ;
	wire _w16914_ ;
	wire _w16913_ ;
	wire _w16912_ ;
	wire _w16911_ ;
	wire _w16910_ ;
	wire _w16909_ ;
	wire _w16908_ ;
	wire _w16907_ ;
	wire _w16906_ ;
	wire _w16905_ ;
	wire _w16904_ ;
	wire _w16903_ ;
	wire _w16902_ ;
	wire _w16901_ ;
	wire _w16900_ ;
	wire _w16899_ ;
	wire _w16898_ ;
	wire _w16897_ ;
	wire _w16896_ ;
	wire _w16895_ ;
	wire _w16894_ ;
	wire _w16893_ ;
	wire _w16892_ ;
	wire _w16891_ ;
	wire _w16890_ ;
	wire _w16889_ ;
	wire _w16888_ ;
	wire _w16887_ ;
	wire _w16886_ ;
	wire _w16885_ ;
	wire _w16884_ ;
	wire _w16883_ ;
	wire _w16882_ ;
	wire _w16881_ ;
	wire _w16880_ ;
	wire _w16879_ ;
	wire _w16878_ ;
	wire _w16877_ ;
	wire _w16876_ ;
	wire _w16875_ ;
	wire _w16874_ ;
	wire _w16873_ ;
	wire _w16872_ ;
	wire _w16871_ ;
	wire _w16870_ ;
	wire _w16869_ ;
	wire _w16868_ ;
	wire _w16867_ ;
	wire _w16866_ ;
	wire _w16865_ ;
	wire _w16864_ ;
	wire _w16863_ ;
	wire _w16862_ ;
	wire _w16861_ ;
	wire _w16860_ ;
	wire _w16859_ ;
	wire _w16858_ ;
	wire _w16857_ ;
	wire _w16856_ ;
	wire _w16855_ ;
	wire _w16854_ ;
	wire _w16853_ ;
	wire _w16852_ ;
	wire _w16851_ ;
	wire _w16850_ ;
	wire _w16849_ ;
	wire _w16848_ ;
	wire _w16847_ ;
	wire _w16846_ ;
	wire _w16845_ ;
	wire _w16844_ ;
	wire _w16843_ ;
	wire _w16842_ ;
	wire _w16841_ ;
	wire _w16840_ ;
	wire _w16839_ ;
	wire _w16838_ ;
	wire _w16837_ ;
	wire _w16836_ ;
	wire _w16835_ ;
	wire _w16834_ ;
	wire _w16833_ ;
	wire _w16832_ ;
	wire _w16831_ ;
	wire _w16830_ ;
	wire _w16829_ ;
	wire _w16828_ ;
	wire _w16827_ ;
	wire _w16826_ ;
	wire _w16825_ ;
	wire _w16824_ ;
	wire _w16823_ ;
	wire _w16822_ ;
	wire _w16821_ ;
	wire _w16820_ ;
	wire _w16819_ ;
	wire _w16818_ ;
	wire _w16817_ ;
	wire _w16816_ ;
	wire _w16815_ ;
	wire _w16814_ ;
	wire _w16813_ ;
	wire _w16812_ ;
	wire _w16811_ ;
	wire _w16810_ ;
	wire _w16809_ ;
	wire _w16808_ ;
	wire _w16807_ ;
	wire _w16806_ ;
	wire _w16805_ ;
	wire _w16804_ ;
	wire _w16803_ ;
	wire _w16802_ ;
	wire _w16801_ ;
	wire _w16800_ ;
	wire _w16799_ ;
	wire _w16798_ ;
	wire _w16797_ ;
	wire _w16796_ ;
	wire _w16795_ ;
	wire _w16794_ ;
	wire _w16793_ ;
	wire _w16792_ ;
	wire _w16791_ ;
	wire _w16790_ ;
	wire _w16789_ ;
	wire _w16788_ ;
	wire _w16787_ ;
	wire _w16786_ ;
	wire _w16785_ ;
	wire _w16784_ ;
	wire _w16783_ ;
	wire _w16782_ ;
	wire _w16781_ ;
	wire _w16780_ ;
	wire _w16779_ ;
	wire _w16778_ ;
	wire _w16777_ ;
	wire _w16776_ ;
	wire _w16775_ ;
	wire _w16774_ ;
	wire _w16773_ ;
	wire _w16772_ ;
	wire _w16771_ ;
	wire _w16770_ ;
	wire _w16769_ ;
	wire _w16768_ ;
	wire _w16767_ ;
	wire _w16766_ ;
	wire _w16765_ ;
	wire _w16764_ ;
	wire _w16763_ ;
	wire _w16762_ ;
	wire _w16761_ ;
	wire _w16760_ ;
	wire _w16759_ ;
	wire _w16758_ ;
	wire _w16757_ ;
	wire _w16756_ ;
	wire _w16755_ ;
	wire _w16754_ ;
	wire _w16753_ ;
	wire _w16752_ ;
	wire _w16751_ ;
	wire _w16750_ ;
	wire _w16749_ ;
	wire _w16748_ ;
	wire _w16747_ ;
	wire _w16746_ ;
	wire _w16745_ ;
	wire _w16744_ ;
	wire _w16743_ ;
	wire _w16742_ ;
	wire _w16741_ ;
	wire _w16740_ ;
	wire _w16739_ ;
	wire _w16738_ ;
	wire _w16737_ ;
	wire _w16736_ ;
	wire _w16735_ ;
	wire _w16734_ ;
	wire _w16733_ ;
	wire _w16732_ ;
	wire _w16731_ ;
	wire _w16730_ ;
	wire _w16729_ ;
	wire _w16728_ ;
	wire _w16727_ ;
	wire _w16726_ ;
	wire _w16725_ ;
	wire _w16724_ ;
	wire _w16723_ ;
	wire _w16722_ ;
	wire _w16721_ ;
	wire _w16720_ ;
	wire _w16719_ ;
	wire _w16718_ ;
	wire _w16717_ ;
	wire _w16716_ ;
	wire _w16715_ ;
	wire _w16714_ ;
	wire _w16713_ ;
	wire _w16712_ ;
	wire _w16711_ ;
	wire _w16710_ ;
	wire _w16709_ ;
	wire _w16708_ ;
	wire _w16707_ ;
	wire _w16706_ ;
	wire _w16705_ ;
	wire _w16704_ ;
	wire _w16703_ ;
	wire _w16702_ ;
	wire _w16701_ ;
	wire _w16700_ ;
	wire _w16699_ ;
	wire _w16698_ ;
	wire _w16697_ ;
	wire _w16696_ ;
	wire _w16695_ ;
	wire _w16694_ ;
	wire _w16693_ ;
	wire _w16692_ ;
	wire _w16691_ ;
	wire _w16690_ ;
	wire _w16689_ ;
	wire _w16688_ ;
	wire _w16687_ ;
	wire _w16686_ ;
	wire _w16685_ ;
	wire _w16684_ ;
	wire _w16683_ ;
	wire _w16682_ ;
	wire _w16681_ ;
	wire _w16680_ ;
	wire _w16679_ ;
	wire _w16678_ ;
	wire _w16677_ ;
	wire _w16676_ ;
	wire _w16675_ ;
	wire _w16674_ ;
	wire _w16673_ ;
	wire _w16672_ ;
	wire _w16671_ ;
	wire _w16670_ ;
	wire _w16669_ ;
	wire _w16668_ ;
	wire _w16667_ ;
	wire _w16666_ ;
	wire _w16665_ ;
	wire _w16664_ ;
	wire _w16663_ ;
	wire _w16662_ ;
	wire _w16661_ ;
	wire _w16660_ ;
	wire _w16659_ ;
	wire _w16658_ ;
	wire _w16657_ ;
	wire _w16656_ ;
	wire _w16655_ ;
	wire _w16654_ ;
	wire _w16653_ ;
	wire _w16652_ ;
	wire _w16651_ ;
	wire _w16650_ ;
	wire _w16649_ ;
	wire _w16648_ ;
	wire _w16647_ ;
	wire _w16646_ ;
	wire _w16645_ ;
	wire _w16644_ ;
	wire _w16643_ ;
	wire _w16642_ ;
	wire _w16641_ ;
	wire _w16640_ ;
	wire _w16639_ ;
	wire _w16638_ ;
	wire _w16637_ ;
	wire _w16636_ ;
	wire _w16635_ ;
	wire _w16634_ ;
	wire _w16633_ ;
	wire _w16632_ ;
	wire _w16631_ ;
	wire _w16630_ ;
	wire _w16629_ ;
	wire _w16628_ ;
	wire _w16627_ ;
	wire _w16626_ ;
	wire _w16625_ ;
	wire _w16624_ ;
	wire _w16623_ ;
	wire _w16622_ ;
	wire _w16621_ ;
	wire _w16620_ ;
	wire _w16619_ ;
	wire _w16618_ ;
	wire _w16617_ ;
	wire _w16616_ ;
	wire _w16615_ ;
	wire _w16614_ ;
	wire _w16613_ ;
	wire _w16612_ ;
	wire _w16611_ ;
	wire _w16610_ ;
	wire _w16609_ ;
	wire _w16608_ ;
	wire _w16607_ ;
	wire _w16606_ ;
	wire _w16605_ ;
	wire _w16604_ ;
	wire _w16603_ ;
	wire _w16602_ ;
	wire _w16601_ ;
	wire _w16600_ ;
	wire _w16599_ ;
	wire _w16598_ ;
	wire _w16597_ ;
	wire _w16596_ ;
	wire _w16595_ ;
	wire _w16594_ ;
	wire _w16593_ ;
	wire _w16592_ ;
	wire _w16591_ ;
	wire _w16590_ ;
	wire _w16589_ ;
	wire _w16588_ ;
	wire _w16587_ ;
	wire _w16586_ ;
	wire _w16585_ ;
	wire _w16584_ ;
	wire _w16583_ ;
	wire _w16582_ ;
	wire _w16581_ ;
	wire _w16580_ ;
	wire _w16579_ ;
	wire _w16578_ ;
	wire _w16577_ ;
	wire _w16576_ ;
	wire _w16575_ ;
	wire _w16574_ ;
	wire _w16573_ ;
	wire _w16572_ ;
	wire _w16571_ ;
	wire _w16570_ ;
	wire _w16569_ ;
	wire _w16568_ ;
	wire _w16567_ ;
	wire _w16566_ ;
	wire _w16565_ ;
	wire _w16564_ ;
	wire _w16563_ ;
	wire _w16562_ ;
	wire _w16561_ ;
	wire _w16560_ ;
	wire _w16559_ ;
	wire _w16558_ ;
	wire _w16557_ ;
	wire _w16556_ ;
	wire _w16555_ ;
	wire _w16554_ ;
	wire _w16553_ ;
	wire _w16552_ ;
	wire _w16551_ ;
	wire _w16550_ ;
	wire _w16549_ ;
	wire _w16548_ ;
	wire _w16547_ ;
	wire _w16546_ ;
	wire _w16545_ ;
	wire _w16544_ ;
	wire _w16543_ ;
	wire _w16542_ ;
	wire _w16541_ ;
	wire _w16540_ ;
	wire _w16539_ ;
	wire _w16538_ ;
	wire _w16537_ ;
	wire _w16536_ ;
	wire _w16535_ ;
	wire _w16534_ ;
	wire _w16533_ ;
	wire _w16532_ ;
	wire _w16531_ ;
	wire _w16530_ ;
	wire _w16529_ ;
	wire _w16528_ ;
	wire _w16527_ ;
	wire _w16526_ ;
	wire _w16525_ ;
	wire _w16524_ ;
	wire _w16523_ ;
	wire _w16522_ ;
	wire _w16521_ ;
	wire _w16520_ ;
	wire _w16519_ ;
	wire _w16518_ ;
	wire _w16517_ ;
	wire _w16516_ ;
	wire _w16515_ ;
	wire _w16514_ ;
	wire _w16513_ ;
	wire _w16512_ ;
	wire _w16511_ ;
	wire _w16510_ ;
	wire _w16509_ ;
	wire _w16508_ ;
	wire _w16507_ ;
	wire _w16506_ ;
	wire _w16505_ ;
	wire _w16504_ ;
	wire _w16503_ ;
	wire _w16502_ ;
	wire _w16501_ ;
	wire _w16500_ ;
	wire _w16499_ ;
	wire _w16498_ ;
	wire _w16497_ ;
	wire _w16496_ ;
	wire _w16495_ ;
	wire _w16494_ ;
	wire _w16493_ ;
	wire _w16492_ ;
	wire _w16491_ ;
	wire _w16490_ ;
	wire _w16489_ ;
	wire _w16488_ ;
	wire _w16487_ ;
	wire _w16486_ ;
	wire _w16485_ ;
	wire _w16484_ ;
	wire _w16483_ ;
	wire _w16482_ ;
	wire _w16481_ ;
	wire _w16480_ ;
	wire _w16479_ ;
	wire _w16478_ ;
	wire _w16477_ ;
	wire _w16476_ ;
	wire _w16475_ ;
	wire _w16474_ ;
	wire _w16473_ ;
	wire _w16472_ ;
	wire _w16471_ ;
	wire _w16470_ ;
	wire _w16469_ ;
	wire _w16468_ ;
	wire _w16467_ ;
	wire _w16466_ ;
	wire _w16465_ ;
	wire _w16464_ ;
	wire _w16463_ ;
	wire _w16462_ ;
	wire _w16461_ ;
	wire _w16460_ ;
	wire _w16459_ ;
	wire _w16458_ ;
	wire _w16457_ ;
	wire _w16456_ ;
	wire _w16455_ ;
	wire _w16454_ ;
	wire _w16453_ ;
	wire _w16452_ ;
	wire _w16451_ ;
	wire _w16450_ ;
	wire _w16449_ ;
	wire _w16448_ ;
	wire _w16447_ ;
	wire _w16446_ ;
	wire _w16445_ ;
	wire _w16444_ ;
	wire _w16443_ ;
	wire _w16442_ ;
	wire _w16441_ ;
	wire _w16440_ ;
	wire _w16439_ ;
	wire _w16438_ ;
	wire _w16437_ ;
	wire _w16436_ ;
	wire _w16435_ ;
	wire _w16434_ ;
	wire _w16433_ ;
	wire _w16432_ ;
	wire _w16431_ ;
	wire _w16430_ ;
	wire _w16429_ ;
	wire _w16428_ ;
	wire _w16427_ ;
	wire _w16426_ ;
	wire _w16425_ ;
	wire _w16424_ ;
	wire _w16423_ ;
	wire _w16422_ ;
	wire _w16421_ ;
	wire _w16420_ ;
	wire _w16419_ ;
	wire _w16418_ ;
	wire _w16417_ ;
	wire _w16416_ ;
	wire _w16415_ ;
	wire _w16414_ ;
	wire _w16413_ ;
	wire _w16412_ ;
	wire _w16411_ ;
	wire _w16410_ ;
	wire _w16409_ ;
	wire _w16408_ ;
	wire _w16407_ ;
	wire _w16406_ ;
	wire _w16405_ ;
	wire _w16404_ ;
	wire _w16403_ ;
	wire _w16402_ ;
	wire _w16401_ ;
	wire _w16400_ ;
	wire _w16399_ ;
	wire _w16398_ ;
	wire _w16397_ ;
	wire _w16396_ ;
	wire _w16395_ ;
	wire _w16394_ ;
	wire _w16393_ ;
	wire _w16392_ ;
	wire _w16391_ ;
	wire _w16390_ ;
	wire _w16389_ ;
	wire _w16388_ ;
	wire _w16387_ ;
	wire _w16386_ ;
	wire _w16385_ ;
	wire _w16384_ ;
	wire _w16383_ ;
	wire _w16382_ ;
	wire _w16381_ ;
	wire _w16380_ ;
	wire _w16379_ ;
	wire _w16378_ ;
	wire _w16377_ ;
	wire _w16376_ ;
	wire _w16375_ ;
	wire _w16374_ ;
	wire _w16373_ ;
	wire _w16372_ ;
	wire _w16371_ ;
	wire _w16370_ ;
	wire _w16369_ ;
	wire _w16368_ ;
	wire _w16367_ ;
	wire _w16366_ ;
	wire _w16365_ ;
	wire _w16364_ ;
	wire _w16363_ ;
	wire _w16362_ ;
	wire _w16361_ ;
	wire _w16360_ ;
	wire _w16359_ ;
	wire _w16358_ ;
	wire _w16357_ ;
	wire _w16356_ ;
	wire _w16355_ ;
	wire _w16354_ ;
	wire _w16353_ ;
	wire _w16352_ ;
	wire _w16351_ ;
	wire _w16350_ ;
	wire _w16349_ ;
	wire _w16348_ ;
	wire _w16347_ ;
	wire _w16346_ ;
	wire _w16345_ ;
	wire _w16344_ ;
	wire _w16343_ ;
	wire _w16342_ ;
	wire _w16341_ ;
	wire _w16340_ ;
	wire _w16339_ ;
	wire _w16338_ ;
	wire _w16337_ ;
	wire _w16336_ ;
	wire _w16335_ ;
	wire _w16334_ ;
	wire _w16333_ ;
	wire _w16332_ ;
	wire _w16331_ ;
	wire _w16330_ ;
	wire _w16329_ ;
	wire _w16328_ ;
	wire _w16327_ ;
	wire _w16326_ ;
	wire _w16325_ ;
	wire _w16324_ ;
	wire _w16323_ ;
	wire _w16322_ ;
	wire _w16321_ ;
	wire _w16320_ ;
	wire _w16319_ ;
	wire _w16318_ ;
	wire _w16317_ ;
	wire _w16316_ ;
	wire _w16315_ ;
	wire _w16314_ ;
	wire _w16313_ ;
	wire _w16312_ ;
	wire _w16311_ ;
	wire _w16310_ ;
	wire _w16309_ ;
	wire _w16308_ ;
	wire _w16307_ ;
	wire _w16306_ ;
	wire _w16305_ ;
	wire _w16304_ ;
	wire _w16303_ ;
	wire _w16302_ ;
	wire _w16301_ ;
	wire _w16300_ ;
	wire _w16299_ ;
	wire _w16298_ ;
	wire _w16297_ ;
	wire _w16296_ ;
	wire _w16295_ ;
	wire _w16294_ ;
	wire _w16293_ ;
	wire _w16292_ ;
	wire _w16291_ ;
	wire _w16290_ ;
	wire _w16289_ ;
	wire _w16288_ ;
	wire _w16287_ ;
	wire _w16286_ ;
	wire _w16285_ ;
	wire _w16284_ ;
	wire _w16283_ ;
	wire _w16282_ ;
	wire _w16281_ ;
	wire _w16280_ ;
	wire _w16279_ ;
	wire _w16278_ ;
	wire _w16277_ ;
	wire _w16276_ ;
	wire _w16275_ ;
	wire _w16274_ ;
	wire _w16273_ ;
	wire _w16272_ ;
	wire _w16271_ ;
	wire _w16270_ ;
	wire _w16269_ ;
	wire _w16268_ ;
	wire _w16267_ ;
	wire _w16266_ ;
	wire _w16265_ ;
	wire _w16264_ ;
	wire _w16263_ ;
	wire _w16262_ ;
	wire _w16261_ ;
	wire _w16260_ ;
	wire _w16259_ ;
	wire _w16258_ ;
	wire _w16257_ ;
	wire _w16256_ ;
	wire _w16255_ ;
	wire _w16254_ ;
	wire _w16253_ ;
	wire _w16252_ ;
	wire _w16251_ ;
	wire _w16250_ ;
	wire _w16249_ ;
	wire _w16248_ ;
	wire _w16247_ ;
	wire _w16246_ ;
	wire _w16245_ ;
	wire _w16244_ ;
	wire _w16243_ ;
	wire _w16242_ ;
	wire _w16241_ ;
	wire _w16240_ ;
	wire _w16239_ ;
	wire _w16238_ ;
	wire _w16237_ ;
	wire _w16236_ ;
	wire _w16235_ ;
	wire _w16234_ ;
	wire _w16233_ ;
	wire _w16232_ ;
	wire _w16231_ ;
	wire _w16230_ ;
	wire _w16229_ ;
	wire _w16228_ ;
	wire _w16227_ ;
	wire _w16226_ ;
	wire _w16225_ ;
	wire _w16224_ ;
	wire _w16223_ ;
	wire _w16222_ ;
	wire _w16221_ ;
	wire _w16220_ ;
	wire _w16219_ ;
	wire _w16218_ ;
	wire _w16217_ ;
	wire _w16216_ ;
	wire _w16215_ ;
	wire _w16214_ ;
	wire _w16213_ ;
	wire _w16212_ ;
	wire _w16211_ ;
	wire _w16210_ ;
	wire _w16209_ ;
	wire _w16208_ ;
	wire _w16207_ ;
	wire _w16206_ ;
	wire _w16205_ ;
	wire _w16204_ ;
	wire _w16203_ ;
	wire _w16202_ ;
	wire _w16201_ ;
	wire _w16200_ ;
	wire _w16199_ ;
	wire _w16198_ ;
	wire _w16197_ ;
	wire _w16196_ ;
	wire _w16195_ ;
	wire _w16194_ ;
	wire _w16193_ ;
	wire _w16192_ ;
	wire _w16191_ ;
	wire _w16190_ ;
	wire _w16189_ ;
	wire _w16188_ ;
	wire _w16187_ ;
	wire _w16186_ ;
	wire _w16185_ ;
	wire _w16184_ ;
	wire _w16183_ ;
	wire _w16182_ ;
	wire _w16181_ ;
	wire _w16180_ ;
	wire _w16179_ ;
	wire _w16178_ ;
	wire _w16177_ ;
	wire _w16176_ ;
	wire _w16175_ ;
	wire _w16174_ ;
	wire _w16173_ ;
	wire _w16172_ ;
	wire _w16171_ ;
	wire _w16170_ ;
	wire _w16169_ ;
	wire _w16168_ ;
	wire _w16167_ ;
	wire _w16166_ ;
	wire _w16165_ ;
	wire _w16164_ ;
	wire _w16163_ ;
	wire _w16162_ ;
	wire _w16161_ ;
	wire _w16160_ ;
	wire _w16159_ ;
	wire _w16158_ ;
	wire _w16157_ ;
	wire _w16156_ ;
	wire _w16155_ ;
	wire _w16154_ ;
	wire _w16153_ ;
	wire _w16152_ ;
	wire _w16151_ ;
	wire _w16150_ ;
	wire _w16149_ ;
	wire _w16148_ ;
	wire _w16147_ ;
	wire _w16146_ ;
	wire _w16145_ ;
	wire _w16144_ ;
	wire _w16143_ ;
	wire _w16142_ ;
	wire _w16141_ ;
	wire _w16140_ ;
	wire _w16139_ ;
	wire _w16138_ ;
	wire _w16137_ ;
	wire _w16136_ ;
	wire _w16135_ ;
	wire _w16134_ ;
	wire _w16133_ ;
	wire _w16132_ ;
	wire _w16131_ ;
	wire _w16130_ ;
	wire _w16129_ ;
	wire _w16128_ ;
	wire _w16127_ ;
	wire _w16126_ ;
	wire _w16125_ ;
	wire _w16124_ ;
	wire _w16123_ ;
	wire _w16122_ ;
	wire _w16121_ ;
	wire _w16120_ ;
	wire _w16119_ ;
	wire _w16118_ ;
	wire _w16117_ ;
	wire _w16116_ ;
	wire _w16115_ ;
	wire _w16114_ ;
	wire _w16113_ ;
	wire _w16112_ ;
	wire _w16111_ ;
	wire _w16110_ ;
	wire _w16109_ ;
	wire _w16108_ ;
	wire _w16107_ ;
	wire _w16106_ ;
	wire _w16105_ ;
	wire _w16104_ ;
	wire _w16103_ ;
	wire _w16102_ ;
	wire _w16101_ ;
	wire _w16100_ ;
	wire _w16099_ ;
	wire _w16098_ ;
	wire _w16097_ ;
	wire _w16096_ ;
	wire _w16095_ ;
	wire _w16094_ ;
	wire _w16093_ ;
	wire _w16092_ ;
	wire _w16091_ ;
	wire _w16090_ ;
	wire _w16089_ ;
	wire _w16088_ ;
	wire _w16087_ ;
	wire _w16086_ ;
	wire _w16085_ ;
	wire _w16084_ ;
	wire _w16083_ ;
	wire _w16082_ ;
	wire _w16081_ ;
	wire _w16080_ ;
	wire _w16079_ ;
	wire _w16078_ ;
	wire _w16077_ ;
	wire _w16076_ ;
	wire _w16075_ ;
	wire _w16074_ ;
	wire _w16073_ ;
	wire _w16072_ ;
	wire _w16071_ ;
	wire _w16070_ ;
	wire _w16069_ ;
	wire _w16068_ ;
	wire _w16067_ ;
	wire _w16066_ ;
	wire _w16065_ ;
	wire _w16064_ ;
	wire _w16063_ ;
	wire _w16062_ ;
	wire _w16061_ ;
	wire _w16060_ ;
	wire _w16059_ ;
	wire _w16058_ ;
	wire _w16057_ ;
	wire _w16056_ ;
	wire _w16055_ ;
	wire _w16054_ ;
	wire _w16053_ ;
	wire _w16052_ ;
	wire _w16051_ ;
	wire _w16050_ ;
	wire _w16049_ ;
	wire _w16048_ ;
	wire _w16047_ ;
	wire _w16046_ ;
	wire _w16045_ ;
	wire _w16044_ ;
	wire _w16043_ ;
	wire _w16042_ ;
	wire _w16041_ ;
	wire _w16040_ ;
	wire _w16039_ ;
	wire _w16038_ ;
	wire _w16037_ ;
	wire _w16036_ ;
	wire _w16035_ ;
	wire _w16034_ ;
	wire _w16033_ ;
	wire _w16032_ ;
	wire _w16031_ ;
	wire _w16030_ ;
	wire _w16029_ ;
	wire _w16028_ ;
	wire _w16027_ ;
	wire _w16026_ ;
	wire _w16025_ ;
	wire _w16024_ ;
	wire _w16023_ ;
	wire _w16022_ ;
	wire _w16021_ ;
	wire _w16020_ ;
	wire _w16019_ ;
	wire _w16018_ ;
	wire _w16017_ ;
	wire _w16016_ ;
	wire _w16015_ ;
	wire _w16014_ ;
	wire _w16013_ ;
	wire _w16012_ ;
	wire _w16011_ ;
	wire _w16010_ ;
	wire _w16009_ ;
	wire _w16008_ ;
	wire _w16007_ ;
	wire _w16006_ ;
	wire _w16005_ ;
	wire _w16004_ ;
	wire _w16003_ ;
	wire _w16002_ ;
	wire _w16001_ ;
	wire _w16000_ ;
	wire _w15999_ ;
	wire _w15998_ ;
	wire _w15997_ ;
	wire _w15996_ ;
	wire _w15995_ ;
	wire _w15994_ ;
	wire _w15993_ ;
	wire _w15992_ ;
	wire _w15991_ ;
	wire _w15990_ ;
	wire _w15989_ ;
	wire _w15988_ ;
	wire _w15987_ ;
	wire _w15986_ ;
	wire _w15985_ ;
	wire _w15984_ ;
	wire _w15983_ ;
	wire _w15982_ ;
	wire _w15981_ ;
	wire _w15980_ ;
	wire _w15979_ ;
	wire _w15978_ ;
	wire _w15977_ ;
	wire _w15976_ ;
	wire _w15975_ ;
	wire _w15974_ ;
	wire _w15973_ ;
	wire _w15972_ ;
	wire _w15971_ ;
	wire _w15970_ ;
	wire _w15969_ ;
	wire _w15968_ ;
	wire _w15967_ ;
	wire _w15966_ ;
	wire _w15965_ ;
	wire _w15964_ ;
	wire _w15963_ ;
	wire _w15962_ ;
	wire _w15961_ ;
	wire _w15960_ ;
	wire _w15959_ ;
	wire _w15958_ ;
	wire _w15957_ ;
	wire _w15956_ ;
	wire _w15955_ ;
	wire _w15954_ ;
	wire _w15953_ ;
	wire _w15952_ ;
	wire _w15951_ ;
	wire _w15950_ ;
	wire _w15949_ ;
	wire _w15948_ ;
	wire _w15947_ ;
	wire _w15946_ ;
	wire _w15945_ ;
	wire _w15944_ ;
	wire _w15943_ ;
	wire _w15942_ ;
	wire _w15941_ ;
	wire _w15940_ ;
	wire _w15939_ ;
	wire _w15938_ ;
	wire _w15937_ ;
	wire _w15936_ ;
	wire _w15935_ ;
	wire _w15934_ ;
	wire _w15933_ ;
	wire _w15932_ ;
	wire _w15931_ ;
	wire _w15930_ ;
	wire _w15929_ ;
	wire _w15928_ ;
	wire _w15927_ ;
	wire _w15926_ ;
	wire _w15925_ ;
	wire _w15924_ ;
	wire _w15923_ ;
	wire _w15922_ ;
	wire _w15921_ ;
	wire _w15920_ ;
	wire _w15919_ ;
	wire _w15918_ ;
	wire _w15917_ ;
	wire _w15916_ ;
	wire _w15915_ ;
	wire _w15914_ ;
	wire _w15913_ ;
	wire _w15912_ ;
	wire _w15911_ ;
	wire _w15910_ ;
	wire _w15909_ ;
	wire _w15908_ ;
	wire _w15907_ ;
	wire _w15906_ ;
	wire _w15905_ ;
	wire _w15904_ ;
	wire _w15903_ ;
	wire _w15902_ ;
	wire _w15901_ ;
	wire _w15900_ ;
	wire _w15899_ ;
	wire _w15898_ ;
	wire _w15897_ ;
	wire _w15896_ ;
	wire _w15895_ ;
	wire _w15894_ ;
	wire _w15893_ ;
	wire _w15892_ ;
	wire _w15891_ ;
	wire _w15890_ ;
	wire _w15889_ ;
	wire _w15888_ ;
	wire _w15887_ ;
	wire _w15886_ ;
	wire _w15885_ ;
	wire _w15884_ ;
	wire _w15883_ ;
	wire _w15882_ ;
	wire _w15881_ ;
	wire _w15880_ ;
	wire _w15879_ ;
	wire _w15878_ ;
	wire _w15877_ ;
	wire _w15876_ ;
	wire _w15875_ ;
	wire _w15874_ ;
	wire _w15873_ ;
	wire _w15872_ ;
	wire _w15871_ ;
	wire _w15870_ ;
	wire _w15869_ ;
	wire _w15868_ ;
	wire _w15867_ ;
	wire _w15866_ ;
	wire _w15865_ ;
	wire _w15864_ ;
	wire _w15863_ ;
	wire _w15862_ ;
	wire _w15861_ ;
	wire _w15860_ ;
	wire _w15859_ ;
	wire _w15858_ ;
	wire _w15857_ ;
	wire _w15856_ ;
	wire _w15855_ ;
	wire _w15854_ ;
	wire _w15853_ ;
	wire _w15852_ ;
	wire _w15851_ ;
	wire _w15850_ ;
	wire _w15849_ ;
	wire _w15848_ ;
	wire _w15847_ ;
	wire _w15846_ ;
	wire _w15845_ ;
	wire _w15844_ ;
	wire _w15843_ ;
	wire _w15842_ ;
	wire _w15841_ ;
	wire _w15840_ ;
	wire _w15839_ ;
	wire _w15838_ ;
	wire _w15837_ ;
	wire _w15836_ ;
	wire _w15835_ ;
	wire _w15834_ ;
	wire _w15833_ ;
	wire _w15832_ ;
	wire _w15831_ ;
	wire _w15830_ ;
	wire _w15829_ ;
	wire _w15828_ ;
	wire _w15827_ ;
	wire _w15826_ ;
	wire _w15825_ ;
	wire _w15824_ ;
	wire _w15823_ ;
	wire _w15822_ ;
	wire _w15821_ ;
	wire _w15820_ ;
	wire _w15819_ ;
	wire _w15818_ ;
	wire _w15817_ ;
	wire _w15816_ ;
	wire _w15815_ ;
	wire _w15814_ ;
	wire _w15813_ ;
	wire _w15812_ ;
	wire _w15811_ ;
	wire _w15810_ ;
	wire _w15809_ ;
	wire _w15808_ ;
	wire _w15807_ ;
	wire _w15806_ ;
	wire _w15805_ ;
	wire _w15804_ ;
	wire _w15803_ ;
	wire _w15802_ ;
	wire _w15801_ ;
	wire _w15800_ ;
	wire _w15799_ ;
	wire _w15798_ ;
	wire _w15797_ ;
	wire _w15796_ ;
	wire _w15795_ ;
	wire _w15794_ ;
	wire _w15793_ ;
	wire _w15792_ ;
	wire _w15791_ ;
	wire _w15790_ ;
	wire _w15789_ ;
	wire _w15788_ ;
	wire _w15787_ ;
	wire _w15786_ ;
	wire _w15785_ ;
	wire _w15784_ ;
	wire _w15783_ ;
	wire _w15782_ ;
	wire _w15781_ ;
	wire _w15780_ ;
	wire _w15779_ ;
	wire _w15778_ ;
	wire _w15777_ ;
	wire _w15776_ ;
	wire _w15775_ ;
	wire _w15774_ ;
	wire _w15773_ ;
	wire _w15772_ ;
	wire _w15771_ ;
	wire _w15770_ ;
	wire _w15769_ ;
	wire _w15768_ ;
	wire _w15767_ ;
	wire _w15766_ ;
	wire _w15765_ ;
	wire _w15764_ ;
	wire _w15763_ ;
	wire _w15762_ ;
	wire _w15761_ ;
	wire _w15760_ ;
	wire _w15759_ ;
	wire _w15758_ ;
	wire _w15757_ ;
	wire _w15756_ ;
	wire _w15755_ ;
	wire _w15754_ ;
	wire _w15753_ ;
	wire _w15752_ ;
	wire _w15751_ ;
	wire _w15750_ ;
	wire _w15749_ ;
	wire _w15748_ ;
	wire _w15747_ ;
	wire _w15746_ ;
	wire _w15745_ ;
	wire _w15744_ ;
	wire _w15743_ ;
	wire _w15742_ ;
	wire _w15741_ ;
	wire _w15740_ ;
	wire _w15739_ ;
	wire _w15738_ ;
	wire _w15737_ ;
	wire _w15736_ ;
	wire _w15735_ ;
	wire _w15734_ ;
	wire _w15733_ ;
	wire _w15732_ ;
	wire _w15731_ ;
	wire _w15730_ ;
	wire _w15729_ ;
	wire _w15728_ ;
	wire _w15727_ ;
	wire _w15726_ ;
	wire _w15725_ ;
	wire _w15724_ ;
	wire _w15723_ ;
	wire _w15722_ ;
	wire _w15721_ ;
	wire _w15720_ ;
	wire _w15719_ ;
	wire _w15718_ ;
	wire _w15717_ ;
	wire _w15716_ ;
	wire _w15715_ ;
	wire _w15714_ ;
	wire _w15713_ ;
	wire _w15712_ ;
	wire _w15711_ ;
	wire _w15710_ ;
	wire _w15709_ ;
	wire _w15708_ ;
	wire _w15707_ ;
	wire _w15706_ ;
	wire _w15705_ ;
	wire _w15704_ ;
	wire _w15703_ ;
	wire _w15702_ ;
	wire _w15701_ ;
	wire _w15700_ ;
	wire _w15699_ ;
	wire _w15698_ ;
	wire _w15697_ ;
	wire _w15696_ ;
	wire _w15695_ ;
	wire _w15694_ ;
	wire _w15693_ ;
	wire _w15692_ ;
	wire _w15691_ ;
	wire _w15690_ ;
	wire _w15689_ ;
	wire _w15688_ ;
	wire _w15687_ ;
	wire _w15686_ ;
	wire _w15685_ ;
	wire _w15684_ ;
	wire _w15683_ ;
	wire _w15682_ ;
	wire _w15681_ ;
	wire _w15680_ ;
	wire _w15679_ ;
	wire _w15678_ ;
	wire _w15677_ ;
	wire _w15676_ ;
	wire _w15675_ ;
	wire _w15674_ ;
	wire _w15673_ ;
	wire _w15672_ ;
	wire _w15671_ ;
	wire _w15670_ ;
	wire _w15669_ ;
	wire _w15668_ ;
	wire _w15667_ ;
	wire _w15666_ ;
	wire _w15665_ ;
	wire _w15664_ ;
	wire _w15663_ ;
	wire _w15662_ ;
	wire _w15661_ ;
	wire _w15660_ ;
	wire _w15659_ ;
	wire _w15658_ ;
	wire _w15657_ ;
	wire _w15656_ ;
	wire _w15655_ ;
	wire _w15654_ ;
	wire _w15653_ ;
	wire _w15652_ ;
	wire _w15651_ ;
	wire _w15650_ ;
	wire _w15649_ ;
	wire _w15648_ ;
	wire _w15647_ ;
	wire _w15646_ ;
	wire _w15645_ ;
	wire _w15644_ ;
	wire _w15643_ ;
	wire _w15642_ ;
	wire _w15641_ ;
	wire _w15640_ ;
	wire _w15639_ ;
	wire _w15638_ ;
	wire _w15637_ ;
	wire _w15636_ ;
	wire _w15635_ ;
	wire _w15634_ ;
	wire _w15633_ ;
	wire _w15632_ ;
	wire _w15631_ ;
	wire _w15630_ ;
	wire _w15629_ ;
	wire _w15628_ ;
	wire _w15627_ ;
	wire _w15626_ ;
	wire _w15625_ ;
	wire _w15624_ ;
	wire _w15623_ ;
	wire _w15622_ ;
	wire _w15621_ ;
	wire _w15620_ ;
	wire _w15619_ ;
	wire _w15618_ ;
	wire _w15617_ ;
	wire _w15616_ ;
	wire _w15615_ ;
	wire _w15614_ ;
	wire _w15613_ ;
	wire _w15612_ ;
	wire _w15611_ ;
	wire _w15610_ ;
	wire _w15609_ ;
	wire _w15608_ ;
	wire _w15607_ ;
	wire _w15606_ ;
	wire _w15605_ ;
	wire _w15604_ ;
	wire _w15603_ ;
	wire _w15602_ ;
	wire _w15601_ ;
	wire _w15600_ ;
	wire _w15599_ ;
	wire _w15598_ ;
	wire _w15597_ ;
	wire _w15596_ ;
	wire _w15595_ ;
	wire _w15594_ ;
	wire _w15593_ ;
	wire _w15592_ ;
	wire _w15591_ ;
	wire _w15590_ ;
	wire _w15589_ ;
	wire _w15588_ ;
	wire _w15587_ ;
	wire _w15586_ ;
	wire _w15585_ ;
	wire _w15584_ ;
	wire _w15583_ ;
	wire _w15582_ ;
	wire _w15581_ ;
	wire _w15580_ ;
	wire _w15579_ ;
	wire _w15578_ ;
	wire _w15577_ ;
	wire _w15576_ ;
	wire _w15575_ ;
	wire _w15574_ ;
	wire _w15573_ ;
	wire _w15572_ ;
	wire _w15571_ ;
	wire _w15570_ ;
	wire _w15569_ ;
	wire _w15568_ ;
	wire _w15567_ ;
	wire _w15566_ ;
	wire _w15565_ ;
	wire _w15564_ ;
	wire _w15563_ ;
	wire _w15562_ ;
	wire _w15561_ ;
	wire _w15560_ ;
	wire _w15559_ ;
	wire _w15558_ ;
	wire _w15557_ ;
	wire _w15556_ ;
	wire _w15555_ ;
	wire _w15554_ ;
	wire _w15553_ ;
	wire _w15552_ ;
	wire _w15551_ ;
	wire _w15550_ ;
	wire _w15549_ ;
	wire _w15548_ ;
	wire _w15547_ ;
	wire _w15546_ ;
	wire _w15545_ ;
	wire _w15544_ ;
	wire _w15543_ ;
	wire _w15542_ ;
	wire _w15541_ ;
	wire _w15540_ ;
	wire _w15539_ ;
	wire _w15538_ ;
	wire _w15537_ ;
	wire _w15536_ ;
	wire _w15535_ ;
	wire _w15534_ ;
	wire _w15533_ ;
	wire _w15532_ ;
	wire _w15531_ ;
	wire _w15530_ ;
	wire _w15529_ ;
	wire _w15528_ ;
	wire _w15527_ ;
	wire _w15526_ ;
	wire _w15525_ ;
	wire _w15524_ ;
	wire _w15523_ ;
	wire _w15522_ ;
	wire _w15521_ ;
	wire _w15520_ ;
	wire _w15519_ ;
	wire _w15518_ ;
	wire _w15517_ ;
	wire _w15516_ ;
	wire _w15515_ ;
	wire _w15514_ ;
	wire _w15513_ ;
	wire _w15512_ ;
	wire _w15511_ ;
	wire _w15510_ ;
	wire _w15509_ ;
	wire _w15508_ ;
	wire _w15507_ ;
	wire _w15506_ ;
	wire _w15505_ ;
	wire _w15504_ ;
	wire _w15503_ ;
	wire _w15502_ ;
	wire _w15501_ ;
	wire _w15500_ ;
	wire _w15499_ ;
	wire _w15498_ ;
	wire _w15497_ ;
	wire _w15496_ ;
	wire _w15495_ ;
	wire _w15494_ ;
	wire _w15493_ ;
	wire _w15492_ ;
	wire _w15491_ ;
	wire _w15490_ ;
	wire _w15489_ ;
	wire _w15488_ ;
	wire _w15487_ ;
	wire _w15486_ ;
	wire _w15485_ ;
	wire _w15484_ ;
	wire _w15483_ ;
	wire _w15482_ ;
	wire _w15481_ ;
	wire _w15480_ ;
	wire _w15479_ ;
	wire _w15478_ ;
	wire _w15477_ ;
	wire _w15476_ ;
	wire _w15475_ ;
	wire _w15474_ ;
	wire _w15473_ ;
	wire _w15472_ ;
	wire _w15471_ ;
	wire _w15470_ ;
	wire _w15469_ ;
	wire _w15468_ ;
	wire _w15467_ ;
	wire _w15466_ ;
	wire _w15465_ ;
	wire _w15464_ ;
	wire _w15463_ ;
	wire _w15462_ ;
	wire _w15461_ ;
	wire _w15460_ ;
	wire _w15459_ ;
	wire _w15458_ ;
	wire _w15457_ ;
	wire _w15456_ ;
	wire _w15455_ ;
	wire _w15454_ ;
	wire _w15453_ ;
	wire _w15452_ ;
	wire _w15451_ ;
	wire _w15450_ ;
	wire _w15449_ ;
	wire _w15448_ ;
	wire _w15447_ ;
	wire _w15446_ ;
	wire _w15445_ ;
	wire _w15444_ ;
	wire _w15443_ ;
	wire _w15442_ ;
	wire _w15441_ ;
	wire _w15440_ ;
	wire _w15439_ ;
	wire _w15438_ ;
	wire _w15437_ ;
	wire _w15436_ ;
	wire _w15435_ ;
	wire _w15434_ ;
	wire _w15433_ ;
	wire _w15432_ ;
	wire _w15431_ ;
	wire _w15430_ ;
	wire _w15429_ ;
	wire _w15428_ ;
	wire _w15427_ ;
	wire _w15426_ ;
	wire _w15425_ ;
	wire _w15424_ ;
	wire _w15423_ ;
	wire _w15422_ ;
	wire _w15421_ ;
	wire _w15420_ ;
	wire _w15419_ ;
	wire _w15418_ ;
	wire _w15417_ ;
	wire _w15416_ ;
	wire _w15415_ ;
	wire _w15414_ ;
	wire _w15413_ ;
	wire _w15412_ ;
	wire _w15411_ ;
	wire _w15410_ ;
	wire _w15409_ ;
	wire _w15408_ ;
	wire _w15407_ ;
	wire _w15406_ ;
	wire _w15405_ ;
	wire _w15404_ ;
	wire _w15403_ ;
	wire _w15402_ ;
	wire _w15401_ ;
	wire _w15400_ ;
	wire _w15399_ ;
	wire _w15398_ ;
	wire _w15397_ ;
	wire _w15396_ ;
	wire _w15395_ ;
	wire _w15394_ ;
	wire _w15393_ ;
	wire _w15392_ ;
	wire _w15391_ ;
	wire _w15390_ ;
	wire _w15389_ ;
	wire _w15388_ ;
	wire _w15387_ ;
	wire _w15386_ ;
	wire _w15385_ ;
	wire _w15384_ ;
	wire _w15383_ ;
	wire _w15382_ ;
	wire _w15381_ ;
	wire _w15380_ ;
	wire _w15379_ ;
	wire _w15378_ ;
	wire _w15377_ ;
	wire _w15376_ ;
	wire _w15375_ ;
	wire _w15374_ ;
	wire _w15373_ ;
	wire _w15372_ ;
	wire _w15371_ ;
	wire _w15370_ ;
	wire _w15369_ ;
	wire _w15368_ ;
	wire _w15367_ ;
	wire _w15366_ ;
	wire _w15365_ ;
	wire _w15364_ ;
	wire _w15363_ ;
	wire _w15362_ ;
	wire _w15361_ ;
	wire _w15360_ ;
	wire _w15359_ ;
	wire _w15358_ ;
	wire _w15357_ ;
	wire _w15356_ ;
	wire _w15355_ ;
	wire _w15354_ ;
	wire _w15353_ ;
	wire _w15352_ ;
	wire _w15351_ ;
	wire _w15350_ ;
	wire _w15349_ ;
	wire _w15348_ ;
	wire _w15347_ ;
	wire _w15346_ ;
	wire _w15345_ ;
	wire _w15344_ ;
	wire _w15343_ ;
	wire _w15342_ ;
	wire _w15341_ ;
	wire _w15340_ ;
	wire _w15339_ ;
	wire _w15338_ ;
	wire _w15337_ ;
	wire _w15336_ ;
	wire _w15335_ ;
	wire _w15334_ ;
	wire _w15333_ ;
	wire _w15332_ ;
	wire _w15331_ ;
	wire _w15330_ ;
	wire _w15329_ ;
	wire _w15328_ ;
	wire _w15327_ ;
	wire _w15326_ ;
	wire _w15325_ ;
	wire _w15324_ ;
	wire _w15323_ ;
	wire _w15322_ ;
	wire _w15321_ ;
	wire _w15320_ ;
	wire _w15319_ ;
	wire _w15318_ ;
	wire _w15317_ ;
	wire _w15316_ ;
	wire _w15315_ ;
	wire _w15314_ ;
	wire _w15313_ ;
	wire _w15312_ ;
	wire _w15311_ ;
	wire _w15310_ ;
	wire _w15309_ ;
	wire _w15308_ ;
	wire _w15307_ ;
	wire _w15306_ ;
	wire _w15305_ ;
	wire _w15304_ ;
	wire _w15303_ ;
	wire _w15302_ ;
	wire _w15301_ ;
	wire _w15300_ ;
	wire _w15299_ ;
	wire _w15298_ ;
	wire _w15297_ ;
	wire _w15296_ ;
	wire _w15295_ ;
	wire _w15294_ ;
	wire _w15293_ ;
	wire _w15292_ ;
	wire _w15291_ ;
	wire _w15290_ ;
	wire _w15289_ ;
	wire _w15288_ ;
	wire _w15287_ ;
	wire _w15286_ ;
	wire _w15285_ ;
	wire _w15284_ ;
	wire _w15283_ ;
	wire _w15282_ ;
	wire _w15281_ ;
	wire _w15280_ ;
	wire _w15279_ ;
	wire _w15278_ ;
	wire _w15277_ ;
	wire _w15276_ ;
	wire _w15275_ ;
	wire _w15274_ ;
	wire _w15273_ ;
	wire _w15272_ ;
	wire _w15271_ ;
	wire _w15270_ ;
	wire _w15269_ ;
	wire _w15268_ ;
	wire _w15267_ ;
	wire _w15266_ ;
	wire _w15265_ ;
	wire _w15264_ ;
	wire _w15263_ ;
	wire _w15262_ ;
	wire _w15261_ ;
	wire _w15260_ ;
	wire _w15259_ ;
	wire _w15258_ ;
	wire _w15257_ ;
	wire _w15256_ ;
	wire _w15255_ ;
	wire _w15254_ ;
	wire _w15253_ ;
	wire _w15252_ ;
	wire _w15251_ ;
	wire _w15250_ ;
	wire _w15249_ ;
	wire _w15248_ ;
	wire _w15247_ ;
	wire _w15246_ ;
	wire _w15245_ ;
	wire _w15244_ ;
	wire _w15243_ ;
	wire _w15242_ ;
	wire _w15241_ ;
	wire _w15240_ ;
	wire _w15239_ ;
	wire _w15238_ ;
	wire _w15237_ ;
	wire _w15236_ ;
	wire _w15235_ ;
	wire _w15234_ ;
	wire _w15233_ ;
	wire _w15232_ ;
	wire _w15231_ ;
	wire _w15230_ ;
	wire _w15229_ ;
	wire _w15228_ ;
	wire _w15227_ ;
	wire _w15226_ ;
	wire _w15225_ ;
	wire _w15224_ ;
	wire _w15223_ ;
	wire _w15222_ ;
	wire _w15221_ ;
	wire _w15220_ ;
	wire _w15219_ ;
	wire _w15218_ ;
	wire _w15217_ ;
	wire _w15216_ ;
	wire _w15215_ ;
	wire _w15214_ ;
	wire _w15213_ ;
	wire _w15212_ ;
	wire _w15211_ ;
	wire _w15210_ ;
	wire _w15209_ ;
	wire _w15208_ ;
	wire _w15207_ ;
	wire _w15206_ ;
	wire _w15205_ ;
	wire _w15204_ ;
	wire _w15203_ ;
	wire _w15202_ ;
	wire _w15201_ ;
	wire _w15200_ ;
	wire _w15199_ ;
	wire _w15198_ ;
	wire _w15197_ ;
	wire _w15196_ ;
	wire _w15195_ ;
	wire _w15194_ ;
	wire _w15193_ ;
	wire _w15192_ ;
	wire _w15191_ ;
	wire _w15190_ ;
	wire _w15189_ ;
	wire _w15188_ ;
	wire _w15187_ ;
	wire _w15186_ ;
	wire _w15185_ ;
	wire _w15184_ ;
	wire _w15183_ ;
	wire _w15182_ ;
	wire _w15181_ ;
	wire _w15180_ ;
	wire _w15179_ ;
	wire _w15178_ ;
	wire _w15177_ ;
	wire _w15176_ ;
	wire _w15175_ ;
	wire _w15174_ ;
	wire _w15173_ ;
	wire _w15172_ ;
	wire _w15171_ ;
	wire _w15170_ ;
	wire _w15169_ ;
	wire _w15168_ ;
	wire _w15167_ ;
	wire _w15166_ ;
	wire _w15165_ ;
	wire _w15164_ ;
	wire _w15163_ ;
	wire _w15162_ ;
	wire _w15161_ ;
	wire _w15160_ ;
	wire _w15159_ ;
	wire _w15158_ ;
	wire _w15157_ ;
	wire _w15156_ ;
	wire _w15155_ ;
	wire _w15154_ ;
	wire _w15153_ ;
	wire _w15152_ ;
	wire _w15151_ ;
	wire _w15150_ ;
	wire _w15149_ ;
	wire _w15148_ ;
	wire _w15147_ ;
	wire _w15146_ ;
	wire _w15145_ ;
	wire _w15144_ ;
	wire _w15143_ ;
	wire _w15142_ ;
	wire _w15141_ ;
	wire _w15140_ ;
	wire _w15139_ ;
	wire _w15138_ ;
	wire _w15137_ ;
	wire _w15136_ ;
	wire _w15135_ ;
	wire _w15134_ ;
	wire _w15133_ ;
	wire _w15132_ ;
	wire _w15131_ ;
	wire _w15130_ ;
	wire _w15129_ ;
	wire _w15128_ ;
	wire _w15127_ ;
	wire _w15126_ ;
	wire _w15125_ ;
	wire _w15124_ ;
	wire _w15123_ ;
	wire _w15122_ ;
	wire _w15121_ ;
	wire _w15120_ ;
	wire _w15119_ ;
	wire _w15118_ ;
	wire _w15117_ ;
	wire _w15116_ ;
	wire _w15115_ ;
	wire _w15114_ ;
	wire _w15113_ ;
	wire _w15112_ ;
	wire _w15111_ ;
	wire _w15110_ ;
	wire _w15109_ ;
	wire _w15108_ ;
	wire _w15107_ ;
	wire _w15106_ ;
	wire _w15105_ ;
	wire _w15104_ ;
	wire _w15103_ ;
	wire _w15102_ ;
	wire _w15101_ ;
	wire _w15100_ ;
	wire _w15099_ ;
	wire _w15098_ ;
	wire _w15097_ ;
	wire _w15096_ ;
	wire _w15095_ ;
	wire _w15094_ ;
	wire _w15093_ ;
	wire _w15092_ ;
	wire _w15091_ ;
	wire _w15090_ ;
	wire _w15089_ ;
	wire _w15088_ ;
	wire _w15087_ ;
	wire _w15086_ ;
	wire _w15085_ ;
	wire _w15084_ ;
	wire _w15083_ ;
	wire _w15082_ ;
	wire _w15081_ ;
	wire _w15080_ ;
	wire _w15079_ ;
	wire _w15078_ ;
	wire _w15077_ ;
	wire _w15076_ ;
	wire _w15075_ ;
	wire _w15074_ ;
	wire _w15073_ ;
	wire _w15072_ ;
	wire _w15071_ ;
	wire _w15070_ ;
	wire _w15069_ ;
	wire _w15068_ ;
	wire _w15067_ ;
	wire _w15066_ ;
	wire _w15065_ ;
	wire _w15064_ ;
	wire _w15063_ ;
	wire _w15062_ ;
	wire _w15061_ ;
	wire _w15060_ ;
	wire _w15059_ ;
	wire _w15058_ ;
	wire _w15057_ ;
	wire _w15056_ ;
	wire _w15055_ ;
	wire _w15054_ ;
	wire _w15053_ ;
	wire _w15052_ ;
	wire _w15051_ ;
	wire _w15050_ ;
	wire _w15049_ ;
	wire _w15048_ ;
	wire _w15047_ ;
	wire _w15046_ ;
	wire _w15045_ ;
	wire _w15044_ ;
	wire _w15043_ ;
	wire _w15042_ ;
	wire _w15041_ ;
	wire _w15040_ ;
	wire _w15039_ ;
	wire _w15038_ ;
	wire _w15037_ ;
	wire _w15036_ ;
	wire _w15035_ ;
	wire _w15034_ ;
	wire _w15033_ ;
	wire _w15032_ ;
	wire _w15031_ ;
	wire _w15030_ ;
	wire _w15029_ ;
	wire _w15028_ ;
	wire _w15027_ ;
	wire _w15026_ ;
	wire _w15025_ ;
	wire _w15024_ ;
	wire _w15023_ ;
	wire _w15022_ ;
	wire _w15021_ ;
	wire _w15020_ ;
	wire _w15019_ ;
	wire _w15018_ ;
	wire _w15017_ ;
	wire _w15016_ ;
	wire _w15015_ ;
	wire _w15014_ ;
	wire _w15013_ ;
	wire _w15012_ ;
	wire _w15011_ ;
	wire _w15010_ ;
	wire _w15009_ ;
	wire _w15008_ ;
	wire _w15007_ ;
	wire _w15006_ ;
	wire _w15005_ ;
	wire _w15004_ ;
	wire _w15003_ ;
	wire _w15002_ ;
	wire _w15001_ ;
	wire _w15000_ ;
	wire _w14999_ ;
	wire _w14998_ ;
	wire _w14997_ ;
	wire _w14996_ ;
	wire _w14995_ ;
	wire _w14994_ ;
	wire _w14993_ ;
	wire _w14992_ ;
	wire _w14991_ ;
	wire _w14990_ ;
	wire _w14989_ ;
	wire _w14988_ ;
	wire _w14987_ ;
	wire _w14986_ ;
	wire _w14985_ ;
	wire _w14984_ ;
	wire _w14983_ ;
	wire _w14982_ ;
	wire _w14981_ ;
	wire _w14980_ ;
	wire _w14979_ ;
	wire _w14978_ ;
	wire _w14977_ ;
	wire _w14976_ ;
	wire _w14975_ ;
	wire _w14974_ ;
	wire _w14973_ ;
	wire _w14972_ ;
	wire _w14971_ ;
	wire _w14970_ ;
	wire _w14969_ ;
	wire _w14968_ ;
	wire _w14967_ ;
	wire _w14966_ ;
	wire _w14965_ ;
	wire _w14964_ ;
	wire _w14963_ ;
	wire _w14962_ ;
	wire _w14961_ ;
	wire _w14960_ ;
	wire _w14959_ ;
	wire _w14958_ ;
	wire _w14957_ ;
	wire _w14956_ ;
	wire _w14955_ ;
	wire _w14954_ ;
	wire _w14953_ ;
	wire _w14952_ ;
	wire _w14951_ ;
	wire _w14950_ ;
	wire _w14949_ ;
	wire _w14948_ ;
	wire _w14947_ ;
	wire _w14946_ ;
	wire _w14945_ ;
	wire _w14944_ ;
	wire _w14943_ ;
	wire _w14942_ ;
	wire _w14941_ ;
	wire _w14940_ ;
	wire _w14939_ ;
	wire _w14938_ ;
	wire _w14937_ ;
	wire _w14936_ ;
	wire _w14935_ ;
	wire _w14934_ ;
	wire _w14933_ ;
	wire _w14932_ ;
	wire _w14931_ ;
	wire _w14930_ ;
	wire _w14929_ ;
	wire _w14928_ ;
	wire _w14927_ ;
	wire _w14926_ ;
	wire _w14925_ ;
	wire _w14924_ ;
	wire _w14923_ ;
	wire _w14922_ ;
	wire _w14921_ ;
	wire _w14920_ ;
	wire _w14919_ ;
	wire _w14918_ ;
	wire _w14917_ ;
	wire _w14916_ ;
	wire _w14915_ ;
	wire _w14914_ ;
	wire _w14913_ ;
	wire _w14912_ ;
	wire _w14911_ ;
	wire _w14910_ ;
	wire _w14909_ ;
	wire _w14908_ ;
	wire _w14907_ ;
	wire _w14906_ ;
	wire _w14905_ ;
	wire _w14904_ ;
	wire _w14903_ ;
	wire _w14902_ ;
	wire _w14901_ ;
	wire _w14900_ ;
	wire _w14899_ ;
	wire _w14898_ ;
	wire _w14897_ ;
	wire _w14896_ ;
	wire _w14895_ ;
	wire _w14894_ ;
	wire _w14893_ ;
	wire _w14892_ ;
	wire _w14891_ ;
	wire _w14890_ ;
	wire _w14889_ ;
	wire _w14888_ ;
	wire _w14887_ ;
	wire _w14886_ ;
	wire _w14885_ ;
	wire _w14884_ ;
	wire _w14883_ ;
	wire _w14882_ ;
	wire _w14881_ ;
	wire _w14880_ ;
	wire _w14879_ ;
	wire _w14878_ ;
	wire _w14877_ ;
	wire _w14876_ ;
	wire _w14875_ ;
	wire _w14874_ ;
	wire _w14873_ ;
	wire _w14872_ ;
	wire _w14871_ ;
	wire _w14870_ ;
	wire _w14869_ ;
	wire _w14868_ ;
	wire _w14867_ ;
	wire _w14866_ ;
	wire _w14865_ ;
	wire _w14864_ ;
	wire _w14863_ ;
	wire _w14862_ ;
	wire _w14861_ ;
	wire _w14860_ ;
	wire _w14859_ ;
	wire _w14858_ ;
	wire _w14857_ ;
	wire _w14856_ ;
	wire _w14855_ ;
	wire _w14854_ ;
	wire _w14853_ ;
	wire _w14852_ ;
	wire _w14851_ ;
	wire _w14850_ ;
	wire _w14849_ ;
	wire _w14848_ ;
	wire _w14847_ ;
	wire _w14846_ ;
	wire _w14845_ ;
	wire _w14844_ ;
	wire _w14843_ ;
	wire _w14842_ ;
	wire _w14841_ ;
	wire _w14840_ ;
	wire _w14839_ ;
	wire _w14838_ ;
	wire _w14837_ ;
	wire _w14836_ ;
	wire _w14835_ ;
	wire _w14834_ ;
	wire _w14833_ ;
	wire _w14832_ ;
	wire _w14831_ ;
	wire _w14830_ ;
	wire _w14829_ ;
	wire _w14828_ ;
	wire _w14827_ ;
	wire _w14826_ ;
	wire _w14825_ ;
	wire _w14824_ ;
	wire _w14823_ ;
	wire _w14822_ ;
	wire _w14821_ ;
	wire _w14820_ ;
	wire _w14819_ ;
	wire _w14818_ ;
	wire _w14817_ ;
	wire _w14816_ ;
	wire _w14815_ ;
	wire _w14814_ ;
	wire _w14813_ ;
	wire _w14812_ ;
	wire _w14811_ ;
	wire _w14810_ ;
	wire _w14809_ ;
	wire _w14808_ ;
	wire _w14807_ ;
	wire _w14806_ ;
	wire _w14805_ ;
	wire _w14804_ ;
	wire _w14803_ ;
	wire _w14802_ ;
	wire _w14801_ ;
	wire _w14800_ ;
	wire _w14799_ ;
	wire _w14798_ ;
	wire _w14797_ ;
	wire _w14796_ ;
	wire _w14795_ ;
	wire _w14794_ ;
	wire _w14793_ ;
	wire _w14792_ ;
	wire _w14791_ ;
	wire _w14790_ ;
	wire _w14789_ ;
	wire _w14788_ ;
	wire _w14787_ ;
	wire _w14786_ ;
	wire _w14785_ ;
	wire _w14784_ ;
	wire _w14783_ ;
	wire _w14782_ ;
	wire _w14781_ ;
	wire _w14780_ ;
	wire _w14779_ ;
	wire _w14778_ ;
	wire _w14777_ ;
	wire _w14776_ ;
	wire _w14775_ ;
	wire _w14774_ ;
	wire _w14773_ ;
	wire _w14772_ ;
	wire _w14771_ ;
	wire _w14770_ ;
	wire _w14769_ ;
	wire _w14768_ ;
	wire _w14767_ ;
	wire _w14766_ ;
	wire _w14765_ ;
	wire _w14764_ ;
	wire _w14763_ ;
	wire _w14762_ ;
	wire _w14761_ ;
	wire _w14760_ ;
	wire _w14759_ ;
	wire _w14758_ ;
	wire _w14757_ ;
	wire _w14756_ ;
	wire _w14755_ ;
	wire _w14754_ ;
	wire _w14753_ ;
	wire _w14752_ ;
	wire _w14751_ ;
	wire _w14750_ ;
	wire _w14749_ ;
	wire _w14748_ ;
	wire _w14747_ ;
	wire _w14746_ ;
	wire _w14745_ ;
	wire _w14744_ ;
	wire _w14743_ ;
	wire _w14742_ ;
	wire _w14741_ ;
	wire _w14740_ ;
	wire _w14739_ ;
	wire _w14738_ ;
	wire _w14737_ ;
	wire _w14736_ ;
	wire _w14735_ ;
	wire _w14734_ ;
	wire _w14733_ ;
	wire _w14732_ ;
	wire _w14731_ ;
	wire _w14730_ ;
	wire _w14729_ ;
	wire _w14728_ ;
	wire _w14727_ ;
	wire _w14726_ ;
	wire _w14725_ ;
	wire _w14724_ ;
	wire _w14723_ ;
	wire _w14722_ ;
	wire _w14721_ ;
	wire _w14720_ ;
	wire _w14719_ ;
	wire _w14718_ ;
	wire _w14717_ ;
	wire _w14716_ ;
	wire _w14715_ ;
	wire _w14714_ ;
	wire _w14713_ ;
	wire _w14712_ ;
	wire _w14711_ ;
	wire _w14710_ ;
	wire _w14709_ ;
	wire _w14708_ ;
	wire _w14707_ ;
	wire _w14706_ ;
	wire _w14705_ ;
	wire _w14704_ ;
	wire _w14703_ ;
	wire _w14702_ ;
	wire _w14701_ ;
	wire _w14700_ ;
	wire _w14699_ ;
	wire _w14698_ ;
	wire _w14697_ ;
	wire _w14696_ ;
	wire _w14695_ ;
	wire _w14694_ ;
	wire _w14693_ ;
	wire _w14692_ ;
	wire _w14691_ ;
	wire _w14690_ ;
	wire _w14689_ ;
	wire _w14688_ ;
	wire _w14687_ ;
	wire _w14686_ ;
	wire _w14685_ ;
	wire _w14684_ ;
	wire _w14683_ ;
	wire _w14682_ ;
	wire _w14681_ ;
	wire _w14680_ ;
	wire _w14679_ ;
	wire _w14678_ ;
	wire _w14677_ ;
	wire _w14676_ ;
	wire _w14675_ ;
	wire _w14674_ ;
	wire _w14673_ ;
	wire _w14672_ ;
	wire _w14671_ ;
	wire _w14670_ ;
	wire _w14669_ ;
	wire _w14668_ ;
	wire _w14667_ ;
	wire _w14666_ ;
	wire _w14665_ ;
	wire _w14664_ ;
	wire _w14663_ ;
	wire _w14662_ ;
	wire _w14661_ ;
	wire _w14660_ ;
	wire _w14659_ ;
	wire _w14658_ ;
	wire _w14657_ ;
	wire _w14656_ ;
	wire _w14655_ ;
	wire _w14654_ ;
	wire _w14653_ ;
	wire _w14652_ ;
	wire _w14651_ ;
	wire _w14650_ ;
	wire _w14649_ ;
	wire _w14648_ ;
	wire _w14647_ ;
	wire _w14646_ ;
	wire _w14645_ ;
	wire _w14644_ ;
	wire _w14643_ ;
	wire _w14642_ ;
	wire _w14641_ ;
	wire _w14640_ ;
	wire _w14639_ ;
	wire _w14638_ ;
	wire _w14637_ ;
	wire _w14636_ ;
	wire _w14635_ ;
	wire _w14634_ ;
	wire _w14633_ ;
	wire _w14632_ ;
	wire _w14631_ ;
	wire _w14630_ ;
	wire _w14629_ ;
	wire _w14628_ ;
	wire _w14627_ ;
	wire _w14626_ ;
	wire _w14625_ ;
	wire _w14624_ ;
	wire _w14623_ ;
	wire _w14622_ ;
	wire _w14621_ ;
	wire _w14620_ ;
	wire _w14619_ ;
	wire _w14618_ ;
	wire _w14617_ ;
	wire _w14616_ ;
	wire _w14615_ ;
	wire _w14614_ ;
	wire _w14613_ ;
	wire _w14612_ ;
	wire _w14611_ ;
	wire _w14610_ ;
	wire _w14609_ ;
	wire _w14608_ ;
	wire _w14607_ ;
	wire _w14606_ ;
	wire _w14605_ ;
	wire _w14604_ ;
	wire _w14603_ ;
	wire _w14602_ ;
	wire _w14601_ ;
	wire _w14600_ ;
	wire _w14599_ ;
	wire _w14598_ ;
	wire _w14597_ ;
	wire _w14596_ ;
	wire _w14595_ ;
	wire _w14594_ ;
	wire _w14593_ ;
	wire _w14592_ ;
	wire _w14591_ ;
	wire _w14590_ ;
	wire _w14589_ ;
	wire _w14588_ ;
	wire _w14587_ ;
	wire _w14586_ ;
	wire _w14585_ ;
	wire _w14584_ ;
	wire _w14583_ ;
	wire _w14582_ ;
	wire _w14581_ ;
	wire _w14580_ ;
	wire _w14579_ ;
	wire _w14578_ ;
	wire _w14577_ ;
	wire _w14576_ ;
	wire _w14575_ ;
	wire _w14574_ ;
	wire _w14573_ ;
	wire _w14572_ ;
	wire _w14571_ ;
	wire _w14570_ ;
	wire _w14569_ ;
	wire _w14568_ ;
	wire _w14567_ ;
	wire _w14566_ ;
	wire _w14565_ ;
	wire _w14564_ ;
	wire _w14563_ ;
	wire _w14562_ ;
	wire _w14561_ ;
	wire _w14560_ ;
	wire _w14559_ ;
	wire _w14558_ ;
	wire _w14557_ ;
	wire _w14556_ ;
	wire _w14555_ ;
	wire _w14554_ ;
	wire _w14553_ ;
	wire _w14552_ ;
	wire _w14551_ ;
	wire _w14550_ ;
	wire _w14549_ ;
	wire _w14548_ ;
	wire _w14547_ ;
	wire _w14546_ ;
	wire _w14545_ ;
	wire _w14544_ ;
	wire _w14543_ ;
	wire _w14542_ ;
	wire _w14541_ ;
	wire _w14540_ ;
	wire _w14539_ ;
	wire _w14538_ ;
	wire _w14537_ ;
	wire _w14536_ ;
	wire _w14535_ ;
	wire _w14534_ ;
	wire _w14533_ ;
	wire _w14532_ ;
	wire _w14531_ ;
	wire _w14530_ ;
	wire _w14529_ ;
	wire _w14528_ ;
	wire _w14527_ ;
	wire _w14526_ ;
	wire _w14525_ ;
	wire _w14524_ ;
	wire _w14523_ ;
	wire _w14522_ ;
	wire _w14521_ ;
	wire _w14520_ ;
	wire _w14519_ ;
	wire _w14518_ ;
	wire _w14517_ ;
	wire _w14516_ ;
	wire _w14515_ ;
	wire _w14514_ ;
	wire _w14513_ ;
	wire _w14512_ ;
	wire _w14511_ ;
	wire _w14510_ ;
	wire _w14509_ ;
	wire _w14508_ ;
	wire _w14507_ ;
	wire _w14506_ ;
	wire _w14505_ ;
	wire _w14504_ ;
	wire _w14503_ ;
	wire _w14502_ ;
	wire _w14501_ ;
	wire _w14500_ ;
	wire _w14499_ ;
	wire _w14498_ ;
	wire _w14497_ ;
	wire _w14496_ ;
	wire _w14495_ ;
	wire _w14494_ ;
	wire _w14493_ ;
	wire _w14492_ ;
	wire _w14491_ ;
	wire _w14490_ ;
	wire _w14489_ ;
	wire _w14488_ ;
	wire _w14487_ ;
	wire _w14486_ ;
	wire _w14485_ ;
	wire _w14484_ ;
	wire _w14483_ ;
	wire _w14482_ ;
	wire _w14481_ ;
	wire _w14480_ ;
	wire _w14479_ ;
	wire _w14478_ ;
	wire _w14477_ ;
	wire _w14476_ ;
	wire _w14475_ ;
	wire _w14474_ ;
	wire _w14473_ ;
	wire _w14472_ ;
	wire _w14471_ ;
	wire _w14470_ ;
	wire _w14469_ ;
	wire _w14468_ ;
	wire _w14467_ ;
	wire _w14466_ ;
	wire _w14465_ ;
	wire _w14464_ ;
	wire _w14463_ ;
	wire _w14462_ ;
	wire _w14461_ ;
	wire _w14460_ ;
	wire _w14459_ ;
	wire _w14458_ ;
	wire _w14457_ ;
	wire _w14456_ ;
	wire _w14455_ ;
	wire _w14454_ ;
	wire _w14453_ ;
	wire _w14452_ ;
	wire _w14451_ ;
	wire _w14450_ ;
	wire _w14449_ ;
	wire _w14448_ ;
	wire _w14447_ ;
	wire _w14446_ ;
	wire _w14445_ ;
	wire _w14444_ ;
	wire _w14443_ ;
	wire _w14442_ ;
	wire _w14441_ ;
	wire _w14440_ ;
	wire _w14439_ ;
	wire _w14438_ ;
	wire _w14437_ ;
	wire _w14436_ ;
	wire _w14435_ ;
	wire _w14434_ ;
	wire _w14433_ ;
	wire _w14432_ ;
	wire _w14431_ ;
	wire _w14430_ ;
	wire _w14429_ ;
	wire _w14428_ ;
	wire _w14427_ ;
	wire _w14426_ ;
	wire _w14425_ ;
	wire _w14424_ ;
	wire _w14423_ ;
	wire _w14422_ ;
	wire _w14421_ ;
	wire _w14420_ ;
	wire _w14419_ ;
	wire _w14418_ ;
	wire _w14417_ ;
	wire _w14416_ ;
	wire _w14415_ ;
	wire _w14414_ ;
	wire _w14413_ ;
	wire _w14412_ ;
	wire _w14411_ ;
	wire _w14410_ ;
	wire _w14409_ ;
	wire _w14408_ ;
	wire _w14407_ ;
	wire _w14406_ ;
	wire _w14405_ ;
	wire _w14404_ ;
	wire _w14403_ ;
	wire _w14402_ ;
	wire _w14401_ ;
	wire _w14400_ ;
	wire _w14399_ ;
	wire _w14398_ ;
	wire _w14397_ ;
	wire _w14396_ ;
	wire _w14395_ ;
	wire _w14394_ ;
	wire _w14393_ ;
	wire _w14392_ ;
	wire _w14391_ ;
	wire _w14390_ ;
	wire _w14389_ ;
	wire _w14388_ ;
	wire _w14387_ ;
	wire _w14386_ ;
	wire _w14385_ ;
	wire _w14384_ ;
	wire _w14383_ ;
	wire _w14382_ ;
	wire _w14381_ ;
	wire _w14380_ ;
	wire _w14379_ ;
	wire _w14378_ ;
	wire _w14377_ ;
	wire _w14376_ ;
	wire _w14375_ ;
	wire _w14374_ ;
	wire _w14373_ ;
	wire _w14372_ ;
	wire _w14371_ ;
	wire _w14370_ ;
	wire _w14369_ ;
	wire _w14368_ ;
	wire _w14367_ ;
	wire _w14366_ ;
	wire _w14365_ ;
	wire _w14364_ ;
	wire _w14363_ ;
	wire _w14362_ ;
	wire _w14361_ ;
	wire _w14360_ ;
	wire _w14359_ ;
	wire _w14358_ ;
	wire _w14357_ ;
	wire _w14356_ ;
	wire _w14355_ ;
	wire _w14354_ ;
	wire _w14353_ ;
	wire _w14352_ ;
	wire _w14351_ ;
	wire _w14350_ ;
	wire _w14349_ ;
	wire _w14348_ ;
	wire _w14347_ ;
	wire _w14346_ ;
	wire _w14345_ ;
	wire _w14344_ ;
	wire _w14343_ ;
	wire _w14342_ ;
	wire _w14341_ ;
	wire _w14340_ ;
	wire _w14339_ ;
	wire _w14338_ ;
	wire _w14337_ ;
	wire _w14336_ ;
	wire _w14335_ ;
	wire _w14334_ ;
	wire _w14333_ ;
	wire _w14332_ ;
	wire _w14331_ ;
	wire _w14330_ ;
	wire _w14329_ ;
	wire _w14328_ ;
	wire _w14327_ ;
	wire _w14326_ ;
	wire _w14325_ ;
	wire _w14324_ ;
	wire _w14323_ ;
	wire _w14322_ ;
	wire _w14321_ ;
	wire _w9134_ ;
	wire _w9133_ ;
	wire _w9132_ ;
	wire _w9131_ ;
	wire _w9130_ ;
	wire _w9129_ ;
	wire _w9128_ ;
	wire _w9127_ ;
	wire _w9126_ ;
	wire _w9125_ ;
	wire _w9124_ ;
	wire _w9123_ ;
	wire _w9122_ ;
	wire _w9121_ ;
	wire _w9120_ ;
	wire _w9119_ ;
	wire _w9118_ ;
	wire _w9117_ ;
	wire _w9116_ ;
	wire _w9115_ ;
	wire _w9114_ ;
	wire _w9113_ ;
	wire _w9112_ ;
	wire _w9111_ ;
	wire _w9110_ ;
	wire _w9109_ ;
	wire _w9108_ ;
	wire _w9107_ ;
	wire _w9106_ ;
	wire _w9105_ ;
	wire _w9104_ ;
	wire _w9103_ ;
	wire _w9102_ ;
	wire _w9101_ ;
	wire _w9100_ ;
	wire _w9099_ ;
	wire _w9098_ ;
	wire _w9097_ ;
	wire _w9096_ ;
	wire _w9095_ ;
	wire _w9094_ ;
	wire _w9093_ ;
	wire _w9092_ ;
	wire _w9091_ ;
	wire _w9090_ ;
	wire _w9089_ ;
	wire _w9088_ ;
	wire _w9087_ ;
	wire _w9086_ ;
	wire _w9085_ ;
	wire _w9084_ ;
	wire _w9083_ ;
	wire _w9082_ ;
	wire _w9081_ ;
	wire _w9080_ ;
	wire _w9079_ ;
	wire _w9078_ ;
	wire _w9077_ ;
	wire _w9076_ ;
	wire _w9075_ ;
	wire _w9074_ ;
	wire _w9073_ ;
	wire _w9072_ ;
	wire _w9071_ ;
	wire _w9070_ ;
	wire _w9069_ ;
	wire _w9068_ ;
	wire _w9067_ ;
	wire _w9066_ ;
	wire _w9065_ ;
	wire _w9064_ ;
	wire _w9063_ ;
	wire _w9062_ ;
	wire _w9061_ ;
	wire _w9060_ ;
	wire _w9059_ ;
	wire _w9058_ ;
	wire _w9057_ ;
	wire _w9056_ ;
	wire _w9055_ ;
	wire _w9054_ ;
	wire _w9053_ ;
	wire _w9052_ ;
	wire _w9051_ ;
	wire _w9050_ ;
	wire _w9049_ ;
	wire _w9048_ ;
	wire _w9047_ ;
	wire _w9046_ ;
	wire _w9045_ ;
	wire _w9044_ ;
	wire _w9043_ ;
	wire _w9042_ ;
	wire _w9041_ ;
	wire _w9040_ ;
	wire _w9039_ ;
	wire _w9038_ ;
	wire _w9037_ ;
	wire _w9036_ ;
	wire _w9035_ ;
	wire _w9034_ ;
	wire _w9033_ ;
	wire _w9032_ ;
	wire _w9031_ ;
	wire _w9030_ ;
	wire _w9029_ ;
	wire _w9028_ ;
	wire _w9027_ ;
	wire _w9026_ ;
	wire _w9025_ ;
	wire _w9024_ ;
	wire _w9023_ ;
	wire _w9022_ ;
	wire _w9021_ ;
	wire _w9020_ ;
	wire _w9019_ ;
	wire _w9018_ ;
	wire _w9017_ ;
	wire _w9016_ ;
	wire _w9015_ ;
	wire _w9014_ ;
	wire _w9013_ ;
	wire _w9012_ ;
	wire _w9011_ ;
	wire _w9010_ ;
	wire _w9009_ ;
	wire _w9008_ ;
	wire _w9007_ ;
	wire _w9006_ ;
	wire _w9005_ ;
	wire _w9004_ ;
	wire _w9003_ ;
	wire _w9002_ ;
	wire _w9001_ ;
	wire _w9000_ ;
	wire _w8999_ ;
	wire _w8998_ ;
	wire _w8997_ ;
	wire _w8996_ ;
	wire _w8995_ ;
	wire _w8994_ ;
	wire _w8993_ ;
	wire _w8992_ ;
	wire _w8991_ ;
	wire _w8990_ ;
	wire _w8989_ ;
	wire _w8988_ ;
	wire _w8987_ ;
	wire _w8986_ ;
	wire _w8985_ ;
	wire _w8984_ ;
	wire _w8983_ ;
	wire _w8982_ ;
	wire _w8981_ ;
	wire _w8980_ ;
	wire _w8979_ ;
	wire _w8978_ ;
	wire _w8977_ ;
	wire _w8976_ ;
	wire _w8975_ ;
	wire _w8974_ ;
	wire _w8973_ ;
	wire _w8972_ ;
	wire _w8971_ ;
	wire _w8970_ ;
	wire _w8969_ ;
	wire _w8968_ ;
	wire _w8967_ ;
	wire _w8966_ ;
	wire _w8965_ ;
	wire _w8964_ ;
	wire _w8963_ ;
	wire _w8962_ ;
	wire _w8961_ ;
	wire _w8960_ ;
	wire _w8959_ ;
	wire _w8958_ ;
	wire _w8957_ ;
	wire _w8956_ ;
	wire _w8955_ ;
	wire _w8954_ ;
	wire _w8953_ ;
	wire _w8952_ ;
	wire _w8951_ ;
	wire _w8950_ ;
	wire _w8949_ ;
	wire _w8948_ ;
	wire _w8947_ ;
	wire _w8946_ ;
	wire _w8945_ ;
	wire _w8944_ ;
	wire _w8943_ ;
	wire _w8942_ ;
	wire _w8941_ ;
	wire _w8940_ ;
	wire _w8939_ ;
	wire _w8938_ ;
	wire _w8937_ ;
	wire _w8936_ ;
	wire _w8935_ ;
	wire _w8934_ ;
	wire _w8933_ ;
	wire _w8932_ ;
	wire _w8931_ ;
	wire _w8930_ ;
	wire _w8929_ ;
	wire _w8928_ ;
	wire _w8927_ ;
	wire _w8926_ ;
	wire _w8925_ ;
	wire _w8924_ ;
	wire _w8923_ ;
	wire _w8922_ ;
	wire _w8921_ ;
	wire _w8920_ ;
	wire _w8919_ ;
	wire _w8918_ ;
	wire _w8917_ ;
	wire _w8916_ ;
	wire _w8915_ ;
	wire _w8914_ ;
	wire _w8913_ ;
	wire _w8912_ ;
	wire _w8911_ ;
	wire _w8910_ ;
	wire _w8909_ ;
	wire _w8908_ ;
	wire _w8907_ ;
	wire _w8906_ ;
	wire _w8905_ ;
	wire _w8904_ ;
	wire _w8903_ ;
	wire _w8902_ ;
	wire _w8901_ ;
	wire _w8900_ ;
	wire _w8899_ ;
	wire _w8898_ ;
	wire _w8897_ ;
	wire _w8896_ ;
	wire _w8895_ ;
	wire _w8894_ ;
	wire _w8893_ ;
	wire _w8892_ ;
	wire _w8891_ ;
	wire _w8890_ ;
	wire _w8889_ ;
	wire _w8888_ ;
	wire _w8887_ ;
	wire _w8886_ ;
	wire _w8885_ ;
	wire _w8884_ ;
	wire _w8883_ ;
	wire _w8882_ ;
	wire _w8881_ ;
	wire _w8880_ ;
	wire _w8879_ ;
	wire _w8878_ ;
	wire _w8877_ ;
	wire _w8876_ ;
	wire _w8875_ ;
	wire _w8874_ ;
	wire _w8873_ ;
	wire _w8872_ ;
	wire _w8871_ ;
	wire _w8870_ ;
	wire _w8869_ ;
	wire _w8868_ ;
	wire _w8867_ ;
	wire _w8866_ ;
	wire _w8865_ ;
	wire _w8864_ ;
	wire _w8863_ ;
	wire _w8862_ ;
	wire _w8861_ ;
	wire _w8860_ ;
	wire _w8859_ ;
	wire _w8858_ ;
	wire _w8857_ ;
	wire _w8856_ ;
	wire _w8855_ ;
	wire _w8854_ ;
	wire _w8853_ ;
	wire _w8852_ ;
	wire _w8851_ ;
	wire _w8850_ ;
	wire _w8849_ ;
	wire _w8848_ ;
	wire _w8847_ ;
	wire _w8846_ ;
	wire _w8845_ ;
	wire _w8844_ ;
	wire _w8843_ ;
	wire _w8842_ ;
	wire _w8841_ ;
	wire _w8840_ ;
	wire _w8839_ ;
	wire _w8838_ ;
	wire _w8837_ ;
	wire _w8836_ ;
	wire _w8835_ ;
	wire _w8834_ ;
	wire _w8833_ ;
	wire _w8832_ ;
	wire _w8831_ ;
	wire _w8830_ ;
	wire _w8829_ ;
	wire _w8828_ ;
	wire _w8827_ ;
	wire _w8826_ ;
	wire _w8825_ ;
	wire _w8824_ ;
	wire _w8823_ ;
	wire _w8822_ ;
	wire _w8821_ ;
	wire _w8820_ ;
	wire _w8819_ ;
	wire _w8818_ ;
	wire _w8817_ ;
	wire _w8816_ ;
	wire _w8815_ ;
	wire _w8814_ ;
	wire _w8813_ ;
	wire _w8812_ ;
	wire _w8811_ ;
	wire _w8810_ ;
	wire _w8809_ ;
	wire _w8808_ ;
	wire _w8807_ ;
	wire _w8806_ ;
	wire _w8805_ ;
	wire _w8804_ ;
	wire _w8803_ ;
	wire _w8802_ ;
	wire _w8801_ ;
	wire _w8800_ ;
	wire _w8799_ ;
	wire _w8798_ ;
	wire _w8797_ ;
	wire _w8796_ ;
	wire _w8795_ ;
	wire _w8794_ ;
	wire _w8793_ ;
	wire _w8792_ ;
	wire _w8791_ ;
	wire _w8790_ ;
	wire _w8789_ ;
	wire _w8788_ ;
	wire _w8787_ ;
	wire _w8786_ ;
	wire _w8785_ ;
	wire _w8784_ ;
	wire _w8783_ ;
	wire _w8782_ ;
	wire _w8781_ ;
	wire _w8780_ ;
	wire _w8779_ ;
	wire _w8778_ ;
	wire _w8777_ ;
	wire _w8776_ ;
	wire _w8775_ ;
	wire _w8774_ ;
	wire _w8773_ ;
	wire _w8772_ ;
	wire _w8771_ ;
	wire _w8770_ ;
	wire _w8769_ ;
	wire _w8768_ ;
	wire _w8767_ ;
	wire _w8766_ ;
	wire _w8765_ ;
	wire _w8764_ ;
	wire _w8763_ ;
	wire _w8762_ ;
	wire _w8761_ ;
	wire _w8760_ ;
	wire _w8759_ ;
	wire _w8758_ ;
	wire _w8757_ ;
	wire _w8756_ ;
	wire _w8755_ ;
	wire _w8754_ ;
	wire _w8753_ ;
	wire _w8752_ ;
	wire _w8751_ ;
	wire _w8750_ ;
	wire _w8749_ ;
	wire _w8748_ ;
	wire _w8747_ ;
	wire _w8746_ ;
	wire _w8745_ ;
	wire _w8744_ ;
	wire _w8743_ ;
	wire _w8742_ ;
	wire _w8741_ ;
	wire _w8740_ ;
	wire _w8739_ ;
	wire _w8738_ ;
	wire _w8737_ ;
	wire _w8736_ ;
	wire _w8735_ ;
	wire _w8734_ ;
	wire _w8733_ ;
	wire _w8732_ ;
	wire _w8731_ ;
	wire _w8730_ ;
	wire _w8729_ ;
	wire _w8728_ ;
	wire _w8727_ ;
	wire _w8726_ ;
	wire _w8725_ ;
	wire _w8724_ ;
	wire _w8723_ ;
	wire _w8722_ ;
	wire _w8721_ ;
	wire _w8720_ ;
	wire _w8719_ ;
	wire _w8718_ ;
	wire _w8717_ ;
	wire _w8716_ ;
	wire _w8715_ ;
	wire _w8714_ ;
	wire _w8713_ ;
	wire _w8712_ ;
	wire _w8711_ ;
	wire _w8710_ ;
	wire _w8709_ ;
	wire _w8708_ ;
	wire _w8707_ ;
	wire _w8706_ ;
	wire _w8705_ ;
	wire _w8704_ ;
	wire _w8703_ ;
	wire _w8702_ ;
	wire _w8701_ ;
	wire _w8700_ ;
	wire _w8699_ ;
	wire _w8698_ ;
	wire _w8697_ ;
	wire _w8696_ ;
	wire _w8695_ ;
	wire _w8694_ ;
	wire _w8693_ ;
	wire _w8692_ ;
	wire _w8691_ ;
	wire _w8690_ ;
	wire _w8689_ ;
	wire _w8688_ ;
	wire _w8687_ ;
	wire _w8686_ ;
	wire _w8685_ ;
	wire _w8684_ ;
	wire _w8683_ ;
	wire _w8682_ ;
	wire _w8681_ ;
	wire _w8680_ ;
	wire _w8679_ ;
	wire _w8678_ ;
	wire _w8677_ ;
	wire _w8676_ ;
	wire _w8675_ ;
	wire _w8674_ ;
	wire _w8673_ ;
	wire _w8672_ ;
	wire _w8671_ ;
	wire _w8670_ ;
	wire _w8669_ ;
	wire _w8668_ ;
	wire _w8667_ ;
	wire _w8666_ ;
	wire _w8665_ ;
	wire _w8664_ ;
	wire _w8663_ ;
	wire _w8662_ ;
	wire _w8661_ ;
	wire _w8660_ ;
	wire _w8659_ ;
	wire _w8658_ ;
	wire _w8657_ ;
	wire _w8656_ ;
	wire _w8655_ ;
	wire _w8654_ ;
	wire _w8653_ ;
	wire _w8652_ ;
	wire _w8651_ ;
	wire _w8650_ ;
	wire _w8649_ ;
	wire _w8648_ ;
	wire _w8647_ ;
	wire _w8646_ ;
	wire _w8645_ ;
	wire _w8644_ ;
	wire _w8643_ ;
	wire _w8642_ ;
	wire _w8641_ ;
	wire _w8640_ ;
	wire _w8639_ ;
	wire _w8638_ ;
	wire _w8637_ ;
	wire _w8636_ ;
	wire _w8635_ ;
	wire _w8634_ ;
	wire _w8633_ ;
	wire _w8632_ ;
	wire _w8631_ ;
	wire _w8630_ ;
	wire _w8629_ ;
	wire _w8628_ ;
	wire _w8627_ ;
	wire _w8626_ ;
	wire _w8625_ ;
	wire _w8624_ ;
	wire _w8623_ ;
	wire _w8622_ ;
	wire _w8621_ ;
	wire _w8620_ ;
	wire _w8619_ ;
	wire _w8618_ ;
	wire _w8617_ ;
	wire _w8616_ ;
	wire _w8615_ ;
	wire _w8614_ ;
	wire _w8613_ ;
	wire _w8612_ ;
	wire _w8611_ ;
	wire _w8610_ ;
	wire _w8609_ ;
	wire _w8608_ ;
	wire _w8607_ ;
	wire _w8606_ ;
	wire _w8605_ ;
	wire _w8604_ ;
	wire _w8603_ ;
	wire _w8602_ ;
	wire _w8601_ ;
	wire _w8600_ ;
	wire _w8599_ ;
	wire _w8598_ ;
	wire _w8597_ ;
	wire _w8596_ ;
	wire _w8595_ ;
	wire _w8594_ ;
	wire _w8593_ ;
	wire _w8592_ ;
	wire _w8591_ ;
	wire _w8590_ ;
	wire _w8589_ ;
	wire _w8588_ ;
	wire _w8587_ ;
	wire _w8586_ ;
	wire _w8585_ ;
	wire _w8584_ ;
	wire _w8583_ ;
	wire _w8582_ ;
	wire _w8581_ ;
	wire _w8580_ ;
	wire _w8579_ ;
	wire _w8578_ ;
	wire _w8577_ ;
	wire _w8576_ ;
	wire _w8575_ ;
	wire _w8574_ ;
	wire _w8573_ ;
	wire _w8572_ ;
	wire _w8571_ ;
	wire _w8570_ ;
	wire _w8569_ ;
	wire _w8568_ ;
	wire _w8567_ ;
	wire _w8566_ ;
	wire _w8565_ ;
	wire _w8564_ ;
	wire _w8563_ ;
	wire _w8562_ ;
	wire _w8561_ ;
	wire _w8560_ ;
	wire _w8559_ ;
	wire _w8558_ ;
	wire _w8557_ ;
	wire _w8556_ ;
	wire _w8555_ ;
	wire _w8554_ ;
	wire _w8553_ ;
	wire _w8552_ ;
	wire _w8551_ ;
	wire _w8550_ ;
	wire _w8549_ ;
	wire _w8548_ ;
	wire _w8547_ ;
	wire _w8546_ ;
	wire _w8545_ ;
	wire _w8544_ ;
	wire _w8543_ ;
	wire _w8542_ ;
	wire _w8541_ ;
	wire _w8540_ ;
	wire _w8539_ ;
	wire _w8538_ ;
	wire _w8537_ ;
	wire _w8536_ ;
	wire _w8535_ ;
	wire _w8534_ ;
	wire _w8533_ ;
	wire _w8532_ ;
	wire _w8531_ ;
	wire _w8530_ ;
	wire _w8529_ ;
	wire _w8528_ ;
	wire _w8527_ ;
	wire _w8526_ ;
	wire _w8525_ ;
	wire _w8524_ ;
	wire _w8523_ ;
	wire _w8522_ ;
	wire _w8521_ ;
	wire _w8520_ ;
	wire _w8519_ ;
	wire _w8518_ ;
	wire _w8517_ ;
	wire _w8516_ ;
	wire _w8515_ ;
	wire _w8514_ ;
	wire _w8513_ ;
	wire _w8512_ ;
	wire _w8511_ ;
	wire _w8510_ ;
	wire _w8509_ ;
	wire _w8508_ ;
	wire _w8507_ ;
	wire _w8506_ ;
	wire _w8505_ ;
	wire _w8504_ ;
	wire _w8503_ ;
	wire _w8502_ ;
	wire _w8501_ ;
	wire _w8500_ ;
	wire _w8499_ ;
	wire _w8498_ ;
	wire _w8497_ ;
	wire _w8496_ ;
	wire _w8495_ ;
	wire _w8494_ ;
	wire _w8493_ ;
	wire _w8492_ ;
	wire _w8491_ ;
	wire _w8490_ ;
	wire _w8489_ ;
	wire _w8488_ ;
	wire _w8487_ ;
	wire _w8486_ ;
	wire _w8485_ ;
	wire _w8484_ ;
	wire _w8483_ ;
	wire _w8482_ ;
	wire _w8481_ ;
	wire _w8480_ ;
	wire _w8479_ ;
	wire _w8478_ ;
	wire _w8477_ ;
	wire _w8476_ ;
	wire _w8475_ ;
	wire _w8474_ ;
	wire _w8473_ ;
	wire _w8472_ ;
	wire _w8471_ ;
	wire _w8470_ ;
	wire _w8469_ ;
	wire _w8468_ ;
	wire _w8467_ ;
	wire _w8466_ ;
	wire _w8465_ ;
	wire _w8464_ ;
	wire _w8463_ ;
	wire _w8462_ ;
	wire _w8461_ ;
	wire _w8460_ ;
	wire _w8459_ ;
	wire _w8458_ ;
	wire _w8457_ ;
	wire _w8456_ ;
	wire _w8455_ ;
	wire _w8454_ ;
	wire _w8453_ ;
	wire _w8452_ ;
	wire _w8451_ ;
	wire _w8450_ ;
	wire _w8449_ ;
	wire _w8448_ ;
	wire _w8447_ ;
	wire _w8446_ ;
	wire _w8445_ ;
	wire _w8444_ ;
	wire _w8443_ ;
	wire _w8442_ ;
	wire _w8441_ ;
	wire _w8440_ ;
	wire _w8439_ ;
	wire _w8438_ ;
	wire _w8437_ ;
	wire _w8436_ ;
	wire _w8435_ ;
	wire _w8434_ ;
	wire _w8433_ ;
	wire _w8432_ ;
	wire _w8431_ ;
	wire _w8430_ ;
	wire _w8429_ ;
	wire _w8428_ ;
	wire _w8427_ ;
	wire _w8426_ ;
	wire _w8425_ ;
	wire _w8424_ ;
	wire _w8423_ ;
	wire _w8422_ ;
	wire _w8421_ ;
	wire _w8420_ ;
	wire _w8419_ ;
	wire _w8418_ ;
	wire _w8417_ ;
	wire _w8416_ ;
	wire _w8415_ ;
	wire _w8414_ ;
	wire _w8413_ ;
	wire _w8412_ ;
	wire _w8411_ ;
	wire _w8410_ ;
	wire _w8409_ ;
	wire _w8408_ ;
	wire _w8407_ ;
	wire _w8406_ ;
	wire _w8405_ ;
	wire _w8404_ ;
	wire _w8403_ ;
	wire _w8402_ ;
	wire _w8401_ ;
	wire _w8400_ ;
	wire _w8399_ ;
	wire _w8398_ ;
	wire _w8397_ ;
	wire _w8396_ ;
	wire _w8395_ ;
	wire _w8394_ ;
	wire _w8393_ ;
	wire _w8392_ ;
	wire _w8391_ ;
	wire _w8390_ ;
	wire _w8389_ ;
	wire _w8388_ ;
	wire _w8387_ ;
	wire _w8386_ ;
	wire _w8385_ ;
	wire _w8384_ ;
	wire _w8383_ ;
	wire _w8382_ ;
	wire _w8381_ ;
	wire _w8380_ ;
	wire _w8379_ ;
	wire _w8378_ ;
	wire _w8377_ ;
	wire _w8376_ ;
	wire _w8375_ ;
	wire _w8374_ ;
	wire _w8373_ ;
	wire _w8372_ ;
	wire _w8371_ ;
	wire _w8370_ ;
	wire _w8369_ ;
	wire _w8368_ ;
	wire _w8367_ ;
	wire _w8366_ ;
	wire _w8365_ ;
	wire _w8364_ ;
	wire _w8363_ ;
	wire _w8362_ ;
	wire _w8361_ ;
	wire _w8360_ ;
	wire _w8359_ ;
	wire _w8358_ ;
	wire _w8357_ ;
	wire _w8356_ ;
	wire _w8355_ ;
	wire _w8354_ ;
	wire _w8353_ ;
	wire _w8352_ ;
	wire _w8351_ ;
	wire _w8350_ ;
	wire _w8349_ ;
	wire _w8348_ ;
	wire _w8347_ ;
	wire _w8346_ ;
	wire _w8345_ ;
	wire _w8344_ ;
	wire _w8343_ ;
	wire _w8342_ ;
	wire _w8341_ ;
	wire _w8340_ ;
	wire _w8339_ ;
	wire _w8338_ ;
	wire _w8337_ ;
	wire _w8336_ ;
	wire _w8335_ ;
	wire _w8334_ ;
	wire _w8333_ ;
	wire _w8332_ ;
	wire _w8331_ ;
	wire _w8330_ ;
	wire _w8329_ ;
	wire _w8328_ ;
	wire _w8327_ ;
	wire _w8326_ ;
	wire _w8325_ ;
	wire _w8324_ ;
	wire _w8323_ ;
	wire _w8322_ ;
	wire _w8321_ ;
	wire _w8320_ ;
	wire _w8319_ ;
	wire _w8318_ ;
	wire _w8317_ ;
	wire _w8316_ ;
	wire _w8315_ ;
	wire _w8314_ ;
	wire _w8313_ ;
	wire _w8312_ ;
	wire _w8311_ ;
	wire _w8310_ ;
	wire _w8309_ ;
	wire _w8308_ ;
	wire _w8307_ ;
	wire _w8306_ ;
	wire _w8305_ ;
	wire _w8304_ ;
	wire _w8303_ ;
	wire _w8302_ ;
	wire _w8301_ ;
	wire _w8300_ ;
	wire _w8299_ ;
	wire _w8298_ ;
	wire _w8297_ ;
	wire _w8296_ ;
	wire _w8295_ ;
	wire _w8294_ ;
	wire _w8293_ ;
	wire _w8292_ ;
	wire _w8291_ ;
	wire _w8290_ ;
	wire _w8289_ ;
	wire _w8288_ ;
	wire _w8287_ ;
	wire _w8286_ ;
	wire _w8285_ ;
	wire _w8284_ ;
	wire _w8283_ ;
	wire _w8282_ ;
	wire _w8281_ ;
	wire _w8280_ ;
	wire _w8279_ ;
	wire _w8278_ ;
	wire _w8277_ ;
	wire _w8276_ ;
	wire _w8275_ ;
	wire _w8274_ ;
	wire _w8273_ ;
	wire _w8272_ ;
	wire _w8271_ ;
	wire _w8270_ ;
	wire _w8269_ ;
	wire _w8268_ ;
	wire _w8267_ ;
	wire _w8266_ ;
	wire _w8265_ ;
	wire _w8264_ ;
	wire _w8263_ ;
	wire _w8262_ ;
	wire _w8261_ ;
	wire _w8260_ ;
	wire _w8259_ ;
	wire _w8258_ ;
	wire _w8257_ ;
	wire _w8256_ ;
	wire _w8255_ ;
	wire _w8254_ ;
	wire _w8253_ ;
	wire _w8252_ ;
	wire _w8251_ ;
	wire _w8250_ ;
	wire _w8249_ ;
	wire _w8248_ ;
	wire _w8247_ ;
	wire _w8246_ ;
	wire _w8245_ ;
	wire _w8244_ ;
	wire _w8243_ ;
	wire _w8242_ ;
	wire _w8241_ ;
	wire _w8240_ ;
	wire _w8239_ ;
	wire _w8238_ ;
	wire _w8237_ ;
	wire _w8236_ ;
	wire _w8235_ ;
	wire _w8234_ ;
	wire _w8233_ ;
	wire _w8232_ ;
	wire _w8231_ ;
	wire _w8230_ ;
	wire _w8229_ ;
	wire _w8228_ ;
	wire _w8227_ ;
	wire _w8226_ ;
	wire _w8225_ ;
	wire _w8224_ ;
	wire _w8223_ ;
	wire _w8222_ ;
	wire _w8221_ ;
	wire _w8220_ ;
	wire _w8219_ ;
	wire _w8218_ ;
	wire _w8217_ ;
	wire _w8216_ ;
	wire _w8215_ ;
	wire _w8214_ ;
	wire _w8213_ ;
	wire _w8212_ ;
	wire _w8211_ ;
	wire _w8210_ ;
	wire _w8209_ ;
	wire _w8208_ ;
	wire _w8207_ ;
	wire _w8206_ ;
	wire _w8205_ ;
	wire _w8204_ ;
	wire _w8203_ ;
	wire _w8202_ ;
	wire _w8201_ ;
	wire _w8200_ ;
	wire _w8199_ ;
	wire _w8198_ ;
	wire _w8197_ ;
	wire _w8196_ ;
	wire _w8195_ ;
	wire _w8194_ ;
	wire _w8193_ ;
	wire _w8192_ ;
	wire _w8191_ ;
	wire _w8190_ ;
	wire _w8189_ ;
	wire _w8188_ ;
	wire _w8187_ ;
	wire _w8186_ ;
	wire _w8185_ ;
	wire _w8184_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4995_ ;
	wire _w4993_ ;
	wire _w4991_ ;
	wire _w4989_ ;
	wire _w4987_ ;
	wire _w4985_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4099_ ;
	wire _w4097_ ;
	wire _w4095_ ;
	wire _w4093_ ;
	wire _w4091_ ;
	wire _w4089_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4059_ ;
	wire _w4090_ ;
	wire _w4244_ ;
	wire _w5082_ ;
	wire _w5360_ ;
	wire _w4433_ ;
	wire _w4075_ ;
	wire _w4068_ ;
	wire _w4100_ ;
	wire _w4116_ ;
	wire _w4069_ ;
	wire _w4098_ ;
	wire _w4114_ ;
	wire _w4067_ ;
	wire _w4096_ ;
	wire _w4112_ ;
	wire _w4065_ ;
	wire _w4094_ ;
	wire _w4236_ ;
	wire _w4574_ ;
	wire _w4110_ ;
	wire _w4063_ ;
	wire _w4087_ ;
	wire _w4221_ ;
	wire _w4383_ ;
	wire _w4066_ ;
	wire _w4092_ ;
	wire _w4108_ ;
	wire _w4061_ ;
	wire _w8038_ ;
	wire _w2951_ ;
	wire _w13224_ ;
	wire _w5308_ ;
	wire _w4060_ ;
	wire _w4132_ ;
	wire _w4088_ ;
	wire _w4062_ ;
	wire _w4064_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4076_ ;
	wire _w4107_ ;
	wire _w4109_ ;
	wire _w4111_ ;
	wire _w4113_ ;
	wire _w4115_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4984_ ;
	wire _w5262_ ;
	wire _w4335_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4986_ ;
	wire _w5264_ ;
	wire _w4337_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4988_ ;
	wire _w5266_ ;
	wire _w4339_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4990_ ;
	wire _w5268_ ;
	wire _w4341_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4992_ ;
	wire _w5270_ ;
	wire _w4343_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4994_ ;
	wire _w5272_ ;
	wire _w4345_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4996_ ;
	wire _w5274_ ;
	wire _w4347_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w5012_ ;
	wire _w5290_ ;
	wire _w4363_ ;
	wire _w4174_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4336_ ;
	wire _w4338_ ;
	wire _w4340_ ;
	wire _w4342_ ;
	wire _w4344_ ;
	wire _w4346_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w5851_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5263_ ;
	wire _w5265_ ;
	wire _w5267_ ;
	wire _w5269_ ;
	wire _w5271_ ;
	wire _w5273_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w21301_ ;
	wire _w548_ ;
	wire _w10821_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w21303_ ;
	wire _w550_ ;
	wire _w10823_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w21305_ ;
	wire _w552_ ;
	wire _w10825_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w21307_ ;
	wire _w554_ ;
	wire _w10827_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w21309_ ;
	wire _w556_ ;
	wire _w10829_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w21311_ ;
	wire _w558_ ;
	wire _w10831_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w21313_ ;
	wire _w560_ ;
	wire _w10833_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w21329_ ;
	wire _w576_ ;
	wire _w10849_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w21399_ ;
	wire _w646_ ;
	wire _w10919_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w21890_ ;
	wire _w1137_ ;
	wire _w11410_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w9135_ ;
	wire _w9136_ ;
	wire _w9137_ ;
	wire _w9138_ ;
	wire _w9139_ ;
	wire _w9140_ ;
	wire _w9141_ ;
	wire _w9142_ ;
	wire _w9143_ ;
	wire _w9144_ ;
	wire _w9145_ ;
	wire _w9146_ ;
	wire _w9147_ ;
	wire _w9148_ ;
	wire _w9149_ ;
	wire _w9150_ ;
	wire _w9151_ ;
	wire _w9152_ ;
	wire _w9153_ ;
	wire _w9154_ ;
	wire _w9155_ ;
	wire _w9156_ ;
	wire _w9157_ ;
	wire _w9158_ ;
	wire _w9159_ ;
	wire _w9160_ ;
	wire _w9161_ ;
	wire _w9162_ ;
	wire _w9163_ ;
	wire _w9164_ ;
	wire _w9165_ ;
	wire _w9166_ ;
	wire _w9167_ ;
	wire _w9168_ ;
	wire _w9169_ ;
	wire _w9170_ ;
	wire _w9171_ ;
	wire _w9172_ ;
	wire _w9173_ ;
	wire _w9174_ ;
	wire _w9175_ ;
	wire _w9176_ ;
	wire _w9177_ ;
	wire _w9178_ ;
	wire _w9179_ ;
	wire _w9180_ ;
	wire _w9181_ ;
	wire _w9182_ ;
	wire _w9183_ ;
	wire _w9184_ ;
	wire _w9185_ ;
	wire _w9186_ ;
	wire _w9187_ ;
	wire _w9188_ ;
	wire _w9189_ ;
	wire _w9190_ ;
	wire _w9191_ ;
	wire _w9192_ ;
	wire _w9193_ ;
	wire _w9194_ ;
	wire _w9195_ ;
	wire _w9196_ ;
	wire _w9197_ ;
	wire _w9198_ ;
	wire _w9199_ ;
	wire _w9200_ ;
	wire _w9201_ ;
	wire _w9202_ ;
	wire _w9203_ ;
	wire _w9204_ ;
	wire _w9205_ ;
	wire _w9206_ ;
	wire _w9207_ ;
	wire _w9208_ ;
	wire _w9209_ ;
	wire _w9210_ ;
	wire _w9211_ ;
	wire _w9212_ ;
	wire _w9213_ ;
	wire _w9214_ ;
	wire _w9215_ ;
	wire _w9216_ ;
	wire _w9217_ ;
	wire _w9218_ ;
	wire _w9219_ ;
	wire _w9220_ ;
	wire _w9221_ ;
	wire _w9222_ ;
	wire _w9223_ ;
	wire _w9224_ ;
	wire _w9225_ ;
	wire _w9226_ ;
	wire _w9227_ ;
	wire _w9228_ ;
	wire _w9229_ ;
	wire _w9230_ ;
	wire _w9231_ ;
	wire _w9232_ ;
	wire _w9233_ ;
	wire _w9234_ ;
	wire _w9235_ ;
	wire _w9236_ ;
	wire _w9237_ ;
	wire _w9238_ ;
	wire _w9239_ ;
	wire _w9240_ ;
	wire _w9241_ ;
	wire _w9242_ ;
	wire _w9243_ ;
	wire _w9244_ ;
	wire _w9245_ ;
	wire _w9246_ ;
	wire _w9247_ ;
	wire _w9248_ ;
	wire _w9249_ ;
	wire _w9250_ ;
	wire _w9251_ ;
	wire _w9252_ ;
	wire _w9253_ ;
	wire _w9254_ ;
	wire _w9255_ ;
	wire _w9256_ ;
	wire _w9257_ ;
	wire _w9258_ ;
	wire _w9259_ ;
	wire _w9260_ ;
	wire _w9261_ ;
	wire _w9262_ ;
	wire _w9263_ ;
	wire _w9264_ ;
	wire _w9265_ ;
	wire _w9266_ ;
	wire _w9267_ ;
	wire _w9268_ ;
	wire _w9269_ ;
	wire _w9270_ ;
	wire _w9271_ ;
	wire _w9272_ ;
	wire _w9273_ ;
	wire _w9274_ ;
	wire _w9275_ ;
	wire _w9276_ ;
	wire _w9277_ ;
	wire _w9278_ ;
	wire _w9279_ ;
	wire _w9280_ ;
	wire _w9281_ ;
	wire _w9282_ ;
	wire _w9283_ ;
	wire _w9284_ ;
	wire _w9285_ ;
	wire _w9286_ ;
	wire _w9287_ ;
	wire _w9288_ ;
	wire _w9289_ ;
	wire _w9290_ ;
	wire _w9291_ ;
	wire _w9292_ ;
	wire _w9293_ ;
	wire _w9294_ ;
	wire _w9295_ ;
	wire _w9296_ ;
	wire _w9297_ ;
	wire _w9298_ ;
	wire _w9299_ ;
	wire _w9300_ ;
	wire _w9301_ ;
	wire _w9302_ ;
	wire _w9303_ ;
	wire _w9304_ ;
	wire _w9305_ ;
	wire _w9306_ ;
	wire _w9307_ ;
	wire _w9308_ ;
	wire _w9309_ ;
	wire _w9310_ ;
	wire _w9311_ ;
	wire _w9312_ ;
	wire _w9313_ ;
	wire _w9314_ ;
	wire _w9315_ ;
	wire _w9316_ ;
	wire _w9317_ ;
	wire _w9318_ ;
	wire _w9319_ ;
	wire _w9320_ ;
	wire _w9321_ ;
	wire _w9322_ ;
	wire _w9323_ ;
	wire _w9324_ ;
	wire _w9325_ ;
	wire _w9326_ ;
	wire _w9327_ ;
	wire _w9328_ ;
	wire _w9329_ ;
	wire _w9330_ ;
	wire _w9331_ ;
	wire _w9332_ ;
	wire _w9333_ ;
	wire _w9334_ ;
	wire _w9335_ ;
	wire _w9336_ ;
	wire _w9337_ ;
	wire _w9338_ ;
	wire _w9339_ ;
	wire _w9340_ ;
	wire _w9341_ ;
	wire _w9342_ ;
	wire _w9343_ ;
	wire _w9344_ ;
	wire _w9345_ ;
	wire _w9346_ ;
	wire _w9347_ ;
	wire _w9348_ ;
	wire _w9349_ ;
	wire _w9350_ ;
	wire _w9351_ ;
	wire _w9352_ ;
	wire _w9353_ ;
	wire _w9354_ ;
	wire _w9355_ ;
	wire _w9356_ ;
	wire _w9357_ ;
	wire _w9358_ ;
	wire _w9359_ ;
	wire _w9360_ ;
	wire _w9361_ ;
	wire _w9362_ ;
	wire _w9363_ ;
	wire _w9364_ ;
	wire _w9365_ ;
	wire _w9366_ ;
	wire _w9367_ ;
	wire _w9368_ ;
	wire _w9369_ ;
	wire _w9370_ ;
	wire _w9371_ ;
	wire _w9372_ ;
	wire _w9373_ ;
	wire _w9374_ ;
	wire _w9375_ ;
	wire _w9376_ ;
	wire _w9377_ ;
	wire _w9378_ ;
	wire _w9379_ ;
	wire _w9380_ ;
	wire _w9381_ ;
	wire _w9382_ ;
	wire _w9383_ ;
	wire _w9384_ ;
	wire _w9385_ ;
	wire _w9386_ ;
	wire _w9387_ ;
	wire _w9388_ ;
	wire _w9389_ ;
	wire _w9390_ ;
	wire _w9391_ ;
	wire _w9392_ ;
	wire _w9393_ ;
	wire _w9394_ ;
	wire _w9395_ ;
	wire _w9396_ ;
	wire _w9397_ ;
	wire _w9398_ ;
	wire _w9399_ ;
	wire _w9400_ ;
	wire _w9401_ ;
	wire _w9402_ ;
	wire _w9403_ ;
	wire _w9404_ ;
	wire _w9405_ ;
	wire _w9406_ ;
	wire _w9407_ ;
	wire _w9408_ ;
	wire _w9409_ ;
	wire _w9410_ ;
	wire _w9411_ ;
	wire _w9412_ ;
	wire _w9413_ ;
	wire _w9414_ ;
	wire _w9415_ ;
	wire _w9416_ ;
	wire _w9417_ ;
	wire _w9418_ ;
	wire _w9419_ ;
	wire _w9420_ ;
	wire _w9421_ ;
	wire _w9422_ ;
	wire _w9423_ ;
	wire _w9424_ ;
	wire _w9425_ ;
	wire _w9426_ ;
	wire _w9427_ ;
	wire _w9428_ ;
	wire _w9429_ ;
	wire _w9430_ ;
	wire _w9431_ ;
	wire _w9432_ ;
	wire _w9433_ ;
	wire _w9434_ ;
	wire _w9435_ ;
	wire _w9436_ ;
	wire _w9437_ ;
	wire _w9438_ ;
	wire _w9439_ ;
	wire _w9440_ ;
	wire _w9441_ ;
	wire _w9442_ ;
	wire _w9443_ ;
	wire _w9444_ ;
	wire _w9445_ ;
	wire _w9446_ ;
	wire _w9447_ ;
	wire _w9448_ ;
	wire _w9449_ ;
	wire _w9450_ ;
	wire _w9451_ ;
	wire _w9452_ ;
	wire _w9453_ ;
	wire _w9454_ ;
	wire _w9455_ ;
	wire _w9456_ ;
	wire _w9457_ ;
	wire _w9458_ ;
	wire _w9459_ ;
	wire _w9460_ ;
	wire _w9461_ ;
	wire _w9462_ ;
	wire _w9463_ ;
	wire _w9464_ ;
	wire _w9465_ ;
	wire _w9466_ ;
	wire _w9467_ ;
	wire _w9468_ ;
	wire _w9469_ ;
	wire _w9470_ ;
	wire _w9471_ ;
	wire _w9472_ ;
	wire _w9473_ ;
	wire _w9474_ ;
	wire _w9475_ ;
	wire _w9476_ ;
	wire _w9477_ ;
	wire _w9478_ ;
	wire _w9479_ ;
	wire _w9480_ ;
	wire _w9481_ ;
	wire _w9482_ ;
	wire _w9483_ ;
	wire _w9484_ ;
	wire _w9485_ ;
	wire _w9486_ ;
	wire _w9487_ ;
	wire _w9488_ ;
	wire _w9489_ ;
	wire _w9490_ ;
	wire _w9491_ ;
	wire _w9492_ ;
	wire _w9493_ ;
	wire _w9494_ ;
	wire _w9495_ ;
	wire _w9496_ ;
	wire _w9497_ ;
	wire _w9498_ ;
	wire _w9499_ ;
	wire _w9500_ ;
	wire _w9501_ ;
	wire _w9502_ ;
	wire _w9503_ ;
	wire _w9504_ ;
	wire _w9505_ ;
	wire _w9506_ ;
	wire _w9507_ ;
	wire _w9508_ ;
	wire _w9509_ ;
	wire _w9510_ ;
	wire _w9511_ ;
	wire _w9512_ ;
	wire _w9513_ ;
	wire _w9514_ ;
	wire _w9515_ ;
	wire _w9516_ ;
	wire _w9517_ ;
	wire _w9518_ ;
	wire _w9519_ ;
	wire _w9520_ ;
	wire _w9521_ ;
	wire _w9522_ ;
	wire _w9523_ ;
	wire _w9524_ ;
	wire _w9525_ ;
	wire _w9526_ ;
	wire _w9527_ ;
	wire _w9528_ ;
	wire _w9529_ ;
	wire _w9530_ ;
	wire _w9531_ ;
	wire _w9532_ ;
	wire _w9533_ ;
	wire _w9534_ ;
	wire _w9535_ ;
	wire _w9536_ ;
	wire _w9537_ ;
	wire _w9538_ ;
	wire _w9539_ ;
	wire _w9540_ ;
	wire _w9541_ ;
	wire _w9542_ ;
	wire _w9543_ ;
	wire _w9544_ ;
	wire _w9545_ ;
	wire _w9546_ ;
	wire _w9547_ ;
	wire _w9548_ ;
	wire _w9549_ ;
	wire _w9550_ ;
	wire _w9551_ ;
	wire _w9552_ ;
	wire _w9553_ ;
	wire _w9554_ ;
	wire _w9555_ ;
	wire _w9556_ ;
	wire _w9557_ ;
	wire _w9558_ ;
	wire _w9559_ ;
	wire _w9560_ ;
	wire _w9561_ ;
	wire _w9562_ ;
	wire _w9563_ ;
	wire _w9564_ ;
	wire _w9565_ ;
	wire _w9566_ ;
	wire _w9567_ ;
	wire _w9568_ ;
	wire _w9569_ ;
	wire _w9570_ ;
	wire _w9571_ ;
	wire _w9572_ ;
	wire _w9573_ ;
	wire _w9574_ ;
	wire _w9575_ ;
	wire _w9576_ ;
	wire _w9577_ ;
	wire _w9578_ ;
	wire _w9579_ ;
	wire _w9580_ ;
	wire _w9581_ ;
	wire _w9582_ ;
	wire _w9583_ ;
	wire _w9584_ ;
	wire _w9585_ ;
	wire _w9586_ ;
	wire _w9587_ ;
	wire _w9588_ ;
	wire _w9589_ ;
	wire _w9590_ ;
	wire _w9591_ ;
	wire _w9592_ ;
	wire _w9593_ ;
	wire _w9594_ ;
	wire _w9595_ ;
	wire _w9596_ ;
	wire _w9597_ ;
	wire _w9598_ ;
	wire _w9599_ ;
	wire _w9600_ ;
	wire _w9601_ ;
	wire _w9602_ ;
	wire _w9603_ ;
	wire _w9604_ ;
	wire _w9605_ ;
	wire _w9606_ ;
	wire _w9607_ ;
	wire _w9608_ ;
	wire _w9609_ ;
	wire _w9610_ ;
	wire _w9611_ ;
	wire _w9612_ ;
	wire _w9613_ ;
	wire _w9614_ ;
	wire _w9615_ ;
	wire _w9616_ ;
	wire _w9617_ ;
	wire _w9618_ ;
	wire _w9619_ ;
	wire _w9620_ ;
	wire _w9621_ ;
	wire _w9622_ ;
	wire _w9623_ ;
	wire _w9624_ ;
	wire _w9625_ ;
	wire _w9626_ ;
	wire _w9627_ ;
	wire _w9628_ ;
	wire _w9629_ ;
	wire _w9630_ ;
	wire _w9631_ ;
	wire _w9632_ ;
	wire _w9633_ ;
	wire _w9634_ ;
	wire _w9635_ ;
	wire _w9636_ ;
	wire _w9637_ ;
	wire _w9638_ ;
	wire _w9639_ ;
	wire _w9640_ ;
	wire _w9641_ ;
	wire _w9642_ ;
	wire _w9643_ ;
	wire _w9644_ ;
	wire _w9645_ ;
	wire _w9646_ ;
	wire _w9647_ ;
	wire _w9648_ ;
	wire _w9649_ ;
	wire _w9650_ ;
	wire _w9651_ ;
	wire _w9652_ ;
	wire _w9653_ ;
	wire _w9654_ ;
	wire _w9655_ ;
	wire _w9656_ ;
	wire _w9657_ ;
	wire _w9658_ ;
	wire _w9659_ ;
	wire _w9660_ ;
	wire _w9661_ ;
	wire _w9662_ ;
	wire _w9663_ ;
	wire _w9664_ ;
	wire _w9665_ ;
	wire _w9666_ ;
	wire _w9667_ ;
	wire _w9668_ ;
	wire _w9669_ ;
	wire _w9670_ ;
	wire _w9671_ ;
	wire _w9672_ ;
	wire _w9673_ ;
	wire _w9674_ ;
	wire _w9675_ ;
	wire _w9676_ ;
	wire _w9677_ ;
	wire _w9678_ ;
	wire _w9679_ ;
	wire _w9680_ ;
	wire _w9681_ ;
	wire _w9682_ ;
	wire _w9683_ ;
	wire _w9684_ ;
	wire _w9685_ ;
	wire _w9686_ ;
	wire _w9687_ ;
	wire _w9688_ ;
	wire _w9689_ ;
	wire _w9690_ ;
	wire _w9691_ ;
	wire _w9692_ ;
	wire _w9693_ ;
	wire _w9694_ ;
	wire _w9695_ ;
	wire _w9696_ ;
	wire _w9697_ ;
	wire _w9698_ ;
	wire _w9699_ ;
	wire _w9700_ ;
	wire _w9701_ ;
	wire _w9702_ ;
	wire _w9703_ ;
	wire _w9704_ ;
	wire _w9705_ ;
	wire _w9706_ ;
	wire _w9707_ ;
	wire _w9708_ ;
	wire _w9709_ ;
	wire _w9710_ ;
	wire _w9711_ ;
	wire _w9712_ ;
	wire _w9713_ ;
	wire _w9714_ ;
	wire _w9715_ ;
	wire _w9716_ ;
	wire _w9717_ ;
	wire _w9718_ ;
	wire _w9719_ ;
	wire _w9720_ ;
	wire _w9721_ ;
	wire _w9722_ ;
	wire _w9723_ ;
	wire _w9724_ ;
	wire _w9725_ ;
	wire _w9726_ ;
	wire _w9727_ ;
	wire _w9728_ ;
	wire _w9729_ ;
	wire _w9730_ ;
	wire _w9731_ ;
	wire _w9732_ ;
	wire _w9733_ ;
	wire _w9734_ ;
	wire _w9735_ ;
	wire _w9736_ ;
	wire _w9737_ ;
	wire _w9738_ ;
	wire _w9739_ ;
	wire _w9740_ ;
	wire _w9741_ ;
	wire _w9742_ ;
	wire _w9743_ ;
	wire _w9744_ ;
	wire _w9745_ ;
	wire _w9746_ ;
	wire _w9747_ ;
	wire _w9748_ ;
	wire _w9749_ ;
	wire _w9750_ ;
	wire _w9751_ ;
	wire _w9752_ ;
	wire _w9753_ ;
	wire _w9754_ ;
	wire _w9755_ ;
	wire _w9756_ ;
	wire _w9757_ ;
	wire _w9758_ ;
	wire _w9759_ ;
	wire _w9760_ ;
	wire _w9761_ ;
	wire _w9762_ ;
	wire _w9763_ ;
	wire _w9764_ ;
	wire _w9765_ ;
	wire _w9766_ ;
	wire _w9767_ ;
	wire _w9768_ ;
	wire _w9769_ ;
	wire _w9770_ ;
	wire _w9771_ ;
	wire _w9772_ ;
	wire _w9773_ ;
	wire _w9774_ ;
	wire _w9775_ ;
	wire _w9776_ ;
	wire _w9777_ ;
	wire _w9778_ ;
	wire _w9779_ ;
	wire _w9780_ ;
	wire _w9781_ ;
	wire _w9782_ ;
	wire _w9783_ ;
	wire _w9784_ ;
	wire _w9785_ ;
	wire _w9786_ ;
	wire _w9787_ ;
	wire _w9788_ ;
	wire _w9789_ ;
	wire _w9790_ ;
	wire _w9791_ ;
	wire _w9792_ ;
	wire _w9793_ ;
	wire _w9794_ ;
	wire _w9795_ ;
	wire _w9796_ ;
	wire _w9797_ ;
	wire _w9798_ ;
	wire _w9799_ ;
	wire _w9800_ ;
	wire _w9801_ ;
	wire _w9802_ ;
	wire _w9803_ ;
	wire _w9804_ ;
	wire _w9805_ ;
	wire _w9806_ ;
	wire _w9807_ ;
	wire _w9808_ ;
	wire _w9809_ ;
	wire _w9810_ ;
	wire _w9811_ ;
	wire _w9812_ ;
	wire _w9813_ ;
	wire _w9814_ ;
	wire _w9815_ ;
	wire _w9816_ ;
	wire _w9817_ ;
	wire _w9818_ ;
	wire _w9819_ ;
	wire _w9820_ ;
	wire _w9821_ ;
	wire _w9822_ ;
	wire _w9823_ ;
	wire _w9824_ ;
	wire _w9825_ ;
	wire _w9826_ ;
	wire _w9827_ ;
	wire _w9828_ ;
	wire _w9829_ ;
	wire _w9830_ ;
	wire _w9831_ ;
	wire _w9832_ ;
	wire _w9833_ ;
	wire _w9834_ ;
	wire _w9835_ ;
	wire _w9836_ ;
	wire _w9837_ ;
	wire _w9838_ ;
	wire _w9839_ ;
	wire _w9840_ ;
	wire _w9841_ ;
	wire _w9842_ ;
	wire _w9843_ ;
	wire _w9844_ ;
	wire _w9845_ ;
	wire _w9846_ ;
	wire _w9847_ ;
	wire _w9848_ ;
	wire _w9849_ ;
	wire _w9850_ ;
	wire _w9851_ ;
	wire _w9852_ ;
	wire _w9853_ ;
	wire _w9854_ ;
	wire _w9855_ ;
	wire _w9856_ ;
	wire _w9857_ ;
	wire _w9858_ ;
	wire _w9859_ ;
	wire _w9860_ ;
	wire _w9861_ ;
	wire _w9862_ ;
	wire _w9863_ ;
	wire _w9864_ ;
	wire _w9865_ ;
	wire _w9866_ ;
	wire _w9867_ ;
	wire _w9868_ ;
	wire _w9869_ ;
	wire _w9870_ ;
	wire _w9871_ ;
	wire _w9872_ ;
	wire _w9873_ ;
	wire _w9874_ ;
	wire _w9875_ ;
	wire _w9876_ ;
	wire _w9877_ ;
	wire _w9878_ ;
	wire _w9879_ ;
	wire _w9880_ ;
	wire _w9881_ ;
	wire _w9882_ ;
	wire _w9883_ ;
	wire _w9884_ ;
	wire _w9885_ ;
	wire _w9886_ ;
	wire _w9887_ ;
	wire _w9888_ ;
	wire _w9889_ ;
	wire _w9890_ ;
	wire _w9891_ ;
	wire _w9892_ ;
	wire _w9893_ ;
	wire _w9894_ ;
	wire _w9895_ ;
	wire _w9896_ ;
	wire _w9897_ ;
	wire _w9898_ ;
	wire _w9899_ ;
	wire _w9900_ ;
	wire _w9901_ ;
	wire _w9902_ ;
	wire _w9903_ ;
	wire _w9904_ ;
	wire _w9905_ ;
	wire _w9906_ ;
	wire _w9907_ ;
	wire _w9908_ ;
	wire _w9909_ ;
	wire _w9910_ ;
	wire _w9911_ ;
	wire _w9912_ ;
	wire _w9913_ ;
	wire _w9914_ ;
	wire _w9915_ ;
	wire _w9916_ ;
	wire _w9917_ ;
	wire _w9918_ ;
	wire _w9919_ ;
	wire _w9920_ ;
	wire _w9921_ ;
	wire _w9922_ ;
	wire _w9923_ ;
	wire _w9924_ ;
	wire _w9925_ ;
	wire _w9926_ ;
	wire _w9927_ ;
	wire _w9928_ ;
	wire _w9929_ ;
	wire _w9930_ ;
	wire _w9931_ ;
	wire _w9932_ ;
	wire _w9933_ ;
	wire _w9934_ ;
	wire _w9935_ ;
	wire _w9936_ ;
	wire _w9937_ ;
	wire _w9938_ ;
	wire _w9939_ ;
	wire _w9940_ ;
	wire _w9941_ ;
	wire _w9942_ ;
	wire _w9943_ ;
	wire _w9944_ ;
	wire _w9945_ ;
	wire _w9946_ ;
	wire _w9947_ ;
	wire _w9948_ ;
	wire _w9949_ ;
	wire _w9950_ ;
	wire _w9951_ ;
	wire _w9952_ ;
	wire _w9953_ ;
	wire _w9954_ ;
	wire _w9955_ ;
	wire _w9956_ ;
	wire _w9957_ ;
	wire _w9958_ ;
	wire _w9959_ ;
	wire _w9960_ ;
	wire _w9961_ ;
	wire _w9962_ ;
	wire _w9963_ ;
	wire _w9964_ ;
	wire _w9965_ ;
	wire _w9966_ ;
	wire _w9967_ ;
	wire _w9968_ ;
	wire _w9969_ ;
	wire _w9970_ ;
	wire _w9971_ ;
	wire _w9972_ ;
	wire _w9973_ ;
	wire _w9974_ ;
	wire _w9975_ ;
	wire _w9976_ ;
	wire _w9977_ ;
	wire _w9978_ ;
	wire _w9979_ ;
	wire _w9980_ ;
	wire _w9981_ ;
	wire _w9982_ ;
	wire _w9983_ ;
	wire _w9984_ ;
	wire _w9985_ ;
	wire _w9986_ ;
	wire _w9987_ ;
	wire _w9988_ ;
	wire _w9989_ ;
	wire _w9990_ ;
	wire _w9991_ ;
	wire _w9992_ ;
	wire _w9993_ ;
	wire _w9994_ ;
	wire _w9995_ ;
	wire _w9996_ ;
	wire _w9997_ ;
	wire _w9998_ ;
	wire _w9999_ ;
	wire _w10000_ ;
	wire _w10001_ ;
	wire _w10002_ ;
	wire _w10003_ ;
	wire _w10004_ ;
	wire _w10005_ ;
	wire _w10006_ ;
	wire _w10007_ ;
	wire _w10008_ ;
	wire _w10009_ ;
	wire _w10010_ ;
	wire _w10011_ ;
	wire _w10012_ ;
	wire _w10013_ ;
	wire _w10014_ ;
	wire _w10015_ ;
	wire _w10016_ ;
	wire _w10017_ ;
	wire _w10018_ ;
	wire _w10019_ ;
	wire _w10020_ ;
	wire _w10021_ ;
	wire _w10022_ ;
	wire _w10023_ ;
	wire _w10024_ ;
	wire _w10025_ ;
	wire _w10026_ ;
	wire _w10027_ ;
	wire _w10028_ ;
	wire _w10029_ ;
	wire _w10030_ ;
	wire _w10031_ ;
	wire _w10032_ ;
	wire _w10033_ ;
	wire _w10034_ ;
	wire _w10035_ ;
	wire _w10036_ ;
	wire _w10037_ ;
	wire _w10038_ ;
	wire _w10039_ ;
	wire _w10040_ ;
	wire _w10041_ ;
	wire _w10042_ ;
	wire _w10043_ ;
	wire _w10044_ ;
	wire _w10045_ ;
	wire _w10046_ ;
	wire _w10047_ ;
	wire _w10048_ ;
	wire _w10049_ ;
	wire _w10050_ ;
	wire _w10051_ ;
	wire _w10052_ ;
	wire _w10053_ ;
	wire _w10054_ ;
	wire _w10055_ ;
	wire _w10056_ ;
	wire _w10057_ ;
	wire _w10058_ ;
	wire _w10059_ ;
	wire _w10060_ ;
	wire _w10061_ ;
	wire _w10062_ ;
	wire _w10063_ ;
	wire _w10064_ ;
	wire _w10065_ ;
	wire _w10066_ ;
	wire _w10067_ ;
	wire _w10068_ ;
	wire _w10069_ ;
	wire _w10070_ ;
	wire _w10071_ ;
	wire _w10072_ ;
	wire _w10073_ ;
	wire _w10074_ ;
	wire _w10075_ ;
	wire _w10076_ ;
	wire _w10077_ ;
	wire _w10078_ ;
	wire _w10079_ ;
	wire _w10080_ ;
	wire _w10081_ ;
	wire _w10082_ ;
	wire _w10083_ ;
	wire _w10084_ ;
	wire _w10085_ ;
	wire _w10086_ ;
	wire _w10087_ ;
	wire _w10088_ ;
	wire _w10089_ ;
	wire _w10090_ ;
	wire _w10091_ ;
	wire _w10092_ ;
	wire _w10093_ ;
	wire _w10094_ ;
	wire _w10095_ ;
	wire _w10096_ ;
	wire _w10097_ ;
	wire _w10098_ ;
	wire _w10099_ ;
	wire _w10100_ ;
	wire _w10101_ ;
	wire _w10102_ ;
	wire _w10103_ ;
	wire _w10104_ ;
	wire _w10105_ ;
	wire _w10106_ ;
	wire _w10107_ ;
	wire _w10108_ ;
	wire _w10109_ ;
	wire _w10110_ ;
	wire _w10111_ ;
	wire _w10112_ ;
	wire _w10113_ ;
	wire _w10114_ ;
	wire _w10115_ ;
	wire _w10116_ ;
	wire _w10117_ ;
	wire _w10118_ ;
	wire _w10119_ ;
	wire _w10120_ ;
	wire _w10121_ ;
	wire _w10122_ ;
	wire _w10123_ ;
	wire _w10124_ ;
	wire _w10125_ ;
	wire _w10126_ ;
	wire _w10127_ ;
	wire _w10128_ ;
	wire _w10129_ ;
	wire _w10130_ ;
	wire _w10131_ ;
	wire _w10132_ ;
	wire _w10133_ ;
	wire _w10134_ ;
	wire _w10135_ ;
	wire _w10136_ ;
	wire _w10137_ ;
	wire _w10138_ ;
	wire _w10139_ ;
	wire _w10140_ ;
	wire _w10141_ ;
	wire _w10142_ ;
	wire _w10143_ ;
	wire _w10144_ ;
	wire _w10145_ ;
	wire _w10146_ ;
	wire _w10147_ ;
	wire _w10148_ ;
	wire _w10149_ ;
	wire _w10150_ ;
	wire _w10151_ ;
	wire _w10152_ ;
	wire _w10153_ ;
	wire _w10154_ ;
	wire _w10155_ ;
	wire _w10156_ ;
	wire _w10157_ ;
	wire _w10158_ ;
	wire _w10159_ ;
	wire _w10160_ ;
	wire _w10161_ ;
	wire _w10162_ ;
	wire _w10163_ ;
	wire _w10164_ ;
	wire _w10165_ ;
	wire _w10166_ ;
	wire _w10167_ ;
	wire _w10168_ ;
	wire _w10169_ ;
	wire _w10170_ ;
	wire _w10171_ ;
	wire _w10172_ ;
	wire _w10173_ ;
	wire _w10174_ ;
	wire _w10175_ ;
	wire _w10176_ ;
	wire _w10177_ ;
	wire _w10178_ ;
	wire _w10179_ ;
	wire _w10180_ ;
	wire _w10181_ ;
	wire _w10182_ ;
	wire _w10183_ ;
	wire _w10184_ ;
	wire _w10185_ ;
	wire _w10186_ ;
	wire _w10187_ ;
	wire _w10188_ ;
	wire _w10189_ ;
	wire _w10190_ ;
	wire _w10191_ ;
	wire _w10192_ ;
	wire _w10193_ ;
	wire _w10194_ ;
	wire _w10195_ ;
	wire _w10196_ ;
	wire _w10197_ ;
	wire _w10198_ ;
	wire _w10199_ ;
	wire _w10200_ ;
	wire _w10201_ ;
	wire _w10202_ ;
	wire _w10203_ ;
	wire _w10204_ ;
	wire _w10205_ ;
	wire _w10206_ ;
	wire _w10207_ ;
	wire _w10208_ ;
	wire _w10209_ ;
	wire _w10210_ ;
	wire _w10211_ ;
	wire _w10212_ ;
	wire _w10213_ ;
	wire _w10214_ ;
	wire _w10215_ ;
	wire _w10216_ ;
	wire _w10217_ ;
	wire _w10218_ ;
	wire _w10219_ ;
	wire _w10220_ ;
	wire _w10221_ ;
	wire _w10222_ ;
	wire _w10223_ ;
	wire _w10224_ ;
	wire _w10225_ ;
	wire _w10226_ ;
	wire _w10227_ ;
	wire _w10228_ ;
	wire _w10229_ ;
	wire _w10230_ ;
	wire _w10231_ ;
	wire _w10232_ ;
	wire _w10233_ ;
	wire _w10234_ ;
	wire _w10235_ ;
	wire _w10236_ ;
	wire _w10237_ ;
	wire _w10238_ ;
	wire _w10239_ ;
	wire _w10240_ ;
	wire _w10241_ ;
	wire _w10242_ ;
	wire _w10243_ ;
	wire _w10244_ ;
	wire _w10245_ ;
	wire _w10246_ ;
	wire _w10247_ ;
	wire _w10248_ ;
	wire _w10249_ ;
	wire _w10250_ ;
	wire _w10251_ ;
	wire _w10252_ ;
	wire _w10253_ ;
	wire _w10254_ ;
	wire _w10255_ ;
	wire _w10256_ ;
	wire _w10257_ ;
	wire _w10258_ ;
	wire _w10259_ ;
	wire _w10260_ ;
	wire _w10261_ ;
	wire _w10262_ ;
	wire _w10263_ ;
	wire _w10264_ ;
	wire _w10265_ ;
	wire _w10266_ ;
	wire _w10267_ ;
	wire _w10268_ ;
	wire _w10269_ ;
	wire _w10270_ ;
	wire _w10271_ ;
	wire _w10272_ ;
	wire _w10273_ ;
	wire _w10274_ ;
	wire _w10275_ ;
	wire _w10276_ ;
	wire _w10277_ ;
	wire _w10278_ ;
	wire _w10279_ ;
	wire _w10280_ ;
	wire _w10281_ ;
	wire _w10282_ ;
	wire _w10283_ ;
	wire _w10284_ ;
	wire _w10285_ ;
	wire _w10286_ ;
	wire _w10287_ ;
	wire _w10288_ ;
	wire _w10289_ ;
	wire _w10290_ ;
	wire _w10291_ ;
	wire _w10292_ ;
	wire _w10293_ ;
	wire _w10294_ ;
	wire _w10295_ ;
	wire _w10296_ ;
	wire _w10297_ ;
	wire _w10298_ ;
	wire _w10299_ ;
	wire _w10300_ ;
	wire _w10301_ ;
	wire _w10302_ ;
	wire _w10303_ ;
	wire _w10304_ ;
	wire _w10305_ ;
	wire _w10306_ ;
	wire _w10307_ ;
	wire _w10308_ ;
	wire _w10309_ ;
	wire _w10310_ ;
	wire _w10311_ ;
	wire _w10312_ ;
	wire _w10313_ ;
	wire _w10314_ ;
	wire _w10315_ ;
	wire _w10316_ ;
	wire _w10317_ ;
	wire _w10318_ ;
	wire _w10319_ ;
	wire _w10320_ ;
	wire _w10321_ ;
	wire _w10322_ ;
	wire _w10323_ ;
	wire _w10324_ ;
	wire _w10325_ ;
	wire _w10326_ ;
	wire _w10327_ ;
	wire _w10328_ ;
	wire _w10329_ ;
	wire _w10330_ ;
	wire _w10331_ ;
	wire _w10332_ ;
	wire _w10333_ ;
	wire _w10334_ ;
	wire _w10335_ ;
	wire _w10336_ ;
	wire _w10337_ ;
	wire _w10338_ ;
	wire _w10339_ ;
	wire _w10340_ ;
	wire _w10341_ ;
	wire _w10342_ ;
	wire _w10343_ ;
	wire _w10344_ ;
	wire _w10345_ ;
	wire _w10346_ ;
	wire _w10347_ ;
	wire _w10348_ ;
	wire _w10349_ ;
	wire _w10350_ ;
	wire _w10351_ ;
	wire _w10352_ ;
	wire _w10353_ ;
	wire _w10354_ ;
	wire _w10355_ ;
	wire _w10356_ ;
	wire _w10357_ ;
	wire _w10358_ ;
	wire _w10359_ ;
	wire _w10360_ ;
	wire _w10361_ ;
	wire _w10362_ ;
	wire _w10363_ ;
	wire _w10364_ ;
	wire _w10365_ ;
	wire _w10366_ ;
	wire _w10367_ ;
	wire _w10368_ ;
	wire _w10369_ ;
	wire _w10370_ ;
	wire _w10371_ ;
	wire _w10372_ ;
	wire _w10373_ ;
	wire _w10374_ ;
	wire _w10375_ ;
	wire _w10376_ ;
	wire _w10377_ ;
	wire _w10378_ ;
	wire _w10379_ ;
	wire _w10380_ ;
	wire _w10381_ ;
	wire _w10382_ ;
	wire _w10383_ ;
	wire _w10384_ ;
	wire _w10385_ ;
	wire _w10386_ ;
	wire _w10387_ ;
	wire _w10388_ ;
	wire _w10389_ ;
	wire _w10390_ ;
	wire _w10391_ ;
	wire _w10392_ ;
	wire _w10393_ ;
	wire _w10394_ ;
	wire _w10395_ ;
	wire _w10396_ ;
	wire _w10397_ ;
	wire _w10398_ ;
	wire _w10399_ ;
	wire _w10400_ ;
	wire _w10401_ ;
	wire _w10402_ ;
	wire _w10403_ ;
	wire _w10404_ ;
	wire _w10405_ ;
	wire _w10406_ ;
	wire _w10407_ ;
	wire _w10408_ ;
	wire _w10409_ ;
	wire _w10410_ ;
	wire _w10411_ ;
	wire _w10412_ ;
	wire _w10413_ ;
	wire _w10414_ ;
	wire _w10415_ ;
	wire _w10416_ ;
	wire _w10417_ ;
	wire _w10418_ ;
	wire _w10419_ ;
	wire _w10420_ ;
	wire _w10421_ ;
	wire _w10422_ ;
	wire _w10423_ ;
	wire _w10424_ ;
	wire _w10425_ ;
	wire _w10426_ ;
	wire _w10427_ ;
	wire _w10428_ ;
	wire _w10429_ ;
	wire _w10430_ ;
	wire _w10431_ ;
	wire _w10432_ ;
	wire _w10433_ ;
	wire _w10434_ ;
	wire _w10435_ ;
	wire _w10436_ ;
	wire _w10437_ ;
	wire _w10438_ ;
	wire _w10439_ ;
	wire _w10440_ ;
	wire _w10441_ ;
	wire _w10442_ ;
	wire _w10443_ ;
	wire _w10444_ ;
	wire _w10445_ ;
	wire _w10446_ ;
	wire _w10447_ ;
	wire _w10448_ ;
	wire _w10449_ ;
	wire _w10450_ ;
	wire _w10451_ ;
	wire _w10452_ ;
	wire _w10453_ ;
	wire _w10454_ ;
	wire _w10455_ ;
	wire _w10456_ ;
	wire _w10457_ ;
	wire _w10458_ ;
	wire _w10459_ ;
	wire _w10460_ ;
	wire _w10461_ ;
	wire _w10462_ ;
	wire _w10463_ ;
	wire _w10464_ ;
	wire _w10465_ ;
	wire _w10466_ ;
	wire _w10467_ ;
	wire _w10468_ ;
	wire _w10469_ ;
	wire _w10470_ ;
	wire _w10471_ ;
	wire _w10472_ ;
	wire _w10473_ ;
	wire _w10474_ ;
	wire _w10475_ ;
	wire _w10476_ ;
	wire _w10477_ ;
	wire _w10478_ ;
	wire _w10479_ ;
	wire _w10480_ ;
	wire _w10481_ ;
	wire _w10482_ ;
	wire _w10483_ ;
	wire _w10484_ ;
	wire _w10485_ ;
	wire _w10486_ ;
	wire _w10487_ ;
	wire _w10488_ ;
	wire _w10489_ ;
	wire _w10490_ ;
	wire _w10491_ ;
	wire _w10492_ ;
	wire _w10493_ ;
	wire _w10494_ ;
	wire _w10495_ ;
	wire _w10496_ ;
	wire _w10497_ ;
	wire _w10498_ ;
	wire _w10499_ ;
	wire _w10500_ ;
	wire _w10501_ ;
	wire _w10502_ ;
	wire _w10503_ ;
	wire _w10504_ ;
	wire _w10505_ ;
	wire _w10506_ ;
	wire _w10507_ ;
	wire _w10508_ ;
	wire _w10509_ ;
	wire _w10510_ ;
	wire _w10511_ ;
	wire _w10512_ ;
	wire _w10513_ ;
	wire _w10514_ ;
	wire _w10515_ ;
	wire _w10516_ ;
	wire _w10517_ ;
	wire _w10518_ ;
	wire _w10519_ ;
	wire _w10520_ ;
	wire _w10521_ ;
	wire _w10522_ ;
	wire _w10523_ ;
	wire _w10524_ ;
	wire _w10525_ ;
	wire _w10526_ ;
	wire _w10527_ ;
	wire _w10528_ ;
	wire _w10529_ ;
	wire _w10530_ ;
	wire _w10531_ ;
	wire _w10532_ ;
	wire _w10533_ ;
	wire _w10534_ ;
	wire _w10535_ ;
	wire _w10536_ ;
	wire _w10537_ ;
	wire _w10538_ ;
	wire _w10539_ ;
	wire _w10540_ ;
	wire _w10541_ ;
	wire _w10542_ ;
	wire _w10543_ ;
	wire _w10544_ ;
	wire _w10545_ ;
	wire _w10546_ ;
	wire _w10547_ ;
	wire _w10548_ ;
	wire _w10549_ ;
	wire _w10550_ ;
	wire _w10551_ ;
	wire _w10552_ ;
	wire _w10553_ ;
	wire _w10554_ ;
	wire _w10555_ ;
	wire _w10556_ ;
	wire _w10557_ ;
	wire _w10558_ ;
	wire _w10559_ ;
	wire _w10560_ ;
	wire _w10561_ ;
	wire _w10562_ ;
	wire _w10563_ ;
	wire _w10564_ ;
	wire _w10565_ ;
	wire _w10566_ ;
	wire _w10567_ ;
	wire _w10568_ ;
	wire _w10569_ ;
	wire _w10570_ ;
	wire _w10571_ ;
	wire _w10572_ ;
	wire _w10573_ ;
	wire _w10574_ ;
	wire _w10575_ ;
	wire _w10576_ ;
	wire _w10577_ ;
	wire _w10578_ ;
	wire _w10579_ ;
	wire _w10580_ ;
	wire _w10581_ ;
	wire _w10582_ ;
	wire _w10583_ ;
	wire _w10584_ ;
	wire _w10585_ ;
	wire _w10586_ ;
	wire _w10587_ ;
	wire _w10588_ ;
	wire _w10589_ ;
	wire _w10590_ ;
	wire _w10591_ ;
	wire _w10592_ ;
	wire _w10593_ ;
	wire _w10594_ ;
	wire _w10595_ ;
	wire _w10596_ ;
	wire _w10597_ ;
	wire _w10598_ ;
	wire _w10599_ ;
	wire _w10600_ ;
	wire _w10601_ ;
	wire _w10602_ ;
	wire _w10603_ ;
	wire _w10604_ ;
	wire _w10605_ ;
	wire _w10606_ ;
	wire _w10607_ ;
	wire _w10608_ ;
	wire _w10609_ ;
	wire _w10610_ ;
	wire _w10611_ ;
	wire _w10612_ ;
	wire _w10613_ ;
	wire _w10614_ ;
	wire _w10615_ ;
	wire _w10616_ ;
	wire _w10617_ ;
	wire _w10618_ ;
	wire _w10619_ ;
	wire _w10620_ ;
	wire _w10621_ ;
	wire _w10622_ ;
	wire _w10623_ ;
	wire _w10624_ ;
	wire _w10625_ ;
	wire _w10626_ ;
	wire _w10627_ ;
	wire _w10628_ ;
	wire _w10629_ ;
	wire _w10630_ ;
	wire _w10631_ ;
	wire _w10632_ ;
	wire _w10633_ ;
	wire _w10634_ ;
	wire _w10635_ ;
	wire _w10636_ ;
	wire _w10637_ ;
	wire _w10638_ ;
	wire _w10639_ ;
	wire _w10640_ ;
	wire _w10641_ ;
	wire _w10642_ ;
	wire _w10643_ ;
	wire _w10644_ ;
	wire _w10645_ ;
	wire _w10646_ ;
	wire _w10647_ ;
	wire _w10648_ ;
	wire _w10649_ ;
	wire _w10650_ ;
	wire _w10651_ ;
	wire _w10652_ ;
	wire _w10653_ ;
	wire _w10654_ ;
	wire _w10655_ ;
	wire _w10656_ ;
	wire _w10657_ ;
	wire _w10658_ ;
	wire _w10659_ ;
	wire _w10660_ ;
	wire _w10661_ ;
	wire _w10662_ ;
	wire _w10663_ ;
	wire _w10664_ ;
	wire _w10665_ ;
	wire _w10666_ ;
	wire _w10667_ ;
	wire _w10668_ ;
	wire _w10669_ ;
	wire _w10670_ ;
	wire _w10671_ ;
	wire _w10672_ ;
	wire _w10673_ ;
	wire _w10674_ ;
	wire _w10675_ ;
	wire _w10676_ ;
	wire _w10677_ ;
	wire _w10678_ ;
	wire _w10679_ ;
	wire _w10680_ ;
	wire _w10681_ ;
	wire _w10682_ ;
	wire _w10683_ ;
	wire _w10684_ ;
	wire _w10685_ ;
	wire _w10686_ ;
	wire _w10687_ ;
	wire _w10688_ ;
	wire _w10689_ ;
	wire _w10690_ ;
	wire _w10691_ ;
	wire _w10692_ ;
	wire _w10693_ ;
	wire _w10694_ ;
	wire _w10695_ ;
	wire _w10696_ ;
	wire _w10697_ ;
	wire _w10698_ ;
	wire _w10699_ ;
	wire _w10700_ ;
	wire _w10701_ ;
	wire _w10702_ ;
	wire _w10703_ ;
	wire _w10704_ ;
	wire _w10705_ ;
	wire _w10706_ ;
	wire _w10707_ ;
	wire _w10708_ ;
	wire _w10709_ ;
	wire _w10710_ ;
	wire _w10711_ ;
	wire _w10712_ ;
	wire _w10713_ ;
	wire _w10714_ ;
	wire _w10715_ ;
	wire _w10716_ ;
	wire _w10717_ ;
	wire _w10718_ ;
	wire _w10719_ ;
	wire _w10720_ ;
	wire _w10721_ ;
	wire _w10722_ ;
	wire _w10723_ ;
	wire _w10724_ ;
	wire _w10725_ ;
	wire _w10726_ ;
	wire _w10727_ ;
	wire _w10728_ ;
	wire _w10729_ ;
	wire _w10730_ ;
	wire _w10731_ ;
	wire _w10732_ ;
	wire _w10733_ ;
	wire _w10734_ ;
	wire _w10735_ ;
	wire _w10736_ ;
	wire _w10737_ ;
	wire _w10738_ ;
	wire _w10739_ ;
	wire _w10740_ ;
	wire _w10741_ ;
	wire _w10742_ ;
	wire _w10743_ ;
	wire _w10744_ ;
	wire _w10745_ ;
	wire _w10746_ ;
	wire _w10747_ ;
	wire _w10748_ ;
	wire _w10749_ ;
	wire _w10750_ ;
	wire _w10751_ ;
	wire _w10752_ ;
	wire _w10753_ ;
	wire _w10754_ ;
	wire _w10755_ ;
	wire _w10756_ ;
	wire _w10757_ ;
	wire _w10758_ ;
	wire _w10759_ ;
	wire _w10760_ ;
	wire _w10761_ ;
	wire _w10762_ ;
	wire _w10763_ ;
	wire _w10764_ ;
	wire _w10765_ ;
	wire _w10766_ ;
	wire _w10767_ ;
	wire _w10768_ ;
	wire _w10769_ ;
	wire _w10770_ ;
	wire _w10771_ ;
	wire _w10772_ ;
	wire _w10773_ ;
	wire _w10774_ ;
	wire _w10775_ ;
	wire _w10776_ ;
	wire _w10777_ ;
	wire _w10778_ ;
	wire _w10779_ ;
	wire _w10780_ ;
	wire _w10781_ ;
	wire _w10782_ ;
	wire _w10783_ ;
	wire _w10784_ ;
	wire _w10785_ ;
	wire _w10786_ ;
	wire _w10787_ ;
	wire _w10788_ ;
	wire _w10789_ ;
	wire _w10790_ ;
	wire _w10791_ ;
	wire _w10792_ ;
	wire _w10793_ ;
	wire _w10794_ ;
	wire _w10795_ ;
	wire _w10796_ ;
	wire _w10797_ ;
	wire _w10798_ ;
	wire _w10799_ ;
	wire _w10800_ ;
	wire _w10801_ ;
	wire _w10802_ ;
	wire _w10803_ ;
	wire _w10804_ ;
	wire _w10805_ ;
	wire _w10806_ ;
	wire _w10807_ ;
	wire _w10808_ ;
	wire _w10809_ ;
	wire _w10810_ ;
	wire _w10811_ ;
	wire _w10812_ ;
	wire _w10813_ ;
	wire _w10814_ ;
	wire _w10815_ ;
	wire _w10816_ ;
	wire _w10817_ ;
	wire _w10818_ ;
	wire _w10819_ ;
	wire _w10820_ ;
	wire _w10822_ ;
	wire _w10824_ ;
	wire _w10826_ ;
	wire _w10828_ ;
	wire _w10830_ ;
	wire _w10832_ ;
	wire _w10834_ ;
	wire _w10835_ ;
	wire _w10836_ ;
	wire _w10837_ ;
	wire _w10838_ ;
	wire _w10839_ ;
	wire _w10840_ ;
	wire _w10841_ ;
	wire _w10842_ ;
	wire _w10843_ ;
	wire _w10844_ ;
	wire _w10845_ ;
	wire _w10846_ ;
	wire _w10847_ ;
	wire _w10848_ ;
	wire _w10850_ ;
	wire _w10851_ ;
	wire _w10852_ ;
	wire _w10853_ ;
	wire _w10854_ ;
	wire _w10855_ ;
	wire _w10856_ ;
	wire _w10857_ ;
	wire _w10858_ ;
	wire _w10859_ ;
	wire _w10860_ ;
	wire _w10861_ ;
	wire _w10862_ ;
	wire _w10863_ ;
	wire _w10864_ ;
	wire _w10865_ ;
	wire _w10866_ ;
	wire _w10867_ ;
	wire _w10868_ ;
	wire _w10869_ ;
	wire _w10870_ ;
	wire _w10871_ ;
	wire _w10872_ ;
	wire _w10873_ ;
	wire _w10874_ ;
	wire _w10875_ ;
	wire _w10876_ ;
	wire _w10877_ ;
	wire _w10878_ ;
	wire _w10879_ ;
	wire _w10880_ ;
	wire _w10881_ ;
	wire _w10882_ ;
	wire _w10883_ ;
	wire _w10884_ ;
	wire _w10885_ ;
	wire _w10886_ ;
	wire _w10887_ ;
	wire _w10888_ ;
	wire _w10889_ ;
	wire _w10890_ ;
	wire _w10891_ ;
	wire _w10892_ ;
	wire _w10893_ ;
	wire _w10894_ ;
	wire _w10895_ ;
	wire _w10896_ ;
	wire _w10897_ ;
	wire _w10898_ ;
	wire _w10899_ ;
	wire _w10900_ ;
	wire _w10901_ ;
	wire _w10902_ ;
	wire _w10903_ ;
	wire _w10904_ ;
	wire _w10905_ ;
	wire _w10906_ ;
	wire _w10907_ ;
	wire _w10908_ ;
	wire _w10909_ ;
	wire _w10910_ ;
	wire _w10911_ ;
	wire _w10912_ ;
	wire _w10913_ ;
	wire _w10914_ ;
	wire _w10915_ ;
	wire _w10916_ ;
	wire _w10917_ ;
	wire _w10918_ ;
	wire _w10920_ ;
	wire _w10921_ ;
	wire _w10922_ ;
	wire _w10923_ ;
	wire _w10924_ ;
	wire _w10925_ ;
	wire _w10926_ ;
	wire _w10927_ ;
	wire _w10928_ ;
	wire _w10929_ ;
	wire _w10930_ ;
	wire _w10931_ ;
	wire _w10932_ ;
	wire _w10933_ ;
	wire _w10934_ ;
	wire _w10935_ ;
	wire _w10936_ ;
	wire _w10937_ ;
	wire _w10938_ ;
	wire _w10939_ ;
	wire _w10940_ ;
	wire _w10941_ ;
	wire _w10942_ ;
	wire _w10943_ ;
	wire _w10944_ ;
	wire _w10945_ ;
	wire _w10946_ ;
	wire _w10947_ ;
	wire _w10948_ ;
	wire _w10949_ ;
	wire _w10950_ ;
	wire _w10951_ ;
	wire _w10952_ ;
	wire _w10953_ ;
	wire _w10954_ ;
	wire _w10955_ ;
	wire _w10956_ ;
	wire _w10957_ ;
	wire _w10958_ ;
	wire _w10959_ ;
	wire _w10960_ ;
	wire _w10961_ ;
	wire _w10962_ ;
	wire _w10963_ ;
	wire _w10964_ ;
	wire _w10965_ ;
	wire _w10966_ ;
	wire _w10967_ ;
	wire _w10968_ ;
	wire _w10969_ ;
	wire _w10970_ ;
	wire _w10971_ ;
	wire _w10972_ ;
	wire _w10973_ ;
	wire _w10974_ ;
	wire _w10975_ ;
	wire _w10976_ ;
	wire _w10977_ ;
	wire _w10978_ ;
	wire _w10979_ ;
	wire _w10980_ ;
	wire _w10981_ ;
	wire _w10982_ ;
	wire _w10983_ ;
	wire _w10984_ ;
	wire _w10985_ ;
	wire _w10986_ ;
	wire _w10987_ ;
	wire _w10988_ ;
	wire _w10989_ ;
	wire _w10990_ ;
	wire _w10991_ ;
	wire _w10992_ ;
	wire _w10993_ ;
	wire _w10994_ ;
	wire _w10995_ ;
	wire _w10996_ ;
	wire _w10997_ ;
	wire _w10998_ ;
	wire _w10999_ ;
	wire _w11000_ ;
	wire _w11001_ ;
	wire _w11002_ ;
	wire _w11003_ ;
	wire _w11004_ ;
	wire _w11005_ ;
	wire _w11006_ ;
	wire _w11007_ ;
	wire _w11008_ ;
	wire _w11009_ ;
	wire _w11010_ ;
	wire _w11011_ ;
	wire _w11012_ ;
	wire _w11013_ ;
	wire _w11014_ ;
	wire _w11015_ ;
	wire _w11016_ ;
	wire _w11017_ ;
	wire _w11018_ ;
	wire _w11019_ ;
	wire _w11020_ ;
	wire _w11021_ ;
	wire _w11022_ ;
	wire _w11023_ ;
	wire _w11024_ ;
	wire _w11025_ ;
	wire _w11026_ ;
	wire _w11027_ ;
	wire _w11028_ ;
	wire _w11029_ ;
	wire _w11030_ ;
	wire _w11031_ ;
	wire _w11032_ ;
	wire _w11033_ ;
	wire _w11034_ ;
	wire _w11035_ ;
	wire _w11036_ ;
	wire _w11037_ ;
	wire _w11038_ ;
	wire _w11039_ ;
	wire _w11040_ ;
	wire _w11041_ ;
	wire _w11042_ ;
	wire _w11043_ ;
	wire _w11044_ ;
	wire _w11045_ ;
	wire _w11046_ ;
	wire _w11047_ ;
	wire _w11048_ ;
	wire _w11049_ ;
	wire _w11050_ ;
	wire _w11051_ ;
	wire _w11052_ ;
	wire _w11053_ ;
	wire _w11054_ ;
	wire _w11055_ ;
	wire _w11056_ ;
	wire _w11057_ ;
	wire _w11058_ ;
	wire _w11059_ ;
	wire _w11060_ ;
	wire _w11061_ ;
	wire _w11062_ ;
	wire _w11063_ ;
	wire _w11064_ ;
	wire _w11065_ ;
	wire _w11066_ ;
	wire _w11067_ ;
	wire _w11068_ ;
	wire _w11069_ ;
	wire _w11070_ ;
	wire _w11071_ ;
	wire _w11072_ ;
	wire _w11073_ ;
	wire _w11074_ ;
	wire _w11075_ ;
	wire _w11076_ ;
	wire _w11077_ ;
	wire _w11078_ ;
	wire _w11079_ ;
	wire _w11080_ ;
	wire _w11081_ ;
	wire _w11082_ ;
	wire _w11083_ ;
	wire _w11084_ ;
	wire _w11085_ ;
	wire _w11086_ ;
	wire _w11087_ ;
	wire _w11088_ ;
	wire _w11089_ ;
	wire _w11090_ ;
	wire _w11091_ ;
	wire _w11092_ ;
	wire _w11093_ ;
	wire _w11094_ ;
	wire _w11095_ ;
	wire _w11096_ ;
	wire _w11097_ ;
	wire _w11098_ ;
	wire _w11099_ ;
	wire _w11100_ ;
	wire _w11101_ ;
	wire _w11102_ ;
	wire _w11103_ ;
	wire _w11104_ ;
	wire _w11105_ ;
	wire _w11106_ ;
	wire _w11107_ ;
	wire _w11108_ ;
	wire _w11109_ ;
	wire _w11110_ ;
	wire _w11111_ ;
	wire _w11112_ ;
	wire _w11113_ ;
	wire _w11114_ ;
	wire _w11115_ ;
	wire _w11116_ ;
	wire _w11117_ ;
	wire _w11118_ ;
	wire _w11119_ ;
	wire _w11120_ ;
	wire _w11121_ ;
	wire _w11122_ ;
	wire _w11123_ ;
	wire _w11124_ ;
	wire _w11125_ ;
	wire _w11126_ ;
	wire _w11127_ ;
	wire _w11128_ ;
	wire _w11129_ ;
	wire _w11130_ ;
	wire _w11131_ ;
	wire _w11132_ ;
	wire _w11133_ ;
	wire _w11134_ ;
	wire _w11135_ ;
	wire _w11136_ ;
	wire _w11137_ ;
	wire _w11138_ ;
	wire _w11139_ ;
	wire _w11140_ ;
	wire _w11141_ ;
	wire _w11142_ ;
	wire _w11143_ ;
	wire _w11144_ ;
	wire _w11145_ ;
	wire _w11146_ ;
	wire _w11147_ ;
	wire _w11148_ ;
	wire _w11149_ ;
	wire _w11150_ ;
	wire _w11151_ ;
	wire _w11152_ ;
	wire _w11153_ ;
	wire _w11154_ ;
	wire _w11155_ ;
	wire _w11156_ ;
	wire _w11157_ ;
	wire _w11158_ ;
	wire _w11159_ ;
	wire _w11160_ ;
	wire _w11161_ ;
	wire _w11162_ ;
	wire _w11163_ ;
	wire _w11164_ ;
	wire _w11165_ ;
	wire _w11166_ ;
	wire _w11167_ ;
	wire _w11168_ ;
	wire _w11169_ ;
	wire _w11170_ ;
	wire _w11171_ ;
	wire _w11172_ ;
	wire _w11173_ ;
	wire _w11174_ ;
	wire _w11175_ ;
	wire _w11176_ ;
	wire _w11177_ ;
	wire _w11178_ ;
	wire _w11179_ ;
	wire _w11180_ ;
	wire _w11181_ ;
	wire _w11182_ ;
	wire _w11183_ ;
	wire _w11184_ ;
	wire _w11185_ ;
	wire _w11186_ ;
	wire _w11187_ ;
	wire _w11188_ ;
	wire _w11189_ ;
	wire _w11190_ ;
	wire _w11191_ ;
	wire _w11192_ ;
	wire _w11193_ ;
	wire _w11194_ ;
	wire _w11195_ ;
	wire _w11196_ ;
	wire _w11197_ ;
	wire _w11198_ ;
	wire _w11199_ ;
	wire _w11200_ ;
	wire _w11201_ ;
	wire _w11202_ ;
	wire _w11203_ ;
	wire _w11204_ ;
	wire _w11205_ ;
	wire _w11206_ ;
	wire _w11207_ ;
	wire _w11208_ ;
	wire _w11209_ ;
	wire _w11210_ ;
	wire _w11211_ ;
	wire _w11212_ ;
	wire _w11213_ ;
	wire _w11214_ ;
	wire _w11215_ ;
	wire _w11216_ ;
	wire _w11217_ ;
	wire _w11218_ ;
	wire _w11219_ ;
	wire _w11220_ ;
	wire _w11221_ ;
	wire _w11222_ ;
	wire _w11223_ ;
	wire _w11224_ ;
	wire _w11225_ ;
	wire _w11226_ ;
	wire _w11227_ ;
	wire _w11228_ ;
	wire _w11229_ ;
	wire _w11230_ ;
	wire _w11231_ ;
	wire _w11232_ ;
	wire _w11233_ ;
	wire _w11234_ ;
	wire _w11235_ ;
	wire _w11236_ ;
	wire _w11237_ ;
	wire _w11238_ ;
	wire _w11239_ ;
	wire _w11240_ ;
	wire _w11241_ ;
	wire _w11242_ ;
	wire _w11243_ ;
	wire _w11244_ ;
	wire _w11245_ ;
	wire _w11246_ ;
	wire _w11247_ ;
	wire _w11248_ ;
	wire _w11249_ ;
	wire _w11250_ ;
	wire _w11251_ ;
	wire _w11252_ ;
	wire _w11253_ ;
	wire _w11254_ ;
	wire _w11255_ ;
	wire _w11256_ ;
	wire _w11257_ ;
	wire _w11258_ ;
	wire _w11259_ ;
	wire _w11260_ ;
	wire _w11261_ ;
	wire _w11262_ ;
	wire _w11263_ ;
	wire _w11264_ ;
	wire _w11265_ ;
	wire _w11266_ ;
	wire _w11267_ ;
	wire _w11268_ ;
	wire _w11269_ ;
	wire _w11270_ ;
	wire _w11271_ ;
	wire _w11272_ ;
	wire _w11273_ ;
	wire _w11274_ ;
	wire _w11275_ ;
	wire _w11276_ ;
	wire _w11277_ ;
	wire _w11278_ ;
	wire _w11279_ ;
	wire _w11280_ ;
	wire _w11281_ ;
	wire _w11282_ ;
	wire _w11283_ ;
	wire _w11284_ ;
	wire _w11285_ ;
	wire _w11286_ ;
	wire _w11287_ ;
	wire _w11288_ ;
	wire _w11289_ ;
	wire _w11290_ ;
	wire _w11291_ ;
	wire _w11292_ ;
	wire _w11293_ ;
	wire _w11294_ ;
	wire _w11295_ ;
	wire _w11296_ ;
	wire _w11297_ ;
	wire _w11298_ ;
	wire _w11299_ ;
	wire _w11300_ ;
	wire _w11301_ ;
	wire _w11302_ ;
	wire _w11303_ ;
	wire _w11304_ ;
	wire _w11305_ ;
	wire _w11306_ ;
	wire _w11307_ ;
	wire _w11308_ ;
	wire _w11309_ ;
	wire _w11310_ ;
	wire _w11311_ ;
	wire _w11312_ ;
	wire _w11313_ ;
	wire _w11314_ ;
	wire _w11315_ ;
	wire _w11316_ ;
	wire _w11317_ ;
	wire _w11318_ ;
	wire _w11319_ ;
	wire _w11320_ ;
	wire _w11321_ ;
	wire _w11322_ ;
	wire _w11323_ ;
	wire _w11324_ ;
	wire _w11325_ ;
	wire _w11326_ ;
	wire _w11327_ ;
	wire _w11328_ ;
	wire _w11329_ ;
	wire _w11330_ ;
	wire _w11331_ ;
	wire _w11332_ ;
	wire _w11333_ ;
	wire _w11334_ ;
	wire _w11335_ ;
	wire _w11336_ ;
	wire _w11337_ ;
	wire _w11338_ ;
	wire _w11339_ ;
	wire _w11340_ ;
	wire _w11341_ ;
	wire _w11342_ ;
	wire _w11343_ ;
	wire _w11344_ ;
	wire _w11345_ ;
	wire _w11346_ ;
	wire _w11347_ ;
	wire _w11348_ ;
	wire _w11349_ ;
	wire _w11350_ ;
	wire _w11351_ ;
	wire _w11352_ ;
	wire _w11353_ ;
	wire _w11354_ ;
	wire _w11355_ ;
	wire _w11356_ ;
	wire _w11357_ ;
	wire _w11358_ ;
	wire _w11359_ ;
	wire _w11360_ ;
	wire _w11361_ ;
	wire _w11362_ ;
	wire _w11363_ ;
	wire _w11364_ ;
	wire _w11365_ ;
	wire _w11366_ ;
	wire _w11367_ ;
	wire _w11368_ ;
	wire _w11369_ ;
	wire _w11370_ ;
	wire _w11371_ ;
	wire _w11372_ ;
	wire _w11373_ ;
	wire _w11374_ ;
	wire _w11375_ ;
	wire _w11376_ ;
	wire _w11377_ ;
	wire _w11378_ ;
	wire _w11379_ ;
	wire _w11380_ ;
	wire _w11381_ ;
	wire _w11382_ ;
	wire _w11383_ ;
	wire _w11384_ ;
	wire _w11385_ ;
	wire _w11386_ ;
	wire _w11387_ ;
	wire _w11388_ ;
	wire _w11389_ ;
	wire _w11390_ ;
	wire _w11391_ ;
	wire _w11392_ ;
	wire _w11393_ ;
	wire _w11394_ ;
	wire _w11395_ ;
	wire _w11396_ ;
	wire _w11397_ ;
	wire _w11398_ ;
	wire _w11399_ ;
	wire _w11400_ ;
	wire _w11401_ ;
	wire _w11402_ ;
	wire _w11403_ ;
	wire _w11404_ ;
	wire _w11405_ ;
	wire _w11406_ ;
	wire _w11407_ ;
	wire _w11408_ ;
	wire _w11409_ ;
	wire _w11411_ ;
	wire _w11412_ ;
	wire _w11413_ ;
	wire _w11414_ ;
	wire _w11415_ ;
	wire _w11416_ ;
	wire _w11417_ ;
	wire _w11418_ ;
	wire _w11419_ ;
	wire _w11420_ ;
	wire _w11421_ ;
	wire _w11422_ ;
	wire _w11423_ ;
	wire _w11424_ ;
	wire _w11425_ ;
	wire _w11426_ ;
	wire _w11427_ ;
	wire _w11428_ ;
	wire _w11429_ ;
	wire _w11430_ ;
	wire _w11431_ ;
	wire _w11432_ ;
	wire _w11433_ ;
	wire _w11434_ ;
	wire _w11435_ ;
	wire _w11436_ ;
	wire _w11437_ ;
	wire _w11438_ ;
	wire _w11439_ ;
	wire _w11440_ ;
	wire _w11441_ ;
	wire _w11442_ ;
	wire _w11443_ ;
	wire _w11444_ ;
	wire _w11445_ ;
	wire _w11446_ ;
	wire _w11447_ ;
	wire _w11448_ ;
	wire _w11449_ ;
	wire _w11450_ ;
	wire _w11451_ ;
	wire _w11452_ ;
	wire _w11453_ ;
	wire _w11454_ ;
	wire _w11455_ ;
	wire _w11456_ ;
	wire _w11457_ ;
	wire _w11458_ ;
	wire _w11459_ ;
	wire _w11460_ ;
	wire _w11461_ ;
	wire _w11462_ ;
	wire _w11463_ ;
	wire _w11464_ ;
	wire _w11465_ ;
	wire _w11466_ ;
	wire _w11467_ ;
	wire _w11468_ ;
	wire _w11469_ ;
	wire _w11470_ ;
	wire _w11471_ ;
	wire _w11472_ ;
	wire _w11473_ ;
	wire _w11474_ ;
	wire _w11475_ ;
	wire _w11476_ ;
	wire _w11477_ ;
	wire _w11478_ ;
	wire _w11479_ ;
	wire _w11480_ ;
	wire _w11481_ ;
	wire _w11482_ ;
	wire _w11483_ ;
	wire _w11484_ ;
	wire _w11485_ ;
	wire _w11486_ ;
	wire _w11487_ ;
	wire _w11488_ ;
	wire _w11489_ ;
	wire _w11490_ ;
	wire _w11491_ ;
	wire _w11492_ ;
	wire _w11493_ ;
	wire _w11494_ ;
	wire _w11495_ ;
	wire _w11496_ ;
	wire _w11497_ ;
	wire _w11498_ ;
	wire _w11499_ ;
	wire _w11500_ ;
	wire _w11501_ ;
	wire _w11502_ ;
	wire _w11503_ ;
	wire _w11504_ ;
	wire _w11505_ ;
	wire _w11506_ ;
	wire _w11507_ ;
	wire _w11508_ ;
	wire _w11509_ ;
	wire _w11510_ ;
	wire _w11511_ ;
	wire _w11512_ ;
	wire _w11513_ ;
	wire _w11514_ ;
	wire _w11515_ ;
	wire _w11516_ ;
	wire _w11517_ ;
	wire _w11518_ ;
	wire _w11519_ ;
	wire _w11520_ ;
	wire _w11521_ ;
	wire _w11522_ ;
	wire _w11523_ ;
	wire _w11524_ ;
	wire _w11525_ ;
	wire _w11526_ ;
	wire _w11527_ ;
	wire _w11528_ ;
	wire _w11529_ ;
	wire _w11530_ ;
	wire _w11531_ ;
	wire _w11532_ ;
	wire _w11533_ ;
	wire _w11534_ ;
	wire _w11535_ ;
	wire _w11536_ ;
	wire _w11537_ ;
	wire _w11538_ ;
	wire _w11539_ ;
	wire _w11540_ ;
	wire _w11541_ ;
	wire _w11542_ ;
	wire _w11543_ ;
	wire _w11544_ ;
	wire _w11545_ ;
	wire _w11546_ ;
	wire _w11547_ ;
	wire _w11548_ ;
	wire _w11549_ ;
	wire _w11550_ ;
	wire _w11551_ ;
	wire _w11552_ ;
	wire _w11553_ ;
	wire _w11554_ ;
	wire _w11555_ ;
	wire _w11556_ ;
	wire _w11557_ ;
	wire _w11558_ ;
	wire _w11559_ ;
	wire _w11560_ ;
	wire _w11561_ ;
	wire _w11562_ ;
	wire _w11563_ ;
	wire _w11564_ ;
	wire _w11565_ ;
	wire _w11566_ ;
	wire _w11567_ ;
	wire _w11568_ ;
	wire _w11569_ ;
	wire _w11570_ ;
	wire _w11571_ ;
	wire _w11572_ ;
	wire _w11573_ ;
	wire _w11574_ ;
	wire _w11575_ ;
	wire _w11576_ ;
	wire _w11577_ ;
	wire _w11578_ ;
	wire _w11579_ ;
	wire _w11580_ ;
	wire _w11581_ ;
	wire _w11582_ ;
	wire _w11583_ ;
	wire _w11584_ ;
	wire _w11585_ ;
	wire _w11586_ ;
	wire _w11587_ ;
	wire _w11588_ ;
	wire _w11589_ ;
	wire _w11590_ ;
	wire _w11591_ ;
	wire _w11592_ ;
	wire _w11593_ ;
	wire _w11594_ ;
	wire _w11595_ ;
	wire _w11596_ ;
	wire _w11597_ ;
	wire _w11598_ ;
	wire _w11599_ ;
	wire _w11600_ ;
	wire _w11601_ ;
	wire _w11602_ ;
	wire _w11603_ ;
	wire _w11604_ ;
	wire _w11605_ ;
	wire _w11606_ ;
	wire _w11607_ ;
	wire _w11608_ ;
	wire _w11609_ ;
	wire _w11610_ ;
	wire _w11611_ ;
	wire _w11612_ ;
	wire _w11613_ ;
	wire _w11614_ ;
	wire _w11615_ ;
	wire _w11616_ ;
	wire _w11617_ ;
	wire _w11618_ ;
	wire _w11619_ ;
	wire _w11620_ ;
	wire _w11621_ ;
	wire _w11622_ ;
	wire _w11623_ ;
	wire _w11624_ ;
	wire _w11625_ ;
	wire _w11626_ ;
	wire _w11627_ ;
	wire _w11628_ ;
	wire _w11629_ ;
	wire _w11630_ ;
	wire _w11631_ ;
	wire _w11632_ ;
	wire _w11633_ ;
	wire _w11634_ ;
	wire _w11635_ ;
	wire _w11636_ ;
	wire _w11637_ ;
	wire _w11638_ ;
	wire _w11639_ ;
	wire _w11640_ ;
	wire _w11641_ ;
	wire _w11642_ ;
	wire _w11643_ ;
	wire _w11644_ ;
	wire _w11645_ ;
	wire _w11646_ ;
	wire _w11647_ ;
	wire _w11648_ ;
	wire _w11649_ ;
	wire _w11650_ ;
	wire _w11651_ ;
	wire _w11652_ ;
	wire _w11653_ ;
	wire _w11654_ ;
	wire _w11655_ ;
	wire _w11656_ ;
	wire _w11657_ ;
	wire _w11658_ ;
	wire _w11659_ ;
	wire _w11660_ ;
	wire _w11661_ ;
	wire _w11662_ ;
	wire _w11663_ ;
	wire _w11664_ ;
	wire _w11665_ ;
	wire _w11666_ ;
	wire _w11667_ ;
	wire _w11668_ ;
	wire _w11669_ ;
	wire _w11670_ ;
	wire _w11671_ ;
	wire _w11672_ ;
	wire _w11673_ ;
	wire _w11674_ ;
	wire _w11675_ ;
	wire _w11676_ ;
	wire _w11677_ ;
	wire _w11678_ ;
	wire _w11679_ ;
	wire _w11680_ ;
	wire _w11681_ ;
	wire _w11682_ ;
	wire _w11683_ ;
	wire _w11684_ ;
	wire _w11685_ ;
	wire _w11686_ ;
	wire _w11687_ ;
	wire _w11688_ ;
	wire _w11689_ ;
	wire _w11690_ ;
	wire _w11691_ ;
	wire _w11692_ ;
	wire _w11693_ ;
	wire _w11694_ ;
	wire _w11695_ ;
	wire _w11696_ ;
	wire _w11697_ ;
	wire _w11698_ ;
	wire _w11699_ ;
	wire _w11700_ ;
	wire _w11701_ ;
	wire _w11702_ ;
	wire _w11703_ ;
	wire _w11704_ ;
	wire _w11705_ ;
	wire _w11706_ ;
	wire _w11707_ ;
	wire _w11708_ ;
	wire _w11709_ ;
	wire _w11710_ ;
	wire _w11711_ ;
	wire _w11712_ ;
	wire _w11713_ ;
	wire _w11714_ ;
	wire _w11715_ ;
	wire _w11716_ ;
	wire _w11717_ ;
	wire _w11718_ ;
	wire _w11719_ ;
	wire _w11720_ ;
	wire _w11721_ ;
	wire _w11722_ ;
	wire _w11723_ ;
	wire _w11724_ ;
	wire _w11725_ ;
	wire _w11726_ ;
	wire _w11727_ ;
	wire _w11728_ ;
	wire _w11729_ ;
	wire _w11730_ ;
	wire _w11731_ ;
	wire _w11732_ ;
	wire _w11733_ ;
	wire _w11734_ ;
	wire _w11735_ ;
	wire _w11736_ ;
	wire _w11737_ ;
	wire _w11738_ ;
	wire _w11739_ ;
	wire _w11740_ ;
	wire _w11741_ ;
	wire _w11742_ ;
	wire _w11743_ ;
	wire _w11744_ ;
	wire _w11745_ ;
	wire _w11746_ ;
	wire _w11747_ ;
	wire _w11748_ ;
	wire _w11749_ ;
	wire _w11750_ ;
	wire _w11751_ ;
	wire _w11752_ ;
	wire _w11753_ ;
	wire _w11754_ ;
	wire _w11755_ ;
	wire _w11756_ ;
	wire _w11757_ ;
	wire _w11758_ ;
	wire _w11759_ ;
	wire _w11760_ ;
	wire _w11761_ ;
	wire _w11762_ ;
	wire _w11763_ ;
	wire _w11764_ ;
	wire _w11765_ ;
	wire _w11766_ ;
	wire _w11767_ ;
	wire _w11768_ ;
	wire _w11769_ ;
	wire _w11770_ ;
	wire _w11771_ ;
	wire _w11772_ ;
	wire _w11773_ ;
	wire _w11774_ ;
	wire _w11775_ ;
	wire _w11776_ ;
	wire _w11777_ ;
	wire _w11778_ ;
	wire _w11779_ ;
	wire _w11780_ ;
	wire _w11781_ ;
	wire _w11782_ ;
	wire _w11783_ ;
	wire _w11784_ ;
	wire _w11785_ ;
	wire _w11786_ ;
	wire _w11787_ ;
	wire _w11788_ ;
	wire _w11789_ ;
	wire _w11790_ ;
	wire _w11791_ ;
	wire _w11792_ ;
	wire _w11793_ ;
	wire _w11794_ ;
	wire _w11795_ ;
	wire _w11796_ ;
	wire _w11797_ ;
	wire _w11798_ ;
	wire _w11799_ ;
	wire _w11800_ ;
	wire _w11801_ ;
	wire _w11802_ ;
	wire _w11803_ ;
	wire _w11804_ ;
	wire _w11805_ ;
	wire _w11806_ ;
	wire _w11807_ ;
	wire _w11808_ ;
	wire _w11809_ ;
	wire _w11810_ ;
	wire _w11811_ ;
	wire _w11812_ ;
	wire _w11813_ ;
	wire _w11814_ ;
	wire _w11815_ ;
	wire _w11816_ ;
	wire _w11817_ ;
	wire _w11818_ ;
	wire _w11819_ ;
	wire _w11820_ ;
	wire _w11821_ ;
	wire _w11822_ ;
	wire _w11823_ ;
	wire _w11824_ ;
	wire _w11825_ ;
	wire _w11826_ ;
	wire _w11827_ ;
	wire _w11828_ ;
	wire _w11829_ ;
	wire _w11830_ ;
	wire _w11831_ ;
	wire _w11832_ ;
	wire _w11833_ ;
	wire _w11834_ ;
	wire _w11835_ ;
	wire _w11836_ ;
	wire _w11837_ ;
	wire _w11838_ ;
	wire _w11839_ ;
	wire _w11840_ ;
	wire _w11841_ ;
	wire _w11842_ ;
	wire _w11843_ ;
	wire _w11844_ ;
	wire _w11845_ ;
	wire _w11846_ ;
	wire _w11847_ ;
	wire _w11848_ ;
	wire _w11849_ ;
	wire _w11850_ ;
	wire _w11851_ ;
	wire _w11852_ ;
	wire _w11853_ ;
	wire _w11854_ ;
	wire _w11855_ ;
	wire _w11856_ ;
	wire _w11857_ ;
	wire _w11858_ ;
	wire _w11859_ ;
	wire _w11860_ ;
	wire _w11861_ ;
	wire _w11862_ ;
	wire _w11863_ ;
	wire _w11864_ ;
	wire _w11865_ ;
	wire _w11866_ ;
	wire _w11867_ ;
	wire _w11868_ ;
	wire _w11869_ ;
	wire _w11870_ ;
	wire _w11871_ ;
	wire _w11872_ ;
	wire _w11873_ ;
	wire _w11874_ ;
	wire _w11875_ ;
	wire _w11876_ ;
	wire _w11877_ ;
	wire _w11878_ ;
	wire _w11879_ ;
	wire _w11880_ ;
	wire _w11881_ ;
	wire _w11882_ ;
	wire _w11883_ ;
	wire _w11884_ ;
	wire _w11885_ ;
	wire _w11886_ ;
	wire _w11887_ ;
	wire _w11888_ ;
	wire _w11889_ ;
	wire _w11890_ ;
	wire _w11891_ ;
	wire _w11892_ ;
	wire _w11893_ ;
	wire _w11894_ ;
	wire _w11895_ ;
	wire _w11896_ ;
	wire _w11897_ ;
	wire _w11898_ ;
	wire _w11899_ ;
	wire _w11900_ ;
	wire _w11901_ ;
	wire _w11902_ ;
	wire _w11903_ ;
	wire _w11904_ ;
	wire _w11905_ ;
	wire _w11906_ ;
	wire _w11907_ ;
	wire _w11908_ ;
	wire _w11909_ ;
	wire _w11910_ ;
	wire _w11911_ ;
	wire _w11912_ ;
	wire _w11913_ ;
	wire _w11914_ ;
	wire _w11915_ ;
	wire _w11916_ ;
	wire _w11917_ ;
	wire _w11918_ ;
	wire _w11919_ ;
	wire _w11920_ ;
	wire _w11921_ ;
	wire _w11922_ ;
	wire _w11923_ ;
	wire _w11924_ ;
	wire _w11925_ ;
	wire _w11926_ ;
	wire _w11927_ ;
	wire _w11928_ ;
	wire _w11929_ ;
	wire _w11930_ ;
	wire _w11931_ ;
	wire _w11932_ ;
	wire _w11933_ ;
	wire _w11934_ ;
	wire _w11935_ ;
	wire _w11936_ ;
	wire _w11937_ ;
	wire _w11938_ ;
	wire _w11939_ ;
	wire _w11940_ ;
	wire _w11941_ ;
	wire _w11942_ ;
	wire _w11943_ ;
	wire _w11944_ ;
	wire _w11945_ ;
	wire _w11946_ ;
	wire _w11947_ ;
	wire _w11948_ ;
	wire _w11949_ ;
	wire _w11950_ ;
	wire _w11951_ ;
	wire _w11952_ ;
	wire _w11953_ ;
	wire _w11954_ ;
	wire _w11955_ ;
	wire _w11956_ ;
	wire _w11957_ ;
	wire _w11958_ ;
	wire _w11959_ ;
	wire _w11960_ ;
	wire _w11961_ ;
	wire _w11962_ ;
	wire _w11963_ ;
	wire _w11964_ ;
	wire _w11965_ ;
	wire _w11966_ ;
	wire _w11967_ ;
	wire _w11968_ ;
	wire _w11969_ ;
	wire _w11970_ ;
	wire _w11971_ ;
	wire _w11972_ ;
	wire _w11973_ ;
	wire _w11974_ ;
	wire _w11975_ ;
	wire _w11976_ ;
	wire _w11977_ ;
	wire _w11978_ ;
	wire _w11979_ ;
	wire _w11980_ ;
	wire _w11981_ ;
	wire _w11982_ ;
	wire _w11983_ ;
	wire _w11984_ ;
	wire _w11985_ ;
	wire _w11986_ ;
	wire _w11987_ ;
	wire _w11988_ ;
	wire _w11989_ ;
	wire _w11990_ ;
	wire _w11991_ ;
	wire _w11992_ ;
	wire _w11993_ ;
	wire _w11994_ ;
	wire _w11995_ ;
	wire _w11996_ ;
	wire _w11997_ ;
	wire _w11998_ ;
	wire _w11999_ ;
	wire _w12000_ ;
	wire _w12001_ ;
	wire _w12002_ ;
	wire _w12003_ ;
	wire _w12004_ ;
	wire _w12005_ ;
	wire _w12006_ ;
	wire _w12007_ ;
	wire _w12008_ ;
	wire _w12009_ ;
	wire _w12010_ ;
	wire _w12011_ ;
	wire _w12012_ ;
	wire _w12013_ ;
	wire _w12014_ ;
	wire _w12015_ ;
	wire _w12016_ ;
	wire _w12017_ ;
	wire _w12018_ ;
	wire _w12019_ ;
	wire _w12020_ ;
	wire _w12021_ ;
	wire _w12022_ ;
	wire _w12023_ ;
	wire _w12024_ ;
	wire _w12025_ ;
	wire _w12026_ ;
	wire _w12027_ ;
	wire _w12028_ ;
	wire _w12029_ ;
	wire _w12030_ ;
	wire _w12031_ ;
	wire _w12032_ ;
	wire _w12033_ ;
	wire _w12034_ ;
	wire _w12035_ ;
	wire _w12036_ ;
	wire _w12037_ ;
	wire _w12038_ ;
	wire _w12039_ ;
	wire _w12040_ ;
	wire _w12041_ ;
	wire _w12042_ ;
	wire _w12043_ ;
	wire _w12044_ ;
	wire _w12045_ ;
	wire _w12046_ ;
	wire _w12047_ ;
	wire _w12048_ ;
	wire _w12049_ ;
	wire _w12050_ ;
	wire _w12051_ ;
	wire _w12052_ ;
	wire _w12053_ ;
	wire _w12054_ ;
	wire _w12055_ ;
	wire _w12056_ ;
	wire _w12057_ ;
	wire _w12058_ ;
	wire _w12059_ ;
	wire _w12060_ ;
	wire _w12061_ ;
	wire _w12062_ ;
	wire _w12063_ ;
	wire _w12064_ ;
	wire _w12065_ ;
	wire _w12066_ ;
	wire _w12067_ ;
	wire _w12068_ ;
	wire _w12069_ ;
	wire _w12070_ ;
	wire _w12071_ ;
	wire _w12072_ ;
	wire _w12073_ ;
	wire _w12074_ ;
	wire _w12075_ ;
	wire _w12076_ ;
	wire _w12077_ ;
	wire _w12078_ ;
	wire _w12079_ ;
	wire _w12080_ ;
	wire _w12081_ ;
	wire _w12082_ ;
	wire _w12083_ ;
	wire _w12084_ ;
	wire _w12085_ ;
	wire _w12086_ ;
	wire _w12087_ ;
	wire _w12088_ ;
	wire _w12089_ ;
	wire _w12090_ ;
	wire _w12091_ ;
	wire _w12092_ ;
	wire _w12093_ ;
	wire _w12094_ ;
	wire _w12095_ ;
	wire _w12096_ ;
	wire _w12097_ ;
	wire _w12098_ ;
	wire _w12099_ ;
	wire _w12100_ ;
	wire _w12101_ ;
	wire _w12102_ ;
	wire _w12103_ ;
	wire _w12104_ ;
	wire _w12105_ ;
	wire _w12106_ ;
	wire _w12107_ ;
	wire _w12108_ ;
	wire _w12109_ ;
	wire _w12110_ ;
	wire _w12111_ ;
	wire _w12112_ ;
	wire _w12113_ ;
	wire _w12114_ ;
	wire _w12115_ ;
	wire _w12116_ ;
	wire _w12117_ ;
	wire _w12118_ ;
	wire _w12119_ ;
	wire _w12120_ ;
	wire _w12121_ ;
	wire _w12122_ ;
	wire _w12123_ ;
	wire _w12124_ ;
	wire _w12125_ ;
	wire _w12126_ ;
	wire _w12127_ ;
	wire _w12128_ ;
	wire _w12129_ ;
	wire _w12130_ ;
	wire _w12131_ ;
	wire _w12132_ ;
	wire _w12133_ ;
	wire _w12134_ ;
	wire _w12135_ ;
	wire _w12136_ ;
	wire _w12137_ ;
	wire _w12138_ ;
	wire _w12139_ ;
	wire _w12140_ ;
	wire _w12141_ ;
	wire _w12142_ ;
	wire _w12143_ ;
	wire _w12144_ ;
	wire _w12145_ ;
	wire _w12146_ ;
	wire _w12147_ ;
	wire _w12148_ ;
	wire _w12149_ ;
	wire _w12150_ ;
	wire _w12151_ ;
	wire _w12152_ ;
	wire _w12153_ ;
	wire _w12154_ ;
	wire _w12155_ ;
	wire _w12156_ ;
	wire _w12157_ ;
	wire _w12158_ ;
	wire _w12159_ ;
	wire _w12160_ ;
	wire _w12161_ ;
	wire _w12162_ ;
	wire _w12163_ ;
	wire _w12164_ ;
	wire _w12165_ ;
	wire _w12166_ ;
	wire _w12167_ ;
	wire _w12168_ ;
	wire _w12169_ ;
	wire _w12170_ ;
	wire _w12171_ ;
	wire _w12172_ ;
	wire _w12173_ ;
	wire _w12174_ ;
	wire _w12175_ ;
	wire _w12176_ ;
	wire _w12177_ ;
	wire _w12178_ ;
	wire _w12179_ ;
	wire _w12180_ ;
	wire _w12181_ ;
	wire _w12182_ ;
	wire _w12183_ ;
	wire _w12184_ ;
	wire _w12185_ ;
	wire _w12186_ ;
	wire _w12187_ ;
	wire _w12188_ ;
	wire _w12189_ ;
	wire _w12190_ ;
	wire _w12191_ ;
	wire _w12192_ ;
	wire _w12193_ ;
	wire _w12194_ ;
	wire _w12195_ ;
	wire _w12196_ ;
	wire _w12197_ ;
	wire _w12198_ ;
	wire _w12199_ ;
	wire _w12200_ ;
	wire _w12201_ ;
	wire _w12202_ ;
	wire _w12203_ ;
	wire _w12204_ ;
	wire _w12205_ ;
	wire _w12206_ ;
	wire _w12207_ ;
	wire _w12208_ ;
	wire _w12209_ ;
	wire _w12210_ ;
	wire _w12211_ ;
	wire _w12212_ ;
	wire _w12213_ ;
	wire _w12214_ ;
	wire _w12215_ ;
	wire _w12216_ ;
	wire _w12217_ ;
	wire _w12218_ ;
	wire _w12219_ ;
	wire _w12220_ ;
	wire _w12221_ ;
	wire _w12222_ ;
	wire _w12223_ ;
	wire _w12224_ ;
	wire _w12225_ ;
	wire _w12226_ ;
	wire _w12227_ ;
	wire _w12228_ ;
	wire _w12229_ ;
	wire _w12230_ ;
	wire _w12231_ ;
	wire _w12232_ ;
	wire _w12233_ ;
	wire _w12234_ ;
	wire _w12235_ ;
	wire _w12236_ ;
	wire _w12237_ ;
	wire _w12238_ ;
	wire _w12239_ ;
	wire _w12240_ ;
	wire _w12241_ ;
	wire _w12242_ ;
	wire _w12243_ ;
	wire _w12244_ ;
	wire _w12245_ ;
	wire _w12246_ ;
	wire _w12247_ ;
	wire _w12248_ ;
	wire _w12249_ ;
	wire _w12250_ ;
	wire _w12251_ ;
	wire _w12252_ ;
	wire _w12253_ ;
	wire _w12254_ ;
	wire _w12255_ ;
	wire _w12256_ ;
	wire _w12257_ ;
	wire _w12258_ ;
	wire _w12259_ ;
	wire _w12260_ ;
	wire _w12261_ ;
	wire _w12262_ ;
	wire _w12263_ ;
	wire _w12264_ ;
	wire _w12265_ ;
	wire _w12266_ ;
	wire _w12267_ ;
	wire _w12268_ ;
	wire _w12269_ ;
	wire _w12270_ ;
	wire _w12271_ ;
	wire _w12272_ ;
	wire _w12273_ ;
	wire _w12274_ ;
	wire _w12275_ ;
	wire _w12276_ ;
	wire _w12277_ ;
	wire _w12278_ ;
	wire _w12279_ ;
	wire _w12280_ ;
	wire _w12281_ ;
	wire _w12282_ ;
	wire _w12283_ ;
	wire _w12284_ ;
	wire _w12285_ ;
	wire _w12286_ ;
	wire _w12287_ ;
	wire _w12288_ ;
	wire _w12289_ ;
	wire _w12290_ ;
	wire _w12291_ ;
	wire _w12292_ ;
	wire _w12293_ ;
	wire _w12294_ ;
	wire _w12295_ ;
	wire _w12296_ ;
	wire _w12297_ ;
	wire _w12298_ ;
	wire _w12299_ ;
	wire _w12300_ ;
	wire _w12301_ ;
	wire _w12302_ ;
	wire _w12303_ ;
	wire _w12304_ ;
	wire _w12305_ ;
	wire _w12306_ ;
	wire _w12307_ ;
	wire _w12308_ ;
	wire _w12309_ ;
	wire _w12310_ ;
	wire _w12311_ ;
	wire _w12312_ ;
	wire _w12313_ ;
	wire _w12314_ ;
	wire _w12315_ ;
	wire _w12316_ ;
	wire _w12317_ ;
	wire _w12318_ ;
	wire _w12319_ ;
	wire _w12320_ ;
	wire _w12321_ ;
	wire _w12322_ ;
	wire _w12323_ ;
	wire _w12324_ ;
	wire _w12325_ ;
	wire _w12326_ ;
	wire _w12327_ ;
	wire _w12328_ ;
	wire _w12329_ ;
	wire _w12330_ ;
	wire _w12331_ ;
	wire _w12332_ ;
	wire _w12333_ ;
	wire _w12334_ ;
	wire _w12335_ ;
	wire _w12336_ ;
	wire _w12337_ ;
	wire _w12338_ ;
	wire _w12339_ ;
	wire _w12340_ ;
	wire _w12341_ ;
	wire _w12342_ ;
	wire _w12343_ ;
	wire _w12344_ ;
	wire _w12345_ ;
	wire _w12346_ ;
	wire _w12347_ ;
	wire _w12348_ ;
	wire _w12349_ ;
	wire _w12350_ ;
	wire _w12351_ ;
	wire _w12352_ ;
	wire _w12353_ ;
	wire _w12354_ ;
	wire _w12355_ ;
	wire _w12356_ ;
	wire _w12357_ ;
	wire _w12358_ ;
	wire _w12359_ ;
	wire _w12360_ ;
	wire _w12361_ ;
	wire _w12362_ ;
	wire _w12363_ ;
	wire _w12364_ ;
	wire _w12365_ ;
	wire _w12366_ ;
	wire _w12367_ ;
	wire _w12368_ ;
	wire _w12369_ ;
	wire _w12370_ ;
	wire _w12371_ ;
	wire _w12372_ ;
	wire _w12373_ ;
	wire _w12374_ ;
	wire _w12375_ ;
	wire _w12376_ ;
	wire _w12377_ ;
	wire _w12378_ ;
	wire _w12379_ ;
	wire _w12380_ ;
	wire _w12381_ ;
	wire _w12382_ ;
	wire _w12383_ ;
	wire _w12384_ ;
	wire _w12385_ ;
	wire _w12386_ ;
	wire _w12387_ ;
	wire _w12388_ ;
	wire _w12389_ ;
	wire _w12390_ ;
	wire _w12391_ ;
	wire _w12392_ ;
	wire _w12393_ ;
	wire _w12394_ ;
	wire _w12395_ ;
	wire _w12396_ ;
	wire _w12397_ ;
	wire _w12398_ ;
	wire _w12399_ ;
	wire _w12400_ ;
	wire _w12401_ ;
	wire _w12402_ ;
	wire _w12403_ ;
	wire _w12404_ ;
	wire _w12405_ ;
	wire _w12406_ ;
	wire _w12407_ ;
	wire _w12408_ ;
	wire _w12409_ ;
	wire _w12410_ ;
	wire _w12411_ ;
	wire _w12412_ ;
	wire _w12413_ ;
	wire _w12414_ ;
	wire _w12415_ ;
	wire _w12416_ ;
	wire _w12417_ ;
	wire _w12418_ ;
	wire _w12419_ ;
	wire _w12420_ ;
	wire _w12421_ ;
	wire _w12422_ ;
	wire _w12423_ ;
	wire _w12424_ ;
	wire _w12425_ ;
	wire _w12426_ ;
	wire _w12427_ ;
	wire _w12428_ ;
	wire _w12429_ ;
	wire _w12430_ ;
	wire _w12431_ ;
	wire _w12432_ ;
	wire _w12433_ ;
	wire _w12434_ ;
	wire _w12435_ ;
	wire _w12436_ ;
	wire _w12437_ ;
	wire _w12438_ ;
	wire _w12439_ ;
	wire _w12440_ ;
	wire _w12441_ ;
	wire _w12442_ ;
	wire _w12443_ ;
	wire _w12444_ ;
	wire _w12445_ ;
	wire _w12446_ ;
	wire _w12447_ ;
	wire _w12448_ ;
	wire _w12449_ ;
	wire _w12450_ ;
	wire _w12451_ ;
	wire _w12452_ ;
	wire _w12453_ ;
	wire _w12454_ ;
	wire _w12455_ ;
	wire _w12456_ ;
	wire _w12457_ ;
	wire _w12458_ ;
	wire _w12459_ ;
	wire _w12460_ ;
	wire _w12461_ ;
	wire _w12462_ ;
	wire _w12463_ ;
	wire _w12464_ ;
	wire _w12465_ ;
	wire _w12466_ ;
	wire _w12467_ ;
	wire _w12468_ ;
	wire _w12469_ ;
	wire _w12470_ ;
	wire _w12471_ ;
	wire _w12472_ ;
	wire _w12473_ ;
	wire _w12474_ ;
	wire _w12475_ ;
	wire _w12476_ ;
	wire _w12477_ ;
	wire _w12478_ ;
	wire _w12479_ ;
	wire _w12480_ ;
	wire _w12481_ ;
	wire _w12482_ ;
	wire _w12483_ ;
	wire _w12484_ ;
	wire _w12485_ ;
	wire _w12486_ ;
	wire _w12487_ ;
	wire _w12488_ ;
	wire _w12489_ ;
	wire _w12490_ ;
	wire _w12491_ ;
	wire _w12492_ ;
	wire _w12493_ ;
	wire _w12494_ ;
	wire _w12495_ ;
	wire _w12496_ ;
	wire _w12497_ ;
	wire _w12498_ ;
	wire _w12499_ ;
	wire _w12500_ ;
	wire _w12501_ ;
	wire _w12502_ ;
	wire _w12503_ ;
	wire _w12504_ ;
	wire _w12505_ ;
	wire _w12506_ ;
	wire _w12507_ ;
	wire _w12508_ ;
	wire _w12509_ ;
	wire _w12510_ ;
	wire _w12511_ ;
	wire _w12512_ ;
	wire _w12513_ ;
	wire _w12514_ ;
	wire _w12515_ ;
	wire _w12516_ ;
	wire _w12517_ ;
	wire _w12518_ ;
	wire _w12519_ ;
	wire _w12520_ ;
	wire _w12521_ ;
	wire _w12522_ ;
	wire _w12523_ ;
	wire _w12524_ ;
	wire _w12525_ ;
	wire _w12526_ ;
	wire _w12527_ ;
	wire _w12528_ ;
	wire _w12529_ ;
	wire _w12530_ ;
	wire _w12531_ ;
	wire _w12532_ ;
	wire _w12533_ ;
	wire _w12534_ ;
	wire _w12535_ ;
	wire _w12536_ ;
	wire _w12537_ ;
	wire _w12538_ ;
	wire _w12539_ ;
	wire _w12540_ ;
	wire _w12541_ ;
	wire _w12542_ ;
	wire _w12543_ ;
	wire _w12544_ ;
	wire _w12545_ ;
	wire _w12546_ ;
	wire _w12547_ ;
	wire _w12548_ ;
	wire _w12549_ ;
	wire _w12550_ ;
	wire _w12551_ ;
	wire _w12552_ ;
	wire _w12553_ ;
	wire _w12554_ ;
	wire _w12555_ ;
	wire _w12556_ ;
	wire _w12557_ ;
	wire _w12558_ ;
	wire _w12559_ ;
	wire _w12560_ ;
	wire _w12561_ ;
	wire _w12562_ ;
	wire _w12563_ ;
	wire _w12564_ ;
	wire _w12565_ ;
	wire _w12566_ ;
	wire _w12567_ ;
	wire _w12568_ ;
	wire _w12569_ ;
	wire _w12570_ ;
	wire _w12571_ ;
	wire _w12572_ ;
	wire _w12573_ ;
	wire _w12574_ ;
	wire _w12575_ ;
	wire _w12576_ ;
	wire _w12577_ ;
	wire _w12578_ ;
	wire _w12579_ ;
	wire _w12580_ ;
	wire _w12581_ ;
	wire _w12582_ ;
	wire _w12583_ ;
	wire _w12584_ ;
	wire _w12585_ ;
	wire _w12586_ ;
	wire _w12587_ ;
	wire _w12588_ ;
	wire _w12589_ ;
	wire _w12590_ ;
	wire _w12591_ ;
	wire _w12592_ ;
	wire _w12593_ ;
	wire _w12594_ ;
	wire _w12595_ ;
	wire _w12596_ ;
	wire _w12597_ ;
	wire _w12598_ ;
	wire _w12599_ ;
	wire _w12600_ ;
	wire _w12601_ ;
	wire _w12602_ ;
	wire _w12603_ ;
	wire _w12604_ ;
	wire _w12605_ ;
	wire _w12606_ ;
	wire _w12607_ ;
	wire _w12608_ ;
	wire _w12609_ ;
	wire _w12610_ ;
	wire _w12611_ ;
	wire _w12612_ ;
	wire _w12613_ ;
	wire _w12614_ ;
	wire _w12615_ ;
	wire _w12616_ ;
	wire _w12617_ ;
	wire _w12618_ ;
	wire _w12619_ ;
	wire _w12620_ ;
	wire _w12621_ ;
	wire _w12622_ ;
	wire _w12623_ ;
	wire _w12624_ ;
	wire _w12625_ ;
	wire _w12626_ ;
	wire _w12627_ ;
	wire _w12628_ ;
	wire _w12629_ ;
	wire _w12630_ ;
	wire _w12631_ ;
	wire _w12632_ ;
	wire _w12633_ ;
	wire _w12634_ ;
	wire _w12635_ ;
	wire _w12636_ ;
	wire _w12637_ ;
	wire _w12638_ ;
	wire _w12639_ ;
	wire _w12640_ ;
	wire _w12641_ ;
	wire _w12642_ ;
	wire _w12643_ ;
	wire _w12644_ ;
	wire _w12645_ ;
	wire _w12646_ ;
	wire _w12647_ ;
	wire _w12648_ ;
	wire _w12649_ ;
	wire _w12650_ ;
	wire _w12651_ ;
	wire _w12652_ ;
	wire _w12653_ ;
	wire _w12654_ ;
	wire _w12655_ ;
	wire _w12656_ ;
	wire _w12657_ ;
	wire _w12658_ ;
	wire _w12659_ ;
	wire _w12660_ ;
	wire _w12661_ ;
	wire _w12662_ ;
	wire _w12663_ ;
	wire _w12664_ ;
	wire _w12665_ ;
	wire _w12666_ ;
	wire _w12667_ ;
	wire _w12668_ ;
	wire _w12669_ ;
	wire _w12670_ ;
	wire _w12671_ ;
	wire _w12672_ ;
	wire _w12673_ ;
	wire _w12674_ ;
	wire _w12675_ ;
	wire _w12676_ ;
	wire _w12677_ ;
	wire _w12678_ ;
	wire _w12679_ ;
	wire _w12680_ ;
	wire _w12681_ ;
	wire _w12682_ ;
	wire _w12683_ ;
	wire _w12684_ ;
	wire _w12685_ ;
	wire _w12686_ ;
	wire _w12687_ ;
	wire _w12688_ ;
	wire _w12689_ ;
	wire _w12690_ ;
	wire _w12691_ ;
	wire _w12692_ ;
	wire _w12693_ ;
	wire _w12694_ ;
	wire _w12695_ ;
	wire _w12696_ ;
	wire _w12697_ ;
	wire _w12698_ ;
	wire _w12699_ ;
	wire _w12700_ ;
	wire _w12701_ ;
	wire _w12702_ ;
	wire _w12703_ ;
	wire _w12704_ ;
	wire _w12705_ ;
	wire _w12706_ ;
	wire _w12707_ ;
	wire _w12708_ ;
	wire _w12709_ ;
	wire _w12710_ ;
	wire _w12711_ ;
	wire _w12712_ ;
	wire _w12713_ ;
	wire _w12714_ ;
	wire _w12715_ ;
	wire _w12716_ ;
	wire _w12717_ ;
	wire _w12718_ ;
	wire _w12719_ ;
	wire _w12720_ ;
	wire _w12721_ ;
	wire _w12722_ ;
	wire _w12723_ ;
	wire _w12724_ ;
	wire _w12725_ ;
	wire _w12726_ ;
	wire _w12727_ ;
	wire _w12728_ ;
	wire _w12729_ ;
	wire _w12730_ ;
	wire _w12731_ ;
	wire _w12732_ ;
	wire _w12733_ ;
	wire _w12734_ ;
	wire _w12735_ ;
	wire _w12736_ ;
	wire _w12737_ ;
	wire _w12738_ ;
	wire _w12739_ ;
	wire _w12740_ ;
	wire _w12741_ ;
	wire _w12742_ ;
	wire _w12743_ ;
	wire _w12744_ ;
	wire _w12745_ ;
	wire _w12746_ ;
	wire _w12747_ ;
	wire _w12748_ ;
	wire _w12749_ ;
	wire _w12750_ ;
	wire _w12751_ ;
	wire _w12752_ ;
	wire _w12753_ ;
	wire _w12754_ ;
	wire _w12755_ ;
	wire _w12756_ ;
	wire _w12757_ ;
	wire _w12758_ ;
	wire _w12759_ ;
	wire _w12760_ ;
	wire _w12761_ ;
	wire _w12762_ ;
	wire _w12763_ ;
	wire _w12764_ ;
	wire _w12765_ ;
	wire _w12766_ ;
	wire _w12767_ ;
	wire _w12768_ ;
	wire _w12769_ ;
	wire _w12770_ ;
	wire _w12771_ ;
	wire _w12772_ ;
	wire _w12773_ ;
	wire _w12774_ ;
	wire _w12775_ ;
	wire _w12776_ ;
	wire _w12777_ ;
	wire _w12778_ ;
	wire _w12779_ ;
	wire _w12780_ ;
	wire _w12781_ ;
	wire _w12782_ ;
	wire _w12783_ ;
	wire _w12784_ ;
	wire _w12785_ ;
	wire _w12786_ ;
	wire _w12787_ ;
	wire _w12788_ ;
	wire _w12789_ ;
	wire _w12790_ ;
	wire _w12791_ ;
	wire _w12792_ ;
	wire _w12793_ ;
	wire _w12794_ ;
	wire _w12795_ ;
	wire _w12796_ ;
	wire _w12797_ ;
	wire _w12798_ ;
	wire _w12799_ ;
	wire _w12800_ ;
	wire _w12801_ ;
	wire _w12802_ ;
	wire _w12803_ ;
	wire _w12804_ ;
	wire _w12805_ ;
	wire _w12806_ ;
	wire _w12807_ ;
	wire _w12808_ ;
	wire _w12809_ ;
	wire _w12810_ ;
	wire _w12811_ ;
	wire _w12812_ ;
	wire _w12813_ ;
	wire _w12814_ ;
	wire _w12815_ ;
	wire _w12816_ ;
	wire _w12817_ ;
	wire _w12818_ ;
	wire _w12819_ ;
	wire _w12820_ ;
	wire _w12821_ ;
	wire _w12822_ ;
	wire _w12823_ ;
	wire _w12824_ ;
	wire _w12825_ ;
	wire _w12826_ ;
	wire _w12827_ ;
	wire _w12828_ ;
	wire _w12829_ ;
	wire _w12830_ ;
	wire _w12831_ ;
	wire _w12832_ ;
	wire _w12833_ ;
	wire _w12834_ ;
	wire _w12835_ ;
	wire _w12836_ ;
	wire _w12837_ ;
	wire _w12838_ ;
	wire _w12839_ ;
	wire _w12840_ ;
	wire _w12841_ ;
	wire _w12842_ ;
	wire _w12843_ ;
	wire _w12844_ ;
	wire _w12845_ ;
	wire _w12846_ ;
	wire _w12847_ ;
	wire _w12848_ ;
	wire _w12849_ ;
	wire _w12850_ ;
	wire _w12851_ ;
	wire _w12852_ ;
	wire _w12853_ ;
	wire _w12854_ ;
	wire _w12855_ ;
	wire _w12856_ ;
	wire _w12857_ ;
	wire _w12858_ ;
	wire _w12859_ ;
	wire _w12860_ ;
	wire _w12861_ ;
	wire _w12862_ ;
	wire _w12863_ ;
	wire _w12864_ ;
	wire _w12865_ ;
	wire _w12866_ ;
	wire _w12867_ ;
	wire _w12868_ ;
	wire _w12869_ ;
	wire _w12870_ ;
	wire _w12871_ ;
	wire _w12872_ ;
	wire _w12873_ ;
	wire _w12874_ ;
	wire _w12875_ ;
	wire _w12876_ ;
	wire _w12877_ ;
	wire _w12878_ ;
	wire _w12879_ ;
	wire _w12880_ ;
	wire _w12881_ ;
	wire _w12882_ ;
	wire _w12883_ ;
	wire _w12884_ ;
	wire _w12885_ ;
	wire _w12886_ ;
	wire _w12887_ ;
	wire _w12888_ ;
	wire _w12889_ ;
	wire _w12890_ ;
	wire _w12891_ ;
	wire _w12892_ ;
	wire _w12893_ ;
	wire _w12894_ ;
	wire _w12895_ ;
	wire _w12896_ ;
	wire _w12897_ ;
	wire _w12898_ ;
	wire _w12899_ ;
	wire _w12900_ ;
	wire _w12901_ ;
	wire _w12902_ ;
	wire _w12903_ ;
	wire _w12904_ ;
	wire _w12905_ ;
	wire _w12906_ ;
	wire _w12907_ ;
	wire _w12908_ ;
	wire _w12909_ ;
	wire _w12910_ ;
	wire _w12911_ ;
	wire _w12912_ ;
	wire _w12913_ ;
	wire _w12914_ ;
	wire _w12915_ ;
	wire _w12916_ ;
	wire _w12917_ ;
	wire _w12918_ ;
	wire _w12919_ ;
	wire _w12920_ ;
	wire _w12921_ ;
	wire _w12922_ ;
	wire _w12923_ ;
	wire _w12924_ ;
	wire _w12925_ ;
	wire _w12926_ ;
	wire _w12927_ ;
	wire _w12928_ ;
	wire _w12929_ ;
	wire _w12930_ ;
	wire _w12931_ ;
	wire _w12932_ ;
	wire _w12933_ ;
	wire _w12934_ ;
	wire _w12935_ ;
	wire _w12936_ ;
	wire _w12937_ ;
	wire _w12938_ ;
	wire _w12939_ ;
	wire _w12940_ ;
	wire _w12941_ ;
	wire _w12942_ ;
	wire _w12943_ ;
	wire _w12944_ ;
	wire _w12945_ ;
	wire _w12946_ ;
	wire _w12947_ ;
	wire _w12948_ ;
	wire _w12949_ ;
	wire _w12950_ ;
	wire _w12951_ ;
	wire _w12952_ ;
	wire _w12953_ ;
	wire _w12954_ ;
	wire _w12955_ ;
	wire _w12956_ ;
	wire _w12957_ ;
	wire _w12958_ ;
	wire _w12959_ ;
	wire _w12960_ ;
	wire _w12961_ ;
	wire _w12962_ ;
	wire _w12963_ ;
	wire _w12964_ ;
	wire _w12965_ ;
	wire _w12966_ ;
	wire _w12967_ ;
	wire _w12968_ ;
	wire _w12969_ ;
	wire _w12970_ ;
	wire _w12971_ ;
	wire _w12972_ ;
	wire _w12973_ ;
	wire _w12974_ ;
	wire _w12975_ ;
	wire _w12976_ ;
	wire _w12977_ ;
	wire _w12978_ ;
	wire _w12979_ ;
	wire _w12980_ ;
	wire _w12981_ ;
	wire _w12982_ ;
	wire _w12983_ ;
	wire _w12984_ ;
	wire _w12985_ ;
	wire _w12986_ ;
	wire _w12987_ ;
	wire _w12988_ ;
	wire _w12989_ ;
	wire _w12990_ ;
	wire _w12991_ ;
	wire _w12992_ ;
	wire _w12993_ ;
	wire _w12994_ ;
	wire _w12995_ ;
	wire _w12996_ ;
	wire _w12997_ ;
	wire _w12998_ ;
	wire _w12999_ ;
	wire _w13000_ ;
	wire _w13001_ ;
	wire _w13002_ ;
	wire _w13003_ ;
	wire _w13004_ ;
	wire _w13005_ ;
	wire _w13006_ ;
	wire _w13007_ ;
	wire _w13008_ ;
	wire _w13009_ ;
	wire _w13010_ ;
	wire _w13011_ ;
	wire _w13012_ ;
	wire _w13013_ ;
	wire _w13014_ ;
	wire _w13015_ ;
	wire _w13016_ ;
	wire _w13017_ ;
	wire _w13018_ ;
	wire _w13019_ ;
	wire _w13020_ ;
	wire _w13021_ ;
	wire _w13022_ ;
	wire _w13023_ ;
	wire _w13024_ ;
	wire _w13025_ ;
	wire _w13026_ ;
	wire _w13027_ ;
	wire _w13028_ ;
	wire _w13029_ ;
	wire _w13030_ ;
	wire _w13031_ ;
	wire _w13032_ ;
	wire _w13033_ ;
	wire _w13034_ ;
	wire _w13035_ ;
	wire _w13036_ ;
	wire _w13037_ ;
	wire _w13038_ ;
	wire _w13039_ ;
	wire _w13040_ ;
	wire _w13041_ ;
	wire _w13042_ ;
	wire _w13043_ ;
	wire _w13044_ ;
	wire _w13045_ ;
	wire _w13046_ ;
	wire _w13047_ ;
	wire _w13048_ ;
	wire _w13049_ ;
	wire _w13050_ ;
	wire _w13051_ ;
	wire _w13052_ ;
	wire _w13053_ ;
	wire _w13054_ ;
	wire _w13055_ ;
	wire _w13056_ ;
	wire _w13057_ ;
	wire _w13058_ ;
	wire _w13059_ ;
	wire _w13060_ ;
	wire _w13061_ ;
	wire _w13062_ ;
	wire _w13063_ ;
	wire _w13064_ ;
	wire _w13065_ ;
	wire _w13066_ ;
	wire _w13067_ ;
	wire _w13068_ ;
	wire _w13069_ ;
	wire _w13070_ ;
	wire _w13071_ ;
	wire _w13072_ ;
	wire _w13073_ ;
	wire _w13074_ ;
	wire _w13075_ ;
	wire _w13076_ ;
	wire _w13077_ ;
	wire _w13078_ ;
	wire _w13079_ ;
	wire _w13080_ ;
	wire _w13081_ ;
	wire _w13082_ ;
	wire _w13083_ ;
	wire _w13084_ ;
	wire _w13085_ ;
	wire _w13086_ ;
	wire _w13087_ ;
	wire _w13088_ ;
	wire _w13089_ ;
	wire _w13090_ ;
	wire _w13091_ ;
	wire _w13092_ ;
	wire _w13093_ ;
	wire _w13094_ ;
	wire _w13095_ ;
	wire _w13096_ ;
	wire _w13097_ ;
	wire _w13098_ ;
	wire _w13099_ ;
	wire _w13100_ ;
	wire _w13101_ ;
	wire _w13102_ ;
	wire _w13103_ ;
	wire _w13104_ ;
	wire _w13105_ ;
	wire _w13106_ ;
	wire _w13107_ ;
	wire _w13108_ ;
	wire _w13109_ ;
	wire _w13110_ ;
	wire _w13111_ ;
	wire _w13112_ ;
	wire _w13113_ ;
	wire _w13114_ ;
	wire _w13115_ ;
	wire _w13116_ ;
	wire _w13117_ ;
	wire _w13118_ ;
	wire _w13119_ ;
	wire _w13120_ ;
	wire _w13121_ ;
	wire _w13122_ ;
	wire _w13123_ ;
	wire _w13124_ ;
	wire _w13125_ ;
	wire _w13126_ ;
	wire _w13127_ ;
	wire _w13128_ ;
	wire _w13129_ ;
	wire _w13130_ ;
	wire _w13131_ ;
	wire _w13132_ ;
	wire _w13133_ ;
	wire _w13134_ ;
	wire _w13135_ ;
	wire _w13136_ ;
	wire _w13137_ ;
	wire _w13138_ ;
	wire _w13139_ ;
	wire _w13140_ ;
	wire _w13141_ ;
	wire _w13142_ ;
	wire _w13143_ ;
	wire _w13144_ ;
	wire _w13145_ ;
	wire _w13146_ ;
	wire _w13147_ ;
	wire _w13148_ ;
	wire _w13149_ ;
	wire _w13150_ ;
	wire _w13151_ ;
	wire _w13152_ ;
	wire _w13153_ ;
	wire _w13154_ ;
	wire _w13155_ ;
	wire _w13156_ ;
	wire _w13157_ ;
	wire _w13158_ ;
	wire _w13159_ ;
	wire _w13160_ ;
	wire _w13161_ ;
	wire _w13162_ ;
	wire _w13163_ ;
	wire _w13164_ ;
	wire _w13165_ ;
	wire _w13166_ ;
	wire _w13167_ ;
	wire _w13168_ ;
	wire _w13169_ ;
	wire _w13170_ ;
	wire _w13171_ ;
	wire _w13172_ ;
	wire _w13173_ ;
	wire _w13174_ ;
	wire _w13175_ ;
	wire _w13176_ ;
	wire _w13177_ ;
	wire _w13178_ ;
	wire _w13179_ ;
	wire _w13180_ ;
	wire _w13181_ ;
	wire _w13182_ ;
	wire _w13183_ ;
	wire _w13184_ ;
	wire _w13185_ ;
	wire _w13186_ ;
	wire _w13187_ ;
	wire _w13188_ ;
	wire _w13189_ ;
	wire _w13190_ ;
	wire _w13191_ ;
	wire _w13192_ ;
	wire _w13193_ ;
	wire _w13194_ ;
	wire _w13195_ ;
	wire _w13196_ ;
	wire _w13197_ ;
	wire _w13198_ ;
	wire _w13199_ ;
	wire _w13200_ ;
	wire _w13201_ ;
	wire _w13202_ ;
	wire _w13203_ ;
	wire _w13204_ ;
	wire _w13205_ ;
	wire _w13206_ ;
	wire _w13207_ ;
	wire _w13208_ ;
	wire _w13209_ ;
	wire _w13210_ ;
	wire _w13211_ ;
	wire _w13212_ ;
	wire _w13213_ ;
	wire _w13214_ ;
	wire _w13215_ ;
	wire _w13216_ ;
	wire _w13217_ ;
	wire _w13218_ ;
	wire _w13219_ ;
	wire _w13220_ ;
	wire _w13221_ ;
	wire _w13222_ ;
	wire _w13223_ ;
	wire _w13225_ ;
	wire _w13226_ ;
	wire _w13227_ ;
	wire _w13228_ ;
	wire _w13229_ ;
	wire _w13230_ ;
	wire _w13231_ ;
	wire _w13232_ ;
	wire _w13233_ ;
	wire _w13234_ ;
	wire _w13235_ ;
	wire _w13236_ ;
	wire _w13237_ ;
	wire _w13238_ ;
	wire _w13239_ ;
	wire _w13240_ ;
	wire _w13241_ ;
	wire _w13242_ ;
	wire _w13243_ ;
	wire _w13244_ ;
	wire _w13245_ ;
	wire _w13246_ ;
	wire _w13247_ ;
	wire _w13248_ ;
	wire _w13249_ ;
	wire _w13250_ ;
	wire _w13251_ ;
	wire _w13252_ ;
	wire _w13253_ ;
	wire _w13254_ ;
	wire _w13255_ ;
	wire _w13256_ ;
	wire _w13257_ ;
	wire _w13258_ ;
	wire _w13259_ ;
	wire _w13260_ ;
	wire _w13261_ ;
	wire _w13262_ ;
	wire _w13263_ ;
	wire _w13264_ ;
	wire _w13265_ ;
	wire _w13266_ ;
	wire _w13267_ ;
	wire _w13268_ ;
	wire _w13269_ ;
	wire _w13270_ ;
	wire _w13271_ ;
	wire _w13272_ ;
	wire _w13273_ ;
	wire _w13274_ ;
	wire _w13275_ ;
	wire _w13276_ ;
	wire _w13277_ ;
	wire _w13278_ ;
	wire _w13279_ ;
	wire _w13280_ ;
	wire _w13281_ ;
	wire _w13282_ ;
	wire _w13283_ ;
	wire _w13284_ ;
	wire _w13285_ ;
	wire _w13286_ ;
	wire _w13287_ ;
	wire _w13288_ ;
	wire _w13289_ ;
	wire _w13290_ ;
	wire _w13291_ ;
	wire _w13292_ ;
	wire _w13293_ ;
	wire _w13294_ ;
	wire _w13295_ ;
	wire _w13296_ ;
	wire _w13297_ ;
	wire _w13298_ ;
	wire _w13299_ ;
	wire _w13300_ ;
	wire _w13301_ ;
	wire _w13302_ ;
	wire _w13303_ ;
	wire _w13304_ ;
	wire _w13305_ ;
	wire _w13306_ ;
	wire _w13307_ ;
	wire _w13308_ ;
	wire _w13309_ ;
	wire _w13310_ ;
	wire _w13311_ ;
	wire _w13312_ ;
	wire _w13313_ ;
	wire _w13314_ ;
	wire _w13315_ ;
	wire _w13316_ ;
	wire _w13317_ ;
	wire _w13318_ ;
	wire _w13319_ ;
	wire _w13320_ ;
	wire _w13321_ ;
	wire _w13322_ ;
	wire _w13323_ ;
	wire _w13324_ ;
	wire _w13325_ ;
	wire _w13326_ ;
	wire _w13327_ ;
	wire _w13328_ ;
	wire _w13329_ ;
	wire _w13330_ ;
	wire _w13331_ ;
	wire _w13332_ ;
	wire _w13333_ ;
	wire _w13334_ ;
	wire _w13335_ ;
	wire _w13336_ ;
	wire _w13337_ ;
	wire _w13338_ ;
	wire _w13339_ ;
	wire _w13340_ ;
	wire _w13341_ ;
	wire _w13342_ ;
	wire _w13343_ ;
	wire _w13344_ ;
	wire _w13345_ ;
	wire _w13346_ ;
	wire _w13347_ ;
	wire _w13348_ ;
	wire _w13349_ ;
	wire _w13350_ ;
	wire _w13351_ ;
	wire _w13352_ ;
	wire _w13353_ ;
	wire _w13354_ ;
	wire _w13355_ ;
	wire _w13356_ ;
	wire _w13357_ ;
	wire _w13358_ ;
	wire _w13359_ ;
	wire _w13360_ ;
	wire _w13361_ ;
	wire _w13362_ ;
	wire _w13363_ ;
	wire _w13364_ ;
	wire _w13365_ ;
	wire _w13366_ ;
	wire _w13367_ ;
	wire _w13368_ ;
	wire _w13369_ ;
	wire _w13370_ ;
	wire _w13371_ ;
	wire _w13372_ ;
	wire _w13373_ ;
	wire _w13374_ ;
	wire _w13375_ ;
	wire _w13376_ ;
	wire _w13377_ ;
	wire _w13378_ ;
	wire _w13379_ ;
	wire _w13380_ ;
	wire _w13381_ ;
	wire _w13382_ ;
	wire _w13383_ ;
	wire _w13384_ ;
	wire _w13385_ ;
	wire _w13386_ ;
	wire _w13387_ ;
	wire _w13388_ ;
	wire _w13389_ ;
	wire _w13390_ ;
	wire _w13391_ ;
	wire _w13392_ ;
	wire _w13393_ ;
	wire _w13394_ ;
	wire _w13395_ ;
	wire _w13396_ ;
	wire _w13397_ ;
	wire _w13398_ ;
	wire _w13399_ ;
	wire _w13400_ ;
	wire _w13401_ ;
	wire _w13402_ ;
	wire _w13403_ ;
	wire _w13404_ ;
	wire _w13405_ ;
	wire _w13406_ ;
	wire _w13407_ ;
	wire _w13408_ ;
	wire _w13409_ ;
	wire _w13410_ ;
	wire _w13411_ ;
	wire _w13412_ ;
	wire _w13413_ ;
	wire _w13414_ ;
	wire _w13415_ ;
	wire _w13416_ ;
	wire _w13417_ ;
	wire _w13418_ ;
	wire _w13419_ ;
	wire _w13420_ ;
	wire _w13421_ ;
	wire _w13422_ ;
	wire _w13423_ ;
	wire _w13424_ ;
	wire _w13425_ ;
	wire _w13426_ ;
	wire _w13427_ ;
	wire _w13428_ ;
	wire _w13429_ ;
	wire _w13430_ ;
	wire _w13431_ ;
	wire _w13432_ ;
	wire _w13433_ ;
	wire _w13434_ ;
	wire _w13435_ ;
	wire _w13436_ ;
	wire _w13437_ ;
	wire _w13438_ ;
	wire _w13439_ ;
	wire _w13440_ ;
	wire _w13441_ ;
	wire _w13442_ ;
	wire _w13443_ ;
	wire _w13444_ ;
	wire _w13445_ ;
	wire _w13446_ ;
	wire _w13447_ ;
	wire _w13448_ ;
	wire _w13449_ ;
	wire _w13450_ ;
	wire _w13451_ ;
	wire _w13452_ ;
	wire _w13453_ ;
	wire _w13454_ ;
	wire _w13455_ ;
	wire _w13456_ ;
	wire _w13457_ ;
	wire _w13458_ ;
	wire _w13459_ ;
	wire _w13460_ ;
	wire _w13461_ ;
	wire _w13462_ ;
	wire _w13463_ ;
	wire _w13464_ ;
	wire _w13465_ ;
	wire _w13466_ ;
	wire _w13467_ ;
	wire _w13468_ ;
	wire _w13469_ ;
	wire _w13470_ ;
	wire _w13471_ ;
	wire _w13472_ ;
	wire _w13473_ ;
	wire _w13474_ ;
	wire _w13475_ ;
	wire _w13476_ ;
	wire _w13477_ ;
	wire _w13478_ ;
	wire _w13479_ ;
	wire _w13480_ ;
	wire _w13481_ ;
	wire _w13482_ ;
	wire _w13483_ ;
	wire _w13484_ ;
	wire _w13485_ ;
	wire _w13486_ ;
	wire _w13487_ ;
	wire _w13488_ ;
	wire _w13489_ ;
	wire _w13490_ ;
	wire _w13491_ ;
	wire _w13492_ ;
	wire _w13493_ ;
	wire _w13494_ ;
	wire _w13495_ ;
	wire _w13496_ ;
	wire _w13497_ ;
	wire _w13498_ ;
	wire _w13499_ ;
	wire _w13500_ ;
	wire _w13501_ ;
	wire _w13502_ ;
	wire _w13503_ ;
	wire _w13504_ ;
	wire _w13505_ ;
	wire _w13506_ ;
	wire _w13507_ ;
	wire _w13508_ ;
	wire _w13509_ ;
	wire _w13510_ ;
	wire _w13511_ ;
	wire _w13512_ ;
	wire _w13513_ ;
	wire _w13514_ ;
	wire _w13515_ ;
	wire _w13516_ ;
	wire _w13517_ ;
	wire _w13518_ ;
	wire _w13519_ ;
	wire _w13520_ ;
	wire _w13521_ ;
	wire _w13522_ ;
	wire _w13523_ ;
	wire _w13524_ ;
	wire _w13525_ ;
	wire _w13526_ ;
	wire _w13527_ ;
	wire _w13528_ ;
	wire _w13529_ ;
	wire _w13530_ ;
	wire _w13531_ ;
	wire _w13532_ ;
	wire _w13533_ ;
	wire _w13534_ ;
	wire _w13535_ ;
	wire _w13536_ ;
	wire _w13537_ ;
	wire _w13538_ ;
	wire _w13539_ ;
	wire _w13540_ ;
	wire _w13541_ ;
	wire _w13542_ ;
	wire _w13543_ ;
	wire _w13544_ ;
	wire _w13545_ ;
	wire _w13546_ ;
	wire _w13547_ ;
	wire _w13548_ ;
	wire _w13549_ ;
	wire _w13550_ ;
	wire _w13551_ ;
	wire _w13552_ ;
	wire _w13553_ ;
	wire _w13554_ ;
	wire _w13555_ ;
	wire _w13556_ ;
	wire _w13557_ ;
	wire _w13558_ ;
	wire _w13559_ ;
	wire _w13560_ ;
	wire _w13561_ ;
	wire _w13562_ ;
	wire _w13563_ ;
	wire _w13564_ ;
	wire _w13565_ ;
	wire _w13566_ ;
	wire _w13567_ ;
	wire _w13568_ ;
	wire _w13569_ ;
	wire _w13570_ ;
	wire _w13571_ ;
	wire _w13572_ ;
	wire _w13573_ ;
	wire _w13574_ ;
	wire _w13575_ ;
	wire _w13576_ ;
	wire _w13577_ ;
	wire _w13578_ ;
	wire _w13579_ ;
	wire _w13580_ ;
	wire _w13581_ ;
	wire _w13582_ ;
	wire _w13583_ ;
	wire _w13584_ ;
	wire _w13585_ ;
	wire _w13586_ ;
	wire _w13587_ ;
	wire _w13588_ ;
	wire _w13589_ ;
	wire _w13590_ ;
	wire _w13591_ ;
	wire _w13592_ ;
	wire _w13593_ ;
	wire _w13594_ ;
	wire _w13595_ ;
	wire _w13596_ ;
	wire _w13597_ ;
	wire _w13598_ ;
	wire _w13599_ ;
	wire _w13600_ ;
	wire _w13601_ ;
	wire _w13602_ ;
	wire _w13603_ ;
	wire _w13604_ ;
	wire _w13605_ ;
	wire _w13606_ ;
	wire _w13607_ ;
	wire _w13608_ ;
	wire _w13609_ ;
	wire _w13610_ ;
	wire _w13611_ ;
	wire _w13612_ ;
	wire _w13613_ ;
	wire _w13614_ ;
	wire _w13615_ ;
	wire _w13616_ ;
	wire _w13617_ ;
	wire _w13618_ ;
	wire _w13619_ ;
	wire _w13620_ ;
	wire _w13621_ ;
	wire _w13622_ ;
	wire _w13623_ ;
	wire _w13624_ ;
	wire _w13625_ ;
	wire _w13626_ ;
	wire _w13627_ ;
	wire _w13628_ ;
	wire _w13629_ ;
	wire _w13630_ ;
	wire _w13631_ ;
	wire _w13632_ ;
	wire _w13633_ ;
	wire _w13634_ ;
	wire _w13635_ ;
	wire _w13636_ ;
	wire _w13637_ ;
	wire _w13638_ ;
	wire _w13639_ ;
	wire _w13640_ ;
	wire _w13641_ ;
	wire _w13642_ ;
	wire _w13643_ ;
	wire _w13644_ ;
	wire _w13645_ ;
	wire _w13646_ ;
	wire _w13647_ ;
	wire _w13648_ ;
	wire _w13649_ ;
	wire _w13650_ ;
	wire _w13651_ ;
	wire _w13652_ ;
	wire _w13653_ ;
	wire _w13654_ ;
	wire _w13655_ ;
	wire _w13656_ ;
	wire _w13657_ ;
	wire _w13658_ ;
	wire _w13659_ ;
	wire _w13660_ ;
	wire _w13661_ ;
	wire _w13662_ ;
	wire _w13663_ ;
	wire _w13664_ ;
	wire _w13665_ ;
	wire _w13666_ ;
	wire _w13667_ ;
	wire _w13668_ ;
	wire _w13669_ ;
	wire _w13670_ ;
	wire _w13671_ ;
	wire _w13672_ ;
	wire _w13673_ ;
	wire _w13674_ ;
	wire _w13675_ ;
	wire _w13676_ ;
	wire _w13677_ ;
	wire _w13678_ ;
	wire _w13679_ ;
	wire _w13680_ ;
	wire _w13681_ ;
	wire _w13682_ ;
	wire _w13683_ ;
	wire _w13684_ ;
	wire _w13685_ ;
	wire _w13686_ ;
	wire _w13687_ ;
	wire _w13688_ ;
	wire _w13689_ ;
	wire _w13690_ ;
	wire _w13691_ ;
	wire _w13692_ ;
	wire _w13693_ ;
	wire _w13694_ ;
	wire _w13695_ ;
	wire _w13696_ ;
	wire _w13697_ ;
	wire _w13698_ ;
	wire _w13699_ ;
	wire _w13700_ ;
	wire _w13701_ ;
	wire _w13702_ ;
	wire _w13703_ ;
	wire _w13704_ ;
	wire _w13705_ ;
	wire _w13706_ ;
	wire _w13707_ ;
	wire _w13708_ ;
	wire _w13709_ ;
	wire _w13710_ ;
	wire _w13711_ ;
	wire _w13712_ ;
	wire _w13713_ ;
	wire _w13714_ ;
	wire _w13715_ ;
	wire _w13716_ ;
	wire _w13717_ ;
	wire _w13718_ ;
	wire _w13719_ ;
	wire _w13720_ ;
	wire _w13721_ ;
	wire _w13722_ ;
	wire _w13723_ ;
	wire _w13724_ ;
	wire _w13725_ ;
	wire _w13726_ ;
	wire _w13727_ ;
	wire _w13728_ ;
	wire _w13729_ ;
	wire _w13730_ ;
	wire _w13731_ ;
	wire _w13732_ ;
	wire _w13733_ ;
	wire _w13734_ ;
	wire _w13735_ ;
	wire _w13736_ ;
	wire _w13737_ ;
	wire _w13738_ ;
	wire _w13739_ ;
	wire _w13740_ ;
	wire _w13741_ ;
	wire _w13742_ ;
	wire _w13743_ ;
	wire _w13744_ ;
	wire _w13745_ ;
	wire _w13746_ ;
	wire _w13747_ ;
	wire _w13748_ ;
	wire _w13749_ ;
	wire _w13750_ ;
	wire _w13751_ ;
	wire _w13752_ ;
	wire _w13753_ ;
	wire _w13754_ ;
	wire _w13755_ ;
	wire _w13756_ ;
	wire _w13757_ ;
	wire _w13758_ ;
	wire _w13759_ ;
	wire _w13760_ ;
	wire _w13761_ ;
	wire _w13762_ ;
	wire _w13763_ ;
	wire _w13764_ ;
	wire _w13765_ ;
	wire _w13766_ ;
	wire _w13767_ ;
	wire _w13768_ ;
	wire _w13769_ ;
	wire _w13770_ ;
	wire _w13771_ ;
	wire _w13772_ ;
	wire _w13773_ ;
	wire _w13774_ ;
	wire _w13775_ ;
	wire _w13776_ ;
	wire _w13777_ ;
	wire _w13778_ ;
	wire _w13779_ ;
	wire _w13780_ ;
	wire _w13781_ ;
	wire _w13782_ ;
	wire _w13783_ ;
	wire _w13784_ ;
	wire _w13785_ ;
	wire _w13786_ ;
	wire _w13787_ ;
	wire _w13788_ ;
	wire _w13789_ ;
	wire _w13790_ ;
	wire _w13791_ ;
	wire _w13792_ ;
	wire _w13793_ ;
	wire _w13794_ ;
	wire _w13795_ ;
	wire _w13796_ ;
	wire _w13797_ ;
	wire _w13798_ ;
	wire _w13799_ ;
	wire _w13800_ ;
	wire _w13801_ ;
	wire _w13802_ ;
	wire _w13803_ ;
	wire _w13804_ ;
	wire _w13805_ ;
	wire _w13806_ ;
	wire _w13807_ ;
	wire _w13808_ ;
	wire _w13809_ ;
	wire _w13810_ ;
	wire _w13811_ ;
	wire _w13812_ ;
	wire _w13813_ ;
	wire _w13814_ ;
	wire _w13815_ ;
	wire _w13816_ ;
	wire _w13817_ ;
	wire _w13818_ ;
	wire _w13819_ ;
	wire _w13820_ ;
	wire _w13821_ ;
	wire _w13822_ ;
	wire _w13823_ ;
	wire _w13824_ ;
	wire _w13825_ ;
	wire _w13826_ ;
	wire _w13827_ ;
	wire _w13828_ ;
	wire _w13829_ ;
	wire _w13830_ ;
	wire _w13831_ ;
	wire _w13832_ ;
	wire _w13833_ ;
	wire _w13834_ ;
	wire _w13835_ ;
	wire _w13836_ ;
	wire _w13837_ ;
	wire _w13838_ ;
	wire _w13839_ ;
	wire _w13840_ ;
	wire _w13841_ ;
	wire _w13842_ ;
	wire _w13843_ ;
	wire _w13844_ ;
	wire _w13845_ ;
	wire _w13846_ ;
	wire _w13847_ ;
	wire _w13848_ ;
	wire _w13849_ ;
	wire _w13850_ ;
	wire _w13851_ ;
	wire _w13852_ ;
	wire _w13853_ ;
	wire _w13854_ ;
	wire _w13855_ ;
	wire _w13856_ ;
	wire _w13857_ ;
	wire _w13858_ ;
	wire _w13859_ ;
	wire _w13860_ ;
	wire _w13861_ ;
	wire _w13862_ ;
	wire _w13863_ ;
	wire _w13864_ ;
	wire _w13865_ ;
	wire _w13866_ ;
	wire _w13867_ ;
	wire _w13868_ ;
	wire _w13869_ ;
	wire _w13870_ ;
	wire _w13871_ ;
	wire _w13872_ ;
	wire _w13873_ ;
	wire _w13874_ ;
	wire _w13875_ ;
	wire _w13876_ ;
	wire _w13877_ ;
	wire _w13878_ ;
	wire _w13879_ ;
	wire _w13880_ ;
	wire _w13881_ ;
	wire _w13882_ ;
	wire _w13883_ ;
	wire _w13884_ ;
	wire _w13885_ ;
	wire _w13886_ ;
	wire _w13887_ ;
	wire _w13888_ ;
	wire _w13889_ ;
	wire _w13890_ ;
	wire _w13891_ ;
	wire _w13892_ ;
	wire _w13893_ ;
	wire _w13894_ ;
	wire _w13895_ ;
	wire _w13896_ ;
	wire _w13897_ ;
	wire _w13898_ ;
	wire _w13899_ ;
	wire _w13900_ ;
	wire _w13901_ ;
	wire _w13902_ ;
	wire _w13903_ ;
	wire _w13904_ ;
	wire _w13905_ ;
	wire _w13906_ ;
	wire _w13907_ ;
	wire _w13908_ ;
	wire _w13909_ ;
	wire _w13910_ ;
	wire _w13911_ ;
	wire _w13912_ ;
	wire _w13913_ ;
	wire _w13914_ ;
	wire _w13915_ ;
	wire _w13916_ ;
	wire _w13917_ ;
	wire _w13918_ ;
	wire _w13919_ ;
	wire _w13920_ ;
	wire _w13921_ ;
	wire _w13922_ ;
	wire _w13923_ ;
	wire _w13924_ ;
	wire _w13925_ ;
	wire _w13926_ ;
	wire _w13927_ ;
	wire _w13928_ ;
	wire _w13929_ ;
	wire _w13930_ ;
	wire _w13931_ ;
	wire _w13932_ ;
	wire _w13933_ ;
	wire _w13934_ ;
	wire _w13935_ ;
	wire _w13936_ ;
	wire _w13937_ ;
	wire _w13938_ ;
	wire _w13939_ ;
	wire _w13940_ ;
	wire _w13941_ ;
	wire _w13942_ ;
	wire _w13943_ ;
	wire _w13944_ ;
	wire _w13945_ ;
	wire _w13946_ ;
	wire _w13947_ ;
	wire _w13948_ ;
	wire _w13949_ ;
	wire _w13950_ ;
	wire _w13951_ ;
	wire _w13952_ ;
	wire _w13953_ ;
	wire _w13954_ ;
	wire _w13955_ ;
	wire _w13956_ ;
	wire _w13957_ ;
	wire _w13958_ ;
	wire _w13959_ ;
	wire _w13960_ ;
	wire _w13961_ ;
	wire _w13962_ ;
	wire _w13963_ ;
	wire _w13964_ ;
	wire _w13965_ ;
	wire _w13966_ ;
	wire _w13967_ ;
	wire _w13968_ ;
	wire _w13969_ ;
	wire _w13970_ ;
	wire _w13971_ ;
	wire _w13972_ ;
	wire _w13973_ ;
	wire _w13974_ ;
	wire _w13975_ ;
	wire _w13976_ ;
	wire _w13977_ ;
	wire _w13978_ ;
	wire _w13979_ ;
	wire _w13980_ ;
	wire _w13981_ ;
	wire _w13982_ ;
	wire _w13983_ ;
	wire _w13984_ ;
	wire _w13985_ ;
	wire _w13986_ ;
	wire _w13987_ ;
	wire _w13988_ ;
	wire _w13989_ ;
	wire _w13990_ ;
	wire _w13991_ ;
	wire _w13992_ ;
	wire _w13993_ ;
	wire _w13994_ ;
	wire _w13995_ ;
	wire _w13996_ ;
	wire _w13997_ ;
	wire _w13998_ ;
	wire _w13999_ ;
	wire _w14000_ ;
	wire _w14001_ ;
	wire _w14002_ ;
	wire _w14003_ ;
	wire _w14004_ ;
	wire _w14005_ ;
	wire _w14006_ ;
	wire _w14007_ ;
	wire _w14008_ ;
	wire _w14009_ ;
	wire _w14010_ ;
	wire _w14011_ ;
	wire _w14012_ ;
	wire _w14013_ ;
	wire _w14014_ ;
	wire _w14015_ ;
	wire _w14016_ ;
	wire _w14017_ ;
	wire _w14018_ ;
	wire _w14019_ ;
	wire _w14020_ ;
	wire _w14021_ ;
	wire _w14022_ ;
	wire _w14023_ ;
	wire _w14024_ ;
	wire _w14025_ ;
	wire _w14026_ ;
	wire _w14027_ ;
	wire _w14028_ ;
	wire _w14029_ ;
	wire _w14030_ ;
	wire _w14031_ ;
	wire _w14032_ ;
	wire _w14033_ ;
	wire _w14034_ ;
	wire _w14035_ ;
	wire _w14036_ ;
	wire _w14037_ ;
	wire _w14038_ ;
	wire _w14039_ ;
	wire _w14040_ ;
	wire _w14041_ ;
	wire _w14042_ ;
	wire _w14043_ ;
	wire _w14044_ ;
	wire _w14045_ ;
	wire _w14046_ ;
	wire _w14047_ ;
	wire _w14048_ ;
	wire _w14049_ ;
	wire _w14050_ ;
	wire _w14051_ ;
	wire _w14052_ ;
	wire _w14053_ ;
	wire _w14054_ ;
	wire _w14055_ ;
	wire _w14056_ ;
	wire _w14057_ ;
	wire _w14058_ ;
	wire _w14059_ ;
	wire _w14060_ ;
	wire _w14061_ ;
	wire _w14062_ ;
	wire _w14063_ ;
	wire _w14064_ ;
	wire _w14065_ ;
	wire _w14066_ ;
	wire _w14067_ ;
	wire _w14068_ ;
	wire _w14069_ ;
	wire _w14070_ ;
	wire _w14071_ ;
	wire _w14072_ ;
	wire _w14073_ ;
	wire _w14074_ ;
	wire _w14075_ ;
	wire _w14076_ ;
	wire _w14077_ ;
	wire _w14078_ ;
	wire _w14079_ ;
	wire _w14080_ ;
	wire _w14081_ ;
	wire _w14082_ ;
	wire _w14083_ ;
	wire _w14084_ ;
	wire _w14085_ ;
	wire _w14086_ ;
	wire _w14087_ ;
	wire _w14088_ ;
	wire _w14089_ ;
	wire _w14090_ ;
	wire _w14091_ ;
	wire _w14092_ ;
	wire _w14093_ ;
	wire _w14094_ ;
	wire _w14095_ ;
	wire _w14096_ ;
	wire _w14097_ ;
	wire _w14098_ ;
	wire _w14099_ ;
	wire _w14100_ ;
	wire _w14101_ ;
	wire _w14102_ ;
	wire _w14103_ ;
	wire _w14104_ ;
	wire _w14105_ ;
	wire _w14106_ ;
	wire _w14107_ ;
	wire _w14108_ ;
	wire _w14109_ ;
	wire _w14110_ ;
	wire _w14111_ ;
	wire _w14112_ ;
	wire _w14113_ ;
	wire _w14114_ ;
	wire _w14115_ ;
	wire _w14116_ ;
	wire _w14117_ ;
	wire _w14118_ ;
	wire _w14119_ ;
	wire _w14120_ ;
	wire _w14121_ ;
	wire _w14122_ ;
	wire _w14123_ ;
	wire _w14124_ ;
	wire _w14125_ ;
	wire _w14126_ ;
	wire _w14127_ ;
	wire _w14128_ ;
	wire _w14129_ ;
	wire _w14130_ ;
	wire _w14131_ ;
	wire _w14132_ ;
	wire _w14133_ ;
	wire _w14134_ ;
	wire _w14135_ ;
	wire _w14136_ ;
	wire _w14137_ ;
	wire _w14138_ ;
	wire _w14139_ ;
	wire _w14140_ ;
	wire _w14141_ ;
	wire _w14142_ ;
	wire _w14143_ ;
	wire _w14144_ ;
	wire _w14145_ ;
	wire _w14146_ ;
	wire _w14147_ ;
	wire _w14148_ ;
	wire _w14149_ ;
	wire _w14150_ ;
	wire _w14151_ ;
	wire _w14152_ ;
	wire _w14153_ ;
	wire _w14154_ ;
	wire _w14155_ ;
	wire _w14156_ ;
	wire _w14157_ ;
	wire _w14158_ ;
	wire _w14159_ ;
	wire _w14160_ ;
	wire _w14161_ ;
	wire _w14162_ ;
	wire _w14163_ ;
	wire _w14164_ ;
	wire _w14165_ ;
	wire _w14166_ ;
	wire _w14167_ ;
	wire _w14168_ ;
	wire _w14169_ ;
	wire _w14170_ ;
	wire _w14171_ ;
	wire _w14172_ ;
	wire _w14173_ ;
	wire _w14174_ ;
	wire _w14175_ ;
	wire _w14176_ ;
	wire _w14177_ ;
	wire _w14178_ ;
	wire _w14179_ ;
	wire _w14180_ ;
	wire _w14181_ ;
	wire _w14182_ ;
	wire _w14183_ ;
	wire _w14184_ ;
	wire _w14185_ ;
	wire _w14186_ ;
	wire _w14187_ ;
	wire _w14188_ ;
	wire _w14189_ ;
	wire _w14190_ ;
	wire _w14191_ ;
	wire _w14192_ ;
	wire _w14193_ ;
	wire _w14194_ ;
	wire _w14195_ ;
	wire _w14196_ ;
	wire _w14197_ ;
	wire _w14198_ ;
	wire _w14199_ ;
	wire _w14200_ ;
	wire _w14201_ ;
	wire _w14202_ ;
	wire _w14203_ ;
	wire _w14204_ ;
	wire _w14205_ ;
	wire _w14206_ ;
	wire _w14207_ ;
	wire _w14208_ ;
	wire _w14209_ ;
	wire _w14210_ ;
	wire _w14211_ ;
	wire _w14212_ ;
	wire _w14213_ ;
	wire _w14214_ ;
	wire _w14215_ ;
	wire _w14216_ ;
	wire _w14217_ ;
	wire _w14218_ ;
	wire _w14219_ ;
	wire _w14220_ ;
	wire _w14221_ ;
	wire _w14222_ ;
	wire _w14223_ ;
	wire _w14224_ ;
	wire _w14225_ ;
	wire _w14226_ ;
	wire _w14227_ ;
	wire _w14228_ ;
	wire _w14229_ ;
	wire _w14230_ ;
	wire _w14231_ ;
	wire _w14232_ ;
	wire _w14233_ ;
	wire _w14234_ ;
	wire _w14235_ ;
	wire _w14236_ ;
	wire _w14237_ ;
	wire _w14238_ ;
	wire _w14239_ ;
	wire _w14240_ ;
	wire _w14241_ ;
	wire _w14242_ ;
	wire _w14243_ ;
	wire _w14244_ ;
	wire _w14245_ ;
	wire _w14246_ ;
	wire _w14247_ ;
	wire _w14248_ ;
	wire _w14249_ ;
	wire _w14250_ ;
	wire _w14251_ ;
	wire _w14252_ ;
	wire _w14253_ ;
	wire _w14254_ ;
	wire _w14255_ ;
	wire _w14256_ ;
	wire _w14257_ ;
	wire _w14258_ ;
	wire _w14259_ ;
	wire _w14260_ ;
	wire _w14261_ ;
	wire _w14262_ ;
	wire _w14263_ ;
	wire _w14264_ ;
	wire _w14265_ ;
	wire _w14266_ ;
	wire _w14267_ ;
	wire _w14268_ ;
	wire _w14269_ ;
	wire _w14270_ ;
	wire _w14271_ ;
	wire _w14272_ ;
	wire _w14273_ ;
	wire _w14274_ ;
	wire _w14275_ ;
	wire _w14276_ ;
	wire _w14277_ ;
	wire _w14278_ ;
	wire _w14279_ ;
	wire _w14280_ ;
	wire _w14281_ ;
	wire _w14282_ ;
	wire _w14283_ ;
	wire _w14284_ ;
	wire _w14285_ ;
	wire _w14286_ ;
	wire _w14287_ ;
	wire _w14288_ ;
	wire _w14289_ ;
	wire _w14290_ ;
	wire _w14291_ ;
	wire _w14292_ ;
	wire _w14293_ ;
	wire _w14294_ ;
	wire _w14295_ ;
	wire _w14296_ ;
	wire _w14297_ ;
	wire _w14298_ ;
	wire _w14299_ ;
	wire _w14300_ ;
	wire _w14301_ ;
	wire _w14302_ ;
	wire _w14303_ ;
	wire _w14304_ ;
	wire _w14305_ ;
	wire _w14306_ ;
	wire _w14307_ ;
	wire _w14308_ ;
	wire _w14309_ ;
	wire _w14310_ ;
	wire _w14311_ ;
	wire _w14312_ ;
	wire _w14313_ ;
	wire _w14314_ ;
	wire _w14315_ ;
	wire _w14316_ ;
	wire _w14317_ ;
	wire _w14318_ ;
	wire _w14319_ ;
	wire _w14320_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\T_IRQ0n_pad ,
		_w548_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\T_IRQ1n_pad ,
		_w550_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\T_IRQ2n_pad ,
		_w552_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\T_IRQE0n_pad ,
		_w554_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\T_IRQE1n_pad ,
		_w556_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\T_IRQL1n_pad ,
		_w558_
	);
	LUT1 #(
		.INIT('h1)
	) name6 (
		T_ISn_pad,
		_w560_
	);
	LUT1 #(
		.INIT('h1)
	) name7 (
		T_PWDn_pad,
		_w576_
	);
	LUT1 #(
		.INIT('h1)
	) name8 (
		\bdma_BM_cyc_reg/P0001 ,
		_w646_
	);
	LUT1 #(
		.INIT('h1)
	) name9 (
		\core_c_psq_MGNT_reg/NET0131 ,
		_w1137_
	);
	LUT1 #(
		.INIT('h1)
	) name10 (
		\emc_ECMcs_reg/NET0131 ,
		_w2951_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\clkc_CLKOUT_reg/NET0131 ,
		\clkc_ckr_reg_DO_reg[15]/NET0131 ,
		_w4059_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\bdma_BSreq_reg/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4060_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport1_rxctl_RSreq_reg/NET0131 ,
		_w4061_
	);
	LUT4 #(
		.INIT('haaab)
	) name14 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		\sport1_txctl_TSreq_reg/NET0131 ,
		_w4062_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		_w4061_,
		_w4062_,
		_w4063_
	);
	LUT4 #(
		.INIT('h0100)
	) name16 (
		\idma_DSreq_reg/NET0131 ,
		_w4060_,
		_w4061_,
		_w4062_,
		_w4064_
	);
	LUT3 #(
		.INIT('h1b)
	) name17 (
		\idma_IDMA_boot_reg/NET0131_reg_syn_10 ,
		\idma_IDMA_boot_reg/NET0131_reg_syn_2 ,
		\idma_IDMA_boot_reg/NET0131_reg_syn_8 ,
		_w4065_
	);
	LUT3 #(
		.INIT('h1b)
	) name18 (
		\bdma_BDMA_boot_reg/NET0131_reg_syn_10 ,
		\bdma_BDMA_boot_reg/NET0131_reg_syn_2 ,
		\bdma_BDMA_boot_reg/NET0131_reg_syn_8 ,
		_w4066_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w4065_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\bdma_BM_cyc_reg/P0001 ,
		\core_c_psq_ECYC_reg/P0001 ,
		_w4068_
	);
	LUT3 #(
		.INIT('h1b)
	) name21 (
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		_w4069_
	);
	LUT3 #(
		.INIT('he4)
	) name22 (
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		_w4070_
	);
	LUT4 #(
		.INIT('h028a)
	) name23 (
		\core_c_psq_PCS_reg[2]/NET0131 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		_w4071_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\core_c_psq_PCS_reg[15]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w4072_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w4071_,
		_w4072_,
		_w4073_
	);
	LUT2 #(
		.INIT('he)
	) name26 (
		_w4071_,
		_w4072_,
		_w4074_
	);
	LUT4 #(
		.INIT('h0001)
	) name27 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_IDLE_Eg_reg/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		\sice_HALT_E_reg/P0001 ,
		_w4075_
	);
	LUT4 #(
		.INIT('h5054)
	) name28 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[12]/NET0131 ,
		\memc_LDaST_Eg_reg/NET0131 ,
		_w4076_
	);
	LUT3 #(
		.INIT('h40)
	) name29 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w4075_,
		_w4076_,
		_w4077_
	);
	LUT3 #(
		.INIT('h10)
	) name30 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		\core_c_psq_MGNT_reg/NET0131 ,
		\core_c_psq_PCS_reg[11]/NET0131 ,
		_w4078_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\core_c_psq_PCS_reg[5]/NET0131 ,
		\core_c_psq_PCS_reg[6]/NET0131 ,
		_w4079_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w4078_,
		_w4079_,
		_w4080_
	);
	LUT4 #(
		.INIT('heee2)
	) name33 (
		\clkc_Awake_reg/NET0131 ,
		\clkc_STBY_reg/NET0131 ,
		\core_c_psq_TRAP_R_L_reg/NET0131 ,
		\sice_GOICE_syn_reg/P0001 ,
		_w4081_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\core_c_psq_PCS_reg[10]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w4082_
	);
	LUT3 #(
		.INIT('h07)
	) name35 (
		\core_c_psq_PCS_reg[4]/NET0131 ,
		_w4081_,
		_w4082_,
		_w4083_
	);
	LUT4 #(
		.INIT('h7500)
	) name36 (
		_w4069_,
		_w4077_,
		_w4080_,
		_w4083_,
		_w4084_
	);
	LUT4 #(
		.INIT('h8aff)
	) name37 (
		_w4069_,
		_w4077_,
		_w4080_,
		_w4083_,
		_w4085_
	);
	LUT2 #(
		.INIT('h7)
	) name38 (
		_w4073_,
		_w4084_,
		_w4086_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\auctl_STEAL_reg/NET0131 ,
		\clkc_STBY_reg/NET0131 ,
		_w4087_
	);
	LUT4 #(
		.INIT('h4000)
	) name40 (
		_w4068_,
		_w4073_,
		_w4084_,
		_w4087_,
		_w4088_
	);
	LUT3 #(
		.INIT('h15)
	) name41 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4089_
	);
	LUT3 #(
		.INIT('h10)
	) name42 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w4090_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sice_CMRW_reg/NET0131 ,
		_w4091_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w4090_,
		_w4091_,
		_w4092_
	);
	LUT3 #(
		.INIT('h15)
	) name45 (
		\core_c_dec_accCM_E_reg/NET0131 ,
		_w4090_,
		_w4091_,
		_w4093_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name46 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		\core_c_psq_SRST_reg/P0001 ,
		_w4065_,
		_w4066_,
		_w4094_
	);
	LUT4 #(
		.INIT('hf400)
	) name47 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[12]/NET0131 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4095_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\core_c_psq_PCS_reg[2]/NET0131 ,
		_w4096_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w4095_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('hb)
	) name50 (
		_w4094_,
		_w4097_,
		_w4098_
	);
	LUT3 #(
		.INIT('h0b)
	) name51 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[11]/NET0131 ,
		_w4099_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		\sice_HALT_E_reg/P0001 ,
		_w4100_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w4099_,
		_w4100_,
		_w4101_
	);
	LUT3 #(
		.INIT('h04)
	) name54 (
		_w4094_,
		_w4097_,
		_w4101_,
		_w4102_
	);
	LUT3 #(
		.INIT('hfb)
	) name55 (
		_w4094_,
		_w4097_,
		_w4101_,
		_w4103_
	);
	LUT3 #(
		.INIT('h40)
	) name56 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4104_
	);
	LUT3 #(
		.INIT('hbf)
	) name57 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4105_
	);
	LUT4 #(
		.INIT('h4000)
	) name58 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4102_,
		_w4106_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w4093_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w4089_,
		_w4107_,
		_w4108_
	);
	LUT3 #(
		.INIT('h01)
	) name61 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		_w4109_
	);
	LUT4 #(
		.INIT('h0100)
	) name62 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4110_
	);
	LUT3 #(
		.INIT('h80)
	) name63 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		_w4111_
	);
	LUT4 #(
		.INIT('h0080)
	) name64 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4112_
	);
	LUT4 #(
		.INIT('h135f)
	) name65 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001 ,
		_w4112_,
		_w4110_,
		_w4113_
	);
	LUT4 #(
		.INIT('h8000)
	) name66 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4114_
	);
	LUT4 #(
		.INIT('h0001)
	) name67 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4115_
	);
	LUT4 #(
		.INIT('h153f)
	) name68 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001 ,
		_w4114_,
		_w4115_,
		_w4116_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w4113_,
		_w4116_,
		_w4117_
	);
	LUT4 #(
		.INIT('h2000)
	) name70 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4118_
	);
	LUT4 #(
		.INIT('h0400)
	) name71 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4119_
	);
	LUT4 #(
		.INIT('h135f)
	) name72 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001 ,
		_w4119_,
		_w4118_,
		_w4120_
	);
	LUT4 #(
		.INIT('h0800)
	) name73 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4121_
	);
	LUT4 #(
		.INIT('h0004)
	) name74 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4122_
	);
	LUT4 #(
		.INIT('h135f)
	) name75 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001 ,
		_w4121_,
		_w4122_,
		_w4123_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w4120_,
		_w4123_,
		_w4124_
	);
	LUT4 #(
		.INIT('h4000)
	) name77 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4125_
	);
	LUT4 #(
		.INIT('h0010)
	) name78 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4126_
	);
	LUT4 #(
		.INIT('h153f)
	) name79 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001 ,
		_w4126_,
		_w4125_,
		_w4127_
	);
	LUT4 #(
		.INIT('h0002)
	) name80 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4128_
	);
	LUT4 #(
		.INIT('h0040)
	) name81 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4129_
	);
	LUT4 #(
		.INIT('h135f)
	) name82 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001 ,
		_w4128_,
		_w4129_,
		_w4130_
	);
	LUT4 #(
		.INIT('h0200)
	) name83 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4131_
	);
	LUT4 #(
		.INIT('h0020)
	) name84 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4132_
	);
	LUT4 #(
		.INIT('h135f)
	) name85 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001 ,
		_w4132_,
		_w4131_,
		_w4133_
	);
	LUT4 #(
		.INIT('h0008)
	) name86 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4134_
	);
	LUT4 #(
		.INIT('h1000)
	) name87 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4135_
	);
	LUT4 #(
		.INIT('h135f)
	) name88 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001 ,
		_w4135_,
		_w4134_,
		_w4136_
	);
	LUT4 #(
		.INIT('h8000)
	) name89 (
		_w4133_,
		_w4136_,
		_w4127_,
		_w4130_,
		_w4137_
	);
	LUT3 #(
		.INIT('h80)
	) name90 (
		_w4124_,
		_w4117_,
		_w4137_,
		_w4138_
	);
	LUT3 #(
		.INIT('h80)
	) name91 (
		\clkc_Cnt4096_reg/NET0131 ,
		\clkc_Cnt4096_s2_reg/NET0131 ,
		\sport0_regs_AUTO_a_reg[12]/NET0131 ,
		_w4139_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\bdma_RST_pin_reg/P0001 ,
		\sice_RCS_reg[1]/NET0131 ,
		_w4140_
	);
	LUT2 #(
		.INIT('he)
	) name93 (
		\bdma_RST_pin_reg/P0001 ,
		\sice_RCS_reg[1]/NET0131 ,
		_w4141_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w4139_,
		_w4140_,
		_w4142_
	);
	LUT2 #(
		.INIT('hb)
	) name95 (
		_w4139_,
		_w4140_,
		_w4143_
	);
	LUT3 #(
		.INIT('hef)
	) name96 (
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4139_,
		_w4140_,
		_w4144_
	);
	LUT4 #(
		.INIT('h0200)
	) name97 (
		\core_eu_ec_cun_MV_reg/P0000_reg_syn_2 ,
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4139_,
		_w4140_,
		_w4145_
	);
	LUT3 #(
		.INIT('h01)
	) name98 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001 ,
		_w4146_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001 ,
		_w4147_
	);
	LUT4 #(
		.INIT('h0001)
	) name100 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001 ,
		_w4148_
	);
	LUT3 #(
		.INIT('h80)
	) name101 (
		_w4147_,
		_w4146_,
		_w4148_,
		_w4149_
	);
	LUT3 #(
		.INIT('h80)
	) name102 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001 ,
		_w4150_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001 ,
		_w4151_
	);
	LUT4 #(
		.INIT('h8000)
	) name104 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001 ,
		_w4152_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name105 (
		\core_eu_ec_cun_updateMV_C_reg/P0001 ,
		_w4151_,
		_w4150_,
		_w4152_,
		_w4153_
	);
	LUT4 #(
		.INIT('h8c88)
	) name106 (
		\core_eu_ec_cun_MVi_pre_C_reg/P0001 ,
		_w4142_,
		_w4149_,
		_w4153_,
		_w4154_
	);
	LUT3 #(
		.INIT('h13)
	) name107 (
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4145_,
		_w4154_,
		_w4155_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[3]/P0001 ,
		_w4156_
	);
	LUT4 #(
		.INIT('h1000)
	) name109 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[2]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[3]/P0001 ,
		_w4157_
	);
	LUT4 #(
		.INIT('hec00)
	) name110 (
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4145_,
		_w4154_,
		_w4157_,
		_w4158_
	);
	LUT4 #(
		.INIT('h2000)
	) name111 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[2]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[3]/P0001 ,
		_w4159_
	);
	LUT4 #(
		.INIT('h1300)
	) name112 (
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4145_,
		_w4154_,
		_w4159_,
		_w4160_
	);
	LUT2 #(
		.INIT('h6)
	) name113 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w4161_
	);
	LUT4 #(
		.INIT('h09f0)
	) name114 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		_w4162_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\core_eu_ec_cun_COND_E_reg[2]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[3]/P0001 ,
		_w4163_
	);
	LUT3 #(
		.INIT('h60)
	) name116 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		_w4162_,
		_w4163_,
		_w4164_
	);
	LUT3 #(
		.INIT('h40)
	) name117 (
		\core_c_psq_CE_reg/NET0131 ,
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[2]/P0001 ,
		_w4165_
	);
	LUT3 #(
		.INIT('h15)
	) name118 (
		\core_eu_ec_cun_condOK_CE_reg/P0001 ,
		_w4156_,
		_w4165_,
		_w4166_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		_w4164_,
		_w4166_,
		_w4167_
	);
	LUT3 #(
		.INIT('h10)
	) name120 (
		_w4160_,
		_w4158_,
		_w4167_,
		_w4168_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		\core_c_dec_IDLE_Eg_reg/P0001 ,
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		_w4169_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\core_eu_ec_cun_TERM_E_reg[2]/P0001 ,
		\core_eu_ec_cun_TERM_E_reg[3]/P0001 ,
		_w4170_
	);
	LUT3 #(
		.INIT('h40)
	) name123 (
		\core_eu_ec_cun_TERM_E_reg[1]/P0001 ,
		\core_eu_ec_cun_TERM_E_reg[2]/P0001 ,
		\core_eu_ec_cun_TERM_E_reg[3]/P0001 ,
		_w4171_
	);
	LUT4 #(
		.INIT('h09f0)
	) name124 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		\core_eu_ec_cun_TERM_E_reg[1]/P0001 ,
		_w4172_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\core_eu_ec_cun_TERM_E_reg[2]/P0001 ,
		\core_eu_ec_cun_TERM_E_reg[3]/P0001 ,
		_w4173_
	);
	LUT3 #(
		.INIT('h90)
	) name126 (
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		_w4172_,
		_w4173_,
		_w4174_
	);
	LUT3 #(
		.INIT('h20)
	) name127 (
		\core_c_psq_CE_reg/NET0131 ,
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		\core_eu_ec_cun_TERM_E_reg[1]/P0001 ,
		_w4175_
	);
	LUT3 #(
		.INIT('h15)
	) name128 (
		\core_eu_ec_cun_termOK_CE_reg/P0001 ,
		_w4170_,
		_w4175_,
		_w4176_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w4174_,
		_w4176_,
		_w4177_
	);
	LUT4 #(
		.INIT('h9f00)
	) name130 (
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		_w4155_,
		_w4171_,
		_w4177_,
		_w4178_
	);
	LUT4 #(
		.INIT('h135f)
	) name131 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001 ,
		_w4112_,
		_w4110_,
		_w4179_
	);
	LUT4 #(
		.INIT('h153f)
	) name132 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001 ,
		_w4114_,
		_w4115_,
		_w4180_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w4179_,
		_w4180_,
		_w4181_
	);
	LUT4 #(
		.INIT('h135f)
	) name134 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001 ,
		_w4119_,
		_w4118_,
		_w4182_
	);
	LUT4 #(
		.INIT('h135f)
	) name135 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001 ,
		_w4128_,
		_w4134_,
		_w4183_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w4182_,
		_w4183_,
		_w4184_
	);
	LUT4 #(
		.INIT('h153f)
	) name137 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001 ,
		_w4126_,
		_w4125_,
		_w4185_
	);
	LUT4 #(
		.INIT('h135f)
	) name138 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001 ,
		_w4121_,
		_w4129_,
		_w4186_
	);
	LUT4 #(
		.INIT('h135f)
	) name139 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001 ,
		_w4132_,
		_w4131_,
		_w4187_
	);
	LUT4 #(
		.INIT('h135f)
	) name140 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001 ,
		_w4135_,
		_w4122_,
		_w4188_
	);
	LUT4 #(
		.INIT('h8000)
	) name141 (
		_w4187_,
		_w4188_,
		_w4185_,
		_w4186_,
		_w4189_
	);
	LUT3 #(
		.INIT('h80)
	) name142 (
		_w4184_,
		_w4181_,
		_w4189_,
		_w4190_
	);
	LUT4 #(
		.INIT('h8000)
	) name143 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w4184_,
		_w4181_,
		_w4189_,
		_w4191_
	);
	LUT4 #(
		.INIT('h153f)
	) name144 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001 ,
		_w4114_,
		_w4115_,
		_w4192_
	);
	LUT4 #(
		.INIT('h135f)
	) name145 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001 ,
		_w4112_,
		_w4110_,
		_w4193_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT4 #(
		.INIT('h135f)
	) name147 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001 ,
		_w4122_,
		_w4131_,
		_w4195_
	);
	LUT4 #(
		.INIT('h135f)
	) name148 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001 ,
		_w4119_,
		_w4118_,
		_w4196_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w4195_,
		_w4196_,
		_w4197_
	);
	LUT4 #(
		.INIT('h135f)
	) name150 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001 ,
		_w4132_,
		_w4129_,
		_w4198_
	);
	LUT4 #(
		.INIT('h135f)
	) name151 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001 ,
		_w4128_,
		_w4134_,
		_w4199_
	);
	LUT4 #(
		.INIT('h153f)
	) name152 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001 ,
		_w4135_,
		_w4121_,
		_w4200_
	);
	LUT4 #(
		.INIT('h153f)
	) name153 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001 ,
		_w4126_,
		_w4125_,
		_w4201_
	);
	LUT4 #(
		.INIT('h8000)
	) name154 (
		_w4200_,
		_w4201_,
		_w4198_,
		_w4199_,
		_w4202_
	);
	LUT3 #(
		.INIT('h80)
	) name155 (
		_w4197_,
		_w4194_,
		_w4202_,
		_w4203_
	);
	LUT4 #(
		.INIT('h1555)
	) name156 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w4197_,
		_w4194_,
		_w4202_,
		_w4204_
	);
	LUT4 #(
		.INIT('h135f)
	) name157 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001 ,
		_w4112_,
		_w4110_,
		_w4205_
	);
	LUT4 #(
		.INIT('h153f)
	) name158 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001 ,
		_w4114_,
		_w4115_,
		_w4206_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w4205_,
		_w4206_,
		_w4207_
	);
	LUT4 #(
		.INIT('h135f)
	) name160 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001 ,
		_w4119_,
		_w4118_,
		_w4208_
	);
	LUT4 #(
		.INIT('h135f)
	) name161 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001 ,
		_w4121_,
		_w4122_,
		_w4209_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		_w4208_,
		_w4209_,
		_w4210_
	);
	LUT4 #(
		.INIT('h153f)
	) name163 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001 ,
		_w4126_,
		_w4125_,
		_w4211_
	);
	LUT4 #(
		.INIT('h135f)
	) name164 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001 ,
		_w4128_,
		_w4129_,
		_w4212_
	);
	LUT4 #(
		.INIT('h135f)
	) name165 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001 ,
		_w4132_,
		_w4131_,
		_w4213_
	);
	LUT4 #(
		.INIT('h135f)
	) name166 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001 ,
		_w4135_,
		_w4134_,
		_w4214_
	);
	LUT4 #(
		.INIT('h8000)
	) name167 (
		_w4213_,
		_w4214_,
		_w4211_,
		_w4212_,
		_w4215_
	);
	LUT3 #(
		.INIT('h80)
	) name168 (
		_w4210_,
		_w4207_,
		_w4215_,
		_w4216_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name169 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		_w4210_,
		_w4207_,
		_w4215_,
		_w4217_
	);
	LUT3 #(
		.INIT('h10)
	) name170 (
		_w4191_,
		_w4204_,
		_w4217_,
		_w4218_
	);
	LUT4 #(
		.INIT('h135f)
	) name171 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001 ,
		_w4114_,
		_w4110_,
		_w4219_
	);
	LUT4 #(
		.INIT('h153f)
	) name172 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001 ,
		_w4112_,
		_w4115_,
		_w4220_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w4219_,
		_w4220_,
		_w4221_
	);
	LUT4 #(
		.INIT('h153f)
	) name174 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001 ,
		_w4128_,
		_w4125_,
		_w4222_
	);
	LUT4 #(
		.INIT('h135f)
	) name175 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001 ,
		_w4134_,
		_w4132_,
		_w4223_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w4222_,
		_w4223_,
		_w4224_
	);
	LUT4 #(
		.INIT('h135f)
	) name177 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001 ,
		_w4121_,
		_w4129_,
		_w4225_
	);
	LUT4 #(
		.INIT('h135f)
	) name178 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001 ,
		_w4126_,
		_w4131_,
		_w4226_
	);
	LUT4 #(
		.INIT('h135f)
	) name179 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001 ,
		_w4119_,
		_w4122_,
		_w4227_
	);
	LUT4 #(
		.INIT('h135f)
	) name180 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001 ,
		_w4135_,
		_w4118_,
		_w4228_
	);
	LUT4 #(
		.INIT('h8000)
	) name181 (
		_w4227_,
		_w4228_,
		_w4225_,
		_w4226_,
		_w4229_
	);
	LUT3 #(
		.INIT('h80)
	) name182 (
		_w4224_,
		_w4221_,
		_w4229_,
		_w4230_
	);
	LUT4 #(
		.INIT('h1555)
	) name183 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w4224_,
		_w4221_,
		_w4229_,
		_w4231_
	);
	LUT4 #(
		.INIT('h53ff)
	) name184 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4111_,
		_w4232_
	);
	LUT4 #(
		.INIT('h35ff)
	) name185 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4109_,
		_w4233_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w4232_,
		_w4233_,
		_w4234_
	);
	LUT4 #(
		.INIT('h153f)
	) name187 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001 ,
		_w4125_,
		_w4118_,
		_w4235_
	);
	LUT4 #(
		.INIT('h135f)
	) name188 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001 ,
		_w4129_,
		_w4131_,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w4235_,
		_w4236_,
		_w4237_
	);
	LUT4 #(
		.INIT('h135f)
	) name190 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001 ,
		_w4119_,
		_w4121_,
		_w4238_
	);
	LUT4 #(
		.INIT('h135f)
	) name191 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001 ,
		_w4122_,
		_w4132_,
		_w4239_
	);
	LUT4 #(
		.INIT('h153f)
	) name192 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001 ,
		_w4128_,
		_w4135_,
		_w4240_
	);
	LUT4 #(
		.INIT('h153f)
	) name193 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001 ,
		_w4126_,
		_w4134_,
		_w4241_
	);
	LUT4 #(
		.INIT('h8000)
	) name194 (
		_w4240_,
		_w4241_,
		_w4238_,
		_w4239_,
		_w4242_
	);
	LUT3 #(
		.INIT('h80)
	) name195 (
		_w4237_,
		_w4234_,
		_w4242_,
		_w4243_
	);
	LUT4 #(
		.INIT('h8000)
	) name196 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4237_,
		_w4234_,
		_w4242_,
		_w4244_
	);
	LUT4 #(
		.INIT('h135f)
	) name197 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001 ,
		_w4112_,
		_w4110_,
		_w4245_
	);
	LUT4 #(
		.INIT('h153f)
	) name198 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001 ,
		_w4114_,
		_w4115_,
		_w4246_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w4245_,
		_w4246_,
		_w4247_
	);
	LUT4 #(
		.INIT('h153f)
	) name200 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001 ,
		_w4128_,
		_w4125_,
		_w4248_
	);
	LUT4 #(
		.INIT('h135f)
	) name201 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001 ,
		_w4134_,
		_w4132_,
		_w4249_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		_w4248_,
		_w4249_,
		_w4250_
	);
	LUT4 #(
		.INIT('h135f)
	) name203 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001 ,
		_w4121_,
		_w4129_,
		_w4251_
	);
	LUT4 #(
		.INIT('h135f)
	) name204 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001 ,
		_w4126_,
		_w4131_,
		_w4252_
	);
	LUT4 #(
		.INIT('h135f)
	) name205 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001 ,
		_w4119_,
		_w4122_,
		_w4253_
	);
	LUT4 #(
		.INIT('h135f)
	) name206 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001 ,
		_w4135_,
		_w4118_,
		_w4254_
	);
	LUT4 #(
		.INIT('h8000)
	) name207 (
		_w4253_,
		_w4254_,
		_w4251_,
		_w4252_,
		_w4255_
	);
	LUT3 #(
		.INIT('h80)
	) name208 (
		_w4250_,
		_w4247_,
		_w4255_,
		_w4256_
	);
	LUT4 #(
		.INIT('h1555)
	) name209 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4250_,
		_w4247_,
		_w4255_,
		_w4257_
	);
	LUT4 #(
		.INIT('h135f)
	) name210 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001 ,
		_w4112_,
		_w4110_,
		_w4258_
	);
	LUT4 #(
		.INIT('h153f)
	) name211 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001 ,
		_w4114_,
		_w4115_,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w4258_,
		_w4259_,
		_w4260_
	);
	LUT4 #(
		.INIT('h135f)
	) name213 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001 ,
		_w4119_,
		_w4118_,
		_w4261_
	);
	LUT4 #(
		.INIT('h153f)
	) name214 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001 ,
		_w4128_,
		_w4125_,
		_w4262_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		_w4261_,
		_w4262_,
		_w4263_
	);
	LUT4 #(
		.INIT('h153f)
	) name216 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001 ,
		_w4126_,
		_w4134_,
		_w4264_
	);
	LUT4 #(
		.INIT('h135f)
	) name217 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001 ,
		_w4132_,
		_w4129_,
		_w4265_
	);
	LUT4 #(
		.INIT('h135f)
	) name218 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001 ,
		_w4121_,
		_w4131_,
		_w4266_
	);
	LUT4 #(
		.INIT('h135f)
	) name219 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001 ,
		_w4135_,
		_w4122_,
		_w4267_
	);
	LUT4 #(
		.INIT('h8000)
	) name220 (
		_w4266_,
		_w4267_,
		_w4264_,
		_w4265_,
		_w4268_
	);
	LUT3 #(
		.INIT('h80)
	) name221 (
		_w4263_,
		_w4260_,
		_w4268_,
		_w4269_
	);
	LUT4 #(
		.INIT('h1555)
	) name222 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4263_,
		_w4260_,
		_w4268_,
		_w4270_
	);
	LUT4 #(
		.INIT('h0001)
	) name223 (
		_w4231_,
		_w4244_,
		_w4257_,
		_w4270_,
		_w4271_
	);
	LUT4 #(
		.INIT('h53ff)
	) name224 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4111_,
		_w4272_
	);
	LUT4 #(
		.INIT('h35ff)
	) name225 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4109_,
		_w4273_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w4272_,
		_w4273_,
		_w4274_
	);
	LUT4 #(
		.INIT('h153f)
	) name227 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001 ,
		_w4125_,
		_w4118_,
		_w4275_
	);
	LUT4 #(
		.INIT('h135f)
	) name228 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001 ,
		_w4129_,
		_w4131_,
		_w4276_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w4275_,
		_w4276_,
		_w4277_
	);
	LUT4 #(
		.INIT('h135f)
	) name230 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001 ,
		_w4119_,
		_w4121_,
		_w4278_
	);
	LUT4 #(
		.INIT('h135f)
	) name231 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001 ,
		_w4122_,
		_w4132_,
		_w4279_
	);
	LUT4 #(
		.INIT('h153f)
	) name232 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001 ,
		_w4128_,
		_w4135_,
		_w4280_
	);
	LUT4 #(
		.INIT('h153f)
	) name233 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001 ,
		_w4126_,
		_w4134_,
		_w4281_
	);
	LUT4 #(
		.INIT('h8000)
	) name234 (
		_w4280_,
		_w4281_,
		_w4278_,
		_w4279_,
		_w4282_
	);
	LUT3 #(
		.INIT('h80)
	) name235 (
		_w4277_,
		_w4274_,
		_w4282_,
		_w4283_
	);
	LUT4 #(
		.INIT('h1555)
	) name236 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4277_,
		_w4274_,
		_w4282_,
		_w4284_
	);
	LUT4 #(
		.INIT('h8000)
	) name237 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4263_,
		_w4260_,
		_w4268_,
		_w4285_
	);
	LUT4 #(
		.INIT('h0006)
	) name238 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w4138_,
		_w4284_,
		_w4285_,
		_w4286_
	);
	LUT3 #(
		.INIT('h80)
	) name239 (
		_w4218_,
		_w4271_,
		_w4286_,
		_w4287_
	);
	LUT4 #(
		.INIT('h8000)
	) name240 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4277_,
		_w4274_,
		_w4282_,
		_w4288_
	);
	LUT4 #(
		.INIT('h8000)
	) name241 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w4197_,
		_w4194_,
		_w4202_,
		_w4289_
	);
	LUT4 #(
		.INIT('h53ff)
	) name242 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4111_,
		_w4290_
	);
	LUT4 #(
		.INIT('h35ff)
	) name243 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4109_,
		_w4291_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT4 #(
		.INIT('h153f)
	) name245 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001 ,
		_w4128_,
		_w4118_,
		_w4293_
	);
	LUT4 #(
		.INIT('h135f)
	) name246 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001 ,
		_w4119_,
		_w4121_,
		_w4294_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w4293_,
		_w4294_,
		_w4295_
	);
	LUT4 #(
		.INIT('h135f)
	) name248 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001 ,
		_w4126_,
		_w4131_,
		_w4296_
	);
	LUT4 #(
		.INIT('h135f)
	) name249 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001 ,
		_w4135_,
		_w4134_,
		_w4297_
	);
	LUT4 #(
		.INIT('h135f)
	) name250 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001 ,
		_w4125_,
		_w4129_,
		_w4298_
	);
	LUT4 #(
		.INIT('h135f)
	) name251 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001 ,
		_w4122_,
		_w4132_,
		_w4299_
	);
	LUT4 #(
		.INIT('h8000)
	) name252 (
		_w4298_,
		_w4299_,
		_w4296_,
		_w4297_,
		_w4300_
	);
	LUT3 #(
		.INIT('h80)
	) name253 (
		_w4295_,
		_w4292_,
		_w4300_,
		_w4301_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name254 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		_w4295_,
		_w4292_,
		_w4300_,
		_w4302_
	);
	LUT3 #(
		.INIT('h10)
	) name255 (
		_w4288_,
		_w4289_,
		_w4302_,
		_w4303_
	);
	LUT4 #(
		.INIT('h135f)
	) name256 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001 ,
		_w4114_,
		_w4110_,
		_w4304_
	);
	LUT4 #(
		.INIT('h153f)
	) name257 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001 ,
		_w4112_,
		_w4115_,
		_w4305_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w4304_,
		_w4305_,
		_w4306_
	);
	LUT4 #(
		.INIT('h135f)
	) name259 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001 ,
		_w4119_,
		_w4132_,
		_w4307_
	);
	LUT4 #(
		.INIT('h135f)
	) name260 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001 ,
		_w4121_,
		_w4129_,
		_w4308_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		_w4307_,
		_w4308_,
		_w4309_
	);
	LUT4 #(
		.INIT('h135f)
	) name262 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001 ,
		_w4135_,
		_w4134_,
		_w4310_
	);
	LUT4 #(
		.INIT('h153f)
	) name263 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001 ,
		_w4122_,
		_w4118_,
		_w4311_
	);
	LUT4 #(
		.INIT('h153f)
	) name264 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001 ,
		_w4128_,
		_w4125_,
		_w4312_
	);
	LUT4 #(
		.INIT('h135f)
	) name265 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001 ,
		_w4126_,
		_w4131_,
		_w4313_
	);
	LUT4 #(
		.INIT('h8000)
	) name266 (
		_w4312_,
		_w4313_,
		_w4310_,
		_w4311_,
		_w4314_
	);
	LUT3 #(
		.INIT('h80)
	) name267 (
		_w4309_,
		_w4306_,
		_w4314_,
		_w4315_
	);
	LUT4 #(
		.INIT('h9555)
	) name268 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w4309_,
		_w4306_,
		_w4314_,
		_w4316_
	);
	LUT4 #(
		.INIT('h53ff)
	) name269 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4111_,
		_w4317_
	);
	LUT4 #(
		.INIT('h35ff)
	) name270 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4109_,
		_w4318_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w4317_,
		_w4318_,
		_w4319_
	);
	LUT4 #(
		.INIT('h153f)
	) name272 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001 ,
		_w4125_,
		_w4118_,
		_w4320_
	);
	LUT4 #(
		.INIT('h135f)
	) name273 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001 ,
		_w4129_,
		_w4131_,
		_w4321_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w4320_,
		_w4321_,
		_w4322_
	);
	LUT4 #(
		.INIT('h135f)
	) name275 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001 ,
		_w4119_,
		_w4121_,
		_w4323_
	);
	LUT4 #(
		.INIT('h135f)
	) name276 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001 ,
		_w4122_,
		_w4132_,
		_w4324_
	);
	LUT4 #(
		.INIT('h153f)
	) name277 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001 ,
		_w4128_,
		_w4135_,
		_w4325_
	);
	LUT4 #(
		.INIT('h153f)
	) name278 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001 ,
		_w4126_,
		_w4134_,
		_w4326_
	);
	LUT4 #(
		.INIT('h8000)
	) name279 (
		_w4325_,
		_w4326_,
		_w4323_,
		_w4324_,
		_w4327_
	);
	LUT3 #(
		.INIT('h80)
	) name280 (
		_w4322_,
		_w4319_,
		_w4327_,
		_w4328_
	);
	LUT4 #(
		.INIT('h8000)
	) name281 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4322_,
		_w4319_,
		_w4327_,
		_w4329_
	);
	LUT4 #(
		.INIT('h8000)
	) name282 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4250_,
		_w4247_,
		_w4255_,
		_w4330_
	);
	LUT3 #(
		.INIT('h01)
	) name283 (
		_w4329_,
		_w4330_,
		_w4316_,
		_w4331_
	);
	LUT4 #(
		.INIT('h1555)
	) name284 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4322_,
		_w4319_,
		_w4327_,
		_w4332_
	);
	LUT4 #(
		.INIT('h8000)
	) name285 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w4224_,
		_w4221_,
		_w4229_,
		_w4333_
	);
	LUT4 #(
		.INIT('h135f)
	) name286 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001 ,
		_w4112_,
		_w4110_,
		_w4334_
	);
	LUT4 #(
		.INIT('h153f)
	) name287 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001 ,
		_w4114_,
		_w4115_,
		_w4335_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w4334_,
		_w4335_,
		_w4336_
	);
	LUT4 #(
		.INIT('h135f)
	) name289 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001 ,
		_w4119_,
		_w4125_,
		_w4337_
	);
	LUT4 #(
		.INIT('h135f)
	) name290 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001 ,
		_w4121_,
		_w4129_,
		_w4338_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w4337_,
		_w4338_,
		_w4339_
	);
	LUT4 #(
		.INIT('h135f)
	) name292 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001 ,
		_w4135_,
		_w4134_,
		_w4340_
	);
	LUT4 #(
		.INIT('h153f)
	) name293 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001 ,
		_w4122_,
		_w4118_,
		_w4341_
	);
	LUT4 #(
		.INIT('h135f)
	) name294 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001 ,
		_w4128_,
		_w4132_,
		_w4342_
	);
	LUT4 #(
		.INIT('h135f)
	) name295 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001 ,
		_w4126_,
		_w4131_,
		_w4343_
	);
	LUT4 #(
		.INIT('h8000)
	) name296 (
		_w4342_,
		_w4343_,
		_w4340_,
		_w4341_,
		_w4344_
	);
	LUT3 #(
		.INIT('h80)
	) name297 (
		_w4339_,
		_w4336_,
		_w4344_,
		_w4345_
	);
	LUT4 #(
		.INIT('h8000)
	) name298 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w4339_,
		_w4336_,
		_w4344_,
		_w4346_
	);
	LUT4 #(
		.INIT('h135f)
	) name299 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001 ,
		_w4112_,
		_w4110_,
		_w4347_
	);
	LUT4 #(
		.INIT('h153f)
	) name300 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001 ,
		_w4114_,
		_w4115_,
		_w4348_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w4347_,
		_w4348_,
		_w4349_
	);
	LUT4 #(
		.INIT('h153f)
	) name302 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001 ,
		_w4128_,
		_w4125_,
		_w4350_
	);
	LUT4 #(
		.INIT('h135f)
	) name303 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001 ,
		_w4134_,
		_w4132_,
		_w4351_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		_w4350_,
		_w4351_,
		_w4352_
	);
	LUT4 #(
		.INIT('h135f)
	) name305 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001 ,
		_w4121_,
		_w4129_,
		_w4353_
	);
	LUT4 #(
		.INIT('h135f)
	) name306 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001 ,
		_w4126_,
		_w4131_,
		_w4354_
	);
	LUT4 #(
		.INIT('h135f)
	) name307 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001 ,
		_w4119_,
		_w4122_,
		_w4355_
	);
	LUT4 #(
		.INIT('h135f)
	) name308 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001 ,
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001 ,
		_w4135_,
		_w4118_,
		_w4356_
	);
	LUT4 #(
		.INIT('h8000)
	) name309 (
		_w4355_,
		_w4356_,
		_w4353_,
		_w4354_,
		_w4357_
	);
	LUT3 #(
		.INIT('h80)
	) name310 (
		_w4352_,
		_w4349_,
		_w4357_,
		_w4358_
	);
	LUT4 #(
		.INIT('h8000)
	) name311 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w4352_,
		_w4349_,
		_w4357_,
		_w4359_
	);
	LUT4 #(
		.INIT('h0001)
	) name312 (
		_w4332_,
		_w4333_,
		_w4346_,
		_w4359_,
		_w4360_
	);
	LUT4 #(
		.INIT('h1555)
	) name313 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w4184_,
		_w4181_,
		_w4189_,
		_w4361_
	);
	LUT4 #(
		.INIT('h1555)
	) name314 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w4352_,
		_w4349_,
		_w4357_,
		_w4362_
	);
	LUT4 #(
		.INIT('h1555)
	) name315 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4237_,
		_w4234_,
		_w4242_,
		_w4363_
	);
	LUT4 #(
		.INIT('h1555)
	) name316 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w4339_,
		_w4336_,
		_w4344_,
		_w4364_
	);
	LUT4 #(
		.INIT('h0001)
	) name317 (
		_w4361_,
		_w4362_,
		_w4363_,
		_w4364_,
		_w4365_
	);
	LUT4 #(
		.INIT('h8000)
	) name318 (
		_w4360_,
		_w4365_,
		_w4303_,
		_w4331_,
		_w4366_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name319 (
		_w4169_,
		_w4178_,
		_w4287_,
		_w4366_,
		_w4367_
	);
	LUT2 #(
		.INIT('h2)
	) name320 (
		_w4168_,
		_w4367_,
		_w4368_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[13]/P0001 ,
		_w4369_
	);
	LUT4 #(
		.INIT('h1555)
	) name322 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4237_,
		_w4234_,
		_w4242_,
		_w4370_
	);
	LUT3 #(
		.INIT('h54)
	) name323 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4369_,
		_w4370_,
		_w4371_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[10]/P0001 ,
		_w4372_
	);
	LUT4 #(
		.INIT('h1555)
	) name325 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4250_,
		_w4247_,
		_w4255_,
		_w4373_
	);
	LUT3 #(
		.INIT('h02)
	) name326 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4372_,
		_w4373_,
		_w4374_
	);
	LUT4 #(
		.INIT('h1555)
	) name327 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4263_,
		_w4260_,
		_w4268_,
		_w4375_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[7]/P0001 ,
		_w4376_
	);
	LUT3 #(
		.INIT('h54)
	) name329 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4375_,
		_w4376_,
		_w4377_
	);
	LUT4 #(
		.INIT('h1555)
	) name330 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4322_,
		_w4319_,
		_w4327_,
		_w4378_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[5]/P0001 ,
		_w4379_
	);
	LUT3 #(
		.INIT('h54)
	) name332 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4378_,
		_w4379_,
		_w4380_
	);
	LUT4 #(
		.INIT('h0001)
	) name333 (
		_w4371_,
		_w4374_,
		_w4377_,
		_w4380_,
		_w4381_
	);
	LUT4 #(
		.INIT('h1555)
	) name334 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4277_,
		_w4274_,
		_w4282_,
		_w4382_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[3]/P0001 ,
		_w4383_
	);
	LUT3 #(
		.INIT('h54)
	) name336 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4382_,
		_w4383_,
		_w4384_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[0]/P0001 ,
		_w4385_
	);
	LUT4 #(
		.INIT('h1555)
	) name338 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4124_,
		_w4117_,
		_w4137_,
		_w4386_
	);
	LUT3 #(
		.INIT('h02)
	) name339 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w4385_,
		_w4386_,
		_w4387_
	);
	LUT3 #(
		.INIT('h02)
	) name340 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4375_,
		_w4376_,
		_w4388_
	);
	LUT3 #(
		.INIT('h02)
	) name341 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4369_,
		_w4370_,
		_w4389_
	);
	LUT4 #(
		.INIT('h0001)
	) name342 (
		_w4384_,
		_w4387_,
		_w4388_,
		_w4389_,
		_w4390_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[6]/P0001 ,
		_w4391_
	);
	LUT4 #(
		.INIT('h1555)
	) name344 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4295_,
		_w4292_,
		_w4300_,
		_w4392_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w4391_,
		_w4392_,
		_w4393_
	);
	LUT4 #(
		.INIT('h1555)
	) name346 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4309_,
		_w4306_,
		_w4314_,
		_w4394_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[11]/P0001 ,
		_w4395_
	);
	LUT3 #(
		.INIT('h54)
	) name348 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w4394_,
		_w4395_,
		_w4396_
	);
	LUT3 #(
		.INIT('h02)
	) name349 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4382_,
		_w4383_,
		_w4397_
	);
	LUT4 #(
		.INIT('h0006)
	) name350 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		_w4393_,
		_w4396_,
		_w4397_,
		_w4398_
	);
	LUT3 #(
		.INIT('h80)
	) name351 (
		_w4381_,
		_w4390_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[4]/P0001 ,
		_w4400_
	);
	LUT4 #(
		.INIT('h4000)
	) name353 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4197_,
		_w4194_,
		_w4202_,
		_w4401_
	);
	LUT3 #(
		.INIT('ha9)
	) name354 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w4400_,
		_w4401_,
		_w4402_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[2]/P0001 ,
		_w4403_
	);
	LUT4 #(
		.INIT('h4000)
	) name356 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4339_,
		_w4336_,
		_w4344_,
		_w4404_
	);
	LUT3 #(
		.INIT('ha9)
	) name357 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w4403_,
		_w4404_,
		_w4405_
	);
	LUT4 #(
		.INIT('h1555)
	) name358 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4352_,
		_w4349_,
		_w4357_,
		_w4406_
	);
	LUT2 #(
		.INIT('h8)
	) name359 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[1]/P0001 ,
		_w4407_
	);
	LUT3 #(
		.INIT('h56)
	) name360 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w4406_,
		_w4407_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[12]/P0001 ,
		_w4409_
	);
	LUT4 #(
		.INIT('h1555)
	) name362 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4210_,
		_w4207_,
		_w4215_,
		_w4410_
	);
	LUT3 #(
		.INIT('h56)
	) name363 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		_w4409_,
		_w4410_,
		_w4411_
	);
	LUT4 #(
		.INIT('h0001)
	) name364 (
		_w4402_,
		_w4405_,
		_w4408_,
		_w4411_,
		_w4412_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[9]/P0001 ,
		_w4413_
	);
	LUT4 #(
		.INIT('h1555)
	) name366 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4224_,
		_w4221_,
		_w4229_,
		_w4414_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w4413_,
		_w4414_,
		_w4415_
	);
	LUT3 #(
		.INIT('h54)
	) name368 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4372_,
		_w4373_,
		_w4416_
	);
	LUT3 #(
		.INIT('h02)
	) name369 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4378_,
		_w4379_,
		_w4417_
	);
	LUT4 #(
		.INIT('h0006)
	) name370 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w4415_,
		_w4416_,
		_w4417_,
		_w4418_
	);
	LUT3 #(
		.INIT('h54)
	) name371 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w4385_,
		_w4386_,
		_w4419_
	);
	LUT3 #(
		.INIT('h02)
	) name372 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w4394_,
		_w4395_,
		_w4420_
	);
	LUT4 #(
		.INIT('h1555)
	) name373 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4184_,
		_w4181_,
		_w4189_,
		_w4421_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[8]/P0001 ,
		_w4422_
	);
	LUT3 #(
		.INIT('ha9)
	) name375 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w4421_,
		_w4422_,
		_w4423_
	);
	LUT3 #(
		.INIT('h10)
	) name376 (
		_w4419_,
		_w4420_,
		_w4423_,
		_w4424_
	);
	LUT4 #(
		.INIT('h8000)
	) name377 (
		_w4178_,
		_w4418_,
		_w4424_,
		_w4412_,
		_w4425_
	);
	LUT4 #(
		.INIT('h3222)
	) name378 (
		\core_c_dec_Nseq_Ed_reg/P0001 ,
		_w4168_,
		_w4399_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		\core_c_dec_Nrti_Ed_reg/P0001 ,
		\core_c_dec_RTI_Ed_reg/P0001 ,
		_w4427_
	);
	LUT4 #(
		.INIT('h0233)
	) name380 (
		_w4169_,
		_w4368_,
		_w4426_,
		_w4427_,
		_w4428_
	);
	LUT4 #(
		.INIT('h1000)
	) name381 (
		\core_c_psq_SRST_reg/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4065_,
		_w4066_,
		_w4429_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name382 (
		\core_c_dec_Nseq_Ed_reg/P0001 ,
		_w4160_,
		_w4158_,
		_w4167_,
		_w4430_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		_w4429_,
		_w4430_,
		_w4431_
	);
	LUT3 #(
		.INIT('h40)
	) name384 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4428_,
		_w4431_,
		_w4432_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w4433_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4434_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4435_
	);
	LUT4 #(
		.INIT('hff35)
	) name388 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4436_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4437_
	);
	LUT2 #(
		.INIT('h4)
	) name390 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4438_
	);
	LUT4 #(
		.INIT('h35ff)
	) name391 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4439_
	);
	LUT3 #(
		.INIT('h95)
	) name392 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w4436_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('hff35)
	) name393 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4441_
	);
	LUT4 #(
		.INIT('h35ff)
	) name394 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4442_
	);
	LUT3 #(
		.INIT('h95)
	) name395 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4441_,
		_w4442_,
		_w4443_
	);
	LUT4 #(
		.INIT('hff35)
	) name396 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4444_
	);
	LUT4 #(
		.INIT('h35ff)
	) name397 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4445_
	);
	LUT3 #(
		.INIT('h95)
	) name398 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4444_,
		_w4445_,
		_w4446_
	);
	LUT4 #(
		.INIT('h35ff)
	) name399 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4447_
	);
	LUT4 #(
		.INIT('hff35)
	) name400 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4448_
	);
	LUT3 #(
		.INIT('h95)
	) name401 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w4447_,
		_w4448_,
		_w4449_
	);
	LUT4 #(
		.INIT('h0001)
	) name402 (
		_w4440_,
		_w4443_,
		_w4446_,
		_w4449_,
		_w4450_
	);
	LUT4 #(
		.INIT('hff35)
	) name403 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4451_
	);
	LUT4 #(
		.INIT('h35ff)
	) name404 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4452_
	);
	LUT4 #(
		.INIT('h1222)
	) name405 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[2]/NET0131 ,
		_w4451_,
		_w4452_,
		_w4453_
	);
	LUT4 #(
		.INIT('hff35)
	) name406 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4454_
	);
	LUT4 #(
		.INIT('h35ff)
	) name407 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4455_
	);
	LUT3 #(
		.INIT('h95)
	) name408 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w4454_,
		_w4455_,
		_w4456_
	);
	LUT4 #(
		.INIT('hff35)
	) name409 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4457_
	);
	LUT4 #(
		.INIT('h35ff)
	) name410 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4458_
	);
	LUT3 #(
		.INIT('h95)
	) name411 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w4457_,
		_w4458_,
		_w4459_
	);
	LUT3 #(
		.INIT('h10)
	) name412 (
		_w4456_,
		_w4459_,
		_w4453_,
		_w4460_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w4450_,
		_w4460_,
		_w4461_
	);
	LUT4 #(
		.INIT('hff35)
	) name414 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4462_
	);
	LUT4 #(
		.INIT('h35ff)
	) name415 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4463_
	);
	LUT3 #(
		.INIT('h95)
	) name416 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w4462_,
		_w4463_,
		_w4464_
	);
	LUT4 #(
		.INIT('hff35)
	) name417 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4465_
	);
	LUT4 #(
		.INIT('h35ff)
	) name418 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4466_
	);
	LUT3 #(
		.INIT('h95)
	) name419 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w4465_,
		_w4466_,
		_w4467_
	);
	LUT4 #(
		.INIT('h35ff)
	) name420 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4468_
	);
	LUT4 #(
		.INIT('hff35)
	) name421 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4469_
	);
	LUT3 #(
		.INIT('h95)
	) name422 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w4468_,
		_w4469_,
		_w4470_
	);
	LUT3 #(
		.INIT('h01)
	) name423 (
		_w4467_,
		_w4470_,
		_w4464_,
		_w4471_
	);
	LUT4 #(
		.INIT('hff35)
	) name424 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4472_
	);
	LUT4 #(
		.INIT('h35ff)
	) name425 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4473_
	);
	LUT3 #(
		.INIT('h95)
	) name426 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w4472_,
		_w4473_,
		_w4474_
	);
	LUT4 #(
		.INIT('hff35)
	) name427 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4475_
	);
	LUT4 #(
		.INIT('h35ff)
	) name428 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4476_
	);
	LUT3 #(
		.INIT('h95)
	) name429 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w4475_,
		_w4476_,
		_w4477_
	);
	LUT4 #(
		.INIT('hff35)
	) name430 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4478_
	);
	LUT4 #(
		.INIT('h35ff)
	) name431 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4479_
	);
	LUT3 #(
		.INIT('h95)
	) name432 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w4478_,
		_w4479_,
		_w4480_
	);
	LUT4 #(
		.INIT('h35ff)
	) name433 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4481_
	);
	LUT4 #(
		.INIT('hff35)
	) name434 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4482_
	);
	LUT3 #(
		.INIT('h95)
	) name435 (
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w4481_,
		_w4482_,
		_w4483_
	);
	LUT4 #(
		.INIT('h0001)
	) name436 (
		_w4474_,
		_w4477_,
		_w4480_,
		_w4483_,
		_w4484_
	);
	LUT4 #(
		.INIT('hff35)
	) name437 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4485_
	);
	LUT4 #(
		.INIT('h35ff)
	) name438 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4486_
	);
	LUT3 #(
		.INIT('h95)
	) name439 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w4485_,
		_w4486_,
		_w4487_
	);
	LUT4 #(
		.INIT('h35ff)
	) name440 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4488_
	);
	LUT4 #(
		.INIT('hff35)
	) name441 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4489_
	);
	LUT3 #(
		.INIT('h95)
	) name442 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w4488_,
		_w4489_,
		_w4490_
	);
	LUT4 #(
		.INIT('hff35)
	) name443 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4491_
	);
	LUT4 #(
		.INIT('h35ff)
	) name444 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4492_
	);
	LUT3 #(
		.INIT('h95)
	) name445 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w4491_,
		_w4492_,
		_w4493_
	);
	LUT4 #(
		.INIT('hff35)
	) name446 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4494_
	);
	LUT4 #(
		.INIT('h35ff)
	) name447 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4495_
	);
	LUT3 #(
		.INIT('h95)
	) name448 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w4494_,
		_w4495_,
		_w4496_
	);
	LUT4 #(
		.INIT('h0001)
	) name449 (
		_w4487_,
		_w4490_,
		_w4493_,
		_w4496_,
		_w4497_
	);
	LUT3 #(
		.INIT('h80)
	) name450 (
		_w4471_,
		_w4484_,
		_w4497_,
		_w4498_
	);
	LUT3 #(
		.INIT('h80)
	) name451 (
		_w4433_,
		_w4461_,
		_w4498_,
		_w4499_
	);
	LUT3 #(
		.INIT('h01)
	) name452 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4428_,
		_w4499_,
		_w4500_
	);
	LUT3 #(
		.INIT('h20)
	) name453 (
		_w4169_,
		_w4430_,
		_w4178_,
		_w4501_
	);
	LUT4 #(
		.INIT('hcc04)
	) name454 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4429_,
		_w4428_,
		_w4501_,
		_w4502_
	);
	LUT4 #(
		.INIT('h4544)
	) name455 (
		_w4138_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4503_
	);
	LUT3 #(
		.INIT('h13)
	) name456 (
		_w4169_,
		_w4430_,
		_w4178_,
		_w4504_
	);
	LUT4 #(
		.INIT('h1131)
	) name457 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w4169_,
		_w4430_,
		_w4505_
	);
	LUT4 #(
		.INIT('h80aa)
	) name458 (
		_w4429_,
		_w4428_,
		_w4504_,
		_w4505_,
		_w4506_
	);
	LUT3 #(
		.INIT('h02)
	) name459 (
		_w4169_,
		_w4430_,
		_w4178_,
		_w4507_
	);
	LUT4 #(
		.INIT('haaa2)
	) name460 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4169_,
		_w4430_,
		_w4178_,
		_w4508_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		_w4429_,
		_w4433_,
		_w4509_
	);
	LUT3 #(
		.INIT('h70)
	) name462 (
		_w4461_,
		_w4498_,
		_w4509_,
		_w4510_
	);
	LUT2 #(
		.INIT('h4)
	) name463 (
		_w4508_,
		_w4510_,
		_w4511_
	);
	LUT3 #(
		.INIT('h10)
	) name464 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w4428_,
		_w4511_,
		_w4512_
	);
	LUT3 #(
		.INIT('h80)
	) name465 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[0]/P0001 ,
		_w4429_,
		_w4513_
	);
	LUT4 #(
		.INIT('h070f)
	) name466 (
		_w4385_,
		_w4428_,
		_w4513_,
		_w4431_,
		_w4514_
	);
	LUT4 #(
		.INIT('h0b00)
	) name467 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		_w4506_,
		_w4512_,
		_w4514_,
		_w4515_
	);
	LUT4 #(
		.INIT('h4555)
	) name468 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4516_
	);
	LUT4 #(
		.INIT('h1000)
	) name469 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4517_
	);
	LUT4 #(
		.INIT('h888b)
	) name470 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w4093_,
		_w4516_,
		_w4517_,
		_w4518_
	);
	LUT4 #(
		.INIT('h0400)
	) name471 (
		\idma_DSreq_reg/NET0131 ,
		_w4060_,
		_w4061_,
		_w4062_,
		_w4519_
	);
	LUT3 #(
		.INIT('h20)
	) name472 (
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4520_
	);
	LUT4 #(
		.INIT('h0800)
	) name473 (
		\idma_DCTL_reg[0]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4521_
	);
	LUT3 #(
		.INIT('h07)
	) name474 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w4519_,
		_w4521_,
		_w4522_
	);
	LUT4 #(
		.INIT('h0015)
	) name475 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4522_,
		_w4523_
	);
	LUT4 #(
		.INIT('h00ef)
	) name476 (
		_w4089_,
		_w4107_,
		_w4518_,
		_w4523_,
		_w4524_
	);
	LUT4 #(
		.INIT('h8aff)
	) name477 (
		_w4108_,
		_w4503_,
		_w4515_,
		_w4524_,
		_w4525_
	);
	LUT4 #(
		.INIT('h4544)
	) name478 (
		_w4256_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4526_
	);
	LUT4 #(
		.INIT('h8000)
	) name479 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_EXA_reg[1]/P0001 ,
		\core_c_psq_EXA_reg[2]/P0001 ,
		\core_c_psq_EXA_reg[3]/P0001 ,
		_w4527_
	);
	LUT4 #(
		.INIT('h8000)
	) name480 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		\core_c_psq_EXA_reg[5]/P0001 ,
		\core_c_psq_EXA_reg[6]/P0001 ,
		_w4527_,
		_w4528_
	);
	LUT4 #(
		.INIT('h8000)
	) name481 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_EXA_reg[9]/P0001 ,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h6)
	) name482 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		_w4529_,
		_w4530_
	);
	LUT3 #(
		.INIT('h80)
	) name483 (
		_w4372_,
		_w4428_,
		_w4431_,
		_w4531_
	);
	LUT4 #(
		.INIT('h8000)
	) name484 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		\core_c_psq_IFA_reg[1]/P0001 ,
		\core_c_psq_IFA_reg[2]/P0001 ,
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w4532_
	);
	LUT4 #(
		.INIT('h8000)
	) name485 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		\core_c_psq_IFA_reg[5]/P0001 ,
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w4532_,
		_w4533_
	);
	LUT4 #(
		.INIT('h8000)
	) name486 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		\core_c_psq_IFA_reg[8]/P0001 ,
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w4533_,
		_w4534_
	);
	LUT2 #(
		.INIT('h6)
	) name487 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w4534_,
		_w4535_
	);
	LUT3 #(
		.INIT('h80)
	) name488 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[10]/P0001 ,
		_w4429_,
		_w4536_
	);
	LUT4 #(
		.INIT('h00bf)
	) name489 (
		_w4428_,
		_w4511_,
		_w4535_,
		_w4536_,
		_w4537_
	);
	LUT4 #(
		.INIT('h0700)
	) name490 (
		_w4506_,
		_w4530_,
		_w4531_,
		_w4537_,
		_w4538_
	);
	LUT4 #(
		.INIT('h4555)
	) name491 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4539_
	);
	LUT4 #(
		.INIT('h1000)
	) name492 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4540_
	);
	LUT4 #(
		.INIT('h888b)
	) name493 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w4093_,
		_w4539_,
		_w4540_,
		_w4541_
	);
	LUT4 #(
		.INIT('h0800)
	) name494 (
		\idma_DCTL_reg[10]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4542_
	);
	LUT3 #(
		.INIT('h07)
	) name495 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w4519_,
		_w4542_,
		_w4543_
	);
	LUT4 #(
		.INIT('h0015)
	) name496 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4543_,
		_w4544_
	);
	LUT4 #(
		.INIT('h00ef)
	) name497 (
		_w4089_,
		_w4107_,
		_w4541_,
		_w4544_,
		_w4545_
	);
	LUT4 #(
		.INIT('h8aff)
	) name498 (
		_w4108_,
		_w4526_,
		_w4538_,
		_w4545_,
		_w4546_
	);
	LUT4 #(
		.INIT('h4544)
	) name499 (
		_w4315_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4547_
	);
	LUT3 #(
		.INIT('h6c)
	) name500 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_EXA_reg[11]/P0001 ,
		_w4529_,
		_w4548_
	);
	LUT3 #(
		.INIT('h80)
	) name501 (
		_w4395_,
		_w4428_,
		_w4431_,
		_w4549_
	);
	LUT3 #(
		.INIT('h6c)
	) name502 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w4534_,
		_w4550_
	);
	LUT3 #(
		.INIT('h80)
	) name503 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[11]/P0001 ,
		_w4429_,
		_w4551_
	);
	LUT4 #(
		.INIT('h00bf)
	) name504 (
		_w4428_,
		_w4511_,
		_w4550_,
		_w4551_,
		_w4552_
	);
	LUT4 #(
		.INIT('h0700)
	) name505 (
		_w4506_,
		_w4548_,
		_w4549_,
		_w4552_,
		_w4553_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name506 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4554_
	);
	LUT4 #(
		.INIT('h2000)
	) name507 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4555_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name508 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w4093_,
		_w4555_,
		_w4554_,
		_w4556_
	);
	LUT4 #(
		.INIT('h0800)
	) name509 (
		\idma_DCTL_reg[11]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4557_
	);
	LUT3 #(
		.INIT('h07)
	) name510 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w4519_,
		_w4557_,
		_w4558_
	);
	LUT4 #(
		.INIT('h0015)
	) name511 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4558_,
		_w4559_
	);
	LUT4 #(
		.INIT('h00ef)
	) name512 (
		_w4089_,
		_w4107_,
		_w4556_,
		_w4559_,
		_w4560_
	);
	LUT4 #(
		.INIT('h8aff)
	) name513 (
		_w4108_,
		_w4547_,
		_w4553_,
		_w4560_,
		_w4561_
	);
	LUT4 #(
		.INIT('h4544)
	) name514 (
		_w4358_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4562_
	);
	LUT2 #(
		.INIT('h6)
	) name515 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_EXA_reg[1]/P0001 ,
		_w4563_
	);
	LUT2 #(
		.INIT('h6)
	) name516 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w4564_
	);
	LUT3 #(
		.INIT('h40)
	) name517 (
		_w4428_,
		_w4511_,
		_w4564_,
		_w4565_
	);
	LUT3 #(
		.INIT('h80)
	) name518 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[1]/P0001 ,
		_w4429_,
		_w4566_
	);
	LUT4 #(
		.INIT('h007f)
	) name519 (
		_w4407_,
		_w4428_,
		_w4431_,
		_w4566_,
		_w4567_
	);
	LUT4 #(
		.INIT('h0700)
	) name520 (
		_w4506_,
		_w4563_,
		_w4565_,
		_w4567_,
		_w4568_
	);
	LUT4 #(
		.INIT('h4555)
	) name521 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4569_
	);
	LUT4 #(
		.INIT('h1000)
	) name522 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4570_
	);
	LUT4 #(
		.INIT('h888b)
	) name523 (
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w4093_,
		_w4569_,
		_w4570_,
		_w4571_
	);
	LUT4 #(
		.INIT('h0800)
	) name524 (
		\idma_DCTL_reg[1]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4572_
	);
	LUT3 #(
		.INIT('h07)
	) name525 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w4519_,
		_w4572_,
		_w4573_
	);
	LUT4 #(
		.INIT('h0015)
	) name526 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4573_,
		_w4574_
	);
	LUT4 #(
		.INIT('h00ef)
	) name527 (
		_w4089_,
		_w4107_,
		_w4571_,
		_w4574_,
		_w4575_
	);
	LUT4 #(
		.INIT('h8aff)
	) name528 (
		_w4108_,
		_w4562_,
		_w4568_,
		_w4575_,
		_w4576_
	);
	LUT3 #(
		.INIT('h10)
	) name529 (
		_w4345_,
		_w4500_,
		_w4502_,
		_w4577_
	);
	LUT3 #(
		.INIT('h78)
	) name530 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_EXA_reg[1]/P0001 ,
		\core_c_psq_EXA_reg[2]/P0001 ,
		_w4578_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name531 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4160_,
		_w4158_,
		_w4167_,
		_w4579_
	);
	LUT3 #(
		.INIT('ha3)
	) name532 (
		\core_c_psq_Taddr_Eb_reg[2]/P0001 ,
		_w4345_,
		_w4579_,
		_w4580_
	);
	LUT3 #(
		.INIT('h80)
	) name533 (
		_w4428_,
		_w4431_,
		_w4580_,
		_w4581_
	);
	LUT3 #(
		.INIT('h78)
	) name534 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		\core_c_psq_IFA_reg[1]/P0001 ,
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w4582_
	);
	LUT3 #(
		.INIT('h80)
	) name535 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[2]/P0001 ,
		_w4429_,
		_w4583_
	);
	LUT4 #(
		.INIT('h4000)
	) name536 (
		\core_c_psq_SRST_reg/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4065_,
		_w4066_,
		_w4584_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		_w4585_
	);
	LUT4 #(
		.INIT('h0001)
	) name538 (
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		\core_c_psq_Iact_E_reg[8]/NET0131 ,
		_w4586_
	);
	LUT2 #(
		.INIT('h8)
	) name539 (
		_w4585_,
		_w4586_,
		_w4587_
	);
	LUT2 #(
		.INIT('h2)
	) name540 (
		_w4584_,
		_w4587_,
		_w4588_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w4583_,
		_w4588_,
		_w4589_
	);
	LUT4 #(
		.INIT('hbf00)
	) name542 (
		_w4428_,
		_w4511_,
		_w4582_,
		_w4589_,
		_w4590_
	);
	LUT4 #(
		.INIT('h1300)
	) name543 (
		_w4506_,
		_w4581_,
		_w4578_,
		_w4590_,
		_w4591_
	);
	LUT4 #(
		.INIT('h4555)
	) name544 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4592_
	);
	LUT4 #(
		.INIT('h1000)
	) name545 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4593_
	);
	LUT4 #(
		.INIT('h888b)
	) name546 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w4093_,
		_w4592_,
		_w4593_,
		_w4594_
	);
	LUT4 #(
		.INIT('h0800)
	) name547 (
		\idma_DCTL_reg[2]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4595_
	);
	LUT3 #(
		.INIT('h07)
	) name548 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w4519_,
		_w4595_,
		_w4596_
	);
	LUT4 #(
		.INIT('h0015)
	) name549 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4596_,
		_w4597_
	);
	LUT4 #(
		.INIT('h00ef)
	) name550 (
		_w4089_,
		_w4107_,
		_w4594_,
		_w4597_,
		_w4598_
	);
	LUT4 #(
		.INIT('h8aff)
	) name551 (
		_w4108_,
		_w4577_,
		_w4591_,
		_w4598_,
		_w4599_
	);
	LUT3 #(
		.INIT('h10)
	) name552 (
		_w4283_,
		_w4500_,
		_w4502_,
		_w4600_
	);
	LUT4 #(
		.INIT('h7f80)
	) name553 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_EXA_reg[1]/P0001 ,
		\core_c_psq_EXA_reg[2]/P0001 ,
		\core_c_psq_EXA_reg[3]/P0001 ,
		_w4601_
	);
	LUT3 #(
		.INIT('ha3)
	) name554 (
		\core_c_psq_Taddr_Eb_reg[3]/P0001 ,
		_w4283_,
		_w4579_,
		_w4602_
	);
	LUT3 #(
		.INIT('h80)
	) name555 (
		_w4428_,
		_w4431_,
		_w4602_,
		_w4603_
	);
	LUT4 #(
		.INIT('h7f80)
	) name556 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		\core_c_psq_IFA_reg[1]/P0001 ,
		\core_c_psq_IFA_reg[2]/P0001 ,
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w4604_
	);
	LUT3 #(
		.INIT('h80)
	) name557 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[3]/P0001 ,
		_w4429_,
		_w4605_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		_w4606_
	);
	LUT4 #(
		.INIT('h0001)
	) name559 (
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		\core_c_psq_Iact_E_reg[9]/NET0131 ,
		_w4607_
	);
	LUT2 #(
		.INIT('h8)
	) name560 (
		_w4606_,
		_w4607_,
		_w4608_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		_w4584_,
		_w4608_,
		_w4609_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w4605_,
		_w4609_,
		_w4610_
	);
	LUT4 #(
		.INIT('hbf00)
	) name563 (
		_w4428_,
		_w4511_,
		_w4604_,
		_w4610_,
		_w4611_
	);
	LUT4 #(
		.INIT('h1300)
	) name564 (
		_w4506_,
		_w4603_,
		_w4601_,
		_w4611_,
		_w4612_
	);
	LUT4 #(
		.INIT('h4555)
	) name565 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4613_
	);
	LUT4 #(
		.INIT('h1000)
	) name566 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4614_
	);
	LUT4 #(
		.INIT('h888b)
	) name567 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w4093_,
		_w4613_,
		_w4614_,
		_w4615_
	);
	LUT4 #(
		.INIT('h0800)
	) name568 (
		\idma_DCTL_reg[3]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4616_
	);
	LUT3 #(
		.INIT('h07)
	) name569 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w4519_,
		_w4616_,
		_w4617_
	);
	LUT4 #(
		.INIT('h0015)
	) name570 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4617_,
		_w4618_
	);
	LUT4 #(
		.INIT('h00ef)
	) name571 (
		_w4089_,
		_w4107_,
		_w4615_,
		_w4618_,
		_w4619_
	);
	LUT4 #(
		.INIT('h8aff)
	) name572 (
		_w4108_,
		_w4600_,
		_w4612_,
		_w4619_,
		_w4620_
	);
	LUT3 #(
		.INIT('h10)
	) name573 (
		_w4203_,
		_w4500_,
		_w4502_,
		_w4621_
	);
	LUT2 #(
		.INIT('h6)
	) name574 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		_w4527_,
		_w4622_
	);
	LUT3 #(
		.INIT('ha3)
	) name575 (
		\core_c_psq_Taddr_Eb_reg[4]/P0001 ,
		_w4203_,
		_w4579_,
		_w4623_
	);
	LUT3 #(
		.INIT('h80)
	) name576 (
		_w4428_,
		_w4431_,
		_w4623_,
		_w4624_
	);
	LUT2 #(
		.INIT('h6)
	) name577 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w4532_,
		_w4625_
	);
	LUT3 #(
		.INIT('h80)
	) name578 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[4]/P0001 ,
		_w4429_,
		_w4626_
	);
	LUT4 #(
		.INIT('h0001)
	) name579 (
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		\core_c_psq_Iact_E_reg[7]/NET0131 ,
		_w4627_
	);
	LUT2 #(
		.INIT('h2)
	) name580 (
		_w4584_,
		_w4627_,
		_w4628_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w4626_,
		_w4628_,
		_w4629_
	);
	LUT4 #(
		.INIT('hbf00)
	) name582 (
		_w4428_,
		_w4511_,
		_w4625_,
		_w4629_,
		_w4630_
	);
	LUT4 #(
		.INIT('h1300)
	) name583 (
		_w4506_,
		_w4624_,
		_w4622_,
		_w4630_,
		_w4631_
	);
	LUT4 #(
		.INIT('h4555)
	) name584 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4632_
	);
	LUT4 #(
		.INIT('h1000)
	) name585 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4633_
	);
	LUT4 #(
		.INIT('h888b)
	) name586 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w4093_,
		_w4632_,
		_w4633_,
		_w4634_
	);
	LUT4 #(
		.INIT('h0800)
	) name587 (
		\idma_DCTL_reg[4]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4635_
	);
	LUT3 #(
		.INIT('h07)
	) name588 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w4519_,
		_w4635_,
		_w4636_
	);
	LUT4 #(
		.INIT('h0015)
	) name589 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4636_,
		_w4637_
	);
	LUT4 #(
		.INIT('h00ef)
	) name590 (
		_w4089_,
		_w4107_,
		_w4634_,
		_w4637_,
		_w4638_
	);
	LUT4 #(
		.INIT('h8aff)
	) name591 (
		_w4108_,
		_w4621_,
		_w4631_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('h4544)
	) name592 (
		_w4328_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4640_
	);
	LUT3 #(
		.INIT('h6c)
	) name593 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		\core_c_psq_EXA_reg[5]/P0001 ,
		_w4527_,
		_w4641_
	);
	LUT3 #(
		.INIT('h6c)
	) name594 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w4532_,
		_w4642_
	);
	LUT3 #(
		.INIT('h40)
	) name595 (
		_w4428_,
		_w4511_,
		_w4642_,
		_w4643_
	);
	LUT4 #(
		.INIT('h0001)
	) name596 (
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		\core_c_psq_Iact_E_reg[3]/NET0131 ,
		_w4644_
	);
	LUT2 #(
		.INIT('h2)
	) name597 (
		_w4584_,
		_w4644_,
		_w4645_
	);
	LUT3 #(
		.INIT('h80)
	) name598 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[5]/P0001 ,
		_w4429_,
		_w4646_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		_w4645_,
		_w4646_,
		_w4647_
	);
	LUT4 #(
		.INIT('h7f00)
	) name600 (
		_w4379_,
		_w4428_,
		_w4431_,
		_w4647_,
		_w4648_
	);
	LUT4 #(
		.INIT('h1300)
	) name601 (
		_w4506_,
		_w4643_,
		_w4641_,
		_w4648_,
		_w4649_
	);
	LUT4 #(
		.INIT('h4555)
	) name602 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4650_
	);
	LUT4 #(
		.INIT('h1000)
	) name603 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4651_
	);
	LUT4 #(
		.INIT('h888b)
	) name604 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w4093_,
		_w4650_,
		_w4651_,
		_w4652_
	);
	LUT4 #(
		.INIT('h0800)
	) name605 (
		\idma_DCTL_reg[5]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4653_
	);
	LUT3 #(
		.INIT('h07)
	) name606 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w4519_,
		_w4653_,
		_w4654_
	);
	LUT4 #(
		.INIT('h0015)
	) name607 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4654_,
		_w4655_
	);
	LUT4 #(
		.INIT('h00ef)
	) name608 (
		_w4089_,
		_w4107_,
		_w4652_,
		_w4655_,
		_w4656_
	);
	LUT4 #(
		.INIT('h8aff)
	) name609 (
		_w4108_,
		_w4640_,
		_w4649_,
		_w4656_,
		_w4657_
	);
	LUT4 #(
		.INIT('h4544)
	) name610 (
		_w4301_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4658_
	);
	LUT4 #(
		.INIT('h78f0)
	) name611 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		\core_c_psq_EXA_reg[5]/P0001 ,
		\core_c_psq_EXA_reg[6]/P0001 ,
		_w4527_,
		_w4659_
	);
	LUT3 #(
		.INIT('h80)
	) name612 (
		_w4391_,
		_w4428_,
		_w4431_,
		_w4660_
	);
	LUT4 #(
		.INIT('h78f0)
	) name613 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		\core_c_psq_IFA_reg[5]/P0001 ,
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w4532_,
		_w4661_
	);
	LUT3 #(
		.INIT('h80)
	) name614 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[6]/P0001 ,
		_w4429_,
		_w4662_
	);
	LUT4 #(
		.INIT('h00bf)
	) name615 (
		_w4428_,
		_w4511_,
		_w4661_,
		_w4662_,
		_w4663_
	);
	LUT4 #(
		.INIT('h0700)
	) name616 (
		_w4506_,
		_w4659_,
		_w4660_,
		_w4663_,
		_w4664_
	);
	LUT4 #(
		.INIT('h4555)
	) name617 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4665_
	);
	LUT4 #(
		.INIT('h1000)
	) name618 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4666_
	);
	LUT4 #(
		.INIT('h888b)
	) name619 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w4093_,
		_w4665_,
		_w4666_,
		_w4667_
	);
	LUT4 #(
		.INIT('h0800)
	) name620 (
		\idma_DCTL_reg[6]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4668_
	);
	LUT3 #(
		.INIT('h07)
	) name621 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w4519_,
		_w4668_,
		_w4669_
	);
	LUT4 #(
		.INIT('h0015)
	) name622 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4669_,
		_w4670_
	);
	LUT4 #(
		.INIT('h00ef)
	) name623 (
		_w4089_,
		_w4107_,
		_w4667_,
		_w4670_,
		_w4671_
	);
	LUT4 #(
		.INIT('h8aff)
	) name624 (
		_w4108_,
		_w4658_,
		_w4664_,
		_w4671_,
		_w4672_
	);
	LUT4 #(
		.INIT('h4544)
	) name625 (
		_w4269_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4673_
	);
	LUT2 #(
		.INIT('h6)
	) name626 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		_w4528_,
		_w4674_
	);
	LUT3 #(
		.INIT('h80)
	) name627 (
		_w4376_,
		_w4428_,
		_w4431_,
		_w4675_
	);
	LUT2 #(
		.INIT('h6)
	) name628 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w4533_,
		_w4676_
	);
	LUT3 #(
		.INIT('h80)
	) name629 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[7]/P0001 ,
		_w4429_,
		_w4677_
	);
	LUT4 #(
		.INIT('h00bf)
	) name630 (
		_w4428_,
		_w4511_,
		_w4676_,
		_w4677_,
		_w4678_
	);
	LUT4 #(
		.INIT('h0700)
	) name631 (
		_w4506_,
		_w4674_,
		_w4675_,
		_w4678_,
		_w4679_
	);
	LUT4 #(
		.INIT('h4555)
	) name632 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4680_
	);
	LUT4 #(
		.INIT('h1000)
	) name633 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4681_
	);
	LUT4 #(
		.INIT('h888b)
	) name634 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w4093_,
		_w4680_,
		_w4681_,
		_w4682_
	);
	LUT4 #(
		.INIT('h0800)
	) name635 (
		\idma_DCTL_reg[7]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4683_
	);
	LUT3 #(
		.INIT('h07)
	) name636 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w4519_,
		_w4683_,
		_w4684_
	);
	LUT4 #(
		.INIT('h0015)
	) name637 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4684_,
		_w4685_
	);
	LUT4 #(
		.INIT('h00ef)
	) name638 (
		_w4089_,
		_w4107_,
		_w4682_,
		_w4685_,
		_w4686_
	);
	LUT4 #(
		.INIT('h8aff)
	) name639 (
		_w4108_,
		_w4673_,
		_w4679_,
		_w4686_,
		_w4687_
	);
	LUT4 #(
		.INIT('h4544)
	) name640 (
		_w4190_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4688_
	);
	LUT3 #(
		.INIT('h6c)
	) name641 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		\core_c_psq_EXA_reg[8]/P0001 ,
		_w4528_,
		_w4689_
	);
	LUT3 #(
		.INIT('h80)
	) name642 (
		_w4422_,
		_w4428_,
		_w4431_,
		_w4690_
	);
	LUT3 #(
		.INIT('h6c)
	) name643 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w4533_,
		_w4691_
	);
	LUT3 #(
		.INIT('h80)
	) name644 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[8]/P0001 ,
		_w4429_,
		_w4692_
	);
	LUT4 #(
		.INIT('h00bf)
	) name645 (
		_w4428_,
		_w4511_,
		_w4691_,
		_w4692_,
		_w4693_
	);
	LUT4 #(
		.INIT('h0700)
	) name646 (
		_w4506_,
		_w4689_,
		_w4690_,
		_w4693_,
		_w4694_
	);
	LUT4 #(
		.INIT('h4555)
	) name647 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4695_
	);
	LUT4 #(
		.INIT('h1000)
	) name648 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4696_
	);
	LUT4 #(
		.INIT('h888b)
	) name649 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w4093_,
		_w4695_,
		_w4696_,
		_w4697_
	);
	LUT4 #(
		.INIT('h0800)
	) name650 (
		\idma_DCTL_reg[8]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4698_
	);
	LUT3 #(
		.INIT('h07)
	) name651 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w4519_,
		_w4698_,
		_w4699_
	);
	LUT4 #(
		.INIT('h0015)
	) name652 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4699_,
		_w4700_
	);
	LUT4 #(
		.INIT('h00ef)
	) name653 (
		_w4089_,
		_w4107_,
		_w4697_,
		_w4700_,
		_w4701_
	);
	LUT4 #(
		.INIT('h8aff)
	) name654 (
		_w4108_,
		_w4688_,
		_w4694_,
		_w4701_,
		_w4702_
	);
	LUT4 #(
		.INIT('h4544)
	) name655 (
		_w4230_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4703_
	);
	LUT4 #(
		.INIT('h78f0)
	) name656 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_EXA_reg[9]/P0001 ,
		_w4528_,
		_w4704_
	);
	LUT3 #(
		.INIT('h80)
	) name657 (
		_w4413_,
		_w4428_,
		_w4431_,
		_w4705_
	);
	LUT4 #(
		.INIT('h78f0)
	) name658 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		\core_c_psq_IFA_reg[8]/P0001 ,
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w4533_,
		_w4706_
	);
	LUT3 #(
		.INIT('h80)
	) name659 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[9]/P0001 ,
		_w4429_,
		_w4707_
	);
	LUT4 #(
		.INIT('h00bf)
	) name660 (
		_w4428_,
		_w4511_,
		_w4706_,
		_w4707_,
		_w4708_
	);
	LUT4 #(
		.INIT('h0700)
	) name661 (
		_w4506_,
		_w4704_,
		_w4705_,
		_w4708_,
		_w4709_
	);
	LUT4 #(
		.INIT('h4555)
	) name662 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4710_
	);
	LUT4 #(
		.INIT('h1000)
	) name663 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4711_
	);
	LUT4 #(
		.INIT('h888b)
	) name664 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w4093_,
		_w4710_,
		_w4711_,
		_w4712_
	);
	LUT4 #(
		.INIT('h0800)
	) name665 (
		\idma_DCTL_reg[9]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4713_
	);
	LUT3 #(
		.INIT('h07)
	) name666 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w4519_,
		_w4713_,
		_w4714_
	);
	LUT4 #(
		.INIT('h0015)
	) name667 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4714_,
		_w4715_
	);
	LUT4 #(
		.INIT('h00ef)
	) name668 (
		_w4089_,
		_w4107_,
		_w4712_,
		_w4715_,
		_w4716_
	);
	LUT4 #(
		.INIT('h8aff)
	) name669 (
		_w4108_,
		_w4703_,
		_w4709_,
		_w4716_,
		_w4717_
	);
	LUT4 #(
		.INIT('h0040)
	) name670 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4718_
	);
	LUT4 #(
		.INIT('h0020)
	) name671 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4719_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		_w4720_
	);
	LUT4 #(
		.INIT('h0002)
	) name673 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4721_
	);
	LUT3 #(
		.INIT('h08)
	) name674 (
		\core_c_dec_Double_E_reg/P0001 ,
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		_w4722_
	);
	LUT4 #(
		.INIT('h0145)
	) name675 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[1]/NET0131 ,
		\emc_WSCRreg_DO_reg[3]/NET0131 ,
		_w4723_
	);
	LUT2 #(
		.INIT('h2)
	) name676 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[11]/NET0131 ,
		_w4724_
	);
	LUT4 #(
		.INIT('h888d)
	) name677 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[7]/NET0131 ,
		_w4723_,
		_w4724_,
		_w4725_
	);
	LUT4 #(
		.INIT('h0415)
	) name678 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[0]/NET0131 ,
		\memc_usysr_DO_reg[14]/NET0131 ,
		_w4726_
	);
	LUT2 #(
		.INIT('h2)
	) name679 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[8]/NET0131 ,
		_w4727_
	);
	LUT4 #(
		.INIT('h888d)
	) name680 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[4]/NET0131 ,
		_w4726_,
		_w4727_,
		_w4728_
	);
	LUT4 #(
		.INIT('ha251)
	) name681 (
		\emc_RWcnt_reg[0]/P0001 ,
		\emc_RWcnt_reg[3]/P0001 ,
		_w4725_,
		_w4728_,
		_w4729_
	);
	LUT2 #(
		.INIT('h2)
	) name682 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[4]/NET0131 ,
		_w4730_
	);
	LUT3 #(
		.INIT('h40)
	) name683 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[2]/NET0131 ,
		_w4731_
	);
	LUT3 #(
		.INIT('h13)
	) name684 (
		\emc_DMcst_reg/NET0131 ,
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[6]/NET0131 ,
		_w4732_
	);
	LUT4 #(
		.INIT('h9a99)
	) name685 (
		\emc_RWcnt_reg[4]/P0001 ,
		_w4730_,
		_w4731_,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h2)
	) name686 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[5]/NET0131 ,
		_w4734_
	);
	LUT3 #(
		.INIT('h40)
	) name687 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[3]/NET0131 ,
		_w4735_
	);
	LUT3 #(
		.INIT('h13)
	) name688 (
		\emc_DMcst_reg/NET0131 ,
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[7]/NET0131 ,
		_w4736_
	);
	LUT4 #(
		.INIT('h6566)
	) name689 (
		\emc_RWcnt_reg[5]/P0001 ,
		_w4734_,
		_w4735_,
		_w4736_,
		_w4737_
	);
	LUT4 #(
		.INIT('h0b00)
	) name690 (
		\emc_RWcnt_reg[3]/P0001 ,
		_w4725_,
		_w4733_,
		_w4737_,
		_w4738_
	);
	LUT4 #(
		.INIT('h0415)
	) name691 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[1]/NET0131 ,
		\memc_usysr_DO_reg[15]/NET0131 ,
		_w4739_
	);
	LUT2 #(
		.INIT('h2)
	) name692 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[9]/NET0131 ,
		_w4740_
	);
	LUT4 #(
		.INIT('h888d)
	) name693 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[5]/NET0131 ,
		_w4739_,
		_w4740_,
		_w4741_
	);
	LUT4 #(
		.INIT('h0145)
	) name694 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[0]/NET0131 ,
		\emc_WSCRreg_DO_reg[2]/NET0131 ,
		_w4742_
	);
	LUT2 #(
		.INIT('h2)
	) name695 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[10]/NET0131 ,
		_w4743_
	);
	LUT4 #(
		.INIT('h888d)
	) name696 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[6]/NET0131 ,
		_w4742_,
		_w4743_,
		_w4744_
	);
	LUT4 #(
		.INIT('h8421)
	) name697 (
		\emc_RWcnt_reg[1]/P0001 ,
		\emc_RWcnt_reg[2]/P0001 ,
		_w4741_,
		_w4744_,
		_w4745_
	);
	LUT4 #(
		.INIT('h4000)
	) name698 (
		_w4722_,
		_w4738_,
		_w4729_,
		_w4745_,
		_w4746_
	);
	LUT2 #(
		.INIT('h2)
	) name699 (
		_w4721_,
		_w4746_,
		_w4747_
	);
	LUT3 #(
		.INIT('h10)
	) name700 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4748_
	);
	LUT4 #(
		.INIT('h8000)
	) name701 (
		_w4738_,
		_w4729_,
		_w4745_,
		_w4748_,
		_w4749_
	);
	LUT4 #(
		.INIT('h0200)
	) name702 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4750_
	);
	LUT4 #(
		.INIT('hfddf)
	) name703 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4751_
	);
	LUT4 #(
		.INIT('h007f)
	) name704 (
		_w4738_,
		_w4729_,
		_w4745_,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4753_
	);
	LUT3 #(
		.INIT('h01)
	) name706 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		\emc_PMcst_reg/NET0131 ,
		_w4754_
	);
	LUT2 #(
		.INIT('h2)
	) name707 (
		\core_c_psq_ECYC_reg/P0001 ,
		\emc_eRDY_reg/NET0131 ,
		_w4755_
	);
	LUT3 #(
		.INIT('h01)
	) name708 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4756_
	);
	LUT4 #(
		.INIT('hba00)
	) name709 (
		\emc_ECS_reg[2]/NET0131 ,
		_w4754_,
		_w4755_,
		_w4756_,
		_w4757_
	);
	LUT4 #(
		.INIT('h27d8)
	) name710 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w4758_
	);
	LUT4 #(
		.INIT('hd827)
	) name711 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		\bdma_BCTL_reg[6]/NET0131 ,
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w4759_
	);
	LUT4 #(
		.INIT('hd827)
	) name712 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[6]/NET0131 ,
		\bdma_BCTL_reg[7]/NET0131 ,
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w4760_
	);
	LUT3 #(
		.INIT('h40)
	) name713 (
		_w4758_,
		_w4759_,
		_w4760_,
		_w4761_
	);
	LUT3 #(
		.INIT('h1e)
	) name714 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BWcnt_reg[0]/NET0131 ,
		_w4762_
	);
	LUT3 #(
		.INIT('h2d)
	) name715 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[7]/NET0131 ,
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w4763_
	);
	LUT4 #(
		.INIT('h1000)
	) name716 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4764_
	);
	LUT3 #(
		.INIT('h10)
	) name717 (
		_w4762_,
		_w4763_,
		_w4764_,
		_w4765_
	);
	LUT2 #(
		.INIT('h8)
	) name718 (
		_w4761_,
		_w4765_,
		_w4766_
	);
	LUT3 #(
		.INIT('h15)
	) name719 (
		_w4757_,
		_w4761_,
		_w4765_,
		_w4767_
	);
	LUT3 #(
		.INIT('h10)
	) name720 (
		_w4752_,
		_w4749_,
		_w4767_,
		_w4768_
	);
	LUT2 #(
		.INIT('hb)
	) name721 (
		_w4747_,
		_w4768_,
		_w4769_
	);
	LUT4 #(
		.INIT('h0001)
	) name722 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		\emc_PMcst_reg/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w4770_
	);
	LUT3 #(
		.INIT('h04)
	) name723 (
		\T_TMODE[1]_pad ,
		\bdma_BDMAmode_reg/NET0131 ,
		\core_c_psq_ECYC_reg/P0001 ,
		_w4771_
	);
	LUT3 #(
		.INIT('h5b)
	) name724 (
		\T_TMODE[1]_pad ,
		\bdma_BDMAmode_reg/NET0131 ,
		\core_c_psq_ECYC_reg/P0001 ,
		_w4772_
	);
	LUT4 #(
		.INIT('h0800)
	) name725 (
		_w4720_,
		_w4753_,
		_w4772_,
		_w4770_,
		_w4773_
	);
	LUT4 #(
		.INIT('h2000)
	) name726 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4774_
	);
	LUT4 #(
		.INIT('h4000)
	) name727 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4775_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name728 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BSreq_reg/NET0131 ,
		_w4774_,
		_w4775_,
		_w4776_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name729 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4777_
	);
	LUT2 #(
		.INIT('h8)
	) name730 (
		\T_TMODE[1]_pad ,
		\emc_ECS_reg[1]/NET0131 ,
		_w4778_
	);
	LUT4 #(
		.INIT('h0020)
	) name731 (
		\T_TMODE[1]_pad ,
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4779_
	);
	LUT3 #(
		.INIT('h10)
	) name732 (
		_w4764_,
		_w4779_,
		_w4777_,
		_w4780_
	);
	LUT3 #(
		.INIT('h20)
	) name733 (
		_w4776_,
		_w4773_,
		_w4780_,
		_w4781_
	);
	LUT3 #(
		.INIT('hdf)
	) name734 (
		_w4776_,
		_w4773_,
		_w4780_,
		_w4782_
	);
	LUT4 #(
		.INIT('hfddd)
	) name735 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4783_
	);
	LUT4 #(
		.INIT('h0080)
	) name736 (
		_w4738_,
		_w4729_,
		_w4745_,
		_w4783_,
		_w4784_
	);
	LUT4 #(
		.INIT('h0400)
	) name737 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4785_
	);
	LUT2 #(
		.INIT('h2)
	) name738 (
		_w4776_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h4)
	) name739 (
		_w4784_,
		_w4786_,
		_w4787_
	);
	LUT2 #(
		.INIT('hb)
	) name740 (
		_w4784_,
		_w4786_,
		_w4788_
	);
	LUT3 #(
		.INIT('h20)
	) name741 (
		_w4781_,
		_w4784_,
		_w4786_,
		_w4789_
	);
	LUT2 #(
		.INIT('h2)
	) name742 (
		_w4753_,
		_w4771_,
		_w4790_
	);
	LUT3 #(
		.INIT('h54)
	) name743 (
		\core_c_psq_ECYC_reg/P0001 ,
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4791_
	);
	LUT3 #(
		.INIT('h08)
	) name744 (
		_w4720_,
		_w4770_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		_w4793_
	);
	LUT4 #(
		.INIT('h0008)
	) name746 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4794_
	);
	LUT4 #(
		.INIT('hefc7)
	) name747 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4795_
	);
	LUT4 #(
		.INIT('h8a00)
	) name748 (
		_w4776_,
		_w4790_,
		_w4792_,
		_w4795_,
		_w4796_
	);
	LUT4 #(
		.INIT('h75ff)
	) name749 (
		_w4776_,
		_w4790_,
		_w4792_,
		_w4795_,
		_w4797_
	);
	LUT4 #(
		.INIT('h0020)
	) name750 (
		_w4781_,
		_w4784_,
		_w4786_,
		_w4796_,
		_w4798_
	);
	LUT4 #(
		.INIT('h1055)
	) name751 (
		_w4719_,
		_w4747_,
		_w4768_,
		_w4798_,
		_w4799_
	);
	LUT3 #(
		.INIT('h75)
	) name752 (
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w4800_
	);
	LUT4 #(
		.INIT('h8088)
	) name753 (
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[14]/NET0131 ,
		_w4718_,
		_w4799_,
		_w4801_
	);
	LUT3 #(
		.INIT('h75)
	) name754 (
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w4802_
	);
	LUT4 #(
		.INIT('h8088)
	) name755 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[13]/NET0131 ,
		_w4718_,
		_w4799_,
		_w4803_
	);
	LUT4 #(
		.INIT('h0004)
	) name756 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w4804_
	);
	LUT4 #(
		.INIT('hb000)
	) name757 (
		_w4747_,
		_w4768_,
		_w4789_,
		_w4796_,
		_w4805_
	);
	LUT3 #(
		.INIT('h01)
	) name758 (
		_w4721_,
		_w4804_,
		_w4805_,
		_w4806_
	);
	LUT4 #(
		.INIT('haaa8)
	) name759 (
		\emc_WSCRreg_DO_reg[12]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w4807_
	);
	LUT3 #(
		.INIT('h01)
	) name760 (
		_w4803_,
		_w4807_,
		_w4801_,
		_w4808_
	);
	LUT4 #(
		.INIT('h4544)
	) name761 (
		_w4216_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4809_
	);
	LUT4 #(
		.INIT('h8000)
	) name762 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_EXA_reg[12]/P0001 ,
		_w4529_,
		_w4810_
	);
	LUT4 #(
		.INIT('h78f0)
	) name763 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_EXA_reg[12]/P0001 ,
		_w4529_,
		_w4811_
	);
	LUT3 #(
		.INIT('h80)
	) name764 (
		_w4409_,
		_w4428_,
		_w4431_,
		_w4812_
	);
	LUT4 #(
		.INIT('h8000)
	) name765 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		\core_c_psq_IFA_reg[11]/P0001 ,
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w4534_,
		_w4813_
	);
	LUT4 #(
		.INIT('h78f0)
	) name766 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		\core_c_psq_IFA_reg[11]/P0001 ,
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w4534_,
		_w4814_
	);
	LUT3 #(
		.INIT('h80)
	) name767 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[12]/P0001 ,
		_w4429_,
		_w4815_
	);
	LUT4 #(
		.INIT('h00bf)
	) name768 (
		_w4428_,
		_w4511_,
		_w4814_,
		_w4815_,
		_w4816_
	);
	LUT4 #(
		.INIT('h0700)
	) name769 (
		_w4506_,
		_w4811_,
		_w4812_,
		_w4816_,
		_w4817_
	);
	LUT4 #(
		.INIT('h4555)
	) name770 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4818_
	);
	LUT4 #(
		.INIT('h1000)
	) name771 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4819_
	);
	LUT4 #(
		.INIT('h888b)
	) name772 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w4093_,
		_w4818_,
		_w4819_,
		_w4820_
	);
	LUT4 #(
		.INIT('h0800)
	) name773 (
		\idma_DCTL_reg[12]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4821_
	);
	LUT3 #(
		.INIT('h07)
	) name774 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w4519_,
		_w4821_,
		_w4822_
	);
	LUT4 #(
		.INIT('h0015)
	) name775 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4822_,
		_w4823_
	);
	LUT4 #(
		.INIT('h00ef)
	) name776 (
		_w4089_,
		_w4107_,
		_w4820_,
		_w4823_,
		_w4824_
	);
	LUT4 #(
		.INIT('h7500)
	) name777 (
		_w4108_,
		_w4809_,
		_w4817_,
		_w4824_,
		_w4825_
	);
	LUT4 #(
		.INIT('h8aff)
	) name778 (
		_w4108_,
		_w4809_,
		_w4817_,
		_w4824_,
		_w4826_
	);
	LUT4 #(
		.INIT('h4544)
	) name779 (
		_w4243_,
		_w4432_,
		_w4500_,
		_w4502_,
		_w4827_
	);
	LUT2 #(
		.INIT('h6)
	) name780 (
		\core_c_psq_EXA_reg[13]/P0001 ,
		_w4810_,
		_w4828_
	);
	LUT2 #(
		.INIT('h6)
	) name781 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w4813_,
		_w4829_
	);
	LUT3 #(
		.INIT('h40)
	) name782 (
		_w4428_,
		_w4511_,
		_w4829_,
		_w4830_
	);
	LUT3 #(
		.INIT('h80)
	) name783 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\sice_IRR_reg[13]/P0001 ,
		_w4429_,
		_w4831_
	);
	LUT4 #(
		.INIT('h007f)
	) name784 (
		_w4369_,
		_w4428_,
		_w4431_,
		_w4831_,
		_w4832_
	);
	LUT4 #(
		.INIT('h0700)
	) name785 (
		_w4506_,
		_w4828_,
		_w4830_,
		_w4832_,
		_w4833_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name786 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4834_
	);
	LUT4 #(
		.INIT('h2000)
	) name787 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4835_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name788 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w4093_,
		_w4835_,
		_w4834_,
		_w4836_
	);
	LUT3 #(
		.INIT('h10)
	) name789 (
		_w4089_,
		_w4107_,
		_w4836_,
		_w4837_
	);
	LUT4 #(
		.INIT('h2a00)
	) name790 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w4067_,
		_w4088_,
		_w4519_,
		_w4838_
	);
	LUT4 #(
		.INIT('h0800)
	) name791 (
		\idma_DCTL_reg[13]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4839_
	);
	LUT4 #(
		.INIT('h1500)
	) name792 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4839_,
		_w4840_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w4838_,
		_w4840_,
		_w4841_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		_w4837_,
		_w4841_,
		_w4842_
	);
	LUT4 #(
		.INIT('h7500)
	) name795 (
		_w4108_,
		_w4827_,
		_w4833_,
		_w4842_,
		_w4843_
	);
	LUT4 #(
		.INIT('h8aff)
	) name796 (
		_w4108_,
		_w4827_,
		_w4833_,
		_w4842_,
		_w4844_
	);
	LUT4 #(
		.INIT('h4000)
	) name797 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4087_,
		_w4845_
	);
	LUT3 #(
		.INIT('h20)
	) name798 (
		_w4067_,
		_w4068_,
		_w4845_,
		_w4846_
	);
	LUT2 #(
		.INIT('h8)
	) name799 (
		\core_c_psq_MGNT_reg/NET0131 ,
		\core_c_psq_PCS_reg[10]/NET0131 ,
		_w4847_
	);
	LUT4 #(
		.INIT('h2000)
	) name800 (
		\core_c_psq_PCS_reg[0]/NET0131 ,
		\core_c_psq_SRST_reg/P0001 ,
		_w4065_,
		_w4066_,
		_w4848_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[13]/NET0131 ,
		_w4849_
	);
	LUT3 #(
		.INIT('h51)
	) name802 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		_w4075_,
		_w4849_,
		_w4850_
	);
	LUT4 #(
		.INIT('h1311)
	) name803 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w4847_,
		_w4848_,
		_w4850_,
		_w4851_
	);
	LUT4 #(
		.INIT('hecee)
	) name804 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w4847_,
		_w4848_,
		_w4850_,
		_w4852_
	);
	LUT2 #(
		.INIT('h4)
	) name805 (
		\core_c_psq_MGNT_reg/NET0131 ,
		\core_c_psq_PCS_reg[10]/NET0131 ,
		_w4853_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[11]/NET0131 ,
		_w4854_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name807 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w4075_,
		_w4853_,
		_w4854_,
		_w4855_
	);
	LUT2 #(
		.INIT('h2)
	) name808 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w4856_
	);
	LUT4 #(
		.INIT('h3323)
	) name809 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[11]/NET0131 ,
		\core_c_psq_PCS_reg[5]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w4857_
	);
	LUT4 #(
		.INIT('hccdc)
	) name810 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[11]/NET0131 ,
		\core_c_psq_PCS_reg[5]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w4858_
	);
	LUT2 #(
		.INIT('h8)
	) name811 (
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\memc_LDaST_Eg_reg/NET0131 ,
		_w4859_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name812 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w4075_,
		_w4857_,
		_w4859_,
		_w4860_
	);
	LUT3 #(
		.INIT('hd0)
	) name813 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w4860_,
		_w4861_
	);
	LUT2 #(
		.INIT('h2)
	) name814 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w4862_
	);
	LUT4 #(
		.INIT('ha820)
	) name815 (
		\core_c_psq_PCS_reg[10]/NET0131 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		_w4863_
	);
	LUT4 #(
		.INIT('h4000)
	) name816 (
		\core_c_psq_SRST_reg/P0001 ,
		_w4065_,
		_w4066_,
		_w4863_,
		_w4864_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w4862_,
		_w4864_,
		_w4865_
	);
	LUT2 #(
		.INIT('he)
	) name818 (
		_w4862_,
		_w4864_,
		_w4866_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_c_psq_PCS_reg[8]/NET0131 ,
		_w4867_
	);
	LUT2 #(
		.INIT('h4)
	) name820 (
		_w4078_,
		_w4867_,
		_w4868_
	);
	LUT3 #(
		.INIT('h45)
	) name821 (
		_w4069_,
		_w4077_,
		_w4868_,
		_w4869_
	);
	LUT4 #(
		.INIT('h0080)
	) name822 (
		_w4861_,
		_w4865_,
		_w4851_,
		_w4869_,
		_w4870_
	);
	LUT3 #(
		.INIT('h0b)
	) name823 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[2]/NET0131 ,
		_w4871_
	);
	LUT3 #(
		.INIT('h02)
	) name824 (
		\core_c_dec_IDLE_Eg_reg/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		\sice_HALT_E_reg/P0001 ,
		_w4872_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name825 (
		\core_c_psq_PCS_reg[6]/NET0131 ,
		_w4081_,
		_w4871_,
		_w4872_,
		_w4873_
	);
	LUT4 #(
		.INIT('h2f22)
	) name826 (
		\core_c_psq_PCS_reg[6]/NET0131 ,
		_w4081_,
		_w4871_,
		_w4872_,
		_w4874_
	);
	LUT4 #(
		.INIT('h0400)
	) name827 (
		_w4094_,
		_w4097_,
		_w4101_,
		_w4873_,
		_w4875_
	);
	LUT2 #(
		.INIT('h8)
	) name828 (
		_w4870_,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('h8)
	) name829 (
		\clkc_Cnt4096_s1_reg/NET0131 ,
		\clkc_Cnt4096_s2_reg/NET0131 ,
		_w4877_
	);
	LUT3 #(
		.INIT('h04)
	) name830 (
		_w4099_,
		_w4100_,
		_w4877_,
		_w4878_
	);
	LUT3 #(
		.INIT('h10)
	) name831 (
		_w4519_,
		_w4520_,
		_w4878_,
		_w4879_
	);
	LUT3 #(
		.INIT('h51)
	) name832 (
		\T_TMODE[1]_pad ,
		_w4093_,
		_w4873_,
		_w4880_
	);
	LUT2 #(
		.INIT('h4)
	) name833 (
		_w4879_,
		_w4880_,
		_w4881_
	);
	LUT3 #(
		.INIT('h70)
	) name834 (
		_w4846_,
		_w4876_,
		_w4881_,
		_w4882_
	);
	LUT4 #(
		.INIT('hd000)
	) name835 (
		PM_bdry_sel_pad,
		_w4825_,
		_w4843_,
		_w4882_,
		_w4883_
	);
	LUT4 #(
		.INIT('h1000)
	) name836 (
		\bdma_BCTL_reg[0]/NET0131 ,
		\bdma_BCTL_reg[1]/NET0131 ,
		\bdma_BDMAmode_reg/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w4884_
	);
	LUT3 #(
		.INIT('he0)
	) name837 (
		PM_bdry_sel_pad,
		\bdma_BIAD_reg[12]/NET0131 ,
		\bdma_BIAD_reg[13]/NET0131 ,
		_w4885_
	);
	LUT2 #(
		.INIT('h4)
	) name838 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		\bdma_CMcnt_reg[1]/NET0131 ,
		_w4886_
	);
	LUT4 #(
		.INIT('h1000)
	) name839 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w4885_,
		_w4884_,
		_w4886_,
		_w4887_
	);
	LUT4 #(
		.INIT('h5333)
	) name840 (
		\bdma_BRdataBUF_reg[0]/P0001 ,
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w4519_,
		_w4887_,
		_w4888_
	);
	LUT3 #(
		.INIT('h8b)
	) name841 (
		\idma_DTMP_L_reg[0]/P0001 ,
		_w4520_,
		_w4888_,
		_w4889_
	);
	LUT4 #(
		.INIT('h5333)
	) name842 (
		\bdma_BRdataBUF_reg[10]/P0001 ,
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w4519_,
		_w4887_,
		_w4890_
	);
	LUT3 #(
		.INIT('h8b)
	) name843 (
		\idma_DTMP_H_reg[2]/P0001 ,
		_w4520_,
		_w4890_,
		_w4891_
	);
	LUT4 #(
		.INIT('h5333)
	) name844 (
		\bdma_BRdataBUF_reg[11]/P0001 ,
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w4519_,
		_w4887_,
		_w4892_
	);
	LUT3 #(
		.INIT('h8b)
	) name845 (
		\idma_DTMP_H_reg[3]/P0001 ,
		_w4520_,
		_w4892_,
		_w4893_
	);
	LUT4 #(
		.INIT('h5333)
	) name846 (
		\bdma_BRdataBUF_reg[12]/P0001 ,
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w4519_,
		_w4887_,
		_w4894_
	);
	LUT3 #(
		.INIT('h8b)
	) name847 (
		\idma_DTMP_H_reg[4]/P0001 ,
		_w4520_,
		_w4894_,
		_w4895_
	);
	LUT4 #(
		.INIT('h5333)
	) name848 (
		\bdma_BRdataBUF_reg[13]/P0001 ,
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w4519_,
		_w4887_,
		_w4896_
	);
	LUT3 #(
		.INIT('h8b)
	) name849 (
		\idma_DTMP_H_reg[5]/P0001 ,
		_w4520_,
		_w4896_,
		_w4897_
	);
	LUT4 #(
		.INIT('h5333)
	) name850 (
		\bdma_BRdataBUF_reg[14]/P0001 ,
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w4519_,
		_w4887_,
		_w4898_
	);
	LUT3 #(
		.INIT('h8b)
	) name851 (
		\idma_DTMP_H_reg[6]/P0001 ,
		_w4520_,
		_w4898_,
		_w4899_
	);
	LUT4 #(
		.INIT('h5333)
	) name852 (
		\bdma_BRdataBUF_reg[15]/P0001 ,
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w4519_,
		_w4887_,
		_w4900_
	);
	LUT3 #(
		.INIT('h8b)
	) name853 (
		\idma_DTMP_H_reg[7]/P0001 ,
		_w4520_,
		_w4900_,
		_w4901_
	);
	LUT4 #(
		.INIT('h5333)
	) name854 (
		\bdma_BRdataBUF_reg[16]/P0001 ,
		\sice_idr1_reg_DO_reg[4]/P0001 ,
		_w4519_,
		_w4887_,
		_w4902_
	);
	LUT3 #(
		.INIT('h8b)
	) name855 (
		\idma_DTMP_H_reg[8]/P0001 ,
		_w4520_,
		_w4902_,
		_w4903_
	);
	LUT4 #(
		.INIT('h5333)
	) name856 (
		\bdma_BRdataBUF_reg[17]/P0001 ,
		\sice_idr1_reg_DO_reg[5]/P0001 ,
		_w4519_,
		_w4887_,
		_w4904_
	);
	LUT3 #(
		.INIT('h8b)
	) name857 (
		\idma_DTMP_H_reg[9]/P0001 ,
		_w4520_,
		_w4904_,
		_w4905_
	);
	LUT4 #(
		.INIT('h5333)
	) name858 (
		\bdma_BRdataBUF_reg[18]/P0001 ,
		\sice_idr1_reg_DO_reg[6]/P0001 ,
		_w4519_,
		_w4887_,
		_w4906_
	);
	LUT3 #(
		.INIT('h8b)
	) name859 (
		\idma_DTMP_H_reg[10]/P0001 ,
		_w4520_,
		_w4906_,
		_w4907_
	);
	LUT4 #(
		.INIT('h5333)
	) name860 (
		\bdma_BRdataBUF_reg[19]/P0001 ,
		\sice_idr1_reg_DO_reg[7]/P0001 ,
		_w4519_,
		_w4887_,
		_w4908_
	);
	LUT3 #(
		.INIT('h8b)
	) name861 (
		\idma_DTMP_H_reg[11]/P0001 ,
		_w4520_,
		_w4908_,
		_w4909_
	);
	LUT4 #(
		.INIT('h5333)
	) name862 (
		\bdma_BRdataBUF_reg[1]/P0001 ,
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w4519_,
		_w4887_,
		_w4910_
	);
	LUT3 #(
		.INIT('h8b)
	) name863 (
		\idma_DTMP_L_reg[1]/P0001 ,
		_w4520_,
		_w4910_,
		_w4911_
	);
	LUT4 #(
		.INIT('h5333)
	) name864 (
		\bdma_BRdataBUF_reg[20]/P0001 ,
		\sice_idr1_reg_DO_reg[8]/P0001 ,
		_w4519_,
		_w4887_,
		_w4912_
	);
	LUT3 #(
		.INIT('h8b)
	) name865 (
		\idma_DTMP_H_reg[12]/P0001 ,
		_w4520_,
		_w4912_,
		_w4913_
	);
	LUT4 #(
		.INIT('h5333)
	) name866 (
		\bdma_BRdataBUF_reg[21]/P0001 ,
		\sice_idr1_reg_DO_reg[9]/P0001 ,
		_w4519_,
		_w4887_,
		_w4914_
	);
	LUT3 #(
		.INIT('h8b)
	) name867 (
		\idma_DTMP_H_reg[13]/P0001 ,
		_w4520_,
		_w4914_,
		_w4915_
	);
	LUT4 #(
		.INIT('h5333)
	) name868 (
		\bdma_BRdataBUF_reg[22]/P0001 ,
		\sice_idr1_reg_DO_reg[10]/P0001 ,
		_w4519_,
		_w4887_,
		_w4916_
	);
	LUT3 #(
		.INIT('h8b)
	) name869 (
		\idma_DTMP_H_reg[14]/P0001 ,
		_w4520_,
		_w4916_,
		_w4917_
	);
	LUT4 #(
		.INIT('h5333)
	) name870 (
		\bdma_BRdataBUF_reg[23]/P0001 ,
		\sice_idr1_reg_DO_reg[11]/P0001 ,
		_w4519_,
		_w4887_,
		_w4918_
	);
	LUT3 #(
		.INIT('h8b)
	) name871 (
		\idma_DTMP_H_reg[15]/P0001 ,
		_w4520_,
		_w4918_,
		_w4919_
	);
	LUT4 #(
		.INIT('h5333)
	) name872 (
		\bdma_BRdataBUF_reg[2]/P0001 ,
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w4519_,
		_w4887_,
		_w4920_
	);
	LUT3 #(
		.INIT('h8b)
	) name873 (
		\idma_DTMP_L_reg[2]/P0001 ,
		_w4520_,
		_w4920_,
		_w4921_
	);
	LUT4 #(
		.INIT('h5333)
	) name874 (
		\bdma_BRdataBUF_reg[3]/P0001 ,
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w4519_,
		_w4887_,
		_w4922_
	);
	LUT3 #(
		.INIT('h8b)
	) name875 (
		\idma_DTMP_L_reg[3]/P0001 ,
		_w4520_,
		_w4922_,
		_w4923_
	);
	LUT4 #(
		.INIT('h5333)
	) name876 (
		\bdma_BRdataBUF_reg[4]/P0001 ,
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w4519_,
		_w4887_,
		_w4924_
	);
	LUT3 #(
		.INIT('h8b)
	) name877 (
		\idma_DTMP_L_reg[4]/P0001 ,
		_w4520_,
		_w4924_,
		_w4925_
	);
	LUT4 #(
		.INIT('h5333)
	) name878 (
		\bdma_BRdataBUF_reg[5]/P0001 ,
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w4519_,
		_w4887_,
		_w4926_
	);
	LUT3 #(
		.INIT('h8b)
	) name879 (
		\idma_DTMP_L_reg[5]/P0001 ,
		_w4520_,
		_w4926_,
		_w4927_
	);
	LUT4 #(
		.INIT('h5333)
	) name880 (
		\bdma_BRdataBUF_reg[6]/P0001 ,
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w4519_,
		_w4887_,
		_w4928_
	);
	LUT3 #(
		.INIT('h8b)
	) name881 (
		\idma_DTMP_L_reg[6]/P0001 ,
		_w4520_,
		_w4928_,
		_w4929_
	);
	LUT4 #(
		.INIT('h5333)
	) name882 (
		\bdma_BRdataBUF_reg[7]/P0001 ,
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w4519_,
		_w4887_,
		_w4930_
	);
	LUT3 #(
		.INIT('h8b)
	) name883 (
		\idma_DTMP_L_reg[7]/P0001 ,
		_w4520_,
		_w4930_,
		_w4931_
	);
	LUT4 #(
		.INIT('h5333)
	) name884 (
		\bdma_BRdataBUF_reg[8]/P0001 ,
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w4519_,
		_w4887_,
		_w4932_
	);
	LUT3 #(
		.INIT('h8b)
	) name885 (
		\idma_DTMP_H_reg[0]/P0001 ,
		_w4520_,
		_w4932_,
		_w4933_
	);
	LUT4 #(
		.INIT('h5333)
	) name886 (
		\bdma_BRdataBUF_reg[9]/P0001 ,
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w4519_,
		_w4887_,
		_w4934_
	);
	LUT3 #(
		.INIT('h8b)
	) name887 (
		\idma_DTMP_H_reg[1]/P0001 ,
		_w4520_,
		_w4934_,
		_w4935_
	);
	LUT4 #(
		.INIT('h0400)
	) name888 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w4936_
	);
	LUT3 #(
		.INIT('he0)
	) name889 (
		PM_bdry_sel_pad,
		\idma_DCTL_reg[12]/NET0131 ,
		\idma_DCTL_reg[13]/NET0131 ,
		_w4937_
	);
	LUT4 #(
		.INIT('h1f00)
	) name890 (
		PM_bdry_sel_pad,
		\idma_DCTL_reg[12]/NET0131 ,
		\idma_DCTL_reg[13]/NET0131 ,
		\idma_WRcyc_reg/NET0131 ,
		_w4938_
	);
	LUT4 #(
		.INIT('h0777)
	) name891 (
		_w4519_,
		_w4887_,
		_w4936_,
		_w4938_,
		_w4939_
	);
	LUT2 #(
		.INIT('h2)
	) name892 (
		_w4873_,
		_w4939_,
		_w4940_
	);
	LUT4 #(
		.INIT('hdf00)
	) name893 (
		_w4067_,
		_w4068_,
		_w4845_,
		_w4940_,
		_w4941_
	);
	LUT4 #(
		.INIT('hbf00)
	) name894 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4092_,
		_w4942_
	);
	LUT2 #(
		.INIT('h2)
	) name895 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w4873_,
		_w4943_
	);
	LUT2 #(
		.INIT('h8)
	) name896 (
		_w4942_,
		_w4943_,
		_w4944_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		_w4941_,
		_w4944_,
		_w4945_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name898 (
		_w4067_,
		_w4068_,
		_w4520_,
		_w4845_,
		_w4946_
	);
	LUT2 #(
		.INIT('h8)
	) name899 (
		\idma_DOVL_reg[3]/NET0131 ,
		_w4946_,
		_w4947_
	);
	LUT3 #(
		.INIT('hac)
	) name900 (
		\bdma_BOVL_reg[3]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4519_,
		_w4948_
	);
	LUT2 #(
		.INIT('h4)
	) name901 (
		_w4946_,
		_w4948_,
		_w4949_
	);
	LUT3 #(
		.INIT('h02)
	) name902 (
		_w4882_,
		_w4949_,
		_w4947_,
		_w4950_
	);
	LUT4 #(
		.INIT('h2400)
	) name903 (
		PM_bdry_sel_pad,
		_w4825_,
		_w4843_,
		_w4950_,
		_w4951_
	);
	LUT3 #(
		.INIT('h53)
	) name904 (
		\bdma_BOVL_reg[2]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4519_,
		_w4952_
	);
	LUT3 #(
		.INIT('h74)
	) name905 (
		\idma_DOVL_reg[2]/NET0131 ,
		_w4946_,
		_w4952_,
		_w4953_
	);
	LUT3 #(
		.INIT('h53)
	) name906 (
		\bdma_BOVL_reg[1]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w4519_,
		_w4954_
	);
	LUT3 #(
		.INIT('h74)
	) name907 (
		\idma_DOVL_reg[1]/NET0131 ,
		_w4946_,
		_w4954_,
		_w4955_
	);
	LUT3 #(
		.INIT('h53)
	) name908 (
		\bdma_BOVL_reg[0]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w4519_,
		_w4956_
	);
	LUT3 #(
		.INIT('h74)
	) name909 (
		\idma_DOVL_reg[0]/NET0131 ,
		_w4946_,
		_w4956_,
		_w4957_
	);
	LUT4 #(
		.INIT('h8000)
	) name910 (
		_w4951_,
		_w4953_,
		_w4955_,
		_w4957_,
		_w4958_
	);
	LUT4 #(
		.INIT('h0080)
	) name911 (
		_w4951_,
		_w4953_,
		_w4955_,
		_w4957_,
		_w4959_
	);
	LUT4 #(
		.INIT('h0800)
	) name912 (
		_w4951_,
		_w4953_,
		_w4955_,
		_w4957_,
		_w4960_
	);
	LUT4 #(
		.INIT('h0008)
	) name913 (
		_w4951_,
		_w4953_,
		_w4955_,
		_w4957_,
		_w4961_
	);
	LUT4 #(
		.INIT('h2000)
	) name914 (
		_w4951_,
		_w4953_,
		_w4955_,
		_w4957_,
		_w4962_
	);
	LUT4 #(
		.INIT('h0020)
	) name915 (
		_w4951_,
		_w4953_,
		_w4955_,
		_w4957_,
		_w4963_
	);
	LUT4 #(
		.INIT('h0200)
	) name916 (
		_w4951_,
		_w4953_,
		_w4955_,
		_w4957_,
		_w4964_
	);
	LUT4 #(
		.INIT('h0002)
	) name917 (
		_w4951_,
		_w4953_,
		_w4955_,
		_w4957_,
		_w4965_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		_w4063_,
		_w4845_,
		_w4966_
	);
	LUT3 #(
		.INIT('h20)
	) name919 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w4967_
	);
	LUT2 #(
		.INIT('h8)
	) name920 (
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w4968_
	);
	LUT4 #(
		.INIT('h5504)
	) name921 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w4090_,
		_w4091_,
		_w4968_,
		_w4969_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w4967_,
		_w4969_,
		_w4970_
	);
	LUT2 #(
		.INIT('h4)
	) name923 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w4971_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_dag_ilm2reg_IL_E_reg[0]/P0001 ,
		_w4972_
	);
	LUT4 #(
		.INIT('h0001)
	) name925 (
		\auctl_R0Sack_reg/NET0131 ,
		\auctl_R1Sack_reg/NET0131 ,
		\auctl_T0Sack_reg/NET0131 ,
		\auctl_T1Sack_reg/NET0131 ,
		_w4973_
	);
	LUT4 #(
		.INIT('h2000)
	) name926 (
		\core_c_dec_Post2_E_reg/P0001 ,
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		_w4972_,
		_w4973_,
		_w4974_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		\core_c_dec_MTIreg_E_reg[4]/P0001 ,
		_w4974_,
		_w4975_
	);
	LUT4 #(
		.INIT('h0045)
	) name928 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w4975_,
		_w4976_
	);
	LUT2 #(
		.INIT('h4)
	) name929 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w4977_
	);
	LUT3 #(
		.INIT('h10)
	) name930 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h1)
	) name931 (
		_w4976_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h8)
	) name932 (
		_w4061_,
		_w4062_,
		_w4980_
	);
	LUT3 #(
		.INIT('h80)
	) name933 (
		\sport1_regs_AUTOreg_DO_reg[5]/NET0131 ,
		_w4061_,
		_w4062_,
		_w4981_
	);
	LUT4 #(
		.INIT('h0100)
	) name934 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		\sport1_txctl_TSreq_reg/NET0131 ,
		_w4982_
	);
	LUT3 #(
		.INIT('h40)
	) name935 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[10]/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w4983_
	);
	LUT3 #(
		.INIT('h04)
	) name936 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w4984_
	);
	LUT4 #(
		.INIT('h0040)
	) name937 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w4985_
	);
	LUT4 #(
		.INIT('h0013)
	) name938 (
		\sport1_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w4983_,
		_w4982_,
		_w4985_,
		_w4986_
	);
	LUT2 #(
		.INIT('h4)
	) name939 (
		_w4981_,
		_w4986_,
		_w4987_
	);
	LUT3 #(
		.INIT('h80)
	) name940 (
		\sport1_regs_AUTOreg_DO_reg[6]/NET0131 ,
		_w4061_,
		_w4062_,
		_w4988_
	);
	LUT3 #(
		.INIT('h40)
	) name941 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[11]/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w4989_
	);
	LUT4 #(
		.INIT('h0040)
	) name942 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[6]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w4990_
	);
	LUT4 #(
		.INIT('h0007)
	) name943 (
		\sport1_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w4982_,
		_w4989_,
		_w4990_,
		_w4991_
	);
	LUT2 #(
		.INIT('h4)
	) name944 (
		_w4988_,
		_w4991_,
		_w4992_
	);
	LUT4 #(
		.INIT('h4044)
	) name945 (
		_w4981_,
		_w4986_,
		_w4988_,
		_w4991_,
		_w4993_
	);
	LUT3 #(
		.INIT('h80)
	) name946 (
		\sport1_regs_AUTOreg_DO_reg[4]/NET0131 ,
		_w4061_,
		_w4062_,
		_w4994_
	);
	LUT3 #(
		.INIT('h40)
	) name947 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[9]/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w4995_
	);
	LUT4 #(
		.INIT('h0040)
	) name948 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w4996_
	);
	LUT4 #(
		.INIT('h0007)
	) name949 (
		\sport1_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w4982_,
		_w4995_,
		_w4996_,
		_w4997_
	);
	LUT2 #(
		.INIT('h4)
	) name950 (
		_w4994_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h8)
	) name951 (
		_w4993_,
		_w4998_,
		_w4999_
	);
	LUT3 #(
		.INIT('he0)
	) name952 (
		_w4976_,
		_w4978_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('h4)
	) name953 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_dag_ilm2reg_IL_E_reg[0]/P0001 ,
		_w5001_
	);
	LUT4 #(
		.INIT('h8000)
	) name954 (
		\core_c_dec_Post2_E_reg/P0001 ,
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		_w4973_,
		_w5001_,
		_w5002_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		\core_c_dec_MTIreg_E_reg[7]/P0001 ,
		_w5002_,
		_w5003_
	);
	LUT4 #(
		.INIT('h0045)
	) name956 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w5003_,
		_w5004_
	);
	LUT2 #(
		.INIT('h8)
	) name957 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w5005_
	);
	LUT3 #(
		.INIT('h20)
	) name958 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w5005_,
		_w5006_
	);
	LUT2 #(
		.INIT('h1)
	) name959 (
		_w5004_,
		_w5006_,
		_w5007_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name960 (
		_w4981_,
		_w4986_,
		_w4988_,
		_w4991_,
		_w5008_
	);
	LUT2 #(
		.INIT('h4)
	) name961 (
		_w4998_,
		_w5008_,
		_w5009_
	);
	LUT3 #(
		.INIT('he0)
	) name962 (
		_w5004_,
		_w5006_,
		_w5009_,
		_w5010_
	);
	LUT4 #(
		.INIT('h8000)
	) name963 (
		\core_c_dec_Post2_E_reg/P0001 ,
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		_w4972_,
		_w4973_,
		_w5011_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		\core_c_dec_MTIreg_E_reg[6]/P0001 ,
		_w5011_,
		_w5012_
	);
	LUT4 #(
		.INIT('h0045)
	) name965 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w5012_,
		_w5013_
	);
	LUT3 #(
		.INIT('h20)
	) name966 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w4977_,
		_w5014_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		_w5013_,
		_w5014_,
		_w5015_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		_w4998_,
		_w5008_,
		_w5016_
	);
	LUT3 #(
		.INIT('he0)
	) name969 (
		_w5013_,
		_w5014_,
		_w5016_,
		_w5017_
	);
	LUT4 #(
		.INIT('h2000)
	) name970 (
		\core_c_dec_Post2_E_reg/P0001 ,
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		_w4973_,
		_w5001_,
		_w5018_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		\core_c_dec_MTIreg_E_reg[5]/P0001 ,
		_w5018_,
		_w5019_
	);
	LUT4 #(
		.INIT('h0045)
	) name972 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w5019_,
		_w5020_
	);
	LUT3 #(
		.INIT('h10)
	) name973 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w5005_,
		_w5021_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		_w5020_,
		_w5021_,
		_w5022_
	);
	LUT2 #(
		.INIT('h2)
	) name975 (
		_w4993_,
		_w4998_,
		_w5023_
	);
	LUT3 #(
		.INIT('he0)
	) name976 (
		_w5020_,
		_w5021_,
		_w5023_,
		_w5024_
	);
	LUT4 #(
		.INIT('h0001)
	) name977 (
		_w5000_,
		_w5010_,
		_w5017_,
		_w5024_,
		_w5025_
	);
	LUT2 #(
		.INIT('h1)
	) name978 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w5026_
	);
	LUT2 #(
		.INIT('h8)
	) name979 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w5027_
	);
	LUT4 #(
		.INIT('h0001)
	) name980 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w5028_
	);
	LUT3 #(
		.INIT('h80)
	) name981 (
		_w5026_,
		_w5027_,
		_w5028_,
		_w5029_
	);
	LUT4 #(
		.INIT('h1555)
	) name982 (
		_w4967_,
		_w5026_,
		_w5027_,
		_w5028_,
		_w5030_
	);
	LUT3 #(
		.INIT('h53)
	) name983 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w5030_,
		_w5031_
	);
	LUT3 #(
		.INIT('h53)
	) name984 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w5030_,
		_w5032_
	);
	LUT2 #(
		.INIT('h8)
	) name985 (
		_w5031_,
		_w5032_,
		_w5033_
	);
	LUT3 #(
		.INIT('he0)
	) name986 (
		_w4976_,
		_w4978_,
		_w5033_,
		_w5034_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		_w5031_,
		_w5032_,
		_w5035_
	);
	LUT3 #(
		.INIT('he0)
	) name988 (
		_w5004_,
		_w5006_,
		_w5035_,
		_w5036_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		_w5031_,
		_w5032_,
		_w5037_
	);
	LUT3 #(
		.INIT('he0)
	) name990 (
		_w5013_,
		_w5014_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h2)
	) name991 (
		_w5031_,
		_w5032_,
		_w5039_
	);
	LUT3 #(
		.INIT('he0)
	) name992 (
		_w5020_,
		_w5021_,
		_w5039_,
		_w5040_
	);
	LUT4 #(
		.INIT('h0001)
	) name993 (
		_w5034_,
		_w5036_,
		_w5038_,
		_w5040_,
		_w5041_
	);
	LUT3 #(
		.INIT('h1b)
	) name994 (
		_w4063_,
		_w5025_,
		_w5041_,
		_w5042_
	);
	LUT4 #(
		.INIT('haa08)
	) name995 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w4090_,
		_w4091_,
		_w4968_,
		_w5043_
	);
	LUT2 #(
		.INIT('h2)
	) name996 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w5044_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w5045_
	);
	LUT4 #(
		.INIT('h0002)
	) name998 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w5046_
	);
	LUT2 #(
		.INIT('h8)
	) name999 (
		_w5045_,
		_w5046_,
		_w5047_
	);
	LUT3 #(
		.INIT('h80)
	) name1000 (
		_w5044_,
		_w5045_,
		_w5046_,
		_w5048_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		_w5043_,
		_w5048_,
		_w5049_
	);
	LUT4 #(
		.INIT('h001b)
	) name1002 (
		_w4063_,
		_w5025_,
		_w5041_,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('h2)
	) name1003 (
		_w4970_,
		_w5050_,
		_w5051_
	);
	LUT3 #(
		.INIT('h80)
	) name1004 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		_w5052_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w5053_
	);
	LUT4 #(
		.INIT('h8000)
	) name1006 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		_w5054_
	);
	LUT2 #(
		.INIT('h2)
	) name1007 (
		\memc_Dwrite_E_reg/NET0131 ,
		\memc_EXTC_E_reg/NET0131 ,
		_w5055_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1008 (
		_w5053_,
		_w5052_,
		_w5054_,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h4)
	) name1009 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w5056_,
		_w5057_
	);
	LUT4 #(
		.INIT('h00ea)
	) name1010 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w5057_,
		_w5058_
	);
	LUT2 #(
		.INIT('h4)
	) name1011 (
		_w4104_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w5060_
	);
	LUT3 #(
		.INIT('h10)
	) name1013 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w5060_,
		_w5061_
	);
	LUT2 #(
		.INIT('h4)
	) name1014 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_Post1_E_reg/P0001 ,
		_w5062_
	);
	LUT4 #(
		.INIT('h1000)
	) name1015 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w4973_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h1)
	) name1016 (
		\core_c_dec_MTIreg_E_reg[0]/P0001 ,
		_w5063_,
		_w5064_
	);
	LUT4 #(
		.INIT('h0045)
	) name1017 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w5064_,
		_w5065_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w5061_,
		_w5065_,
		_w5066_
	);
	LUT4 #(
		.INIT('h0400)
	) name1019 (
		_w4981_,
		_w4986_,
		_w4988_,
		_w4991_,
		_w5067_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		_w4998_,
		_w5067_,
		_w5068_
	);
	LUT4 #(
		.INIT('h0155)
	) name1021 (
		_w4063_,
		_w5061_,
		_w5065_,
		_w5068_,
		_w5069_
	);
	LUT3 #(
		.INIT('h20)
	) name1022 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w5060_,
		_w5070_
	);
	LUT2 #(
		.INIT('h4)
	) name1023 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w5071_
	);
	LUT4 #(
		.INIT('h1555)
	) name1024 (
		\core_c_dec_MTIreg_E_reg[2]/P0001 ,
		_w4973_,
		_w5062_,
		_w5071_,
		_w5072_
	);
	LUT4 #(
		.INIT('h0045)
	) name1025 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w5072_,
		_w5073_
	);
	LUT2 #(
		.INIT('h1)
	) name1026 (
		_w5070_,
		_w5073_,
		_w5074_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1027 (
		_w4981_,
		_w4986_,
		_w4988_,
		_w4991_,
		_w5075_
	);
	LUT2 #(
		.INIT('h8)
	) name1028 (
		_w4998_,
		_w5075_,
		_w5076_
	);
	LUT3 #(
		.INIT('he0)
	) name1029 (
		_w5070_,
		_w5073_,
		_w5076_,
		_w5077_
	);
	LUT2 #(
		.INIT('h2)
	) name1030 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w5078_
	);
	LUT3 #(
		.INIT('h10)
	) name1031 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w5078_,
		_w5079_
	);
	LUT4 #(
		.INIT('h2000)
	) name1032 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w4973_,
		_w5062_,
		_w5080_
	);
	LUT2 #(
		.INIT('h1)
	) name1033 (
		\core_c_dec_MTIreg_E_reg[1]/P0001 ,
		_w5080_,
		_w5081_
	);
	LUT4 #(
		.INIT('h0045)
	) name1034 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w5081_,
		_w5082_
	);
	LUT2 #(
		.INIT('h1)
	) name1035 (
		_w5079_,
		_w5082_,
		_w5083_
	);
	LUT2 #(
		.INIT('he)
	) name1036 (
		_w5079_,
		_w5082_,
		_w5084_
	);
	LUT2 #(
		.INIT('h4)
	) name1037 (
		_w4998_,
		_w5067_,
		_w5085_
	);
	LUT3 #(
		.INIT('he0)
	) name1038 (
		_w5079_,
		_w5082_,
		_w5085_,
		_w5086_
	);
	LUT3 #(
		.INIT('h20)
	) name1039 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w5078_,
		_w5087_
	);
	LUT2 #(
		.INIT('h8)
	) name1040 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w5088_
	);
	LUT4 #(
		.INIT('h1555)
	) name1041 (
		\core_c_dec_MTIreg_E_reg[3]/P0001 ,
		_w4973_,
		_w5062_,
		_w5088_,
		_w5089_
	);
	LUT4 #(
		.INIT('h0045)
	) name1042 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		_w5087_,
		_w5090_,
		_w5091_
	);
	LUT2 #(
		.INIT('he)
	) name1044 (
		_w5087_,
		_w5090_,
		_w5092_
	);
	LUT2 #(
		.INIT('h4)
	) name1045 (
		_w4998_,
		_w5075_,
		_w5093_
	);
	LUT3 #(
		.INIT('he0)
	) name1046 (
		_w5087_,
		_w5090_,
		_w5093_,
		_w5094_
	);
	LUT4 #(
		.INIT('h0100)
	) name1047 (
		_w5086_,
		_w5094_,
		_w5077_,
		_w5069_,
		_w5095_
	);
	LUT2 #(
		.INIT('h2)
	) name1048 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w5096_
	);
	LUT3 #(
		.INIT('he0)
	) name1049 (
		_w5079_,
		_w5082_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h1)
	) name1050 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w5098_
	);
	LUT3 #(
		.INIT('he0)
	) name1051 (
		_w5061_,
		_w5065_,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h4)
	) name1052 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w5100_
	);
	LUT3 #(
		.INIT('he0)
	) name1053 (
		_w5070_,
		_w5073_,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w5102_
	);
	LUT3 #(
		.INIT('he0)
	) name1055 (
		_w5087_,
		_w5090_,
		_w5102_,
		_w5103_
	);
	LUT4 #(
		.INIT('h0001)
	) name1056 (
		_w5097_,
		_w5099_,
		_w5101_,
		_w5103_,
		_w5104_
	);
	LUT3 #(
		.INIT('h13)
	) name1057 (
		_w4063_,
		_w5095_,
		_w5104_,
		_w5105_
	);
	LUT2 #(
		.INIT('h1)
	) name1058 (
		_w5042_,
		_w5105_,
		_w5106_
	);
	LUT2 #(
		.INIT('h4)
	) name1059 (
		\core_c_dec_Post1_E_reg/P0001 ,
		_w4973_,
		_w5107_
	);
	LUT3 #(
		.INIT('ha8)
	) name1060 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w4967_,
		_w4969_,
		_w5108_
	);
	LUT4 #(
		.INIT('ha080)
	) name1061 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w4967_,
		_w5107_,
		_w4969_,
		_w5109_
	);
	LUT4 #(
		.INIT('h00a8)
	) name1062 (
		_w5059_,
		_w5042_,
		_w5105_,
		_w5109_,
		_w5110_
	);
	LUT3 #(
		.INIT('h54)
	) name1063 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w4967_,
		_w4969_,
		_w5111_
	);
	LUT4 #(
		.INIT('h0f01)
	) name1064 (
		_w4063_,
		_w4845_,
		_w5107_,
		_w5111_,
		_w5112_
	);
	LUT4 #(
		.INIT('h1300)
	) name1065 (
		_w4063_,
		_w5095_,
		_w5104_,
		_w5112_,
		_w5113_
	);
	LUT3 #(
		.INIT('h04)
	) name1066 (
		_w4104_,
		_w5058_,
		_w4970_,
		_w5114_
	);
	LUT4 #(
		.INIT('h1b00)
	) name1067 (
		_w4063_,
		_w5025_,
		_w5041_,
		_w5114_,
		_w5115_
	);
	LUT3 #(
		.INIT('h23)
	) name1068 (
		_w5105_,
		_w5113_,
		_w5115_,
		_w5116_
	);
	LUT4 #(
		.INIT('hba00)
	) name1069 (
		_w4966_,
		_w5051_,
		_w5110_,
		_w5116_,
		_w5117_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		_w5118_
	);
	LUT2 #(
		.INIT('h1)
	) name1071 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w5119_
	);
	LUT3 #(
		.INIT('h01)
	) name1072 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w5120_
	);
	LUT2 #(
		.INIT('h1)
	) name1073 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w5121_
	);
	LUT3 #(
		.INIT('h01)
	) name1074 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w5122_
	);
	LUT2 #(
		.INIT('h8)
	) name1075 (
		_w5120_,
		_w5122_,
		_w5123_
	);
	LUT3 #(
		.INIT('h80)
	) name1076 (
		_w5118_,
		_w5120_,
		_w5122_,
		_w5124_
	);
	LUT2 #(
		.INIT('h1)
	) name1077 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w5125_
	);
	LUT3 #(
		.INIT('h01)
	) name1078 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w5126_
	);
	LUT4 #(
		.INIT('h8000)
	) name1079 (
		_w5118_,
		_w5120_,
		_w5122_,
		_w5126_,
		_w5127_
	);
	LUT2 #(
		.INIT('h1)
	) name1080 (
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w5128_
	);
	LUT2 #(
		.INIT('h8)
	) name1081 (
		_w5127_,
		_w5128_,
		_w5129_
	);
	LUT3 #(
		.INIT('h2a)
	) name1082 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		_w5127_,
		_w5128_,
		_w5130_
	);
	LUT3 #(
		.INIT('h01)
	) name1083 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		_w5131_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		_w5132_
	);
	LUT4 #(
		.INIT('h0001)
	) name1085 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w5133_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w5133_,
		_w5134_
	);
	LUT3 #(
		.INIT('h40)
	) name1087 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w5132_,
		_w5133_,
		_w5135_
	);
	LUT4 #(
		.INIT('h2333)
	) name1088 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w5131_,
		_w5132_,
		_w5133_,
		_w5136_
	);
	LUT3 #(
		.INIT('h23)
	) name1089 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w5132_,
		_w5133_,
		_w5137_
	);
	LUT3 #(
		.INIT('he0)
	) name1090 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		_w5138_
	);
	LUT3 #(
		.INIT('ha8)
	) name1091 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w5139_
	);
	LUT4 #(
		.INIT('h0777)
	) name1092 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w5140_
	);
	LUT3 #(
		.INIT('h10)
	) name1093 (
		_w5139_,
		_w5138_,
		_w5140_,
		_w5141_
	);
	LUT2 #(
		.INIT('h8)
	) name1094 (
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w5142_
	);
	LUT4 #(
		.INIT('h153f)
	) name1095 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w5143_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1096 (
		_w5120_,
		_w5121_,
		_w5142_,
		_w5143_,
		_w5144_
	);
	LUT4 #(
		.INIT('h1000)
	) name1097 (
		_w5136_,
		_w5137_,
		_w5141_,
		_w5144_,
		_w5145_
	);
	LUT4 #(
		.INIT('hd540)
	) name1098 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		_w5124_,
		_w5125_,
		_w5128_,
		_w5146_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1099 (
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w5130_,
		_w5145_,
		_w5146_,
		_w5147_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		_w5148_
	);
	LUT3 #(
		.INIT('h01)
	) name1101 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w5149_
	);
	LUT4 #(
		.INIT('h0001)
	) name1102 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		_w5150_
	);
	LUT2 #(
		.INIT('h8)
	) name1103 (
		_w5125_,
		_w5150_,
		_w5151_
	);
	LUT3 #(
		.INIT('h80)
	) name1104 (
		_w5118_,
		_w5125_,
		_w5150_,
		_w5152_
	);
	LUT4 #(
		.INIT('h4000)
	) name1105 (
		_w5130_,
		_w5145_,
		_w5146_,
		_w5152_,
		_w5153_
	);
	LUT4 #(
		.INIT('h070f)
	) name1106 (
		_w5120_,
		_w5122_,
		_w5147_,
		_w5153_,
		_w5154_
	);
	LUT2 #(
		.INIT('h2)
	) name1107 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		_w5154_,
		_w5155_
	);
	LUT4 #(
		.INIT('hc0e2)
	) name1108 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5154_,
		_w5156_
	);
	LUT2 #(
		.INIT('h6)
	) name1109 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5157_
	);
	LUT4 #(
		.INIT('h0040)
	) name1110 (
		_w5130_,
		_w5145_,
		_w5146_,
		_w5150_,
		_w5158_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1111 (
		_w5127_,
		_w5130_,
		_w5145_,
		_w5146_,
		_w5159_
	);
	LUT3 #(
		.INIT('h02)
	) name1112 (
		\core_dag_ilm1reg_I_reg[3]/NET0131 ,
		_w5158_,
		_w5159_,
		_w5160_
	);
	LUT4 #(
		.INIT('h0008)
	) name1113 (
		\core_dag_ilm1reg_I_reg[3]/NET0131 ,
		\core_dag_ilm1reg_M_reg[3]/NET0131 ,
		_w5158_,
		_w5159_,
		_w5161_
	);
	LUT4 #(
		.INIT('h3331)
	) name1114 (
		\core_dag_ilm1reg_I_reg[3]/NET0131 ,
		\core_dag_ilm1reg_M_reg[3]/NET0131 ,
		_w5158_,
		_w5159_,
		_w5162_
	);
	LUT4 #(
		.INIT('hccc6)
	) name1115 (
		\core_dag_ilm1reg_I_reg[3]/NET0131 ,
		\core_dag_ilm1reg_M_reg[3]/NET0131 ,
		_w5158_,
		_w5159_,
		_w5163_
	);
	LUT2 #(
		.INIT('h9)
	) name1116 (
		_w5157_,
		_w5163_,
		_w5164_
	);
	LUT4 #(
		.INIT('h0040)
	) name1117 (
		_w5130_,
		_w5145_,
		_w5146_,
		_w5149_,
		_w5165_
	);
	LUT2 #(
		.INIT('h4)
	) name1118 (
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w5127_,
		_w5166_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1119 (
		_w5130_,
		_w5145_,
		_w5146_,
		_w5166_,
		_w5167_
	);
	LUT3 #(
		.INIT('h02)
	) name1120 (
		\core_dag_ilm1reg_I_reg[2]/NET0131 ,
		_w5165_,
		_w5167_,
		_w5168_
	);
	LUT2 #(
		.INIT('h6)
	) name1121 (
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5169_
	);
	LUT3 #(
		.INIT('h71)
	) name1122 (
		\core_dag_ilm1reg_M_reg[2]/NET0131 ,
		_w5168_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h2)
	) name1123 (
		_w5164_,
		_w5170_,
		_w5171_
	);
	LUT2 #(
		.INIT('h4)
	) name1124 (
		_w5164_,
		_w5170_,
		_w5172_
	);
	LUT4 #(
		.INIT('h0040)
	) name1125 (
		_w5130_,
		_w5145_,
		_w5146_,
		_w5148_,
		_w5173_
	);
	LUT4 #(
		.INIT('ha222)
	) name1126 (
		\core_dag_ilm1reg_I_reg[1]/NET0131 ,
		_w5129_,
		_w5145_,
		_w5146_,
		_w5174_
	);
	LUT2 #(
		.INIT('h4)
	) name1127 (
		_w5173_,
		_w5174_,
		_w5175_
	);
	LUT2 #(
		.INIT('h6)
	) name1128 (
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5176_
	);
	LUT4 #(
		.INIT('hdf45)
	) name1129 (
		\core_dag_ilm1reg_M_reg[1]/NET0131 ,
		_w5173_,
		_w5174_,
		_w5176_,
		_w5177_
	);
	LUT4 #(
		.INIT('hccc6)
	) name1130 (
		\core_dag_ilm1reg_I_reg[2]/NET0131 ,
		\core_dag_ilm1reg_M_reg[2]/NET0131 ,
		_w5165_,
		_w5167_,
		_w5178_
	);
	LUT3 #(
		.INIT('h21)
	) name1131 (
		_w5169_,
		_w5177_,
		_w5178_,
		_w5179_
	);
	LUT3 #(
		.INIT('h48)
	) name1132 (
		_w5169_,
		_w5177_,
		_w5178_,
		_w5180_
	);
	LUT4 #(
		.INIT('h8000)
	) name1133 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		_w5129_,
		_w5145_,
		_w5146_,
		_w5181_
	);
	LUT4 #(
		.INIT('h002a)
	) name1134 (
		\core_dag_ilm1reg_I_reg[0]/NET0131 ,
		_w5148_,
		_w5167_,
		_w5181_,
		_w5182_
	);
	LUT2 #(
		.INIT('h6)
	) name1135 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5183_
	);
	LUT3 #(
		.INIT('h8e)
	) name1136 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w5182_,
		_w5183_,
		_w5184_
	);
	LUT3 #(
		.INIT('h9a)
	) name1137 (
		\core_dag_ilm1reg_M_reg[1]/NET0131 ,
		_w5173_,
		_w5174_,
		_w5185_
	);
	LUT4 #(
		.INIT('h9a65)
	) name1138 (
		\core_dag_ilm1reg_M_reg[1]/NET0131 ,
		_w5173_,
		_w5174_,
		_w5176_,
		_w5186_
	);
	LUT4 #(
		.INIT('h0071)
	) name1139 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w5182_,
		_w5183_,
		_w5186_,
		_w5187_
	);
	LUT4 #(
		.INIT('h8e00)
	) name1140 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w5182_,
		_w5183_,
		_w5186_,
		_w5188_
	);
	LUT2 #(
		.INIT('h6)
	) name1141 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w5182_,
		_w5189_
	);
	LUT3 #(
		.INIT('h69)
	) name1142 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w5182_,
		_w5183_,
		_w5190_
	);
	LUT4 #(
		.INIT('h0609)
	) name1143 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5182_,
		_w5191_
	);
	LUT4 #(
		.INIT('h5440)
	) name1144 (
		_w5180_,
		_w5184_,
		_w5186_,
		_w5191_,
		_w5192_
	);
	LUT4 #(
		.INIT('h4445)
	) name1145 (
		_w5171_,
		_w5172_,
		_w5179_,
		_w5192_,
		_w5193_
	);
	LUT4 #(
		.INIT('h1000)
	) name1146 (
		_w5130_,
		_w5131_,
		_w5145_,
		_w5146_,
		_w5194_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1147 (
		_w5124_,
		_w5130_,
		_w5145_,
		_w5146_,
		_w5195_
	);
	LUT4 #(
		.INIT('h0002)
	) name1148 (
		\core_dag_ilm1reg_I_reg[6]/NET0131 ,
		_w5195_,
		_w5158_,
		_w5194_,
		_w5196_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		\core_dag_ilm1reg_M_reg[6]/NET0131 ,
		_w5196_,
		_w5197_
	);
	LUT2 #(
		.INIT('h6)
	) name1150 (
		\core_dag_ilm1reg_M_reg[6]/NET0131 ,
		_w5196_,
		_w5198_
	);
	LUT2 #(
		.INIT('h6)
	) name1151 (
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5199_
	);
	LUT3 #(
		.INIT('h69)
	) name1152 (
		\core_dag_ilm1reg_M_reg[6]/NET0131 ,
		_w5196_,
		_w5199_,
		_w5200_
	);
	LUT4 #(
		.INIT('h0040)
	) name1153 (
		_w5130_,
		_w5145_,
		_w5146_,
		_w5151_,
		_w5201_
	);
	LUT4 #(
		.INIT('h008a)
	) name1154 (
		\core_dag_ilm1reg_I_reg[5]/NET0131 ,
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w5195_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('h6)
	) name1155 (
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5203_
	);
	LUT3 #(
		.INIT('h71)
	) name1156 (
		\core_dag_ilm1reg_M_reg[5]/NET0131 ,
		_w5202_,
		_w5203_,
		_w5204_
	);
	LUT2 #(
		.INIT('h4)
	) name1157 (
		_w5200_,
		_w5204_,
		_w5205_
	);
	LUT4 #(
		.INIT('h2333)
	) name1158 (
		_w5130_,
		_w5135_,
		_w5145_,
		_w5146_,
		_w5206_
	);
	LUT3 #(
		.INIT('ha8)
	) name1159 (
		\core_dag_ilm1reg_I_reg[7]/NET0131 ,
		_w5153_,
		_w5206_,
		_w5207_
	);
	LUT4 #(
		.INIT('h1113)
	) name1160 (
		\core_dag_ilm1reg_I_reg[7]/NET0131 ,
		\core_dag_ilm1reg_M_reg[7]/NET0131 ,
		_w5153_,
		_w5206_,
		_w5208_
	);
	LUT4 #(
		.INIT('h8880)
	) name1161 (
		\core_dag_ilm1reg_I_reg[7]/NET0131 ,
		\core_dag_ilm1reg_M_reg[7]/NET0131 ,
		_w5153_,
		_w5206_,
		_w5209_
	);
	LUT4 #(
		.INIT('h666c)
	) name1162 (
		\core_dag_ilm1reg_I_reg[7]/NET0131 ,
		\core_dag_ilm1reg_M_reg[7]/NET0131 ,
		_w5153_,
		_w5206_,
		_w5210_
	);
	LUT2 #(
		.INIT('h6)
	) name1163 (
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5211_
	);
	LUT2 #(
		.INIT('h9)
	) name1164 (
		_w5210_,
		_w5211_,
		_w5212_
	);
	LUT3 #(
		.INIT('h71)
	) name1165 (
		\core_dag_ilm1reg_M_reg[6]/NET0131 ,
		_w5196_,
		_w5199_,
		_w5213_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1166 (
		_w5200_,
		_w5204_,
		_w5212_,
		_w5213_,
		_w5214_
	);
	LUT2 #(
		.INIT('h4)
	) name1167 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		_w5150_,
		_w5215_
	);
	LUT4 #(
		.INIT('h0040)
	) name1168 (
		_w5130_,
		_w5145_,
		_w5146_,
		_w5215_,
		_w5216_
	);
	LUT4 #(
		.INIT('h002a)
	) name1169 (
		\core_dag_ilm1reg_I_reg[4]/NET0131 ,
		_w5125_,
		_w5195_,
		_w5216_,
		_w5217_
	);
	LUT2 #(
		.INIT('h6)
	) name1170 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5218_
	);
	LUT3 #(
		.INIT('h71)
	) name1171 (
		\core_dag_ilm1reg_M_reg[4]/NET0131 ,
		_w5217_,
		_w5218_,
		_w5219_
	);
	LUT2 #(
		.INIT('h6)
	) name1172 (
		\core_dag_ilm1reg_M_reg[5]/NET0131 ,
		_w5202_,
		_w5220_
	);
	LUT3 #(
		.INIT('h69)
	) name1173 (
		\core_dag_ilm1reg_M_reg[5]/NET0131 ,
		_w5202_,
		_w5203_,
		_w5221_
	);
	LUT3 #(
		.INIT('h71)
	) name1174 (
		\core_dag_ilm1reg_M_reg[3]/NET0131 ,
		_w5160_,
		_w5157_,
		_w5222_
	);
	LUT2 #(
		.INIT('h6)
	) name1175 (
		\core_dag_ilm1reg_M_reg[4]/NET0131 ,
		_w5217_,
		_w5223_
	);
	LUT3 #(
		.INIT('h69)
	) name1176 (
		\core_dag_ilm1reg_M_reg[4]/NET0131 ,
		_w5217_,
		_w5218_,
		_w5224_
	);
	LUT2 #(
		.INIT('h2)
	) name1177 (
		_w5222_,
		_w5224_,
		_w5225_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1178 (
		_w5219_,
		_w5221_,
		_w5222_,
		_w5224_,
		_w5226_
	);
	LUT2 #(
		.INIT('h8)
	) name1179 (
		_w5214_,
		_w5226_,
		_w5227_
	);
	LUT2 #(
		.INIT('h4)
	) name1180 (
		_w5222_,
		_w5224_,
		_w5228_
	);
	LUT4 #(
		.INIT('hb2bb)
	) name1181 (
		_w5219_,
		_w5221_,
		_w5222_,
		_w5224_,
		_w5229_
	);
	LUT2 #(
		.INIT('h2)
	) name1182 (
		_w5200_,
		_w5204_,
		_w5230_
	);
	LUT4 #(
		.INIT('hdf0d)
	) name1183 (
		_w5200_,
		_w5204_,
		_w5212_,
		_w5213_,
		_w5231_
	);
	LUT3 #(
		.INIT('hd0)
	) name1184 (
		_w5214_,
		_w5229_,
		_w5231_,
		_w5232_
	);
	LUT4 #(
		.INIT('h2333)
	) name1185 (
		_w5130_,
		_w5134_,
		_w5145_,
		_w5146_,
		_w5233_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1186 (
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w5153_,
		_w5233_,
		_w5234_
	);
	LUT2 #(
		.INIT('h2)
	) name1187 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		_w5234_,
		_w5235_
	);
	LUT3 #(
		.INIT('h31)
	) name1188 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w5234_,
		_w5236_
	);
	LUT3 #(
		.INIT('hc6)
	) name1189 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w5234_,
		_w5237_
	);
	LUT2 #(
		.INIT('h6)
	) name1190 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5238_
	);
	LUT4 #(
		.INIT('hc639)
	) name1191 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w5234_,
		_w5238_,
		_w5239_
	);
	LUT4 #(
		.INIT('h4555)
	) name1192 (
		_w5123_,
		_w5130_,
		_w5145_,
		_w5146_,
		_w5240_
	);
	LUT4 #(
		.INIT('haa20)
	) name1193 (
		\core_dag_ilm1reg_I_reg[8]/NET0131 ,
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		_w5153_,
		_w5240_,
		_w5241_
	);
	LUT2 #(
		.INIT('h8)
	) name1194 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('h1)
	) name1195 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w5241_,
		_w5243_
	);
	LUT2 #(
		.INIT('h6)
	) name1196 (
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5244_
	);
	LUT3 #(
		.INIT('h71)
	) name1197 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w5241_,
		_w5244_,
		_w5245_
	);
	LUT3 #(
		.INIT('h71)
	) name1198 (
		\core_dag_ilm1reg_M_reg[7]/NET0131 ,
		_w5207_,
		_w5211_,
		_w5246_
	);
	LUT2 #(
		.INIT('h6)
	) name1199 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w5241_,
		_w5247_
	);
	LUT3 #(
		.INIT('h69)
	) name1200 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w5241_,
		_w5244_,
		_w5248_
	);
	LUT2 #(
		.INIT('h2)
	) name1201 (
		_w5246_,
		_w5248_,
		_w5249_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name1202 (
		_w5239_,
		_w5245_,
		_w5246_,
		_w5248_,
		_w5250_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1203 (
		_w5193_,
		_w5227_,
		_w5232_,
		_w5250_,
		_w5251_
	);
	LUT4 #(
		.INIT('hf731)
	) name1204 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w5234_,
		_w5238_,
		_w5252_
	);
	LUT4 #(
		.INIT('h2333)
	) name1205 (
		_w5130_,
		_w5133_,
		_w5145_,
		_w5146_,
		_w5253_
	);
	LUT4 #(
		.INIT('haa80)
	) name1206 (
		\core_dag_ilm1reg_I_reg[10]/NET0131 ,
		_w5122_,
		_w5153_,
		_w5253_,
		_w5254_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		_w5254_,
		_w5255_
	);
	LUT2 #(
		.INIT('h8)
	) name1208 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		_w5254_,
		_w5256_
	);
	LUT2 #(
		.INIT('h6)
	) name1209 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		_w5254_,
		_w5257_
	);
	LUT2 #(
		.INIT('h6)
	) name1210 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5258_
	);
	LUT3 #(
		.INIT('h69)
	) name1211 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		_w5254_,
		_w5258_,
		_w5259_
	);
	LUT2 #(
		.INIT('h2)
	) name1212 (
		_w5252_,
		_w5259_,
		_w5260_
	);
	LUT3 #(
		.INIT('h71)
	) name1213 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		_w5254_,
		_w5258_,
		_w5261_
	);
	LUT4 #(
		.INIT('h0001)
	) name1214 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w5262_
	);
	LUT4 #(
		.INIT('h8000)
	) name1215 (
		_w5118_,
		_w5125_,
		_w5150_,
		_w5262_,
		_w5263_
	);
	LUT4 #(
		.INIT('h0040)
	) name1216 (
		_w5130_,
		_w5145_,
		_w5146_,
		_w5263_,
		_w5264_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1217 (
		_w5119_,
		_w5130_,
		_w5145_,
		_w5146_,
		_w5265_
	);
	LUT4 #(
		.INIT('h080a)
	) name1218 (
		\core_dag_ilm1reg_I_reg[11]/NET0131 ,
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		_w5264_,
		_w5265_,
		_w5266_
	);
	LUT2 #(
		.INIT('h6)
	) name1219 (
		\core_dag_ilm1reg_M_reg[11]/NET0131 ,
		_w5266_,
		_w5267_
	);
	LUT2 #(
		.INIT('h6)
	) name1220 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5268_
	);
	LUT3 #(
		.INIT('h69)
	) name1221 (
		\core_dag_ilm1reg_M_reg[11]/NET0131 ,
		_w5266_,
		_w5268_,
		_w5269_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1222 (
		_w5252_,
		_w5259_,
		_w5261_,
		_w5269_,
		_w5270_
	);
	LUT2 #(
		.INIT('h4)
	) name1223 (
		_w5261_,
		_w5269_,
		_w5271_
	);
	LUT2 #(
		.INIT('h4)
	) name1224 (
		_w5252_,
		_w5259_,
		_w5272_
	);
	LUT2 #(
		.INIT('h4)
	) name1225 (
		_w5246_,
		_w5248_,
		_w5273_
	);
	LUT4 #(
		.INIT('hd4dd)
	) name1226 (
		_w5239_,
		_w5245_,
		_w5246_,
		_w5248_,
		_w5274_
	);
	LUT4 #(
		.INIT('h1311)
	) name1227 (
		_w5270_,
		_w5271_,
		_w5272_,
		_w5274_,
		_w5275_
	);
	LUT3 #(
		.INIT('hc6)
	) name1228 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w5154_,
		_w5276_
	);
	LUT4 #(
		.INIT('h2000)
	) name1229 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		_w5130_,
		_w5145_,
		_w5146_,
		_w5277_
	);
	LUT4 #(
		.INIT('h0002)
	) name1230 (
		\core_dag_ilm1reg_I_reg[12]/NET0131 ,
		_w5264_,
		_w5265_,
		_w5277_,
		_w5278_
	);
	LUT2 #(
		.INIT('h6)
	) name1231 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5279_
	);
	LUT3 #(
		.INIT('h8e)
	) name1232 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w5278_,
		_w5279_,
		_w5280_
	);
	LUT3 #(
		.INIT('h71)
	) name1233 (
		\core_dag_ilm1reg_M_reg[11]/NET0131 ,
		_w5266_,
		_w5268_,
		_w5281_
	);
	LUT2 #(
		.INIT('h6)
	) name1234 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w5278_,
		_w5282_
	);
	LUT3 #(
		.INIT('h69)
	) name1235 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w5278_,
		_w5279_,
		_w5283_
	);
	LUT2 #(
		.INIT('h2)
	) name1236 (
		_w5281_,
		_w5283_,
		_w5284_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1237 (
		_w5276_,
		_w5280_,
		_w5281_,
		_w5283_,
		_w5285_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1238 (
		_w5251_,
		_w5270_,
		_w5275_,
		_w5285_,
		_w5286_
	);
	LUT2 #(
		.INIT('h4)
	) name1239 (
		_w5281_,
		_w5283_,
		_w5287_
	);
	LUT4 #(
		.INIT('hb2bb)
	) name1240 (
		_w5276_,
		_w5280_,
		_w5281_,
		_w5283_,
		_w5288_
	);
	LUT3 #(
		.INIT('h65)
	) name1241 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w5289_
	);
	LUT2 #(
		.INIT('h9)
	) name1242 (
		_w5276_,
		_w5280_,
		_w5290_
	);
	LUT4 #(
		.INIT('h008f)
	) name1243 (
		_w5251_,
		_w5270_,
		_w5275_,
		_w5284_,
		_w5291_
	);
	LUT3 #(
		.INIT('h36)
	) name1244 (
		_w5287_,
		_w5290_,
		_w5291_,
		_w5292_
	);
	LUT3 #(
		.INIT('hc4)
	) name1245 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5154_,
		_w5293_
	);
	LUT3 #(
		.INIT('h02)
	) name1246 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5154_,
		_w5294_
	);
	LUT3 #(
		.INIT('h39)
	) name1247 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5154_,
		_w5295_
	);
	LUT4 #(
		.INIT('he8c0)
	) name1248 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		\core_dag_ilm1reg_M_reg[1]/NET0131 ,
		_w5175_,
		_w5182_,
		_w5296_
	);
	LUT4 #(
		.INIT('h0113)
	) name1249 (
		\core_dag_ilm1reg_M_reg[2]/NET0131 ,
		_w5161_,
		_w5168_,
		_w5296_,
		_w5297_
	);
	LUT4 #(
		.INIT('hfca8)
	) name1250 (
		\core_dag_ilm1reg_M_reg[4]/NET0131 ,
		\core_dag_ilm1reg_M_reg[5]/NET0131 ,
		_w5202_,
		_w5217_,
		_w5298_
	);
	LUT4 #(
		.INIT('h173f)
	) name1251 (
		\core_dag_ilm1reg_M_reg[4]/NET0131 ,
		\core_dag_ilm1reg_M_reg[5]/NET0131 ,
		_w5202_,
		_w5217_,
		_w5299_
	);
	LUT4 #(
		.INIT('hef00)
	) name1252 (
		_w5162_,
		_w5297_,
		_w5298_,
		_w5299_,
		_w5300_
	);
	LUT3 #(
		.INIT('h07)
	) name1253 (
		\core_dag_ilm1reg_M_reg[6]/NET0131 ,
		_w5196_,
		_w5209_,
		_w5301_
	);
	LUT4 #(
		.INIT('h0133)
	) name1254 (
		_w5197_,
		_w5208_,
		_w5300_,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		_w5236_,
		_w5243_,
		_w5303_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1256 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		\core_dag_ilm1reg_M_reg[11]/NET0131 ,
		_w5254_,
		_w5266_,
		_w5304_
	);
	LUT3 #(
		.INIT('he8)
	) name1257 (
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w5235_,
		_w5242_,
		_w5305_
	);
	LUT4 #(
		.INIT('he800)
	) name1258 (
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w5235_,
		_w5242_,
		_w5304_,
		_w5306_
	);
	LUT4 #(
		.INIT('h137f)
	) name1259 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		\core_dag_ilm1reg_M_reg[11]/NET0131 ,
		_w5254_,
		_w5266_,
		_w5307_
	);
	LUT2 #(
		.INIT('h4)
	) name1260 (
		_w5306_,
		_w5307_,
		_w5308_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1261 (
		_w5302_,
		_w5303_,
		_w5304_,
		_w5308_,
		_w5309_
	);
	LUT3 #(
		.INIT('h71)
	) name1262 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w5278_,
		_w5309_,
		_w5310_
	);
	LUT4 #(
		.INIT('h87e1)
	) name1263 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w5278_,
		_w5295_,
		_w5309_,
		_w5311_
	);
	LUT4 #(
		.INIT('h5410)
	) name1264 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5289_,
		_w5311_,
		_w5292_,
		_w5312_
	);
	LUT4 #(
		.INIT('h5041)
	) name1265 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		_w5287_,
		_w5290_,
		_w5291_,
		_w5313_
	);
	LUT2 #(
		.INIT('h8)
	) name1266 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		_w5154_,
		_w5314_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1267 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5311_,
		_w5313_,
		_w5314_,
		_w5315_
	);
	LUT4 #(
		.INIT('h0200)
	) name1268 (
		\core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w5316_
	);
	LUT4 #(
		.INIT('h0200)
	) name1269 (
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w5317_
	);
	LUT4 #(
		.INIT('h0200)
	) name1270 (
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w5318_
	);
	LUT4 #(
		.INIT('h0200)
	) name1271 (
		\core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w5319_
	);
	LUT3 #(
		.INIT('h01)
	) name1272 (
		_w5318_,
		_w5319_,
		_w5317_,
		_w5320_
	);
	LUT4 #(
		.INIT('h0200)
	) name1273 (
		\core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w5321_
	);
	LUT4 #(
		.INIT('h0200)
	) name1274 (
		\core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w5322_
	);
	LUT4 #(
		.INIT('h0200)
	) name1275 (
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w5323_
	);
	LUT4 #(
		.INIT('h0200)
	) name1276 (
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w5324_
	);
	LUT4 #(
		.INIT('h0001)
	) name1277 (
		_w5321_,
		_w5322_,
		_w5323_,
		_w5324_,
		_w5325_
	);
	LUT4 #(
		.INIT('h45ef)
	) name1278 (
		_w4063_,
		_w5316_,
		_w5320_,
		_w5325_,
		_w5326_
	);
	LUT2 #(
		.INIT('h4)
	) name1279 (
		\core_c_dec_Post2_E_reg/P0001 ,
		_w4973_,
		_w5327_
	);
	LUT3 #(
		.INIT('he0)
	) name1280 (
		_w5043_,
		_w5048_,
		_w5327_,
		_w5328_
	);
	LUT4 #(
		.INIT('h1b00)
	) name1281 (
		_w4063_,
		_w5025_,
		_w5041_,
		_w5328_,
		_w5329_
	);
	LUT2 #(
		.INIT('h2)
	) name1282 (
		_w4970_,
		_w5329_,
		_w5330_
	);
	LUT4 #(
		.INIT('h1300)
	) name1283 (
		_w4063_,
		_w5095_,
		_w5104_,
		_w5109_,
		_w5331_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1284 (
		_w5059_,
		_w4970_,
		_w5331_,
		_w5329_,
		_w5332_
	);
	LUT4 #(
		.INIT('hfb00)
	) name1285 (
		_w4104_,
		_w5058_,
		_w4970_,
		_w5327_,
		_w5333_
	);
	LUT4 #(
		.INIT('h00ec)
	) name1286 (
		_w4063_,
		_w5095_,
		_w5104_,
		_w5333_,
		_w5334_
	);
	LUT4 #(
		.INIT('h0020)
	) name1287 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w4104_,
		_w5058_,
		_w4970_,
		_w5335_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		_w5334_,
		_w5335_,
		_w5336_
	);
	LUT4 #(
		.INIT('h0072)
	) name1289 (
		_w4966_,
		_w5106_,
		_w5332_,
		_w5336_,
		_w5337_
	);
	LUT3 #(
		.INIT('hb0)
	) name1290 (
		_w5117_,
		_w5326_,
		_w5337_,
		_w5338_
	);
	LUT4 #(
		.INIT('h7500)
	) name1291 (
		_w5117_,
		_w5312_,
		_w5315_,
		_w5338_,
		_w5339_
	);
	LUT2 #(
		.INIT('h1)
	) name1292 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		_w5340_
	);
	LUT3 #(
		.INIT('h01)
	) name1293 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w5341_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5342_
	);
	LUT2 #(
		.INIT('h1)
	) name1295 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		_w5343_
	);
	LUT4 #(
		.INIT('h0001)
	) name1296 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5344_
	);
	LUT2 #(
		.INIT('h1)
	) name1297 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		_w5345_
	);
	LUT3 #(
		.INIT('h01)
	) name1298 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w5346_
	);
	LUT2 #(
		.INIT('h1)
	) name1299 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w5347_
	);
	LUT3 #(
		.INIT('h01)
	) name1300 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w5348_
	);
	LUT3 #(
		.INIT('h80)
	) name1301 (
		_w5344_,
		_w5346_,
		_w5348_,
		_w5349_
	);
	LUT4 #(
		.INIT('h4000)
	) name1302 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		_w5344_,
		_w5346_,
		_w5348_,
		_w5350_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		_w5341_,
		_w5350_,
		_w5351_
	);
	LUT3 #(
		.INIT('ha8)
	) name1304 (
		_w5344_,
		_w5346_,
		_w5347_,
		_w5352_
	);
	LUT3 #(
		.INIT('h01)
	) name1305 (
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5353_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1306 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5354_
	);
	LUT3 #(
		.INIT('h01)
	) name1307 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w5355_
	);
	LUT2 #(
		.INIT('h4)
	) name1308 (
		_w5354_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h4)
	) name1309 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w5344_,
		_w5357_
	);
	LUT3 #(
		.INIT('h0b)
	) name1310 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w5344_,
		_w5345_,
		_w5358_
	);
	LUT2 #(
		.INIT('h8)
	) name1311 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w5359_
	);
	LUT4 #(
		.INIT('h0777)
	) name1312 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		_w5360_
	);
	LUT3 #(
		.INIT('ha8)
	) name1313 (
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5361_
	);
	LUT3 #(
		.INIT('ha8)
	) name1314 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w5362_
	);
	LUT4 #(
		.INIT('h0100)
	) name1315 (
		_w5361_,
		_w5362_,
		_w5359_,
		_w5360_,
		_w5363_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1316 (
		_w5352_,
		_w5356_,
		_w5358_,
		_w5363_,
		_w5364_
	);
	LUT3 #(
		.INIT('h80)
	) name1317 (
		_w5344_,
		_w5346_,
		_w5347_,
		_w5365_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1318 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		_w5344_,
		_w5346_,
		_w5347_,
		_w5366_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1319 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		_w5344_,
		_w5346_,
		_w5348_,
		_w5367_
	);
	LUT2 #(
		.INIT('h1)
	) name1320 (
		_w5366_,
		_w5367_,
		_w5368_
	);
	LUT2 #(
		.INIT('h8)
	) name1321 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w5369_
	);
	LUT4 #(
		.INIT('h0040)
	) name1322 (
		_w5351_,
		_w5364_,
		_w5368_,
		_w5369_,
		_w5370_
	);
	LUT3 #(
		.INIT('h2a)
	) name1323 (
		\core_dag_ilm2reg_I_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		_w5370_,
		_w5371_
	);
	LUT4 #(
		.INIT('h20a0)
	) name1324 (
		\core_dag_ilm2reg_I_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_M_reg[0]/NET0131 ,
		_w5370_,
		_w5372_
	);
	LUT4 #(
		.INIT('hd25a)
	) name1325 (
		\core_dag_ilm2reg_I_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_M_reg[0]/NET0131 ,
		_w5370_,
		_w5373_
	);
	LUT4 #(
		.INIT('h0001)
	) name1326 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		_w5374_
	);
	LUT2 #(
		.INIT('h8)
	) name1327 (
		_w5348_,
		_w5374_,
		_w5375_
	);
	LUT3 #(
		.INIT('h80)
	) name1328 (
		_w5345_,
		_w5348_,
		_w5374_,
		_w5376_
	);
	LUT2 #(
		.INIT('h8)
	) name1329 (
		_w5357_,
		_w5376_,
		_w5377_
	);
	LUT4 #(
		.INIT('ha808)
	) name1330 (
		\core_dag_ilm2reg_I_reg[13]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5370_,
		_w5377_,
		_w5378_
	);
	LUT2 #(
		.INIT('h8)
	) name1331 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5378_,
		_w5379_
	);
	LUT4 #(
		.INIT('h4000)
	) name1332 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w5345_,
		_w5348_,
		_w5374_,
		_w5380_
	);
	LUT2 #(
		.INIT('h8)
	) name1333 (
		_w5343_,
		_w5380_,
		_w5381_
	);
	LUT4 #(
		.INIT('h5e0e)
	) name1334 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5370_,
		_w5381_,
		_w5382_
	);
	LUT3 #(
		.INIT('h80)
	) name1335 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M_reg[12]/NET0131 ,
		_w5382_,
		_w5383_
	);
	LUT3 #(
		.INIT('h13)
	) name1336 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M_reg[12]/NET0131 ,
		_w5382_,
		_w5384_
	);
	LUT2 #(
		.INIT('h4)
	) name1337 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		_w5380_,
		_w5385_
	);
	LUT4 #(
		.INIT('hf707)
	) name1338 (
		_w5342_,
		_w5343_,
		_w5370_,
		_w5385_,
		_w5386_
	);
	LUT2 #(
		.INIT('h8)
	) name1339 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		_w5386_,
		_w5387_
	);
	LUT3 #(
		.INIT('h13)
	) name1340 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w5386_,
		_w5388_
	);
	LUT4 #(
		.INIT('ha202)
	) name1341 (
		\core_dag_ilm2reg_I_reg[11]/NET0131 ,
		_w5353_,
		_w5370_,
		_w5381_,
		_w5389_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		\core_dag_ilm2reg_M_reg[11]/NET0131 ,
		_w5389_,
		_w5390_
	);
	LUT2 #(
		.INIT('h1)
	) name1343 (
		_w5388_,
		_w5390_,
		_w5391_
	);
	LUT2 #(
		.INIT('h2)
	) name1344 (
		_w5370_,
		_w5380_,
		_w5392_
	);
	LUT4 #(
		.INIT('h0040)
	) name1345 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w5342_,
		_w5343_,
		_w5370_,
		_w5393_
	);
	LUT3 #(
		.INIT('h02)
	) name1346 (
		\core_dag_ilm2reg_I_reg[9]/NET0131 ,
		_w5392_,
		_w5393_,
		_w5394_
	);
	LUT4 #(
		.INIT('h3331)
	) name1347 (
		\core_dag_ilm2reg_I_reg[9]/NET0131 ,
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w5392_,
		_w5393_,
		_w5395_
	);
	LUT2 #(
		.INIT('h2)
	) name1348 (
		_w5370_,
		_w5376_,
		_w5396_
	);
	LUT4 #(
		.INIT('h008a)
	) name1349 (
		\core_dag_ilm2reg_I_reg[8]/NET0131 ,
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		_w5393_,
		_w5396_,
		_w5397_
	);
	LUT2 #(
		.INIT('h1)
	) name1350 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		_w5397_,
		_w5398_
	);
	LUT4 #(
		.INIT('h0080)
	) name1351 (
		_w5342_,
		_w5343_,
		_w5346_,
		_w5370_,
		_w5399_
	);
	LUT2 #(
		.INIT('h2)
	) name1352 (
		_w5370_,
		_w5375_,
		_w5400_
	);
	LUT3 #(
		.INIT('h73)
	) name1353 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		_w5370_,
		_w5375_,
		_w5401_
	);
	LUT3 #(
		.INIT('h20)
	) name1354 (
		\core_dag_ilm2reg_I_reg[7]/NET0131 ,
		_w5399_,
		_w5401_,
		_w5402_
	);
	LUT4 #(
		.INIT('h3133)
	) name1355 (
		\core_dag_ilm2reg_I_reg[7]/NET0131 ,
		\core_dag_ilm2reg_M_reg[7]/NET0131 ,
		_w5399_,
		_w5401_,
		_w5403_
	);
	LUT4 #(
		.INIT('h0800)
	) name1356 (
		\core_dag_ilm2reg_I_reg[7]/NET0131 ,
		\core_dag_ilm2reg_M_reg[7]/NET0131 ,
		_w5399_,
		_w5401_,
		_w5404_
	);
	LUT4 #(
		.INIT('h008a)
	) name1357 (
		\core_dag_ilm2reg_I_reg[6]/NET0131 ,
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w5399_,
		_w5400_,
		_w5405_
	);
	LUT4 #(
		.INIT('haa2a)
	) name1358 (
		_w5350_,
		_w5364_,
		_w5368_,
		_w5369_,
		_w5406_
	);
	LUT4 #(
		.INIT('h00a2)
	) name1359 (
		\core_dag_ilm2reg_I_reg[3]/NET0131 ,
		_w5370_,
		_w5374_,
		_w5406_,
		_w5407_
	);
	LUT2 #(
		.INIT('h1)
	) name1360 (
		\core_dag_ilm2reg_M_reg[3]/NET0131 ,
		_w5407_,
		_w5408_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		\core_dag_ilm2reg_M_reg[3]/NET0131 ,
		_w5407_,
		_w5409_
	);
	LUT2 #(
		.INIT('h4)
	) name1362 (
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w5350_,
		_w5410_
	);
	LUT3 #(
		.INIT('h70)
	) name1363 (
		_w5364_,
		_w5368_,
		_w5410_,
		_w5411_
	);
	LUT4 #(
		.INIT('h008a)
	) name1364 (
		\core_dag_ilm2reg_I_reg[2]/NET0131 ,
		_w5341_,
		_w5370_,
		_w5411_,
		_w5412_
	);
	LUT4 #(
		.INIT('h1500)
	) name1365 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		_w5364_,
		_w5368_,
		_w5410_,
		_w5413_
	);
	LUT4 #(
		.INIT('h008a)
	) name1366 (
		\core_dag_ilm2reg_I_reg[1]/NET0131 ,
		_w5340_,
		_w5370_,
		_w5413_,
		_w5414_
	);
	LUT3 #(
		.INIT('he8)
	) name1367 (
		\core_dag_ilm2reg_M_reg[1]/NET0131 ,
		_w5372_,
		_w5414_,
		_w5415_
	);
	LUT4 #(
		.INIT('h0113)
	) name1368 (
		\core_dag_ilm2reg_M_reg[2]/NET0131 ,
		_w5409_,
		_w5412_,
		_w5415_,
		_w5416_
	);
	LUT2 #(
		.INIT('h4)
	) name1369 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		_w5374_,
		_w5417_
	);
	LUT4 #(
		.INIT('hacfc)
	) name1370 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		_w5365_,
		_w5370_,
		_w5417_,
		_w5418_
	);
	LUT2 #(
		.INIT('h2)
	) name1371 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		_w5418_,
		_w5419_
	);
	LUT3 #(
		.INIT('h31)
	) name1372 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M_reg[5]/NET0131 ,
		_w5418_,
		_w5420_
	);
	LUT4 #(
		.INIT('ha202)
	) name1373 (
		\core_dag_ilm2reg_I_reg[4]/NET0131 ,
		_w5349_,
		_w5370_,
		_w5417_,
		_w5421_
	);
	LUT2 #(
		.INIT('h1)
	) name1374 (
		\core_dag_ilm2reg_M_reg[4]/NET0131 ,
		_w5421_,
		_w5422_
	);
	LUT2 #(
		.INIT('h1)
	) name1375 (
		_w5420_,
		_w5422_,
		_w5423_
	);
	LUT2 #(
		.INIT('h8)
	) name1376 (
		\core_dag_ilm2reg_M_reg[4]/NET0131 ,
		_w5421_,
		_w5424_
	);
	LUT3 #(
		.INIT('h17)
	) name1377 (
		\core_dag_ilm2reg_M_reg[5]/NET0131 ,
		_w5419_,
		_w5424_,
		_w5425_
	);
	LUT4 #(
		.INIT('hef00)
	) name1378 (
		_w5408_,
		_w5416_,
		_w5423_,
		_w5425_,
		_w5426_
	);
	LUT4 #(
		.INIT('h1301)
	) name1379 (
		\core_dag_ilm2reg_M_reg[6]/NET0131 ,
		_w5404_,
		_w5405_,
		_w5426_,
		_w5427_
	);
	LUT4 #(
		.INIT('h0001)
	) name1380 (
		_w5395_,
		_w5398_,
		_w5403_,
		_w5427_,
		_w5428_
	);
	LUT2 #(
		.INIT('h8)
	) name1381 (
		\core_dag_ilm2reg_M_reg[11]/NET0131 ,
		_w5389_,
		_w5429_
	);
	LUT3 #(
		.INIT('h80)
	) name1382 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w5386_,
		_w5430_
	);
	LUT4 #(
		.INIT('he8c0)
	) name1383 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w5394_,
		_w5397_,
		_w5431_
	);
	LUT4 #(
		.INIT('h1113)
	) name1384 (
		_w5391_,
		_w5429_,
		_w5430_,
		_w5431_,
		_w5432_
	);
	LUT4 #(
		.INIT('h4055)
	) name1385 (
		_w5384_,
		_w5391_,
		_w5428_,
		_w5432_,
		_w5433_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1386 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5378_,
		_w5383_,
		_w5433_,
		_w5434_
	);
	LUT4 #(
		.INIT('h4442)
	) name1387 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5378_,
		_w5383_,
		_w5433_,
		_w5435_
	);
	LUT2 #(
		.INIT('h6)
	) name1388 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5436_
	);
	LUT2 #(
		.INIT('h9)
	) name1389 (
		_w5373_,
		_w5436_,
		_w5437_
	);
	LUT4 #(
		.INIT('h0100)
	) name1390 (
		_w5379_,
		_w5383_,
		_w5433_,
		_w5437_,
		_w5438_
	);
	LUT4 #(
		.INIT('haa08)
	) name1391 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5373_,
		_w5435_,
		_w5438_,
		_w5439_
	);
	LUT3 #(
		.INIT('h80)
	) name1392 (
		\core_dag_ilm2reg_I_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		_w5370_,
		_w5440_
	);
	LUT4 #(
		.INIT('h1333)
	) name1393 (
		\core_dag_ilm2reg_I_reg[13]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5370_,
		_w5377_,
		_w5441_
	);
	LUT2 #(
		.INIT('h2)
	) name1394 (
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5442_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		_w5441_,
		_w5442_,
		_w5443_
	);
	LUT4 #(
		.INIT('hc6cc)
	) name1396 (
		\core_dag_ilm2reg_I_reg[7]/NET0131 ,
		\core_dag_ilm2reg_M_reg[7]/NET0131 ,
		_w5399_,
		_w5401_,
		_w5444_
	);
	LUT2 #(
		.INIT('h6)
	) name1397 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5445_
	);
	LUT2 #(
		.INIT('h9)
	) name1398 (
		_w5444_,
		_w5445_,
		_w5446_
	);
	LUT2 #(
		.INIT('h6)
	) name1399 (
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5447_
	);
	LUT3 #(
		.INIT('h71)
	) name1400 (
		\core_dag_ilm2reg_M_reg[6]/NET0131 ,
		_w5405_,
		_w5447_,
		_w5448_
	);
	LUT2 #(
		.INIT('h4)
	) name1401 (
		_w5446_,
		_w5448_,
		_w5449_
	);
	LUT2 #(
		.INIT('h6)
	) name1402 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5450_
	);
	LUT4 #(
		.INIT('hf731)
	) name1403 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M_reg[5]/NET0131 ,
		_w5418_,
		_w5450_,
		_w5451_
	);
	LUT2 #(
		.INIT('h6)
	) name1404 (
		\core_dag_ilm2reg_M_reg[6]/NET0131 ,
		_w5405_,
		_w5452_
	);
	LUT4 #(
		.INIT('h9600)
	) name1405 (
		\core_dag_ilm2reg_M_reg[6]/NET0131 ,
		_w5405_,
		_w5447_,
		_w5451_,
		_w5453_
	);
	LUT2 #(
		.INIT('h6)
	) name1406 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5454_
	);
	LUT3 #(
		.INIT('h71)
	) name1407 (
		\core_dag_ilm2reg_M_reg[4]/NET0131 ,
		_w5421_,
		_w5454_,
		_w5455_
	);
	LUT3 #(
		.INIT('hc6)
	) name1408 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M_reg[5]/NET0131 ,
		_w5418_,
		_w5456_
	);
	LUT4 #(
		.INIT('hc639)
	) name1409 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M_reg[5]/NET0131 ,
		_w5418_,
		_w5450_,
		_w5457_
	);
	LUT2 #(
		.INIT('h6)
	) name1410 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5458_
	);
	LUT3 #(
		.INIT('h71)
	) name1411 (
		\core_dag_ilm2reg_M_reg[3]/NET0131 ,
		_w5407_,
		_w5458_,
		_w5459_
	);
	LUT2 #(
		.INIT('h6)
	) name1412 (
		\core_dag_ilm2reg_M_reg[4]/NET0131 ,
		_w5421_,
		_w5460_
	);
	LUT3 #(
		.INIT('h69)
	) name1413 (
		\core_dag_ilm2reg_M_reg[4]/NET0131 ,
		_w5421_,
		_w5454_,
		_w5461_
	);
	LUT2 #(
		.INIT('h4)
	) name1414 (
		_w5459_,
		_w5461_,
		_w5462_
	);
	LUT4 #(
		.INIT('hb2bb)
	) name1415 (
		_w5455_,
		_w5457_,
		_w5459_,
		_w5461_,
		_w5463_
	);
	LUT2 #(
		.INIT('h1)
	) name1416 (
		_w5453_,
		_w5463_,
		_w5464_
	);
	LUT4 #(
		.INIT('h0069)
	) name1417 (
		\core_dag_ilm2reg_M_reg[6]/NET0131 ,
		_w5405_,
		_w5447_,
		_w5451_,
		_w5465_
	);
	LUT3 #(
		.INIT('h0d)
	) name1418 (
		_w5446_,
		_w5448_,
		_w5465_,
		_w5466_
	);
	LUT3 #(
		.INIT('h45)
	) name1419 (
		_w5449_,
		_w5464_,
		_w5466_,
		_w5467_
	);
	LUT2 #(
		.INIT('h6)
	) name1420 (
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5468_
	);
	LUT3 #(
		.INIT('h71)
	) name1421 (
		\core_dag_ilm2reg_M_reg[2]/NET0131 ,
		_w5412_,
		_w5468_,
		_w5469_
	);
	LUT2 #(
		.INIT('h6)
	) name1422 (
		\core_dag_ilm2reg_M_reg[3]/NET0131 ,
		_w5407_,
		_w5470_
	);
	LUT3 #(
		.INIT('h69)
	) name1423 (
		\core_dag_ilm2reg_M_reg[3]/NET0131 ,
		_w5407_,
		_w5458_,
		_w5471_
	);
	LUT2 #(
		.INIT('h2)
	) name1424 (
		_w5469_,
		_w5471_,
		_w5472_
	);
	LUT2 #(
		.INIT('h4)
	) name1425 (
		_w5469_,
		_w5471_,
		_w5473_
	);
	LUT2 #(
		.INIT('h6)
	) name1426 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5474_
	);
	LUT3 #(
		.INIT('h71)
	) name1427 (
		\core_dag_ilm2reg_M_reg[1]/NET0131 ,
		_w5414_,
		_w5474_,
		_w5475_
	);
	LUT2 #(
		.INIT('h6)
	) name1428 (
		\core_dag_ilm2reg_M_reg[2]/NET0131 ,
		_w5412_,
		_w5476_
	);
	LUT3 #(
		.INIT('h69)
	) name1429 (
		\core_dag_ilm2reg_M_reg[2]/NET0131 ,
		_w5412_,
		_w5468_,
		_w5477_
	);
	LUT2 #(
		.INIT('h2)
	) name1430 (
		_w5475_,
		_w5477_,
		_w5478_
	);
	LUT2 #(
		.INIT('h4)
	) name1431 (
		_w5475_,
		_w5477_,
		_w5479_
	);
	LUT3 #(
		.INIT('h8e)
	) name1432 (
		\core_dag_ilm2reg_M_reg[0]/NET0131 ,
		_w5371_,
		_w5436_,
		_w5480_
	);
	LUT3 #(
		.INIT('h69)
	) name1433 (
		\core_dag_ilm2reg_M_reg[1]/NET0131 ,
		_w5414_,
		_w5474_,
		_w5481_
	);
	LUT3 #(
		.INIT('h21)
	) name1434 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5373_,
		_w5482_
	);
	LUT3 #(
		.INIT('he8)
	) name1435 (
		_w5480_,
		_w5481_,
		_w5482_,
		_w5483_
	);
	LUT4 #(
		.INIT('h0445)
	) name1436 (
		_w5473_,
		_w5475_,
		_w5477_,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h2)
	) name1437 (
		_w5459_,
		_w5461_,
		_w5485_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1438 (
		_w5455_,
		_w5457_,
		_w5459_,
		_w5461_,
		_w5486_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1439 (
		_w5446_,
		_w5448_,
		_w5453_,
		_w5486_,
		_w5487_
	);
	LUT3 #(
		.INIT('h10)
	) name1440 (
		_w5472_,
		_w5484_,
		_w5487_,
		_w5488_
	);
	LUT4 #(
		.INIT('hccc6)
	) name1441 (
		\core_dag_ilm2reg_I_reg[9]/NET0131 ,
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w5392_,
		_w5393_,
		_w5489_
	);
	LUT2 #(
		.INIT('h6)
	) name1442 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5490_
	);
	LUT2 #(
		.INIT('h9)
	) name1443 (
		_w5489_,
		_w5490_,
		_w5491_
	);
	LUT2 #(
		.INIT('h6)
	) name1444 (
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5492_
	);
	LUT3 #(
		.INIT('h71)
	) name1445 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		_w5397_,
		_w5492_,
		_w5493_
	);
	LUT3 #(
		.INIT('h71)
	) name1446 (
		\core_dag_ilm2reg_M_reg[7]/NET0131 ,
		_w5402_,
		_w5445_,
		_w5494_
	);
	LUT2 #(
		.INIT('h6)
	) name1447 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		_w5397_,
		_w5495_
	);
	LUT3 #(
		.INIT('h69)
	) name1448 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		_w5397_,
		_w5492_,
		_w5496_
	);
	LUT2 #(
		.INIT('h2)
	) name1449 (
		_w5494_,
		_w5496_,
		_w5497_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name1450 (
		_w5491_,
		_w5493_,
		_w5494_,
		_w5496_,
		_w5498_
	);
	LUT3 #(
		.INIT('h6c)
	) name1451 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w5386_,
		_w5499_
	);
	LUT2 #(
		.INIT('h6)
	) name1452 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5500_
	);
	LUT4 #(
		.INIT('h6c93)
	) name1453 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w5386_,
		_w5500_,
		_w5501_
	);
	LUT4 #(
		.INIT('h0071)
	) name1454 (
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w5394_,
		_w5490_,
		_w5501_,
		_w5502_
	);
	LUT4 #(
		.INIT('h7f13)
	) name1455 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w5386_,
		_w5500_,
		_w5503_
	);
	LUT2 #(
		.INIT('h6)
	) name1456 (
		\core_dag_ilm2reg_M_reg[11]/NET0131 ,
		_w5389_,
		_w5504_
	);
	LUT2 #(
		.INIT('h6)
	) name1457 (
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5505_
	);
	LUT3 #(
		.INIT('h69)
	) name1458 (
		\core_dag_ilm2reg_M_reg[11]/NET0131 ,
		_w5389_,
		_w5505_,
		_w5506_
	);
	LUT2 #(
		.INIT('h2)
	) name1459 (
		_w5503_,
		_w5506_,
		_w5507_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w5502_,
		_w5507_,
		_w5508_
	);
	LUT4 #(
		.INIT('he000)
	) name1461 (
		_w5467_,
		_w5488_,
		_w5498_,
		_w5508_,
		_w5509_
	);
	LUT2 #(
		.INIT('h4)
	) name1462 (
		_w5494_,
		_w5496_,
		_w5510_
	);
	LUT4 #(
		.INIT('hd4dd)
	) name1463 (
		_w5491_,
		_w5493_,
		_w5494_,
		_w5496_,
		_w5511_
	);
	LUT4 #(
		.INIT('h8e00)
	) name1464 (
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w5394_,
		_w5490_,
		_w5501_,
		_w5512_
	);
	LUT3 #(
		.INIT('h2b)
	) name1465 (
		_w5503_,
		_w5506_,
		_w5512_,
		_w5513_
	);
	LUT3 #(
		.INIT('hd0)
	) name1466 (
		_w5508_,
		_w5511_,
		_w5513_,
		_w5514_
	);
	LUT4 #(
		.INIT('h64c4)
	) name1467 (
		\core_dag_ilm2reg_I_reg[13]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5370_,
		_w5377_,
		_w5515_
	);
	LUT2 #(
		.INIT('h6)
	) name1468 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5516_
	);
	LUT4 #(
		.INIT('h80ec)
	) name1469 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M_reg[12]/NET0131 ,
		_w5382_,
		_w5516_,
		_w5517_
	);
	LUT3 #(
		.INIT('h71)
	) name1470 (
		\core_dag_ilm2reg_M_reg[11]/NET0131 ,
		_w5389_,
		_w5505_,
		_w5518_
	);
	LUT3 #(
		.INIT('h6c)
	) name1471 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M_reg[12]/NET0131 ,
		_w5382_,
		_w5519_
	);
	LUT4 #(
		.INIT('h6c93)
	) name1472 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M_reg[12]/NET0131 ,
		_w5382_,
		_w5516_,
		_w5520_
	);
	LUT2 #(
		.INIT('h2)
	) name1473 (
		_w5518_,
		_w5520_,
		_w5521_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1474 (
		_w5515_,
		_w5517_,
		_w5518_,
		_w5520_,
		_w5522_
	);
	LUT2 #(
		.INIT('h4)
	) name1475 (
		_w5518_,
		_w5520_,
		_w5523_
	);
	LUT4 #(
		.INIT('hb2bb)
	) name1476 (
		_w5515_,
		_w5517_,
		_w5518_,
		_w5520_,
		_w5524_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1477 (
		_w5509_,
		_w5514_,
		_w5522_,
		_w5524_,
		_w5525_
	);
	LUT2 #(
		.INIT('h9)
	) name1478 (
		_w5443_,
		_w5525_,
		_w5526_
	);
	LUT3 #(
		.INIT('h14)
	) name1479 (
		_w5373_,
		_w5443_,
		_w5525_,
		_w5527_
	);
	LUT4 #(
		.INIT('h1551)
	) name1480 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5437_,
		_w5443_,
		_w5525_,
		_w5528_
	);
	LUT3 #(
		.INIT('h45)
	) name1481 (
		_w5440_,
		_w5527_,
		_w5528_,
		_w5529_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name1482 (
		_w4067_,
		_w4068_,
		_w4519_,
		_w4845_,
		_w5530_
	);
	LUT4 #(
		.INIT('he000)
	) name1483 (
		\bdma_BCTL_reg[0]/NET0131 ,
		\bdma_BCTL_reg[1]/NET0131 ,
		\bdma_BDMAmode_reg/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w5531_
	);
	LUT2 #(
		.INIT('h1)
	) name1484 (
		\bdma_BCTL_reg[1]/NET0131 ,
		\bdma_DM_2nd_reg/NET0131 ,
		_w5532_
	);
	LUT3 #(
		.INIT('h32)
	) name1485 (
		\bdma_BCTL_reg[1]/NET0131 ,
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_DM_2nd_reg/NET0131 ,
		_w5533_
	);
	LUT2 #(
		.INIT('h8)
	) name1486 (
		_w5531_,
		_w5533_,
		_w5534_
	);
	LUT3 #(
		.INIT('h8c)
	) name1487 (
		\bdma_BCTL_reg[1]/NET0131 ,
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_DM_2nd_reg/NET0131 ,
		_w5535_
	);
	LUT2 #(
		.INIT('h8)
	) name1488 (
		_w5531_,
		_w5535_,
		_w5536_
	);
	LUT2 #(
		.INIT('h8)
	) name1489 (
		_w4519_,
		_w5536_,
		_w5537_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1490 (
		_w4067_,
		_w4068_,
		_w4845_,
		_w5537_,
		_w5538_
	);
	LUT3 #(
		.INIT('h07)
	) name1491 (
		_w5530_,
		_w5534_,
		_w5538_,
		_w5539_
	);
	LUT4 #(
		.INIT('h0200)
	) name1492 (
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w5540_
	);
	LUT4 #(
		.INIT('h0200)
	) name1493 (
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w5541_
	);
	LUT4 #(
		.INIT('h0200)
	) name1494 (
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w5542_
	);
	LUT4 #(
		.INIT('h0200)
	) name1495 (
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w5543_
	);
	LUT4 #(
		.INIT('h0001)
	) name1496 (
		_w5540_,
		_w5541_,
		_w5542_,
		_w5543_,
		_w5544_
	);
	LUT4 #(
		.INIT('h0200)
	) name1497 (
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w5545_
	);
	LUT4 #(
		.INIT('h0200)
	) name1498 (
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w5546_
	);
	LUT4 #(
		.INIT('h0200)
	) name1499 (
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w5547_
	);
	LUT4 #(
		.INIT('h0200)
	) name1500 (
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w5548_
	);
	LUT4 #(
		.INIT('h0001)
	) name1501 (
		_w5545_,
		_w5546_,
		_w5547_,
		_w5548_,
		_w5549_
	);
	LUT3 #(
		.INIT('h1b)
	) name1502 (
		_w4063_,
		_w5544_,
		_w5549_,
		_w5550_
	);
	LUT4 #(
		.INIT('h0123)
	) name1503 (
		_w4063_,
		_w5049_,
		_w5544_,
		_w5549_,
		_w5551_
	);
	LUT3 #(
		.INIT('h02)
	) name1504 (
		\core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5552_
	);
	LUT4 #(
		.INIT('h0200)
	) name1505 (
		\core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w5553_
	);
	LUT4 #(
		.INIT('h0200)
	) name1506 (
		\core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w5554_
	);
	LUT4 #(
		.INIT('h0200)
	) name1507 (
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w5555_
	);
	LUT4 #(
		.INIT('h0200)
	) name1508 (
		\core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w5556_
	);
	LUT3 #(
		.INIT('h01)
	) name1509 (
		_w5555_,
		_w5556_,
		_w5554_,
		_w5557_
	);
	LUT4 #(
		.INIT('h0200)
	) name1510 (
		\core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w5558_
	);
	LUT4 #(
		.INIT('h0200)
	) name1511 (
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w5559_
	);
	LUT4 #(
		.INIT('h0200)
	) name1512 (
		\core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w5560_
	);
	LUT4 #(
		.INIT('h0200)
	) name1513 (
		\core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w5561_
	);
	LUT4 #(
		.INIT('h0001)
	) name1514 (
		_w5558_,
		_w5559_,
		_w5560_,
		_w5561_,
		_w5562_
	);
	LUT4 #(
		.INIT('h45ef)
	) name1515 (
		_w4063_,
		_w5553_,
		_w5557_,
		_w5562_,
		_w5563_
	);
	LUT3 #(
		.INIT('h08)
	) name1516 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w5564_
	);
	LUT4 #(
		.INIT('h0800)
	) name1517 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w5565_
	);
	LUT4 #(
		.INIT('h000b)
	) name1518 (
		_w4970_,
		_w5563_,
		_w5565_,
		_w5551_,
		_w5566_
	);
	LUT3 #(
		.INIT('h23)
	) name1519 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\core_c_psq_PCS_reg[5]/NET0131 ,
		\core_c_psq_PCS_reg[6]/NET0131 ,
		_w5567_
	);
	LUT3 #(
		.INIT('hdc)
	) name1520 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\core_c_psq_PCS_reg[5]/NET0131 ,
		\core_c_psq_PCS_reg[6]/NET0131 ,
		_w5568_
	);
	LUT2 #(
		.INIT('h8)
	) name1521 (
		_w4870_,
		_w5567_,
		_w5569_
	);
	LUT4 #(
		.INIT('h4555)
	) name1522 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w5570_
	);
	LUT4 #(
		.INIT('hea00)
	) name1523 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w5056_,
		_w5571_
	);
	LUT4 #(
		.INIT('ha222)
	) name1524 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w5572_
	);
	LUT4 #(
		.INIT('h0800)
	) name1525 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w5573_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1526 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w5574_
	);
	LUT3 #(
		.INIT('h40)
	) name1527 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w5575_
	);
	LUT4 #(
		.INIT('h4000)
	) name1528 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[0]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w5576_
	);
	LUT2 #(
		.INIT('h1)
	) name1529 (
		_w5574_,
		_w5576_,
		_w5577_
	);
	LUT2 #(
		.INIT('h4)
	) name1530 (
		_w5572_,
		_w5577_,
		_w5578_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1531 (
		_w5059_,
		_w5539_,
		_w5566_,
		_w5578_,
		_w5579_
	);
	LUT4 #(
		.INIT('haa80)
	) name1532 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w5580_
	);
	LUT4 #(
		.INIT('h2223)
	) name1533 (
		_w5117_,
		_w5337_,
		_w5579_,
		_w5580_,
		_w5581_
	);
	LUT4 #(
		.INIT('h7500)
	) name1534 (
		_w5117_,
		_w5439_,
		_w5529_,
		_w5581_,
		_w5582_
	);
	LUT4 #(
		.INIT('h0a08)
	) name1535 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w4967_,
		_w5107_,
		_w4969_,
		_w5583_
	);
	LUT4 #(
		.INIT('h00a8)
	) name1536 (
		_w5059_,
		_w5042_,
		_w5105_,
		_w5583_,
		_w5584_
	);
	LUT2 #(
		.INIT('h8)
	) name1537 (
		_w5042_,
		_w5334_,
		_w5585_
	);
	LUT4 #(
		.INIT('h00ba)
	) name1538 (
		_w4966_,
		_w5330_,
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		\memc_DMo_oe1_reg/P0001 ,
		\memc_DMo_oe2_reg/P0001 ,
		_w5587_
	);
	LUT2 #(
		.INIT('h1)
	) name1540 (
		\memc_DMo_oe4_reg/P0001 ,
		\memc_DMo_oe5_reg/P0001 ,
		_w5588_
	);
	LUT4 #(
		.INIT('h0001)
	) name1541 (
		\memc_DMo_oe3_reg/P0001 ,
		\memc_DMo_oe4_reg/P0001 ,
		\memc_DMo_oe5_reg/P0001 ,
		\memc_DMo_oe6_reg/P0001 ,
		_w5589_
	);
	LUT2 #(
		.INIT('h4)
	) name1542 (
		\memc_DM_oe_reg/P0001 ,
		\memc_DMo_oe7_reg/P0001 ,
		_w5590_
	);
	LUT4 #(
		.INIT('h4000)
	) name1543 (
		\memc_DMo_oe0_reg/P0001 ,
		_w5587_,
		_w5589_,
		_w5590_,
		_w5591_
	);
	LUT2 #(
		.INIT('h2)
	) name1544 (
		\memc_DM_oe_reg/P0001 ,
		\memc_DMo_oe7_reg/P0001 ,
		_w5592_
	);
	LUT4 #(
		.INIT('h4000)
	) name1545 (
		\memc_DMo_oe0_reg/P0001 ,
		_w5587_,
		_w5589_,
		_w5592_,
		_w5593_
	);
	LUT3 #(
		.INIT('h01)
	) name1546 (
		\memc_DM_oe_reg/P0001 ,
		\memc_DMo_oe0_reg/P0001 ,
		\memc_DMo_oe7_reg/P0001 ,
		_w5594_
	);
	LUT3 #(
		.INIT('h10)
	) name1547 (
		\memc_DMo_oe4_reg/P0001 ,
		\memc_DMo_oe5_reg/P0001 ,
		\memc_DMo_oe6_reg/P0001 ,
		_w5595_
	);
	LUT4 #(
		.INIT('h4000)
	) name1548 (
		\memc_DMo_oe3_reg/P0001 ,
		_w5587_,
		_w5594_,
		_w5595_,
		_w5596_
	);
	LUT3 #(
		.INIT('h01)
	) name1549 (
		_w5593_,
		_w5596_,
		_w5591_,
		_w5597_
	);
	LUT4 #(
		.INIT('h1000)
	) name1550 (
		\memc_DMo_oe3_reg/P0001 ,
		\memc_DMo_oe6_reg/P0001 ,
		_w5587_,
		_w5594_,
		_w5598_
	);
	LUT2 #(
		.INIT('h4)
	) name1551 (
		\memc_DMo_oe4_reg/P0001 ,
		\memc_DMo_oe5_reg/P0001 ,
		_w5599_
	);
	LUT2 #(
		.INIT('h8)
	) name1552 (
		_w5598_,
		_w5599_,
		_w5600_
	);
	LUT2 #(
		.INIT('h2)
	) name1553 (
		\memc_DMo_oe4_reg/P0001 ,
		\memc_DMo_oe5_reg/P0001 ,
		_w5601_
	);
	LUT2 #(
		.INIT('h8)
	) name1554 (
		_w5598_,
		_w5601_,
		_w5602_
	);
	LUT2 #(
		.INIT('h4)
	) name1555 (
		\memc_DMo_oe1_reg/P0001 ,
		\memc_DMo_oe2_reg/P0001 ,
		_w5603_
	);
	LUT3 #(
		.INIT('h80)
	) name1556 (
		_w5589_,
		_w5594_,
		_w5603_,
		_w5604_
	);
	LUT2 #(
		.INIT('h2)
	) name1557 (
		\memc_DMo_oe1_reg/P0001 ,
		\memc_DMo_oe2_reg/P0001 ,
		_w5605_
	);
	LUT3 #(
		.INIT('h80)
	) name1558 (
		_w5589_,
		_w5594_,
		_w5605_,
		_w5606_
	);
	LUT4 #(
		.INIT('h0002)
	) name1559 (
		\memc_DMo_oe3_reg/P0001 ,
		\memc_DMo_oe4_reg/P0001 ,
		\memc_DMo_oe5_reg/P0001 ,
		\memc_DMo_oe6_reg/P0001 ,
		_w5607_
	);
	LUT3 #(
		.INIT('h80)
	) name1560 (
		_w5587_,
		_w5594_,
		_w5607_,
		_w5608_
	);
	LUT3 #(
		.INIT('h01)
	) name1561 (
		_w5606_,
		_w5608_,
		_w5604_,
		_w5609_
	);
	LUT4 #(
		.INIT('h1000)
	) name1562 (
		_w5602_,
		_w5600_,
		_w5609_,
		_w5597_,
		_w5610_
	);
	LUT3 #(
		.INIT('h04)
	) name1563 (
		\memc_DM_oe_reg/P0001 ,
		\memc_DMo_oe0_reg/P0001 ,
		\memc_DMo_oe7_reg/P0001 ,
		_w5611_
	);
	LUT3 #(
		.INIT('h80)
	) name1564 (
		_w5587_,
		_w5589_,
		_w5611_,
		_w5612_
	);
	LUT3 #(
		.INIT('ha8)
	) name1565 (
		\DM_rd0[13]_pad ,
		_w5610_,
		_w5612_,
		_w5613_
	);
	LUT4 #(
		.INIT('h153f)
	) name1566 (
		\DM_rd6[13]_pad ,
		\DM_rdm[13]_pad ,
		_w5593_,
		_w5596_,
		_w5614_
	);
	LUT4 #(
		.INIT('h153f)
	) name1567 (
		\DM_rd7[13]_pad ,
		_w5588_,
		_w5598_,
		_w5591_,
		_w5615_
	);
	LUT2 #(
		.INIT('h8)
	) name1568 (
		_w5614_,
		_w5615_,
		_w5616_
	);
	LUT3 #(
		.INIT('h80)
	) name1569 (
		\DM_rd5[13]_pad ,
		_w5598_,
		_w5599_,
		_w5617_
	);
	LUT3 #(
		.INIT('h80)
	) name1570 (
		\DM_rd4[13]_pad ,
		_w5598_,
		_w5601_,
		_w5618_
	);
	LUT4 #(
		.INIT('h8000)
	) name1571 (
		\DM_rd2[13]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w5619_
	);
	LUT4 #(
		.INIT('h8000)
	) name1572 (
		\DM_rd1[13]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w5620_
	);
	LUT4 #(
		.INIT('h8000)
	) name1573 (
		\DM_rd3[13]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w5621_
	);
	LUT3 #(
		.INIT('h01)
	) name1574 (
		_w5620_,
		_w5621_,
		_w5619_,
		_w5622_
	);
	LUT3 #(
		.INIT('h10)
	) name1575 (
		_w5618_,
		_w5617_,
		_w5622_,
		_w5623_
	);
	LUT2 #(
		.INIT('h8)
	) name1576 (
		_w5616_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h4)
	) name1577 (
		_w5613_,
		_w5624_,
		_w5625_
	);
	LUT4 #(
		.INIT('h4000)
	) name1578 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[13]/P0001 ,
		_w5626_
	);
	LUT4 #(
		.INIT('h0800)
	) name1579 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5627_
	);
	LUT2 #(
		.INIT('h1)
	) name1580 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w5628_
	);
	LUT4 #(
		.INIT('h8000)
	) name1581 (
		_w5053_,
		_w5052_,
		_w5054_,
		_w5628_,
		_w5629_
	);
	LUT3 #(
		.INIT('h80)
	) name1582 (
		\bdma_BCTL_reg[13]/NET0131 ,
		_w5627_,
		_w5629_,
		_w5630_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w5631_
	);
	LUT4 #(
		.INIT('h4000)
	) name1584 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5632_
	);
	LUT3 #(
		.INIT('h80)
	) name1585 (
		\emc_WSCRreg_DO_reg[13]/NET0131 ,
		_w5631_,
		_w5632_,
		_w5633_
	);
	LUT2 #(
		.INIT('h4)
	) name1586 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w5634_
	);
	LUT4 #(
		.INIT('h2000)
	) name1587 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5635_
	);
	LUT3 #(
		.INIT('h80)
	) name1588 (
		\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w5634_,
		_w5635_,
		_w5636_
	);
	LUT4 #(
		.INIT('h1000)
	) name1589 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5637_
	);
	LUT3 #(
		.INIT('h80)
	) name1590 (
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w5634_,
		_w5637_,
		_w5638_
	);
	LUT4 #(
		.INIT('h0100)
	) name1591 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5639_
	);
	LUT3 #(
		.INIT('he2)
	) name1592 (
		\sport1_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_rxctl_SLOT1_EXT_reg[3]/NET0131 ,
		_w5640_
	);
	LUT3 #(
		.INIT('h80)
	) name1593 (
		_w5631_,
		_w5639_,
		_w5640_,
		_w5641_
	);
	LUT4 #(
		.INIT('h0001)
	) name1594 (
		_w5633_,
		_w5636_,
		_w5638_,
		_w5641_,
		_w5642_
	);
	LUT2 #(
		.INIT('h4)
	) name1595 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w5643_
	);
	LUT4 #(
		.INIT('h0400)
	) name1596 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5644_
	);
	LUT3 #(
		.INIT('h80)
	) name1597 (
		\clkc_ckr_reg_DO_reg[13]/NET0131 ,
		_w5631_,
		_w5644_,
		_w5645_
	);
	LUT3 #(
		.INIT('h80)
	) name1598 (
		\PIO_oe[9]_pad ,
		_w5628_,
		_w5632_,
		_w5646_
	);
	LUT2 #(
		.INIT('h2)
	) name1599 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w5647_
	);
	LUT4 #(
		.INIT('h0200)
	) name1600 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5648_
	);
	LUT3 #(
		.INIT('h80)
	) name1601 (
		\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w5648_,
		_w5634_,
		_w5649_
	);
	LUT3 #(
		.INIT('h80)
	) name1602 (
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w5632_,
		_w5634_,
		_w5650_
	);
	LUT4 #(
		.INIT('h0001)
	) name1603 (
		_w5645_,
		_w5646_,
		_w5649_,
		_w5650_,
		_w5651_
	);
	LUT3 #(
		.INIT('h40)
	) name1604 (
		_w5630_,
		_w5642_,
		_w5651_,
		_w5652_
	);
	LUT3 #(
		.INIT('h80)
	) name1605 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w5629_,
		_w5648_,
		_w5653_
	);
	LUT3 #(
		.INIT('h80)
	) name1606 (
		\bdma_BEAD_reg[13]/NET0131 ,
		_w5629_,
		_w5644_,
		_w5654_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w5653_,
		_w5654_,
		_w5655_
	);
	LUT2 #(
		.INIT('h2)
	) name1608 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5656_
	);
	LUT4 #(
		.INIT('h0010)
	) name1609 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5657_
	);
	LUT4 #(
		.INIT('h4000)
	) name1610 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w5053_,
		_w5052_,
		_w5054_,
		_w5658_
	);
	LUT4 #(
		.INIT('h8000)
	) name1611 (
		\bdma_BWCOUNT_reg[13]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w5659_
	);
	LUT4 #(
		.INIT('h8000)
	) name1612 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5660_
	);
	LUT3 #(
		.INIT('h80)
	) name1613 (
		\memc_usysr_DO_reg[13]/NET0131 ,
		_w5631_,
		_w5660_,
		_w5661_
	);
	LUT3 #(
		.INIT('h80)
	) name1614 (
		\pio_pmask_reg_DO_reg[9]/NET0131 ,
		_w5628_,
		_w5660_,
		_w5662_
	);
	LUT3 #(
		.INIT('h80)
	) name1615 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w5628_,
		_w5639_,
		_w5663_
	);
	LUT3 #(
		.INIT('h01)
	) name1616 (
		_w5662_,
		_w5663_,
		_w5661_,
		_w5664_
	);
	LUT3 #(
		.INIT('h80)
	) name1617 (
		\tm_TCR_TMP_reg[13]/NET0131 ,
		_w5631_,
		_w5637_,
		_w5665_
	);
	LUT3 #(
		.INIT('h80)
	) name1618 (
		\PIO_out[9]_pad ,
		_w5628_,
		_w5635_,
		_w5666_
	);
	LUT3 #(
		.INIT('h80)
	) name1619 (
		\tm_tpr_reg_DO_reg[13]/NET0131 ,
		_w5631_,
		_w5635_,
		_w5667_
	);
	LUT3 #(
		.INIT('h80)
	) name1620 (
		\sport0_regs_AUTO_a_reg[13]/NET0131 ,
		_w5627_,
		_w5634_,
		_w5668_
	);
	LUT4 #(
		.INIT('h0001)
	) name1621 (
		_w5665_,
		_w5666_,
		_w5667_,
		_w5668_,
		_w5669_
	);
	LUT2 #(
		.INIT('h4)
	) name1622 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5670_
	);
	LUT2 #(
		.INIT('h4)
	) name1623 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5671_
	);
	LUT4 #(
		.INIT('h0100)
	) name1624 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5672_
	);
	LUT3 #(
		.INIT('h80)
	) name1625 (
		\pio_PINT_reg[9]/NET0131 ,
		_w5670_,
		_w5672_,
		_w5673_
	);
	LUT3 #(
		.INIT('h80)
	) name1626 (
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w5634_,
		_w5639_,
		_w5674_
	);
	LUT3 #(
		.INIT('he2)
	) name1627 (
		\sport0_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_rxctl_SLOT1_EXT_reg[3]/NET0131 ,
		_w5675_
	);
	LUT3 #(
		.INIT('h80)
	) name1628 (
		_w5634_,
		_w5660_,
		_w5675_,
		_w5676_
	);
	LUT3 #(
		.INIT('h80)
	) name1629 (
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w5644_,
		_w5634_,
		_w5677_
	);
	LUT4 #(
		.INIT('h0001)
	) name1630 (
		_w5673_,
		_w5674_,
		_w5676_,
		_w5677_,
		_w5678_
	);
	LUT4 #(
		.INIT('h4000)
	) name1631 (
		_w5659_,
		_w5664_,
		_w5669_,
		_w5678_,
		_w5679_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1632 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w5652_,
		_w5655_,
		_w5679_,
		_w5680_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1633 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_MFPSQ_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w5681_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1634 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4237_,
		_w4234_,
		_w4242_,
		_w5682_
	);
	LUT3 #(
		.INIT('ha8)
	) name1635 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w5683_
	);
	LUT4 #(
		.INIT('h135f)
	) name1636 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w5684_
	);
	LUT2 #(
		.INIT('h4)
	) name1637 (
		_w5683_,
		_w5684_,
		_w5685_
	);
	LUT3 #(
		.INIT('h8a)
	) name1638 (
		_w5681_,
		_w5682_,
		_w5685_,
		_w5686_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1639 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_MFDAG2_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w5687_
	);
	LUT4 #(
		.INIT('h135f)
	) name1640 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131 ,
		_w5688_
	);
	LUT4 #(
		.INIT('h135f)
	) name1641 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131 ,
		_w5689_
	);
	LUT2 #(
		.INIT('h8)
	) name1642 (
		_w5688_,
		_w5689_,
		_w5690_
	);
	LUT4 #(
		.INIT('h135f)
	) name1643 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131 ,
		_w5691_
	);
	LUT4 #(
		.INIT('h135f)
	) name1644 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131 ,
		_w5692_
	);
	LUT4 #(
		.INIT('h135f)
	) name1645 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131 ,
		_w5693_
	);
	LUT4 #(
		.INIT('h135f)
	) name1646 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131 ,
		_w5694_
	);
	LUT4 #(
		.INIT('h8000)
	) name1647 (
		_w5693_,
		_w5694_,
		_w5691_,
		_w5692_,
		_w5695_
	);
	LUT3 #(
		.INIT('h2a)
	) name1648 (
		_w5687_,
		_w5690_,
		_w5695_,
		_w5696_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1649 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_MFDAG1_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w5697_
	);
	LUT4 #(
		.INIT('h135f)
	) name1650 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131 ,
		_w5698_
	);
	LUT4 #(
		.INIT('h135f)
	) name1651 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131 ,
		_w5699_
	);
	LUT2 #(
		.INIT('h8)
	) name1652 (
		_w5698_,
		_w5699_,
		_w5700_
	);
	LUT4 #(
		.INIT('h135f)
	) name1653 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131 ,
		_w5701_
	);
	LUT4 #(
		.INIT('h135f)
	) name1654 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131 ,
		_w5702_
	);
	LUT4 #(
		.INIT('h135f)
	) name1655 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131 ,
		_w5703_
	);
	LUT4 #(
		.INIT('h135f)
	) name1656 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131 ,
		_w5704_
	);
	LUT4 #(
		.INIT('h8000)
	) name1657 (
		_w5703_,
		_w5704_,
		_w5701_,
		_w5702_,
		_w5705_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1658 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_MFSPT_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w5706_
	);
	LUT4 #(
		.INIT('h135f)
	) name1659 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[13]/P0001 ,
		\sport1_txctl_TX_reg[13]/P0001 ,
		_w5707_
	);
	LUT4 #(
		.INIT('h135f)
	) name1660 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[13]/P0001 ,
		\sport1_rxctl_RX_reg[13]/P0001 ,
		_w5708_
	);
	LUT3 #(
		.INIT('h2a)
	) name1661 (
		_w5706_,
		_w5707_,
		_w5708_,
		_w5709_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1662 (
		_w5697_,
		_w5700_,
		_w5705_,
		_w5709_,
		_w5710_
	);
	LUT2 #(
		.INIT('h4)
	) name1663 (
		_w5696_,
		_w5710_,
		_w5711_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1664 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_MFMAC_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w5712_
	);
	LUT3 #(
		.INIT('h1b)
	) name1665 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 ,
		_w5713_
	);
	LUT4 #(
		.INIT('ha820)
	) name1666 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 ,
		_w5714_
	);
	LUT3 #(
		.INIT('h1b)
	) name1667 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001 ,
		_w5715_
	);
	LUT4 #(
		.INIT('ha820)
	) name1668 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001 ,
		_w5716_
	);
	LUT3 #(
		.INIT('h1b)
	) name1669 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 ,
		_w5717_
	);
	LUT4 #(
		.INIT('ha820)
	) name1670 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 ,
		_w5718_
	);
	LUT3 #(
		.INIT('h01)
	) name1671 (
		_w5716_,
		_w5718_,
		_w5714_,
		_w5719_
	);
	LUT3 #(
		.INIT('h1b)
	) name1672 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001 ,
		_w5720_
	);
	LUT4 #(
		.INIT('ha820)
	) name1673 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001 ,
		_w5721_
	);
	LUT3 #(
		.INIT('h1b)
	) name1674 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001 ,
		_w5722_
	);
	LUT4 #(
		.INIT('ha820)
	) name1675 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001 ,
		_w5723_
	);
	LUT3 #(
		.INIT('h1b)
	) name1676 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001 ,
		_w5724_
	);
	LUT4 #(
		.INIT('ha820)
	) name1677 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001 ,
		_w5725_
	);
	LUT3 #(
		.INIT('h1b)
	) name1678 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001 ,
		_w5726_
	);
	LUT4 #(
		.INIT('ha820)
	) name1679 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001 ,
		_w5727_
	);
	LUT4 #(
		.INIT('h0001)
	) name1680 (
		_w5721_,
		_w5723_,
		_w5725_,
		_w5727_,
		_w5728_
	);
	LUT3 #(
		.INIT('h2a)
	) name1681 (
		_w5712_,
		_w5719_,
		_w5728_,
		_w5729_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1682 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_MFALU_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w5730_
	);
	LUT4 #(
		.INIT('ha820)
	) name1683 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001 ,
		_w5731_
	);
	LUT4 #(
		.INIT('ha820)
	) name1684 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001 ,
		_w5732_
	);
	LUT2 #(
		.INIT('h1)
	) name1685 (
		_w5731_,
		_w5732_,
		_w5733_
	);
	LUT3 #(
		.INIT('h1b)
	) name1686 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001 ,
		_w5734_
	);
	LUT4 #(
		.INIT('ha820)
	) name1687 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001 ,
		_w5735_
	);
	LUT3 #(
		.INIT('h1b)
	) name1688 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001 ,
		_w5736_
	);
	LUT4 #(
		.INIT('ha820)
	) name1689 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001 ,
		_w5737_
	);
	LUT4 #(
		.INIT('ha820)
	) name1690 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001 ,
		_w5738_
	);
	LUT3 #(
		.INIT('h01)
	) name1691 (
		_w5737_,
		_w5738_,
		_w5735_,
		_w5739_
	);
	LUT3 #(
		.INIT('h2a)
	) name1692 (
		_w5730_,
		_w5733_,
		_w5739_,
		_w5740_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1693 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_MFSHT_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w5741_
	);
	LUT3 #(
		.INIT('h1b)
	) name1694 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[4]/P0001 ,
		_w5742_
	);
	LUT4 #(
		.INIT('ha820)
	) name1695 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[4]/P0001 ,
		_w5743_
	);
	LUT3 #(
		.INIT('h1b)
	) name1696 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001 ,
		_w5744_
	);
	LUT4 #(
		.INIT('ha820)
	) name1697 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001 ,
		_w5745_
	);
	LUT2 #(
		.INIT('h1)
	) name1698 (
		_w5743_,
		_w5745_,
		_w5746_
	);
	LUT3 #(
		.INIT('h1b)
	) name1699 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001 ,
		_w5747_
	);
	LUT4 #(
		.INIT('ha820)
	) name1700 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001 ,
		_w5748_
	);
	LUT3 #(
		.INIT('h1b)
	) name1701 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001 ,
		_w5749_
	);
	LUT4 #(
		.INIT('ha820)
	) name1702 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001 ,
		_w5750_
	);
	LUT3 #(
		.INIT('h1b)
	) name1703 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001 ,
		_w5751_
	);
	LUT4 #(
		.INIT('ha820)
	) name1704 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001 ,
		_w5752_
	);
	LUT3 #(
		.INIT('h01)
	) name1705 (
		_w5750_,
		_w5752_,
		_w5748_,
		_w5753_
	);
	LUT3 #(
		.INIT('h2a)
	) name1706 (
		_w5741_,
		_w5746_,
		_w5753_,
		_w5754_
	);
	LUT3 #(
		.INIT('h01)
	) name1707 (
		_w5740_,
		_w5754_,
		_w5729_,
		_w5755_
	);
	LUT2 #(
		.INIT('h8)
	) name1708 (
		_w5711_,
		_w5755_,
		_w5756_
	);
	LUT4 #(
		.INIT('h0100)
	) name1709 (
		_w5626_,
		_w5686_,
		_w5680_,
		_w5756_,
		_w5757_
	);
	LUT2 #(
		.INIT('h8)
	) name1710 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[13]/P0001 ,
		_w5758_
	);
	LUT3 #(
		.INIT('h08)
	) name1711 (
		_w5588_,
		_w5598_,
		_w5758_,
		_w5759_
	);
	LUT4 #(
		.INIT('h0133)
	) name1712 (
		\emc_DMDoe_reg/NET0131 ,
		_w5625_,
		_w5757_,
		_w5759_,
		_w5760_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		_w5563_,
		_w5550_,
		_w5761_
	);
	LUT4 #(
		.INIT('h2031)
	) name1714 (
		_w5117_,
		_w5337_,
		_w5761_,
		_w5760_,
		_w5762_
	);
	LUT4 #(
		.INIT('h4844)
	) name1715 (
		_w5156_,
		_w5190_,
		_w5286_,
		_w5288_,
		_w5763_
	);
	LUT4 #(
		.INIT('h2122)
	) name1716 (
		_w5156_,
		_w5189_,
		_w5286_,
		_w5288_,
		_w5764_
	);
	LUT3 #(
		.INIT('h01)
	) name1717 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5764_,
		_w5763_,
		_w5765_
	);
	LUT2 #(
		.INIT('h8)
	) name1718 (
		\core_dag_ilm1reg_I_reg[0]/NET0131 ,
		_w5181_,
		_w5766_
	);
	LUT4 #(
		.INIT('h7010)
	) name1719 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w5278_,
		_w5293_,
		_w5309_,
		_w5767_
	);
	LUT4 #(
		.INIT('h80e0)
	) name1720 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w5278_,
		_w5294_,
		_w5309_,
		_w5768_
	);
	LUT3 #(
		.INIT('h54)
	) name1721 (
		_w5190_,
		_w5767_,
		_w5768_,
		_w5769_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name1722 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5155_,
		_w5189_,
		_w5310_,
		_w5770_
	);
	LUT4 #(
		.INIT('h0045)
	) name1723 (
		_w5766_,
		_w5769_,
		_w5770_,
		_w5765_,
		_w5771_
	);
	LUT3 #(
		.INIT('ha8)
	) name1724 (
		\DM_rd0[0]_pad ,
		_w5610_,
		_w5612_,
		_w5772_
	);
	LUT4 #(
		.INIT('h135f)
	) name1725 (
		\DM_rdm[0]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w5773_
	);
	LUT4 #(
		.INIT('h135f)
	) name1726 (
		\DM_rd6[0]_pad ,
		\DM_rd7[0]_pad ,
		_w5596_,
		_w5591_,
		_w5774_
	);
	LUT2 #(
		.INIT('h8)
	) name1727 (
		_w5773_,
		_w5774_,
		_w5775_
	);
	LUT3 #(
		.INIT('h80)
	) name1728 (
		\DM_rd4[0]_pad ,
		_w5598_,
		_w5601_,
		_w5776_
	);
	LUT3 #(
		.INIT('h80)
	) name1729 (
		\DM_rd5[0]_pad ,
		_w5598_,
		_w5599_,
		_w5777_
	);
	LUT4 #(
		.INIT('h8000)
	) name1730 (
		\DM_rd2[0]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w5778_
	);
	LUT4 #(
		.INIT('h8000)
	) name1731 (
		\DM_rd1[0]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w5779_
	);
	LUT4 #(
		.INIT('h8000)
	) name1732 (
		\DM_rd3[0]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w5780_
	);
	LUT3 #(
		.INIT('h01)
	) name1733 (
		_w5779_,
		_w5780_,
		_w5778_,
		_w5781_
	);
	LUT3 #(
		.INIT('h10)
	) name1734 (
		_w5777_,
		_w5776_,
		_w5781_,
		_w5782_
	);
	LUT2 #(
		.INIT('h8)
	) name1735 (
		_w5775_,
		_w5782_,
		_w5783_
	);
	LUT2 #(
		.INIT('h4)
	) name1736 (
		_w5772_,
		_w5783_,
		_w5784_
	);
	LUT4 #(
		.INIT('h4000)
	) name1737 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[0]/P0001 ,
		_w5785_
	);
	LUT3 #(
		.INIT('h80)
	) name1738 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w5629_,
		_w5648_,
		_w5786_
	);
	LUT3 #(
		.INIT('h80)
	) name1739 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w5632_,
		_w5634_,
		_w5787_
	);
	LUT3 #(
		.INIT('h80)
	) name1740 (
		\PIO_oe[0]_pad ,
		_w5628_,
		_w5632_,
		_w5788_
	);
	LUT3 #(
		.INIT('h80)
	) name1741 (
		\sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w5634_,
		_w5635_,
		_w5789_
	);
	LUT4 #(
		.INIT('h0800)
	) name1742 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5790_
	);
	LUT3 #(
		.INIT('h80)
	) name1743 (
		\emc_WSCRext_reg_DO_reg[0]/NET0131 ,
		_w5670_,
		_w5790_,
		_w5791_
	);
	LUT4 #(
		.INIT('h0001)
	) name1744 (
		_w5787_,
		_w5788_,
		_w5789_,
		_w5791_,
		_w5792_
	);
	LUT3 #(
		.INIT('h80)
	) name1745 (
		\emc_WSCRreg_DO_reg[0]/NET0131 ,
		_w5631_,
		_w5632_,
		_w5793_
	);
	LUT4 #(
		.INIT('h0400)
	) name1746 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5794_
	);
	LUT2 #(
		.INIT('h8)
	) name1747 (
		_w5671_,
		_w5794_,
		_w5795_
	);
	LUT3 #(
		.INIT('h80)
	) name1748 (
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w5634_,
		_w5637_,
		_w5796_
	);
	LUT3 #(
		.INIT('h80)
	) name1749 (
		\sport1_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w5631_,
		_w5639_,
		_w5797_
	);
	LUT4 #(
		.INIT('h0001)
	) name1750 (
		_w5793_,
		_w5796_,
		_w5797_,
		_w5795_,
		_w5798_
	);
	LUT3 #(
		.INIT('h40)
	) name1751 (
		_w5786_,
		_w5792_,
		_w5798_,
		_w5799_
	);
	LUT3 #(
		.INIT('h80)
	) name1752 (
		\bdma_BEAD_reg[0]/NET0131 ,
		_w5629_,
		_w5644_,
		_w5800_
	);
	LUT3 #(
		.INIT('h80)
	) name1753 (
		\bdma_BCTL_reg[0]/NET0131 ,
		_w5627_,
		_w5629_,
		_w5801_
	);
	LUT2 #(
		.INIT('h1)
	) name1754 (
		_w5800_,
		_w5801_,
		_w5802_
	);
	LUT2 #(
		.INIT('h8)
	) name1755 (
		_w5799_,
		_w5802_,
		_w5803_
	);
	LUT4 #(
		.INIT('h0200)
	) name1756 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5804_
	);
	LUT4 #(
		.INIT('h8000)
	) name1757 (
		\bdma_BOVL_reg[0]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w5805_
	);
	LUT4 #(
		.INIT('h8000)
	) name1758 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w5806_
	);
	LUT3 #(
		.INIT('h80)
	) name1759 (
		\tm_TCR_TMP_reg[0]/NET0131 ,
		_w5631_,
		_w5637_,
		_w5807_
	);
	LUT3 #(
		.INIT('h80)
	) name1760 (
		\pio_pmask_reg_DO_reg[0]/NET0131 ,
		_w5628_,
		_w5660_,
		_w5808_
	);
	LUT2 #(
		.INIT('h8)
	) name1761 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5809_
	);
	LUT4 #(
		.INIT('h8000)
	) name1762 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5810_
	);
	LUT3 #(
		.INIT('h80)
	) name1763 (
		\sport1_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w5670_,
		_w5810_,
		_w5811_
	);
	LUT3 #(
		.INIT('h80)
	) name1764 (
		\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w5648_,
		_w5634_,
		_w5812_
	);
	LUT4 #(
		.INIT('h0001)
	) name1765 (
		_w5807_,
		_w5808_,
		_w5811_,
		_w5812_,
		_w5813_
	);
	LUT3 #(
		.INIT('h80)
	) name1766 (
		\memc_usysr_DO_reg[0]/NET0131 ,
		_w5631_,
		_w5660_,
		_w5814_
	);
	LUT3 #(
		.INIT('h80)
	) name1767 (
		\sport0_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w5627_,
		_w5634_,
		_w5815_
	);
	LUT3 #(
		.INIT('h80)
	) name1768 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w5628_,
		_w5639_,
		_w5816_
	);
	LUT3 #(
		.INIT('h80)
	) name1769 (
		\pio_PINT_reg[0]/NET0131 ,
		_w5670_,
		_w5672_,
		_w5817_
	);
	LUT4 #(
		.INIT('h0001)
	) name1770 (
		_w5814_,
		_w5815_,
		_w5816_,
		_w5817_,
		_w5818_
	);
	LUT3 #(
		.INIT('h80)
	) name1771 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w5644_,
		_w5634_,
		_w5819_
	);
	LUT3 #(
		.INIT('h80)
	) name1772 (
		\clkc_ckr_reg_DO_reg[0]/NET0131 ,
		_w5631_,
		_w5644_,
		_w5820_
	);
	LUT3 #(
		.INIT('h80)
	) name1773 (
		\sport0_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w5634_,
		_w5660_,
		_w5821_
	);
	LUT3 #(
		.INIT('h80)
	) name1774 (
		\PIO_out[0]_pad ,
		_w5628_,
		_w5635_,
		_w5822_
	);
	LUT4 #(
		.INIT('h0001)
	) name1775 (
		_w5819_,
		_w5820_,
		_w5821_,
		_w5822_,
		_w5823_
	);
	LUT2 #(
		.INIT('h8)
	) name1776 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5824_
	);
	LUT3 #(
		.INIT('h80)
	) name1777 (
		\idma_DOVL_reg[0]/NET0131 ,
		_w5804_,
		_w5824_,
		_w5825_
	);
	LUT3 #(
		.INIT('h80)
	) name1778 (
		\tm_tpr_reg_DO_reg[0]/NET0131 ,
		_w5631_,
		_w5635_,
		_w5826_
	);
	LUT3 #(
		.INIT('h80)
	) name1779 (
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w5634_,
		_w5639_,
		_w5827_
	);
	LUT3 #(
		.INIT('h80)
	) name1780 (
		\tm_tsr_reg_DO_reg[0]/NET0131 ,
		_w5627_,
		_w5631_,
		_w5828_
	);
	LUT4 #(
		.INIT('h0001)
	) name1781 (
		_w5825_,
		_w5826_,
		_w5827_,
		_w5828_,
		_w5829_
	);
	LUT4 #(
		.INIT('h8000)
	) name1782 (
		_w5823_,
		_w5829_,
		_w5813_,
		_w5818_,
		_w5830_
	);
	LUT3 #(
		.INIT('h10)
	) name1783 (
		_w5806_,
		_w5805_,
		_w5830_,
		_w5831_
	);
	LUT3 #(
		.INIT('h2a)
	) name1784 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w5803_,
		_w5831_,
		_w5832_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1785 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4124_,
		_w4117_,
		_w4137_,
		_w5833_
	);
	LUT4 #(
		.INIT('h135f)
	) name1786 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w5834_
	);
	LUT4 #(
		.INIT('h135f)
	) name1787 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_ICNTL_reg_DO_reg[0]/NET0131 ,
		_w5835_
	);
	LUT2 #(
		.INIT('h8)
	) name1788 (
		_w5834_,
		_w5835_,
		_w5836_
	);
	LUT3 #(
		.INIT('ha8)
	) name1789 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w5837_
	);
	LUT4 #(
		.INIT('h135f)
	) name1790 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w5838_
	);
	LUT4 #(
		.INIT('h135f)
	) name1791 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\core_c_psq_SSTAT_reg[0]/NET0131 ,
		_w5839_
	);
	LUT3 #(
		.INIT('h40)
	) name1792 (
		_w5837_,
		_w5838_,
		_w5839_,
		_w5840_
	);
	LUT2 #(
		.INIT('h8)
	) name1793 (
		_w5836_,
		_w5840_,
		_w5841_
	);
	LUT3 #(
		.INIT('h8a)
	) name1794 (
		_w5681_,
		_w5833_,
		_w5841_,
		_w5842_
	);
	LUT4 #(
		.INIT('h135f)
	) name1795 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131 ,
		_w5843_
	);
	LUT4 #(
		.INIT('h135f)
	) name1796 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131 ,
		_w5844_
	);
	LUT2 #(
		.INIT('h8)
	) name1797 (
		_w5843_,
		_w5844_,
		_w5845_
	);
	LUT4 #(
		.INIT('h135f)
	) name1798 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131 ,
		_w5846_
	);
	LUT4 #(
		.INIT('h135f)
	) name1799 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w5847_
	);
	LUT4 #(
		.INIT('h135f)
	) name1800 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 ,
		_w5848_
	);
	LUT4 #(
		.INIT('h135f)
	) name1801 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131 ,
		_w5849_
	);
	LUT4 #(
		.INIT('h8000)
	) name1802 (
		_w5848_,
		_w5849_,
		_w5846_,
		_w5847_,
		_w5850_
	);
	LUT3 #(
		.INIT('h2a)
	) name1803 (
		_w5697_,
		_w5845_,
		_w5850_,
		_w5851_
	);
	LUT4 #(
		.INIT('h135f)
	) name1804 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w5852_
	);
	LUT4 #(
		.INIT('h135f)
	) name1805 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131 ,
		_w5853_
	);
	LUT2 #(
		.INIT('h8)
	) name1806 (
		_w5852_,
		_w5853_,
		_w5854_
	);
	LUT4 #(
		.INIT('h135f)
	) name1807 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w5855_
	);
	LUT4 #(
		.INIT('h135f)
	) name1808 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131 ,
		_w5856_
	);
	LUT4 #(
		.INIT('h135f)
	) name1809 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131 ,
		_w5857_
	);
	LUT4 #(
		.INIT('h135f)
	) name1810 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131 ,
		_w5858_
	);
	LUT4 #(
		.INIT('h8000)
	) name1811 (
		_w5857_,
		_w5858_,
		_w5855_,
		_w5856_,
		_w5859_
	);
	LUT4 #(
		.INIT('h135f)
	) name1812 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport1_txctl_TX_reg[0]/P0001 ,
		_w5860_
	);
	LUT4 #(
		.INIT('h135f)
	) name1813 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport1_rxctl_RX_reg[0]/P0001 ,
		_w5861_
	);
	LUT3 #(
		.INIT('h2a)
	) name1814 (
		_w5706_,
		_w5860_,
		_w5861_,
		_w5862_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1815 (
		_w5687_,
		_w5854_,
		_w5859_,
		_w5862_,
		_w5863_
	);
	LUT2 #(
		.INIT('h4)
	) name1816 (
		_w5851_,
		_w5863_,
		_w5864_
	);
	LUT3 #(
		.INIT('h1b)
	) name1817 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 ,
		_w5865_
	);
	LUT4 #(
		.INIT('ha820)
	) name1818 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 ,
		_w5866_
	);
	LUT3 #(
		.INIT('h1b)
	) name1819 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001 ,
		_w5867_
	);
	LUT4 #(
		.INIT('ha820)
	) name1820 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001 ,
		_w5868_
	);
	LUT3 #(
		.INIT('h1b)
	) name1821 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001 ,
		_w5869_
	);
	LUT4 #(
		.INIT('ha820)
	) name1822 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001 ,
		_w5870_
	);
	LUT3 #(
		.INIT('h01)
	) name1823 (
		_w5868_,
		_w5870_,
		_w5866_,
		_w5871_
	);
	LUT3 #(
		.INIT('h1b)
	) name1824 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 ,
		_w5872_
	);
	LUT4 #(
		.INIT('ha820)
	) name1825 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 ,
		_w5873_
	);
	LUT3 #(
		.INIT('h1b)
	) name1826 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001 ,
		_w5874_
	);
	LUT4 #(
		.INIT('ha820)
	) name1827 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001 ,
		_w5875_
	);
	LUT3 #(
		.INIT('h1b)
	) name1828 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001 ,
		_w5876_
	);
	LUT4 #(
		.INIT('ha820)
	) name1829 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001 ,
		_w5877_
	);
	LUT3 #(
		.INIT('h1b)
	) name1830 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001 ,
		_w5878_
	);
	LUT4 #(
		.INIT('ha820)
	) name1831 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001 ,
		_w5879_
	);
	LUT4 #(
		.INIT('h0001)
	) name1832 (
		_w5873_,
		_w5875_,
		_w5877_,
		_w5879_,
		_w5880_
	);
	LUT3 #(
		.INIT('h2a)
	) name1833 (
		_w5712_,
		_w5871_,
		_w5880_,
		_w5881_
	);
	LUT3 #(
		.INIT('h1b)
	) name1834 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[0]/P0001 ,
		_w5882_
	);
	LUT4 #(
		.INIT('ha820)
	) name1835 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[0]/P0001 ,
		_w5883_
	);
	LUT3 #(
		.INIT('h1b)
	) name1836 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001 ,
		_w5884_
	);
	LUT4 #(
		.INIT('ha820)
	) name1837 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001 ,
		_w5885_
	);
	LUT2 #(
		.INIT('h1)
	) name1838 (
		_w5883_,
		_w5885_,
		_w5886_
	);
	LUT3 #(
		.INIT('h1b)
	) name1839 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001 ,
		_w5887_
	);
	LUT4 #(
		.INIT('ha820)
	) name1840 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001 ,
		_w5888_
	);
	LUT3 #(
		.INIT('h1b)
	) name1841 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001 ,
		_w5889_
	);
	LUT4 #(
		.INIT('ha820)
	) name1842 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001 ,
		_w5890_
	);
	LUT3 #(
		.INIT('h1b)
	) name1843 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001 ,
		_w5891_
	);
	LUT4 #(
		.INIT('ha820)
	) name1844 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001 ,
		_w5892_
	);
	LUT3 #(
		.INIT('h01)
	) name1845 (
		_w5890_,
		_w5892_,
		_w5888_,
		_w5893_
	);
	LUT3 #(
		.INIT('h2a)
	) name1846 (
		_w5741_,
		_w5886_,
		_w5893_,
		_w5894_
	);
	LUT3 #(
		.INIT('h1b)
	) name1847 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001 ,
		_w5895_
	);
	LUT4 #(
		.INIT('ha820)
	) name1848 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001 ,
		_w5896_
	);
	LUT2 #(
		.INIT('h8)
	) name1849 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w5897_
	);
	LUT2 #(
		.INIT('h1)
	) name1850 (
		_w5896_,
		_w5897_,
		_w5898_
	);
	LUT3 #(
		.INIT('h1b)
	) name1851 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001 ,
		_w5899_
	);
	LUT4 #(
		.INIT('ha820)
	) name1852 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001 ,
		_w5900_
	);
	LUT3 #(
		.INIT('h1b)
	) name1853 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001 ,
		_w5901_
	);
	LUT4 #(
		.INIT('ha820)
	) name1854 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001 ,
		_w5902_
	);
	LUT4 #(
		.INIT('ha820)
	) name1855 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001 ,
		_w5903_
	);
	LUT4 #(
		.INIT('ha820)
	) name1856 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001 ,
		_w5904_
	);
	LUT4 #(
		.INIT('h0001)
	) name1857 (
		_w5900_,
		_w5902_,
		_w5903_,
		_w5904_,
		_w5905_
	);
	LUT3 #(
		.INIT('h2a)
	) name1858 (
		_w5730_,
		_w5898_,
		_w5905_,
		_w5906_
	);
	LUT3 #(
		.INIT('h01)
	) name1859 (
		_w5894_,
		_w5906_,
		_w5881_,
		_w5907_
	);
	LUT2 #(
		.INIT('h8)
	) name1860 (
		_w5864_,
		_w5907_,
		_w5908_
	);
	LUT2 #(
		.INIT('h4)
	) name1861 (
		_w5842_,
		_w5908_,
		_w5909_
	);
	LUT3 #(
		.INIT('h10)
	) name1862 (
		_w5785_,
		_w5832_,
		_w5909_,
		_w5910_
	);
	LUT4 #(
		.INIT('h5455)
	) name1863 (
		\emc_DMDoe_reg/NET0131 ,
		_w5785_,
		_w5832_,
		_w5909_,
		_w5911_
	);
	LUT2 #(
		.INIT('h8)
	) name1864 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[0]/P0001 ,
		_w5912_
	);
	LUT3 #(
		.INIT('h08)
	) name1865 (
		_w5588_,
		_w5598_,
		_w5912_,
		_w5913_
	);
	LUT3 #(
		.INIT('h45)
	) name1866 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w5914_
	);
	LUT3 #(
		.INIT('h4c)
	) name1867 (
		_w5117_,
		_w5337_,
		_w5914_,
		_w5915_
	);
	LUT4 #(
		.INIT('h0133)
	) name1868 (
		_w5117_,
		_w5762_,
		_w5771_,
		_w5915_,
		_w5916_
	);
	LUT4 #(
		.INIT('hf101)
	) name1869 (
		_w5339_,
		_w5582_,
		_w5586_,
		_w5916_,
		_w5917_
	);
	LUT4 #(
		.INIT('h1411)
	) name1870 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5156_,
		_w5286_,
		_w5288_,
		_w5918_
	);
	LUT4 #(
		.INIT('h556a)
	) name1871 (
		_w5257_,
		_w5302_,
		_w5303_,
		_w5305_,
		_w5919_
	);
	LUT3 #(
		.INIT('h10)
	) name1872 (
		_w5767_,
		_w5918_,
		_w5919_,
		_w5920_
	);
	LUT4 #(
		.INIT('h002a)
	) name1873 (
		\core_dag_ilm1reg_I_reg[10]/NET0131 ,
		_w5122_,
		_w5153_,
		_w5253_,
		_w5921_
	);
	LUT2 #(
		.INIT('h9)
	) name1874 (
		_w5252_,
		_w5259_,
		_w5922_
	);
	LUT3 #(
		.INIT('h4b)
	) name1875 (
		_w5251_,
		_w5274_,
		_w5922_,
		_w5923_
	);
	LUT4 #(
		.INIT('h0133)
	) name1876 (
		_w5767_,
		_w5921_,
		_w5918_,
		_w5923_,
		_w5924_
	);
	LUT3 #(
		.INIT('ha8)
	) name1877 (
		\DM_rd0[10]_pad ,
		_w5610_,
		_w5612_,
		_w5925_
	);
	LUT4 #(
		.INIT('h135f)
	) name1878 (
		\DM_rdm[10]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w5926_
	);
	LUT4 #(
		.INIT('h135f)
	) name1879 (
		\DM_rd6[10]_pad ,
		\DM_rd7[10]_pad ,
		_w5596_,
		_w5591_,
		_w5927_
	);
	LUT2 #(
		.INIT('h8)
	) name1880 (
		_w5926_,
		_w5927_,
		_w5928_
	);
	LUT3 #(
		.INIT('h80)
	) name1881 (
		\DM_rd5[10]_pad ,
		_w5598_,
		_w5599_,
		_w5929_
	);
	LUT3 #(
		.INIT('h80)
	) name1882 (
		\DM_rd4[10]_pad ,
		_w5598_,
		_w5601_,
		_w5930_
	);
	LUT4 #(
		.INIT('h8000)
	) name1883 (
		\DM_rd2[10]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w5931_
	);
	LUT4 #(
		.INIT('h8000)
	) name1884 (
		\DM_rd1[10]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w5932_
	);
	LUT4 #(
		.INIT('h8000)
	) name1885 (
		\DM_rd3[10]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w5933_
	);
	LUT3 #(
		.INIT('h01)
	) name1886 (
		_w5932_,
		_w5933_,
		_w5931_,
		_w5934_
	);
	LUT3 #(
		.INIT('h10)
	) name1887 (
		_w5930_,
		_w5929_,
		_w5934_,
		_w5935_
	);
	LUT2 #(
		.INIT('h8)
	) name1888 (
		_w5928_,
		_w5935_,
		_w5936_
	);
	LUT2 #(
		.INIT('h4)
	) name1889 (
		_w5925_,
		_w5936_,
		_w5937_
	);
	LUT4 #(
		.INIT('h4000)
	) name1890 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[10]/P0001 ,
		_w5938_
	);
	LUT3 #(
		.INIT('h80)
	) name1891 (
		\bdma_BCTL_reg[10]/NET0131 ,
		_w5627_,
		_w5629_,
		_w5939_
	);
	LUT3 #(
		.INIT('h80)
	) name1892 (
		\emc_WSCRreg_DO_reg[10]/NET0131 ,
		_w5631_,
		_w5632_,
		_w5940_
	);
	LUT3 #(
		.INIT('h80)
	) name1893 (
		\tm_tpr_reg_DO_reg[10]/NET0131 ,
		_w5631_,
		_w5635_,
		_w5941_
	);
	LUT3 #(
		.INIT('h80)
	) name1894 (
		\sport0_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w5632_,
		_w5634_,
		_w5942_
	);
	LUT3 #(
		.INIT('h80)
	) name1895 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		_w5631_,
		_w5637_,
		_w5943_
	);
	LUT4 #(
		.INIT('h0001)
	) name1896 (
		_w5940_,
		_w5941_,
		_w5942_,
		_w5943_,
		_w5944_
	);
	LUT3 #(
		.INIT('h80)
	) name1897 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w5631_,
		_w5639_,
		_w5945_
	);
	LUT4 #(
		.INIT('h8000)
	) name1898 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		_w5631_,
		_w5639_,
		_w5946_
	);
	LUT3 #(
		.INIT('h80)
	) name1899 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w5634_,
		_w5660_,
		_w5947_
	);
	LUT4 #(
		.INIT('h8000)
	) name1900 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		_w5634_,
		_w5660_,
		_w5948_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w5946_,
		_w5948_,
		_w5949_
	);
	LUT3 #(
		.INIT('h40)
	) name1902 (
		_w5939_,
		_w5944_,
		_w5949_,
		_w5950_
	);
	LUT3 #(
		.INIT('h80)
	) name1903 (
		\bdma_BEAD_reg[10]/NET0131 ,
		_w5629_,
		_w5644_,
		_w5951_
	);
	LUT3 #(
		.INIT('h80)
	) name1904 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w5629_,
		_w5648_,
		_w5952_
	);
	LUT2 #(
		.INIT('h1)
	) name1905 (
		_w5951_,
		_w5952_,
		_w5953_
	);
	LUT4 #(
		.INIT('h8000)
	) name1906 (
		\bdma_BOVL_reg[10]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w5954_
	);
	LUT4 #(
		.INIT('h8000)
	) name1907 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w5955_
	);
	LUT3 #(
		.INIT('h80)
	) name1908 (
		\sport0_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w5627_,
		_w5634_,
		_w5956_
	);
	LUT3 #(
		.INIT('h80)
	) name1909 (
		\sport1_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w5670_,
		_w5810_,
		_w5957_
	);
	LUT3 #(
		.INIT('h80)
	) name1910 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w5628_,
		_w5639_,
		_w5958_
	);
	LUT3 #(
		.INIT('h01)
	) name1911 (
		_w5957_,
		_w5958_,
		_w5956_,
		_w5959_
	);
	LUT3 #(
		.INIT('h80)
	) name1912 (
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w5634_,
		_w5637_,
		_w5960_
	);
	LUT3 #(
		.INIT('h80)
	) name1913 (
		\memc_usysr_DO_reg[10]/NET0131 ,
		_w5631_,
		_w5660_,
		_w5961_
	);
	LUT3 #(
		.INIT('h80)
	) name1914 (
		\sport1_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w5644_,
		_w5634_,
		_w5962_
	);
	LUT3 #(
		.INIT('h80)
	) name1915 (
		\clkc_ckr_reg_DO_reg[10]/NET0131 ,
		_w5631_,
		_w5644_,
		_w5963_
	);
	LUT4 #(
		.INIT('h0001)
	) name1916 (
		_w5960_,
		_w5961_,
		_w5962_,
		_w5963_,
		_w5964_
	);
	LUT3 #(
		.INIT('h80)
	) name1917 (
		\idma_DOVL_reg[10]/NET0131 ,
		_w5804_,
		_w5824_,
		_w5965_
	);
	LUT3 #(
		.INIT('h80)
	) name1918 (
		\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w5634_,
		_w5635_,
		_w5966_
	);
	LUT3 #(
		.INIT('h80)
	) name1919 (
		\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w5648_,
		_w5634_,
		_w5967_
	);
	LUT3 #(
		.INIT('h80)
	) name1920 (
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w5634_,
		_w5639_,
		_w5968_
	);
	LUT4 #(
		.INIT('h0001)
	) name1921 (
		_w5965_,
		_w5966_,
		_w5967_,
		_w5968_,
		_w5969_
	);
	LUT4 #(
		.INIT('h4000)
	) name1922 (
		_w5955_,
		_w5959_,
		_w5964_,
		_w5969_,
		_w5970_
	);
	LUT4 #(
		.INIT('h4000)
	) name1923 (
		_w5954_,
		_w5950_,
		_w5953_,
		_w5970_,
		_w5971_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1924 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4250_,
		_w4247_,
		_w4255_,
		_w5972_
	);
	LUT3 #(
		.INIT('ha8)
	) name1925 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w5973_
	);
	LUT4 #(
		.INIT('h135f)
	) name1926 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w5974_
	);
	LUT2 #(
		.INIT('h4)
	) name1927 (
		_w5973_,
		_w5974_,
		_w5975_
	);
	LUT3 #(
		.INIT('h8a)
	) name1928 (
		_w5681_,
		_w5972_,
		_w5975_,
		_w5976_
	);
	LUT4 #(
		.INIT('h135f)
	) name1929 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131 ,
		_w5977_
	);
	LUT4 #(
		.INIT('h135f)
	) name1930 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 ,
		_w5978_
	);
	LUT2 #(
		.INIT('h8)
	) name1931 (
		_w5977_,
		_w5978_,
		_w5979_
	);
	LUT4 #(
		.INIT('h135f)
	) name1932 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131 ,
		_w5980_
	);
	LUT4 #(
		.INIT('h135f)
	) name1933 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131 ,
		_w5981_
	);
	LUT4 #(
		.INIT('h135f)
	) name1934 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131 ,
		_w5982_
	);
	LUT4 #(
		.INIT('h135f)
	) name1935 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131 ,
		_w5983_
	);
	LUT4 #(
		.INIT('h8000)
	) name1936 (
		_w5982_,
		_w5983_,
		_w5980_,
		_w5981_,
		_w5984_
	);
	LUT3 #(
		.INIT('h2a)
	) name1937 (
		_w5687_,
		_w5979_,
		_w5984_,
		_w5985_
	);
	LUT4 #(
		.INIT('h135f)
	) name1938 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131 ,
		_w5986_
	);
	LUT4 #(
		.INIT('h135f)
	) name1939 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131 ,
		_w5987_
	);
	LUT2 #(
		.INIT('h8)
	) name1940 (
		_w5986_,
		_w5987_,
		_w5988_
	);
	LUT4 #(
		.INIT('h135f)
	) name1941 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 ,
		_w5989_
	);
	LUT4 #(
		.INIT('h135f)
	) name1942 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131 ,
		_w5990_
	);
	LUT4 #(
		.INIT('h135f)
	) name1943 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131 ,
		_w5991_
	);
	LUT4 #(
		.INIT('h135f)
	) name1944 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131 ,
		_w5992_
	);
	LUT4 #(
		.INIT('h8000)
	) name1945 (
		_w5991_,
		_w5992_,
		_w5989_,
		_w5990_,
		_w5993_
	);
	LUT4 #(
		.INIT('h135f)
	) name1946 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[10]/P0001 ,
		\sport1_txctl_TX_reg[10]/P0001 ,
		_w5994_
	);
	LUT4 #(
		.INIT('h153f)
	) name1947 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[10]/P0001 ,
		\sport1_rxctl_RX_reg[10]/P0001 ,
		_w5995_
	);
	LUT3 #(
		.INIT('h2a)
	) name1948 (
		_w5706_,
		_w5994_,
		_w5995_,
		_w5996_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1949 (
		_w5697_,
		_w5988_,
		_w5993_,
		_w5996_,
		_w5997_
	);
	LUT2 #(
		.INIT('h4)
	) name1950 (
		_w5985_,
		_w5997_,
		_w5998_
	);
	LUT3 #(
		.INIT('h1b)
	) name1951 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001 ,
		_w5999_
	);
	LUT4 #(
		.INIT('ha820)
	) name1952 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001 ,
		_w6000_
	);
	LUT3 #(
		.INIT('h1b)
	) name1953 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001 ,
		_w6001_
	);
	LUT4 #(
		.INIT('ha820)
	) name1954 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001 ,
		_w6002_
	);
	LUT3 #(
		.INIT('h1b)
	) name1955 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001 ,
		_w6003_
	);
	LUT4 #(
		.INIT('ha820)
	) name1956 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001 ,
		_w6004_
	);
	LUT3 #(
		.INIT('h01)
	) name1957 (
		_w6002_,
		_w6004_,
		_w6000_,
		_w6005_
	);
	LUT3 #(
		.INIT('h2a)
	) name1958 (
		_w5741_,
		_w5746_,
		_w6005_,
		_w6006_
	);
	LUT3 #(
		.INIT('h1b)
	) name1959 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001 ,
		_w6007_
	);
	LUT4 #(
		.INIT('ha820)
	) name1960 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001 ,
		_w6008_
	);
	LUT3 #(
		.INIT('h1b)
	) name1961 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001 ,
		_w6009_
	);
	LUT4 #(
		.INIT('ha820)
	) name1962 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001 ,
		_w6010_
	);
	LUT3 #(
		.INIT('h1b)
	) name1963 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001 ,
		_w6011_
	);
	LUT4 #(
		.INIT('ha820)
	) name1964 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001 ,
		_w6012_
	);
	LUT3 #(
		.INIT('h01)
	) name1965 (
		_w6010_,
		_w6012_,
		_w6008_,
		_w6013_
	);
	LUT3 #(
		.INIT('h1b)
	) name1966 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 ,
		_w6014_
	);
	LUT4 #(
		.INIT('ha820)
	) name1967 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 ,
		_w6015_
	);
	LUT3 #(
		.INIT('h1b)
	) name1968 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001 ,
		_w6016_
	);
	LUT4 #(
		.INIT('ha820)
	) name1969 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001 ,
		_w6017_
	);
	LUT3 #(
		.INIT('h1b)
	) name1970 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001 ,
		_w6018_
	);
	LUT4 #(
		.INIT('ha820)
	) name1971 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001 ,
		_w6019_
	);
	LUT4 #(
		.INIT('h0001)
	) name1972 (
		_w5714_,
		_w6015_,
		_w6017_,
		_w6019_,
		_w6020_
	);
	LUT3 #(
		.INIT('h2a)
	) name1973 (
		_w5712_,
		_w6013_,
		_w6020_,
		_w6021_
	);
	LUT4 #(
		.INIT('ha820)
	) name1974 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001 ,
		_w6022_
	);
	LUT3 #(
		.INIT('h1b)
	) name1975 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001 ,
		_w6023_
	);
	LUT4 #(
		.INIT('ha820)
	) name1976 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001 ,
		_w6024_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		_w6022_,
		_w6024_,
		_w6025_
	);
	LUT3 #(
		.INIT('h1b)
	) name1978 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001 ,
		_w6026_
	);
	LUT4 #(
		.INIT('ha820)
	) name1979 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001 ,
		_w6027_
	);
	LUT3 #(
		.INIT('h1b)
	) name1980 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001 ,
		_w6028_
	);
	LUT4 #(
		.INIT('ha820)
	) name1981 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001 ,
		_w6029_
	);
	LUT4 #(
		.INIT('ha820)
	) name1982 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001 ,
		_w6030_
	);
	LUT3 #(
		.INIT('h01)
	) name1983 (
		_w6029_,
		_w6030_,
		_w6027_,
		_w6031_
	);
	LUT3 #(
		.INIT('h2a)
	) name1984 (
		_w5730_,
		_w6025_,
		_w6031_,
		_w6032_
	);
	LUT3 #(
		.INIT('h01)
	) name1985 (
		_w6021_,
		_w6032_,
		_w6006_,
		_w6033_
	);
	LUT2 #(
		.INIT('h8)
	) name1986 (
		_w5998_,
		_w6033_,
		_w6034_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1987 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w5971_,
		_w5976_,
		_w6034_,
		_w6035_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[10]/P0001 ,
		_w6036_
	);
	LUT3 #(
		.INIT('h08)
	) name1989 (
		_w5588_,
		_w5598_,
		_w6036_,
		_w6037_
	);
	LUT4 #(
		.INIT('hba00)
	) name1990 (
		\emc_DMDoe_reg/NET0131 ,
		_w5938_,
		_w6035_,
		_w6037_,
		_w6038_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		_w5937_,
		_w6038_,
		_w6039_
	);
	LUT3 #(
		.INIT('hc4)
	) name1992 (
		_w5117_,
		_w5337_,
		_w6039_,
		_w6040_
	);
	LUT4 #(
		.INIT('hef00)
	) name1993 (
		_w5117_,
		_w5920_,
		_w5924_,
		_w6040_,
		_w6041_
	);
	LUT3 #(
		.INIT('ha8)
	) name1994 (
		\DM_rd0[3]_pad ,
		_w5610_,
		_w5612_,
		_w6042_
	);
	LUT4 #(
		.INIT('h135f)
	) name1995 (
		\DM_rdm[3]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w6043_
	);
	LUT4 #(
		.INIT('h135f)
	) name1996 (
		\DM_rd6[3]_pad ,
		\DM_rd7[3]_pad ,
		_w5596_,
		_w5591_,
		_w6044_
	);
	LUT2 #(
		.INIT('h8)
	) name1997 (
		_w6043_,
		_w6044_,
		_w6045_
	);
	LUT3 #(
		.INIT('h80)
	) name1998 (
		\DM_rd5[3]_pad ,
		_w5598_,
		_w5599_,
		_w6046_
	);
	LUT3 #(
		.INIT('h80)
	) name1999 (
		\DM_rd4[3]_pad ,
		_w5598_,
		_w5601_,
		_w6047_
	);
	LUT4 #(
		.INIT('h8000)
	) name2000 (
		\DM_rd2[3]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w6048_
	);
	LUT4 #(
		.INIT('h8000)
	) name2001 (
		\DM_rd1[3]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w6049_
	);
	LUT4 #(
		.INIT('h8000)
	) name2002 (
		\DM_rd3[3]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w6050_
	);
	LUT3 #(
		.INIT('h01)
	) name2003 (
		_w6049_,
		_w6050_,
		_w6048_,
		_w6051_
	);
	LUT3 #(
		.INIT('h10)
	) name2004 (
		_w6047_,
		_w6046_,
		_w6051_,
		_w6052_
	);
	LUT2 #(
		.INIT('h8)
	) name2005 (
		_w6045_,
		_w6052_,
		_w6053_
	);
	LUT2 #(
		.INIT('h4)
	) name2006 (
		_w6042_,
		_w6053_,
		_w6054_
	);
	LUT4 #(
		.INIT('h4000)
	) name2007 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[3]/P0001 ,
		_w6055_
	);
	LUT3 #(
		.INIT('h80)
	) name2008 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w5629_,
		_w5648_,
		_w6056_
	);
	LUT3 #(
		.INIT('h80)
	) name2009 (
		\emc_WSCRreg_DO_reg[3]/NET0131 ,
		_w5631_,
		_w5632_,
		_w6057_
	);
	LUT3 #(
		.INIT('h80)
	) name2010 (
		\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w5634_,
		_w5635_,
		_w6058_
	);
	LUT3 #(
		.INIT('h80)
	) name2011 (
		\sport1_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w5631_,
		_w5639_,
		_w6059_
	);
	LUT3 #(
		.INIT('h80)
	) name2012 (
		\tm_tsr_reg_DO_reg[3]/NET0131 ,
		_w5627_,
		_w5631_,
		_w6060_
	);
	LUT4 #(
		.INIT('h0001)
	) name2013 (
		_w6057_,
		_w6058_,
		_w6059_,
		_w6060_,
		_w6061_
	);
	LUT3 #(
		.INIT('h80)
	) name2014 (
		\idma_DOVL_reg[3]/NET0131 ,
		_w5804_,
		_w5824_,
		_w6062_
	);
	LUT3 #(
		.INIT('h80)
	) name2015 (
		\sport0_regs_AUTOreg_DO_reg[3]/NET0131 ,
		_w5627_,
		_w5634_,
		_w6063_
	);
	LUT3 #(
		.INIT('h80)
	) name2016 (
		\tm_tpr_reg_DO_reg[3]/NET0131 ,
		_w5631_,
		_w5635_,
		_w6064_
	);
	LUT4 #(
		.INIT('h0001)
	) name2017 (
		_w5795_,
		_w6062_,
		_w6063_,
		_w6064_,
		_w6065_
	);
	LUT3 #(
		.INIT('h40)
	) name2018 (
		_w6056_,
		_w6061_,
		_w6065_,
		_w6066_
	);
	LUT3 #(
		.INIT('h80)
	) name2019 (
		\bdma_BEAD_reg[3]/NET0131 ,
		_w5629_,
		_w5644_,
		_w6067_
	);
	LUT3 #(
		.INIT('h80)
	) name2020 (
		\bdma_BCTL_reg[3]/NET0131 ,
		_w5627_,
		_w5629_,
		_w6068_
	);
	LUT2 #(
		.INIT('h1)
	) name2021 (
		_w6067_,
		_w6068_,
		_w6069_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		_w6066_,
		_w6069_,
		_w6070_
	);
	LUT4 #(
		.INIT('h8000)
	) name2023 (
		\bdma_BOVL_reg[3]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w6071_
	);
	LUT4 #(
		.INIT('h8000)
	) name2024 (
		\bdma_BWCOUNT_reg[3]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w6072_
	);
	LUT3 #(
		.INIT('h80)
	) name2025 (
		\pio_pmask_reg_DO_reg[3]/NET0131 ,
		_w5628_,
		_w5660_,
		_w6073_
	);
	LUT3 #(
		.INIT('h80)
	) name2026 (
		\sport0_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w5634_,
		_w5660_,
		_w6074_
	);
	LUT3 #(
		.INIT('h80)
	) name2027 (
		\sport1_regs_AUTOreg_DO_reg[3]/NET0131 ,
		_w5670_,
		_w5810_,
		_w6075_
	);
	LUT3 #(
		.INIT('h80)
	) name2028 (
		\tm_TCR_TMP_reg[3]/NET0131 ,
		_w5631_,
		_w5637_,
		_w6076_
	);
	LUT4 #(
		.INIT('h0001)
	) name2029 (
		_w6073_,
		_w6074_,
		_w6075_,
		_w6076_,
		_w6077_
	);
	LUT3 #(
		.INIT('h80)
	) name2030 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w5632_,
		_w5634_,
		_w6078_
	);
	LUT3 #(
		.INIT('h80)
	) name2031 (
		\emc_WSCRext_reg_DO_reg[3]/NET0131 ,
		_w5670_,
		_w5790_,
		_w6079_
	);
	LUT3 #(
		.INIT('h80)
	) name2032 (
		\sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w5648_,
		_w5634_,
		_w6080_
	);
	LUT3 #(
		.INIT('h80)
	) name2033 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w5644_,
		_w5634_,
		_w6081_
	);
	LUT4 #(
		.INIT('h0001)
	) name2034 (
		_w6078_,
		_w6079_,
		_w6080_,
		_w6081_,
		_w6082_
	);
	LUT3 #(
		.INIT('h80)
	) name2035 (
		\idma_DCTL_reg[3]/NET0131 ,
		_w5628_,
		_w5639_,
		_w6083_
	);
	LUT3 #(
		.INIT('h80)
	) name2036 (
		\PIO_out[3]_pad ,
		_w5628_,
		_w5635_,
		_w6084_
	);
	LUT3 #(
		.INIT('h80)
	) name2037 (
		\PIO_oe[3]_pad ,
		_w5628_,
		_w5632_,
		_w6085_
	);
	LUT3 #(
		.INIT('h80)
	) name2038 (
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w5634_,
		_w5639_,
		_w6086_
	);
	LUT4 #(
		.INIT('h0001)
	) name2039 (
		_w6083_,
		_w6084_,
		_w6085_,
		_w6086_,
		_w6087_
	);
	LUT3 #(
		.INIT('h80)
	) name2040 (
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w5634_,
		_w5637_,
		_w6088_
	);
	LUT3 #(
		.INIT('h80)
	) name2041 (
		\clkc_ckr_reg_DO_reg[3]/NET0131 ,
		_w5631_,
		_w5644_,
		_w6089_
	);
	LUT3 #(
		.INIT('h80)
	) name2042 (
		\memc_usysr_DO_reg[3]/NET0131 ,
		_w5631_,
		_w5660_,
		_w6090_
	);
	LUT3 #(
		.INIT('h80)
	) name2043 (
		\pio_PINT_reg[3]/NET0131 ,
		_w5670_,
		_w5672_,
		_w6091_
	);
	LUT4 #(
		.INIT('h0001)
	) name2044 (
		_w6088_,
		_w6089_,
		_w6090_,
		_w6091_,
		_w6092_
	);
	LUT4 #(
		.INIT('h8000)
	) name2045 (
		_w6087_,
		_w6092_,
		_w6077_,
		_w6082_,
		_w6093_
	);
	LUT3 #(
		.INIT('h10)
	) name2046 (
		_w6072_,
		_w6071_,
		_w6093_,
		_w6094_
	);
	LUT3 #(
		.INIT('h2a)
	) name2047 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w6070_,
		_w6094_,
		_w6095_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2048 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4277_,
		_w4274_,
		_w4282_,
		_w6096_
	);
	LUT2 #(
		.INIT('h8)
	) name2049 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w6097_
	);
	LUT4 #(
		.INIT('h153f)
	) name2050 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w6098_
	);
	LUT2 #(
		.INIT('h4)
	) name2051 (
		_w6097_,
		_w6098_,
		_w6099_
	);
	LUT3 #(
		.INIT('ha8)
	) name2052 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w6100_
	);
	LUT4 #(
		.INIT('h135f)
	) name2053 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_SSTAT_reg[3]/NET0131 ,
		_w6101_
	);
	LUT4 #(
		.INIT('h135f)
	) name2054 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w6102_
	);
	LUT3 #(
		.INIT('h40)
	) name2055 (
		_w6100_,
		_w6101_,
		_w6102_,
		_w6103_
	);
	LUT2 #(
		.INIT('h8)
	) name2056 (
		_w6099_,
		_w6103_,
		_w6104_
	);
	LUT3 #(
		.INIT('h8a)
	) name2057 (
		_w5681_,
		_w6096_,
		_w6104_,
		_w6105_
	);
	LUT4 #(
		.INIT('h135f)
	) name2058 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131 ,
		_w6106_
	);
	LUT4 #(
		.INIT('h135f)
	) name2059 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131 ,
		_w6107_
	);
	LUT2 #(
		.INIT('h8)
	) name2060 (
		_w6106_,
		_w6107_,
		_w6108_
	);
	LUT4 #(
		.INIT('h135f)
	) name2061 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w6109_
	);
	LUT4 #(
		.INIT('h135f)
	) name2062 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131 ,
		_w6110_
	);
	LUT4 #(
		.INIT('h135f)
	) name2063 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131 ,
		_w6111_
	);
	LUT4 #(
		.INIT('h135f)
	) name2064 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131 ,
		_w6112_
	);
	LUT4 #(
		.INIT('h8000)
	) name2065 (
		_w6111_,
		_w6112_,
		_w6109_,
		_w6110_,
		_w6113_
	);
	LUT3 #(
		.INIT('h2a)
	) name2066 (
		_w5687_,
		_w6108_,
		_w6113_,
		_w6114_
	);
	LUT4 #(
		.INIT('h135f)
	) name2067 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131 ,
		_w6115_
	);
	LUT4 #(
		.INIT('h135f)
	) name2068 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131 ,
		_w6116_
	);
	LUT2 #(
		.INIT('h8)
	) name2069 (
		_w6115_,
		_w6116_,
		_w6117_
	);
	LUT4 #(
		.INIT('h135f)
	) name2070 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131 ,
		_w6118_
	);
	LUT4 #(
		.INIT('h135f)
	) name2071 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131 ,
		_w6119_
	);
	LUT4 #(
		.INIT('h135f)
	) name2072 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 ,
		_w6120_
	);
	LUT4 #(
		.INIT('h135f)
	) name2073 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 ,
		_w6121_
	);
	LUT4 #(
		.INIT('h8000)
	) name2074 (
		_w6120_,
		_w6121_,
		_w6118_,
		_w6119_,
		_w6122_
	);
	LUT4 #(
		.INIT('h135f)
	) name2075 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[3]/P0001 ,
		\sport1_txctl_TX_reg[3]/P0001 ,
		_w6123_
	);
	LUT4 #(
		.INIT('h135f)
	) name2076 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		\sport1_rxctl_RX_reg[3]/P0001 ,
		_w6124_
	);
	LUT3 #(
		.INIT('h2a)
	) name2077 (
		_w5706_,
		_w6123_,
		_w6124_,
		_w6125_
	);
	LUT4 #(
		.INIT('h00d5)
	) name2078 (
		_w5697_,
		_w6117_,
		_w6122_,
		_w6125_,
		_w6126_
	);
	LUT2 #(
		.INIT('h4)
	) name2079 (
		_w6114_,
		_w6126_,
		_w6127_
	);
	LUT3 #(
		.INIT('h1b)
	) name2080 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001 ,
		_w6128_
	);
	LUT4 #(
		.INIT('ha820)
	) name2081 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001 ,
		_w6129_
	);
	LUT3 #(
		.INIT('h1b)
	) name2082 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[3]/P0001 ,
		_w6130_
	);
	LUT4 #(
		.INIT('ha820)
	) name2083 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[3]/P0001 ,
		_w6131_
	);
	LUT2 #(
		.INIT('h1)
	) name2084 (
		_w6129_,
		_w6131_,
		_w6132_
	);
	LUT3 #(
		.INIT('h1b)
	) name2085 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001 ,
		_w6133_
	);
	LUT4 #(
		.INIT('ha820)
	) name2086 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001 ,
		_w6134_
	);
	LUT3 #(
		.INIT('h1b)
	) name2087 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001 ,
		_w6135_
	);
	LUT4 #(
		.INIT('ha820)
	) name2088 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001 ,
		_w6136_
	);
	LUT3 #(
		.INIT('h1b)
	) name2089 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001 ,
		_w6137_
	);
	LUT4 #(
		.INIT('ha820)
	) name2090 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001 ,
		_w6138_
	);
	LUT3 #(
		.INIT('h01)
	) name2091 (
		_w6136_,
		_w6138_,
		_w6134_,
		_w6139_
	);
	LUT3 #(
		.INIT('h2a)
	) name2092 (
		_w5741_,
		_w6132_,
		_w6139_,
		_w6140_
	);
	LUT3 #(
		.INIT('h1b)
	) name2093 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001 ,
		_w6141_
	);
	LUT4 #(
		.INIT('ha820)
	) name2094 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001 ,
		_w6142_
	);
	LUT3 #(
		.INIT('h1b)
	) name2095 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001 ,
		_w6143_
	);
	LUT4 #(
		.INIT('ha820)
	) name2096 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001 ,
		_w6144_
	);
	LUT3 #(
		.INIT('h1b)
	) name2097 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001 ,
		_w6145_
	);
	LUT4 #(
		.INIT('ha820)
	) name2098 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001 ,
		_w6146_
	);
	LUT3 #(
		.INIT('h01)
	) name2099 (
		_w6144_,
		_w6146_,
		_w6142_,
		_w6147_
	);
	LUT3 #(
		.INIT('h1b)
	) name2100 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 ,
		_w6148_
	);
	LUT4 #(
		.INIT('ha820)
	) name2101 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 ,
		_w6149_
	);
	LUT3 #(
		.INIT('h1b)
	) name2102 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001 ,
		_w6150_
	);
	LUT4 #(
		.INIT('ha820)
	) name2103 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001 ,
		_w6151_
	);
	LUT3 #(
		.INIT('h1b)
	) name2104 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001 ,
		_w6152_
	);
	LUT4 #(
		.INIT('ha820)
	) name2105 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001 ,
		_w6153_
	);
	LUT3 #(
		.INIT('h1b)
	) name2106 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001 ,
		_w6154_
	);
	LUT4 #(
		.INIT('ha820)
	) name2107 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001 ,
		_w6155_
	);
	LUT4 #(
		.INIT('h0001)
	) name2108 (
		_w6149_,
		_w6151_,
		_w6153_,
		_w6155_,
		_w6156_
	);
	LUT3 #(
		.INIT('h2a)
	) name2109 (
		_w5712_,
		_w6147_,
		_w6156_,
		_w6157_
	);
	LUT3 #(
		.INIT('h1b)
	) name2110 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001 ,
		_w6158_
	);
	LUT4 #(
		.INIT('ha820)
	) name2111 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001 ,
		_w6159_
	);
	LUT2 #(
		.INIT('h8)
	) name2112 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w6160_
	);
	LUT2 #(
		.INIT('h1)
	) name2113 (
		_w6159_,
		_w6160_,
		_w6161_
	);
	LUT4 #(
		.INIT('ha820)
	) name2114 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001 ,
		_w6162_
	);
	LUT3 #(
		.INIT('h1b)
	) name2115 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001 ,
		_w6163_
	);
	LUT4 #(
		.INIT('ha820)
	) name2116 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001 ,
		_w6164_
	);
	LUT4 #(
		.INIT('ha820)
	) name2117 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001 ,
		_w6165_
	);
	LUT4 #(
		.INIT('ha820)
	) name2118 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001 ,
		_w6166_
	);
	LUT4 #(
		.INIT('h0001)
	) name2119 (
		_w6162_,
		_w6164_,
		_w6165_,
		_w6166_,
		_w6167_
	);
	LUT3 #(
		.INIT('h2a)
	) name2120 (
		_w5730_,
		_w6161_,
		_w6167_,
		_w6168_
	);
	LUT3 #(
		.INIT('h01)
	) name2121 (
		_w6157_,
		_w6168_,
		_w6140_,
		_w6169_
	);
	LUT2 #(
		.INIT('h8)
	) name2122 (
		_w6127_,
		_w6169_,
		_w6170_
	);
	LUT2 #(
		.INIT('h4)
	) name2123 (
		_w6105_,
		_w6170_,
		_w6171_
	);
	LUT3 #(
		.INIT('h10)
	) name2124 (
		_w6055_,
		_w6095_,
		_w6171_,
		_w6172_
	);
	LUT4 #(
		.INIT('h5455)
	) name2125 (
		\emc_DMDoe_reg/NET0131 ,
		_w6055_,
		_w6095_,
		_w6171_,
		_w6173_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[3]/P0001 ,
		_w6174_
	);
	LUT3 #(
		.INIT('h08)
	) name2127 (
		_w5588_,
		_w5598_,
		_w6174_,
		_w6175_
	);
	LUT3 #(
		.INIT('h45)
	) name2128 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w6176_
	);
	LUT4 #(
		.INIT('h0200)
	) name2129 (
		\core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w6177_
	);
	LUT4 #(
		.INIT('h0200)
	) name2130 (
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w6178_
	);
	LUT4 #(
		.INIT('h0200)
	) name2131 (
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w6179_
	);
	LUT4 #(
		.INIT('h0200)
	) name2132 (
		\core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w6180_
	);
	LUT4 #(
		.INIT('h0001)
	) name2133 (
		_w6177_,
		_w6178_,
		_w6179_,
		_w6180_,
		_w6181_
	);
	LUT4 #(
		.INIT('h0200)
	) name2134 (
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w6182_
	);
	LUT4 #(
		.INIT('h0200)
	) name2135 (
		\core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w6183_
	);
	LUT4 #(
		.INIT('h0200)
	) name2136 (
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w6184_
	);
	LUT4 #(
		.INIT('h0200)
	) name2137 (
		\core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w6185_
	);
	LUT4 #(
		.INIT('h0001)
	) name2138 (
		_w6182_,
		_w6183_,
		_w6184_,
		_w6185_,
		_w6186_
	);
	LUT3 #(
		.INIT('hd0)
	) name2139 (
		_w4063_,
		_w6181_,
		_w6186_,
		_w6187_
	);
	LUT4 #(
		.INIT('h0200)
	) name2140 (
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w6188_
	);
	LUT4 #(
		.INIT('h0200)
	) name2141 (
		\core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w6189_
	);
	LUT4 #(
		.INIT('h0200)
	) name2142 (
		\core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w6190_
	);
	LUT4 #(
		.INIT('h0200)
	) name2143 (
		\core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w6191_
	);
	LUT3 #(
		.INIT('h01)
	) name2144 (
		_w6190_,
		_w6191_,
		_w6189_,
		_w6192_
	);
	LUT4 #(
		.INIT('h0200)
	) name2145 (
		\core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w6193_
	);
	LUT4 #(
		.INIT('h0200)
	) name2146 (
		\core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w6194_
	);
	LUT4 #(
		.INIT('h0200)
	) name2147 (
		\core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w6195_
	);
	LUT4 #(
		.INIT('h0200)
	) name2148 (
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w6196_
	);
	LUT4 #(
		.INIT('h0001)
	) name2149 (
		_w6193_,
		_w6194_,
		_w6195_,
		_w6196_,
		_w6197_
	);
	LUT4 #(
		.INIT('h45ef)
	) name2150 (
		_w4063_,
		_w6188_,
		_w6192_,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h2)
	) name2151 (
		_w6187_,
		_w6198_,
		_w6199_
	);
	LUT4 #(
		.INIT('hefcd)
	) name2152 (
		_w5117_,
		_w5337_,
		_w6176_,
		_w6199_,
		_w6200_
	);
	LUT3 #(
		.INIT('h8a)
	) name2153 (
		_w5586_,
		_w6041_,
		_w6200_,
		_w6201_
	);
	LUT2 #(
		.INIT('h9)
	) name2154 (
		_w5164_,
		_w5170_,
		_w6202_
	);
	LUT3 #(
		.INIT('h1e)
	) name2155 (
		_w5179_,
		_w5192_,
		_w6202_,
		_w6203_
	);
	LUT3 #(
		.INIT('he0)
	) name2156 (
		_w5767_,
		_w5918_,
		_w6203_,
		_w6204_
	);
	LUT3 #(
		.INIT('ha8)
	) name2157 (
		\core_dag_ilm1reg_I_reg[3]/NET0131 ,
		_w5158_,
		_w5159_,
		_w6205_
	);
	LUT4 #(
		.INIT('h366c)
	) name2158 (
		\core_dag_ilm1reg_M_reg[2]/NET0131 ,
		_w5163_,
		_w5168_,
		_w5296_,
		_w6206_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2159 (
		_w5767_,
		_w5918_,
		_w6205_,
		_w6206_,
		_w6207_
	);
	LUT3 #(
		.INIT('h8a)
	) name2160 (
		_w5337_,
		_w6204_,
		_w6207_,
		_w6208_
	);
	LUT2 #(
		.INIT('h2)
	) name2161 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		_w5386_,
		_w6209_
	);
	LUT3 #(
		.INIT('h14)
	) name2162 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5443_,
		_w5525_,
		_w6210_
	);
	LUT3 #(
		.INIT('he1)
	) name2163 (
		_w5428_,
		_w5431_,
		_w5499_,
		_w6211_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2164 (
		_w5467_,
		_w5488_,
		_w5498_,
		_w5511_,
		_w6212_
	);
	LUT4 #(
		.INIT('h718e)
	) name2165 (
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w5394_,
		_w5490_,
		_w5501_,
		_w6213_
	);
	LUT2 #(
		.INIT('h6)
	) name2166 (
		_w6212_,
		_w6213_,
		_w6214_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2167 (
		_w5434_,
		_w6210_,
		_w6211_,
		_w6214_,
		_w6215_
	);
	LUT4 #(
		.INIT('h888a)
	) name2168 (
		_w5117_,
		_w5337_,
		_w6209_,
		_w6215_,
		_w6216_
	);
	LUT4 #(
		.INIT('h0233)
	) name2169 (
		_w4063_,
		_w5049_,
		_w6181_,
		_w6186_,
		_w6217_
	);
	LUT4 #(
		.INIT('h0080)
	) name2170 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w6218_
	);
	LUT4 #(
		.INIT('h000b)
	) name2171 (
		_w4970_,
		_w6198_,
		_w6217_,
		_w6218_,
		_w6219_
	);
	LUT4 #(
		.INIT('ha222)
	) name2172 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w6220_
	);
	LUT4 #(
		.INIT('h2a00)
	) name2173 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w6221_
	);
	LUT4 #(
		.INIT('h4000)
	) name2174 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w6222_
	);
	LUT2 #(
		.INIT('h1)
	) name2175 (
		_w6221_,
		_w6222_,
		_w6223_
	);
	LUT3 #(
		.INIT('h20)
	) name2176 (
		_w5539_,
		_w6220_,
		_w6223_,
		_w6224_
	);
	LUT3 #(
		.INIT('hd0)
	) name2177 (
		_w5059_,
		_w6219_,
		_w6224_,
		_w6225_
	);
	LUT4 #(
		.INIT('h5540)
	) name2178 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w6226_
	);
	LUT3 #(
		.INIT('h01)
	) name2179 (
		_w5337_,
		_w6226_,
		_w6225_,
		_w6227_
	);
	LUT4 #(
		.INIT('h0200)
	) name2180 (
		\core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w6228_
	);
	LUT4 #(
		.INIT('h0200)
	) name2181 (
		\core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w6229_
	);
	LUT4 #(
		.INIT('h0200)
	) name2182 (
		\core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w6230_
	);
	LUT4 #(
		.INIT('h0200)
	) name2183 (
		\core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w6231_
	);
	LUT3 #(
		.INIT('h01)
	) name2184 (
		_w6230_,
		_w6231_,
		_w6229_,
		_w6232_
	);
	LUT4 #(
		.INIT('h0200)
	) name2185 (
		\core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w6233_
	);
	LUT4 #(
		.INIT('h0200)
	) name2186 (
		\core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w6234_
	);
	LUT4 #(
		.INIT('h0200)
	) name2187 (
		\core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w6235_
	);
	LUT4 #(
		.INIT('h0200)
	) name2188 (
		\core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w6236_
	);
	LUT4 #(
		.INIT('h0001)
	) name2189 (
		_w6233_,
		_w6234_,
		_w6235_,
		_w6236_,
		_w6237_
	);
	LUT4 #(
		.INIT('h45ef)
	) name2190 (
		_w4063_,
		_w6228_,
		_w6232_,
		_w6237_,
		_w6238_
	);
	LUT3 #(
		.INIT('h15)
	) name2191 (
		_w5117_,
		_w5337_,
		_w6238_,
		_w6239_
	);
	LUT3 #(
		.INIT('h45)
	) name2192 (
		_w5586_,
		_w6227_,
		_w6239_,
		_w6240_
	);
	LUT4 #(
		.INIT('h1055)
	) name2193 (
		_w6201_,
		_w6208_,
		_w6216_,
		_w6240_,
		_w6241_
	);
	LUT4 #(
		.INIT('hefaa)
	) name2194 (
		_w6201_,
		_w6208_,
		_w6216_,
		_w6240_,
		_w6242_
	);
	LUT4 #(
		.INIT('h5540)
	) name2195 (
		_w5255_,
		_w5302_,
		_w5303_,
		_w5305_,
		_w6243_
	);
	LUT3 #(
		.INIT('h36)
	) name2196 (
		_w5256_,
		_w5267_,
		_w6243_,
		_w6244_
	);
	LUT3 #(
		.INIT('h10)
	) name2197 (
		_w5767_,
		_w5918_,
		_w6244_,
		_w6245_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name2198 (
		\core_dag_ilm1reg_I_reg[11]/NET0131 ,
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		_w5264_,
		_w5265_,
		_w6246_
	);
	LUT2 #(
		.INIT('h9)
	) name2199 (
		_w5261_,
		_w5269_,
		_w6247_
	);
	LUT4 #(
		.INIT('h3233)
	) name2200 (
		_w5251_,
		_w5260_,
		_w5272_,
		_w5274_,
		_w6248_
	);
	LUT2 #(
		.INIT('h6)
	) name2201 (
		_w6247_,
		_w6248_,
		_w6249_
	);
	LUT4 #(
		.INIT('h010f)
	) name2202 (
		_w5767_,
		_w5918_,
		_w6246_,
		_w6249_,
		_w6250_
	);
	LUT3 #(
		.INIT('ha8)
	) name2203 (
		\DM_rd0[11]_pad ,
		_w5610_,
		_w5612_,
		_w6251_
	);
	LUT4 #(
		.INIT('h135f)
	) name2204 (
		\DM_rdm[11]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w6252_
	);
	LUT4 #(
		.INIT('h135f)
	) name2205 (
		\DM_rd6[11]_pad ,
		\DM_rd7[11]_pad ,
		_w5596_,
		_w5591_,
		_w6253_
	);
	LUT2 #(
		.INIT('h8)
	) name2206 (
		_w6252_,
		_w6253_,
		_w6254_
	);
	LUT3 #(
		.INIT('h80)
	) name2207 (
		\DM_rd5[11]_pad ,
		_w5598_,
		_w5599_,
		_w6255_
	);
	LUT3 #(
		.INIT('h80)
	) name2208 (
		\DM_rd4[11]_pad ,
		_w5598_,
		_w5601_,
		_w6256_
	);
	LUT4 #(
		.INIT('h8000)
	) name2209 (
		\DM_rd2[11]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w6257_
	);
	LUT4 #(
		.INIT('h8000)
	) name2210 (
		\DM_rd1[11]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w6258_
	);
	LUT4 #(
		.INIT('h8000)
	) name2211 (
		\DM_rd3[11]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w6259_
	);
	LUT3 #(
		.INIT('h01)
	) name2212 (
		_w6258_,
		_w6259_,
		_w6257_,
		_w6260_
	);
	LUT3 #(
		.INIT('h10)
	) name2213 (
		_w6256_,
		_w6255_,
		_w6260_,
		_w6261_
	);
	LUT2 #(
		.INIT('h8)
	) name2214 (
		_w6254_,
		_w6261_,
		_w6262_
	);
	LUT2 #(
		.INIT('h4)
	) name2215 (
		_w6251_,
		_w6262_,
		_w6263_
	);
	LUT4 #(
		.INIT('h4000)
	) name2216 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[11]/P0001 ,
		_w6264_
	);
	LUT3 #(
		.INIT('h80)
	) name2217 (
		\bdma_BCTL_reg[11]/NET0131 ,
		_w5627_,
		_w5629_,
		_w6265_
	);
	LUT3 #(
		.INIT('h80)
	) name2218 (
		\tm_tpr_reg_DO_reg[11]/NET0131 ,
		_w5631_,
		_w5635_,
		_w6266_
	);
	LUT3 #(
		.INIT('h80)
	) name2219 (
		\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w5648_,
		_w5634_,
		_w6267_
	);
	LUT3 #(
		.INIT('h80)
	) name2220 (
		\idma_DCTL_reg[11]/NET0131 ,
		_w5628_,
		_w5639_,
		_w6268_
	);
	LUT4 #(
		.INIT('h0001)
	) name2221 (
		_w5795_,
		_w6266_,
		_w6267_,
		_w6268_,
		_w6269_
	);
	LUT4 #(
		.INIT('h8000)
	) name2222 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_txctl_Wcnt_reg[3]/NET0131 ,
		_w5631_,
		_w5639_,
		_w6270_
	);
	LUT4 #(
		.INIT('h8000)
	) name2223 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_txctl_Wcnt_reg[3]/NET0131 ,
		_w5634_,
		_w5660_,
		_w6271_
	);
	LUT2 #(
		.INIT('h1)
	) name2224 (
		_w6270_,
		_w6271_,
		_w6272_
	);
	LUT3 #(
		.INIT('h40)
	) name2225 (
		_w6265_,
		_w6269_,
		_w6272_,
		_w6273_
	);
	LUT3 #(
		.INIT('h80)
	) name2226 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w5629_,
		_w5648_,
		_w6274_
	);
	LUT3 #(
		.INIT('h80)
	) name2227 (
		\bdma_BEAD_reg[11]/NET0131 ,
		_w5629_,
		_w5644_,
		_w6275_
	);
	LUT2 #(
		.INIT('h1)
	) name2228 (
		_w6274_,
		_w6275_,
		_w6276_
	);
	LUT4 #(
		.INIT('h8000)
	) name2229 (
		\bdma_BWCOUNT_reg[11]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w6277_
	);
	LUT4 #(
		.INIT('h8000)
	) name2230 (
		\bdma_BOVL_reg[11]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w6278_
	);
	LUT3 #(
		.INIT('h80)
	) name2231 (
		\sport1_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w5670_,
		_w5810_,
		_w6279_
	);
	LUT3 #(
		.INIT('h80)
	) name2232 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w5631_,
		_w5660_,
		_w6280_
	);
	LUT3 #(
		.INIT('h80)
	) name2233 (
		\clkc_ckr_reg_DO_reg[11]/NET0131 ,
		_w5631_,
		_w5644_,
		_w6281_
	);
	LUT3 #(
		.INIT('h80)
	) name2234 (
		\sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w5634_,
		_w5635_,
		_w6282_
	);
	LUT4 #(
		.INIT('h0001)
	) name2235 (
		_w6279_,
		_w6280_,
		_w6281_,
		_w6282_,
		_w6283_
	);
	LUT3 #(
		.INIT('h80)
	) name2236 (
		\sport0_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w5627_,
		_w5634_,
		_w6284_
	);
	LUT3 #(
		.INIT('h80)
	) name2237 (
		\emc_WSCRreg_DO_reg[11]/NET0131 ,
		_w5631_,
		_w5632_,
		_w6285_
	);
	LUT3 #(
		.INIT('h80)
	) name2238 (
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w5634_,
		_w5639_,
		_w6286_
	);
	LUT3 #(
		.INIT('h80)
	) name2239 (
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w5644_,
		_w5634_,
		_w6287_
	);
	LUT4 #(
		.INIT('h0001)
	) name2240 (
		_w6284_,
		_w6285_,
		_w6286_,
		_w6287_,
		_w6288_
	);
	LUT3 #(
		.INIT('h80)
	) name2241 (
		\idma_DOVL_reg[11]/NET0131 ,
		_w5804_,
		_w5824_,
		_w6289_
	);
	LUT3 #(
		.INIT('h80)
	) name2242 (
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w5634_,
		_w5637_,
		_w6290_
	);
	LUT3 #(
		.INIT('h80)
	) name2243 (
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w5632_,
		_w5634_,
		_w6291_
	);
	LUT3 #(
		.INIT('h80)
	) name2244 (
		\tm_TCR_TMP_reg[11]/NET0131 ,
		_w5631_,
		_w5637_,
		_w6292_
	);
	LUT4 #(
		.INIT('h0001)
	) name2245 (
		_w6289_,
		_w6290_,
		_w6291_,
		_w6292_,
		_w6293_
	);
	LUT4 #(
		.INIT('h4000)
	) name2246 (
		_w6278_,
		_w6283_,
		_w6288_,
		_w6293_,
		_w6294_
	);
	LUT4 #(
		.INIT('h4000)
	) name2247 (
		_w6277_,
		_w6273_,
		_w6276_,
		_w6294_,
		_w6295_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2248 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4309_,
		_w4306_,
		_w4314_,
		_w6296_
	);
	LUT3 #(
		.INIT('ha8)
	) name2249 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w6297_
	);
	LUT4 #(
		.INIT('h135f)
	) name2250 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w6298_
	);
	LUT2 #(
		.INIT('h4)
	) name2251 (
		_w6297_,
		_w6298_,
		_w6299_
	);
	LUT3 #(
		.INIT('h8a)
	) name2252 (
		_w5681_,
		_w6296_,
		_w6299_,
		_w6300_
	);
	LUT4 #(
		.INIT('h135f)
	) name2253 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131 ,
		_w6301_
	);
	LUT4 #(
		.INIT('h135f)
	) name2254 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131 ,
		_w6302_
	);
	LUT2 #(
		.INIT('h8)
	) name2255 (
		_w6301_,
		_w6302_,
		_w6303_
	);
	LUT4 #(
		.INIT('h135f)
	) name2256 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131 ,
		_w6304_
	);
	LUT4 #(
		.INIT('h135f)
	) name2257 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131 ,
		_w6305_
	);
	LUT4 #(
		.INIT('h135f)
	) name2258 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131 ,
		_w6306_
	);
	LUT4 #(
		.INIT('h135f)
	) name2259 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131 ,
		_w6307_
	);
	LUT4 #(
		.INIT('h8000)
	) name2260 (
		_w6306_,
		_w6307_,
		_w6304_,
		_w6305_,
		_w6308_
	);
	LUT3 #(
		.INIT('h2a)
	) name2261 (
		_w5697_,
		_w6303_,
		_w6308_,
		_w6309_
	);
	LUT4 #(
		.INIT('h135f)
	) name2262 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131 ,
		_w6310_
	);
	LUT4 #(
		.INIT('h135f)
	) name2263 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131 ,
		_w6311_
	);
	LUT2 #(
		.INIT('h8)
	) name2264 (
		_w6310_,
		_w6311_,
		_w6312_
	);
	LUT4 #(
		.INIT('h135f)
	) name2265 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131 ,
		_w6313_
	);
	LUT4 #(
		.INIT('h135f)
	) name2266 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131 ,
		_w6314_
	);
	LUT4 #(
		.INIT('h135f)
	) name2267 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131 ,
		_w6315_
	);
	LUT4 #(
		.INIT('h135f)
	) name2268 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131 ,
		_w6316_
	);
	LUT4 #(
		.INIT('h8000)
	) name2269 (
		_w6315_,
		_w6316_,
		_w6313_,
		_w6314_,
		_w6317_
	);
	LUT4 #(
		.INIT('h135f)
	) name2270 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[11]/P0001 ,
		\sport1_txctl_TX_reg[11]/P0001 ,
		_w6318_
	);
	LUT4 #(
		.INIT('h135f)
	) name2271 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[11]/P0001 ,
		\sport1_rxctl_RX_reg[11]/P0001 ,
		_w6319_
	);
	LUT3 #(
		.INIT('h2a)
	) name2272 (
		_w5706_,
		_w6318_,
		_w6319_,
		_w6320_
	);
	LUT4 #(
		.INIT('h00d5)
	) name2273 (
		_w5687_,
		_w6312_,
		_w6317_,
		_w6320_,
		_w6321_
	);
	LUT2 #(
		.INIT('h4)
	) name2274 (
		_w6309_,
		_w6321_,
		_w6322_
	);
	LUT3 #(
		.INIT('h1b)
	) name2275 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001 ,
		_w6323_
	);
	LUT4 #(
		.INIT('ha820)
	) name2276 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001 ,
		_w6324_
	);
	LUT3 #(
		.INIT('h1b)
	) name2277 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001 ,
		_w6325_
	);
	LUT4 #(
		.INIT('ha820)
	) name2278 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001 ,
		_w6326_
	);
	LUT3 #(
		.INIT('h1b)
	) name2279 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001 ,
		_w6327_
	);
	LUT4 #(
		.INIT('ha820)
	) name2280 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001 ,
		_w6328_
	);
	LUT3 #(
		.INIT('h01)
	) name2281 (
		_w6326_,
		_w6328_,
		_w6324_,
		_w6329_
	);
	LUT3 #(
		.INIT('h2a)
	) name2282 (
		_w5741_,
		_w5746_,
		_w6329_,
		_w6330_
	);
	LUT3 #(
		.INIT('h1b)
	) name2283 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 ,
		_w6331_
	);
	LUT4 #(
		.INIT('ha820)
	) name2284 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 ,
		_w6332_
	);
	LUT3 #(
		.INIT('h1b)
	) name2285 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001 ,
		_w6333_
	);
	LUT4 #(
		.INIT('ha820)
	) name2286 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001 ,
		_w6334_
	);
	LUT3 #(
		.INIT('h1b)
	) name2287 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001 ,
		_w6335_
	);
	LUT4 #(
		.INIT('ha820)
	) name2288 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001 ,
		_w6336_
	);
	LUT3 #(
		.INIT('h01)
	) name2289 (
		_w6334_,
		_w6336_,
		_w6332_,
		_w6337_
	);
	LUT3 #(
		.INIT('h1b)
	) name2290 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001 ,
		_w6338_
	);
	LUT4 #(
		.INIT('ha820)
	) name2291 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001 ,
		_w6339_
	);
	LUT3 #(
		.INIT('h1b)
	) name2292 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001 ,
		_w6340_
	);
	LUT4 #(
		.INIT('ha820)
	) name2293 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001 ,
		_w6341_
	);
	LUT3 #(
		.INIT('h1b)
	) name2294 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001 ,
		_w6342_
	);
	LUT4 #(
		.INIT('ha820)
	) name2295 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001 ,
		_w6343_
	);
	LUT4 #(
		.INIT('h0001)
	) name2296 (
		_w5714_,
		_w6339_,
		_w6341_,
		_w6343_,
		_w6344_
	);
	LUT3 #(
		.INIT('h2a)
	) name2297 (
		_w5712_,
		_w6337_,
		_w6344_,
		_w6345_
	);
	LUT4 #(
		.INIT('ha820)
	) name2298 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001 ,
		_w6346_
	);
	LUT4 #(
		.INIT('ha820)
	) name2299 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001 ,
		_w6347_
	);
	LUT2 #(
		.INIT('h1)
	) name2300 (
		_w6346_,
		_w6347_,
		_w6348_
	);
	LUT3 #(
		.INIT('h1b)
	) name2301 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001 ,
		_w6349_
	);
	LUT4 #(
		.INIT('ha820)
	) name2302 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001 ,
		_w6350_
	);
	LUT3 #(
		.INIT('h1b)
	) name2303 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001 ,
		_w6351_
	);
	LUT4 #(
		.INIT('ha820)
	) name2304 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001 ,
		_w6352_
	);
	LUT3 #(
		.INIT('h1b)
	) name2305 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001 ,
		_w6353_
	);
	LUT4 #(
		.INIT('ha820)
	) name2306 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001 ,
		_w6354_
	);
	LUT3 #(
		.INIT('h01)
	) name2307 (
		_w6352_,
		_w6354_,
		_w6350_,
		_w6355_
	);
	LUT3 #(
		.INIT('h2a)
	) name2308 (
		_w5730_,
		_w6348_,
		_w6355_,
		_w6356_
	);
	LUT3 #(
		.INIT('h01)
	) name2309 (
		_w6345_,
		_w6356_,
		_w6330_,
		_w6357_
	);
	LUT2 #(
		.INIT('h8)
	) name2310 (
		_w6322_,
		_w6357_,
		_w6358_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2311 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w6295_,
		_w6300_,
		_w6358_,
		_w6359_
	);
	LUT2 #(
		.INIT('h8)
	) name2312 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[11]/P0001 ,
		_w6360_
	);
	LUT3 #(
		.INIT('h08)
	) name2313 (
		_w5588_,
		_w5598_,
		_w6360_,
		_w6361_
	);
	LUT4 #(
		.INIT('hba00)
	) name2314 (
		\emc_DMDoe_reg/NET0131 ,
		_w6264_,
		_w6359_,
		_w6361_,
		_w6362_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w6263_,
		_w6362_,
		_w6363_
	);
	LUT3 #(
		.INIT('hc4)
	) name2316 (
		_w5117_,
		_w5337_,
		_w6363_,
		_w6364_
	);
	LUT4 #(
		.INIT('hef00)
	) name2317 (
		_w5117_,
		_w6245_,
		_w6250_,
		_w6364_,
		_w6365_
	);
	LUT3 #(
		.INIT('ha8)
	) name2318 (
		\DM_rd0[2]_pad ,
		_w5610_,
		_w5612_,
		_w6366_
	);
	LUT4 #(
		.INIT('h135f)
	) name2319 (
		\DM_rdm[2]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w6367_
	);
	LUT4 #(
		.INIT('h135f)
	) name2320 (
		\DM_rd6[2]_pad ,
		\DM_rd7[2]_pad ,
		_w5596_,
		_w5591_,
		_w6368_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		_w6367_,
		_w6368_,
		_w6369_
	);
	LUT3 #(
		.INIT('h80)
	) name2322 (
		\DM_rd4[2]_pad ,
		_w5598_,
		_w5601_,
		_w6370_
	);
	LUT3 #(
		.INIT('h80)
	) name2323 (
		\DM_rd5[2]_pad ,
		_w5598_,
		_w5599_,
		_w6371_
	);
	LUT4 #(
		.INIT('h8000)
	) name2324 (
		\DM_rd2[2]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w6372_
	);
	LUT4 #(
		.INIT('h8000)
	) name2325 (
		\DM_rd1[2]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w6373_
	);
	LUT4 #(
		.INIT('h8000)
	) name2326 (
		\DM_rd3[2]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w6374_
	);
	LUT3 #(
		.INIT('h01)
	) name2327 (
		_w6373_,
		_w6374_,
		_w6372_,
		_w6375_
	);
	LUT3 #(
		.INIT('h10)
	) name2328 (
		_w6371_,
		_w6370_,
		_w6375_,
		_w6376_
	);
	LUT2 #(
		.INIT('h8)
	) name2329 (
		_w6369_,
		_w6376_,
		_w6377_
	);
	LUT2 #(
		.INIT('h4)
	) name2330 (
		_w6366_,
		_w6377_,
		_w6378_
	);
	LUT4 #(
		.INIT('h4000)
	) name2331 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[2]/P0001 ,
		_w6379_
	);
	LUT3 #(
		.INIT('h80)
	) name2332 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w5629_,
		_w5648_,
		_w6380_
	);
	LUT3 #(
		.INIT('h80)
	) name2333 (
		\emc_WSCRreg_DO_reg[2]/NET0131 ,
		_w5631_,
		_w5632_,
		_w6381_
	);
	LUT3 #(
		.INIT('h80)
	) name2334 (
		\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w5634_,
		_w5635_,
		_w6382_
	);
	LUT3 #(
		.INIT('h80)
	) name2335 (
		\sport1_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w5631_,
		_w5639_,
		_w6383_
	);
	LUT3 #(
		.INIT('h80)
	) name2336 (
		\tm_tsr_reg_DO_reg[2]/NET0131 ,
		_w5627_,
		_w5631_,
		_w6384_
	);
	LUT4 #(
		.INIT('h0001)
	) name2337 (
		_w6381_,
		_w6382_,
		_w6383_,
		_w6384_,
		_w6385_
	);
	LUT3 #(
		.INIT('h80)
	) name2338 (
		\idma_DOVL_reg[2]/NET0131 ,
		_w5804_,
		_w5824_,
		_w6386_
	);
	LUT3 #(
		.INIT('h80)
	) name2339 (
		\sport0_regs_AUTOreg_DO_reg[2]/NET0131 ,
		_w5627_,
		_w5634_,
		_w6387_
	);
	LUT3 #(
		.INIT('h80)
	) name2340 (
		\tm_tpr_reg_DO_reg[2]/NET0131 ,
		_w5631_,
		_w5635_,
		_w6388_
	);
	LUT4 #(
		.INIT('h0001)
	) name2341 (
		_w5795_,
		_w6386_,
		_w6387_,
		_w6388_,
		_w6389_
	);
	LUT3 #(
		.INIT('h40)
	) name2342 (
		_w6380_,
		_w6385_,
		_w6389_,
		_w6390_
	);
	LUT3 #(
		.INIT('h80)
	) name2343 (
		\bdma_BEAD_reg[2]/NET0131 ,
		_w5629_,
		_w5644_,
		_w6391_
	);
	LUT3 #(
		.INIT('h80)
	) name2344 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w5627_,
		_w5629_,
		_w6392_
	);
	LUT2 #(
		.INIT('h1)
	) name2345 (
		_w6391_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h8)
	) name2346 (
		_w6390_,
		_w6393_,
		_w6394_
	);
	LUT4 #(
		.INIT('h8000)
	) name2347 (
		\bdma_BOVL_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w6395_
	);
	LUT4 #(
		.INIT('h8000)
	) name2348 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w6396_
	);
	LUT3 #(
		.INIT('h80)
	) name2349 (
		\pio_pmask_reg_DO_reg[2]/NET0131 ,
		_w5628_,
		_w5660_,
		_w6397_
	);
	LUT3 #(
		.INIT('h80)
	) name2350 (
		\sport0_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w5634_,
		_w5660_,
		_w6398_
	);
	LUT3 #(
		.INIT('h80)
	) name2351 (
		\sport1_regs_AUTOreg_DO_reg[2]/NET0131 ,
		_w5670_,
		_w5810_,
		_w6399_
	);
	LUT3 #(
		.INIT('h80)
	) name2352 (
		\tm_TCR_TMP_reg[2]/NET0131 ,
		_w5631_,
		_w5637_,
		_w6400_
	);
	LUT4 #(
		.INIT('h0001)
	) name2353 (
		_w6397_,
		_w6398_,
		_w6399_,
		_w6400_,
		_w6401_
	);
	LUT3 #(
		.INIT('h80)
	) name2354 (
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w5632_,
		_w5634_,
		_w6402_
	);
	LUT3 #(
		.INIT('h80)
	) name2355 (
		\emc_WSCRext_reg_DO_reg[2]/NET0131 ,
		_w5670_,
		_w5790_,
		_w6403_
	);
	LUT3 #(
		.INIT('h80)
	) name2356 (
		\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w5648_,
		_w5634_,
		_w6404_
	);
	LUT3 #(
		.INIT('h80)
	) name2357 (
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w5644_,
		_w5634_,
		_w6405_
	);
	LUT4 #(
		.INIT('h0001)
	) name2358 (
		_w6402_,
		_w6403_,
		_w6404_,
		_w6405_,
		_w6406_
	);
	LUT3 #(
		.INIT('h80)
	) name2359 (
		\idma_DCTL_reg[2]/NET0131 ,
		_w5628_,
		_w5639_,
		_w6407_
	);
	LUT3 #(
		.INIT('h80)
	) name2360 (
		\PIO_out[2]_pad ,
		_w5628_,
		_w5635_,
		_w6408_
	);
	LUT3 #(
		.INIT('h80)
	) name2361 (
		\PIO_oe[2]_pad ,
		_w5628_,
		_w5632_,
		_w6409_
	);
	LUT3 #(
		.INIT('h80)
	) name2362 (
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w5634_,
		_w5639_,
		_w6410_
	);
	LUT4 #(
		.INIT('h0001)
	) name2363 (
		_w6407_,
		_w6408_,
		_w6409_,
		_w6410_,
		_w6411_
	);
	LUT3 #(
		.INIT('h80)
	) name2364 (
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w5634_,
		_w5637_,
		_w6412_
	);
	LUT3 #(
		.INIT('h80)
	) name2365 (
		\clkc_ckr_reg_DO_reg[2]/NET0131 ,
		_w5631_,
		_w5644_,
		_w6413_
	);
	LUT3 #(
		.INIT('h80)
	) name2366 (
		\memc_usysr_DO_reg[2]/NET0131 ,
		_w5631_,
		_w5660_,
		_w6414_
	);
	LUT3 #(
		.INIT('h80)
	) name2367 (
		\pio_PINT_reg[2]/NET0131 ,
		_w5670_,
		_w5672_,
		_w6415_
	);
	LUT4 #(
		.INIT('h0001)
	) name2368 (
		_w6412_,
		_w6413_,
		_w6414_,
		_w6415_,
		_w6416_
	);
	LUT4 #(
		.INIT('h8000)
	) name2369 (
		_w6411_,
		_w6416_,
		_w6401_,
		_w6406_,
		_w6417_
	);
	LUT3 #(
		.INIT('h10)
	) name2370 (
		_w6396_,
		_w6395_,
		_w6417_,
		_w6418_
	);
	LUT3 #(
		.INIT('h2a)
	) name2371 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w6394_,
		_w6418_,
		_w6419_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2372 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4339_,
		_w4336_,
		_w4344_,
		_w6420_
	);
	LUT4 #(
		.INIT('h135f)
	) name2373 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_SSTAT_reg[2]/NET0131 ,
		_w6421_
	);
	LUT4 #(
		.INIT('h135f)
	) name2374 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		_w6422_
	);
	LUT2 #(
		.INIT('h8)
	) name2375 (
		_w6421_,
		_w6422_,
		_w6423_
	);
	LUT3 #(
		.INIT('ha8)
	) name2376 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w6424_
	);
	LUT4 #(
		.INIT('h153f)
	) name2377 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w6425_
	);
	LUT4 #(
		.INIT('h135f)
	) name2378 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w6426_
	);
	LUT3 #(
		.INIT('h40)
	) name2379 (
		_w6424_,
		_w6425_,
		_w6426_,
		_w6427_
	);
	LUT2 #(
		.INIT('h8)
	) name2380 (
		_w6423_,
		_w6427_,
		_w6428_
	);
	LUT3 #(
		.INIT('h8a)
	) name2381 (
		_w5681_,
		_w6420_,
		_w6428_,
		_w6429_
	);
	LUT4 #(
		.INIT('h135f)
	) name2382 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w6430_
	);
	LUT4 #(
		.INIT('h135f)
	) name2383 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w6431_
	);
	LUT2 #(
		.INIT('h8)
	) name2384 (
		_w6430_,
		_w6431_,
		_w6432_
	);
	LUT4 #(
		.INIT('h135f)
	) name2385 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131 ,
		_w6433_
	);
	LUT4 #(
		.INIT('h135f)
	) name2386 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131 ,
		_w6434_
	);
	LUT4 #(
		.INIT('h135f)
	) name2387 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131 ,
		_w6435_
	);
	LUT4 #(
		.INIT('h135f)
	) name2388 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131 ,
		_w6436_
	);
	LUT4 #(
		.INIT('h8000)
	) name2389 (
		_w6435_,
		_w6436_,
		_w6433_,
		_w6434_,
		_w6437_
	);
	LUT3 #(
		.INIT('h2a)
	) name2390 (
		_w5687_,
		_w6432_,
		_w6437_,
		_w6438_
	);
	LUT4 #(
		.INIT('h135f)
	) name2391 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131 ,
		_w6439_
	);
	LUT4 #(
		.INIT('h135f)
	) name2392 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131 ,
		_w6440_
	);
	LUT2 #(
		.INIT('h8)
	) name2393 (
		_w6439_,
		_w6440_,
		_w6441_
	);
	LUT4 #(
		.INIT('h135f)
	) name2394 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131 ,
		_w6442_
	);
	LUT4 #(
		.INIT('h135f)
	) name2395 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 ,
		_w6443_
	);
	LUT4 #(
		.INIT('h135f)
	) name2396 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 ,
		_w6444_
	);
	LUT4 #(
		.INIT('h135f)
	) name2397 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131 ,
		_w6445_
	);
	LUT4 #(
		.INIT('h8000)
	) name2398 (
		_w6444_,
		_w6445_,
		_w6442_,
		_w6443_,
		_w6446_
	);
	LUT4 #(
		.INIT('h135f)
	) name2399 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[2]/P0001 ,
		\sport1_txctl_TX_reg[2]/P0001 ,
		_w6447_
	);
	LUT4 #(
		.INIT('h135f)
	) name2400 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport1_rxctl_RX_reg[2]/P0001 ,
		_w6448_
	);
	LUT3 #(
		.INIT('h2a)
	) name2401 (
		_w5706_,
		_w6447_,
		_w6448_,
		_w6449_
	);
	LUT4 #(
		.INIT('h00d5)
	) name2402 (
		_w5697_,
		_w6441_,
		_w6446_,
		_w6449_,
		_w6450_
	);
	LUT2 #(
		.INIT('h4)
	) name2403 (
		_w6438_,
		_w6450_,
		_w6451_
	);
	LUT3 #(
		.INIT('h1b)
	) name2404 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001 ,
		_w6452_
	);
	LUT4 #(
		.INIT('ha820)
	) name2405 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001 ,
		_w6453_
	);
	LUT2 #(
		.INIT('h8)
	) name2406 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w6454_
	);
	LUT2 #(
		.INIT('h1)
	) name2407 (
		_w6453_,
		_w6454_,
		_w6455_
	);
	LUT3 #(
		.INIT('h1b)
	) name2408 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001 ,
		_w6456_
	);
	LUT4 #(
		.INIT('ha820)
	) name2409 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001 ,
		_w6457_
	);
	LUT3 #(
		.INIT('h1b)
	) name2410 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001 ,
		_w6458_
	);
	LUT4 #(
		.INIT('ha820)
	) name2411 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001 ,
		_w6459_
	);
	LUT4 #(
		.INIT('ha820)
	) name2412 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001 ,
		_w6460_
	);
	LUT4 #(
		.INIT('ha820)
	) name2413 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001 ,
		_w6461_
	);
	LUT4 #(
		.INIT('h0001)
	) name2414 (
		_w6457_,
		_w6459_,
		_w6460_,
		_w6461_,
		_w6462_
	);
	LUT3 #(
		.INIT('h2a)
	) name2415 (
		_w5730_,
		_w6455_,
		_w6462_,
		_w6463_
	);
	LUT3 #(
		.INIT('h1b)
	) name2416 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001 ,
		_w6464_
	);
	LUT4 #(
		.INIT('ha820)
	) name2417 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001 ,
		_w6465_
	);
	LUT3 #(
		.INIT('h1b)
	) name2418 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[2]/P0001 ,
		_w6466_
	);
	LUT4 #(
		.INIT('ha820)
	) name2419 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[2]/P0001 ,
		_w6467_
	);
	LUT2 #(
		.INIT('h1)
	) name2420 (
		_w6465_,
		_w6467_,
		_w6468_
	);
	LUT3 #(
		.INIT('h1b)
	) name2421 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001 ,
		_w6469_
	);
	LUT4 #(
		.INIT('ha820)
	) name2422 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001 ,
		_w6470_
	);
	LUT3 #(
		.INIT('h1b)
	) name2423 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001 ,
		_w6471_
	);
	LUT4 #(
		.INIT('ha820)
	) name2424 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001 ,
		_w6472_
	);
	LUT3 #(
		.INIT('h1b)
	) name2425 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001 ,
		_w6473_
	);
	LUT4 #(
		.INIT('ha820)
	) name2426 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001 ,
		_w6474_
	);
	LUT3 #(
		.INIT('h01)
	) name2427 (
		_w6472_,
		_w6474_,
		_w6470_,
		_w6475_
	);
	LUT3 #(
		.INIT('h2a)
	) name2428 (
		_w5741_,
		_w6468_,
		_w6475_,
		_w6476_
	);
	LUT3 #(
		.INIT('h1b)
	) name2429 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 ,
		_w6477_
	);
	LUT4 #(
		.INIT('ha820)
	) name2430 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 ,
		_w6478_
	);
	LUT3 #(
		.INIT('h1b)
	) name2431 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001 ,
		_w6479_
	);
	LUT4 #(
		.INIT('ha820)
	) name2432 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001 ,
		_w6480_
	);
	LUT3 #(
		.INIT('h1b)
	) name2433 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001 ,
		_w6481_
	);
	LUT4 #(
		.INIT('ha820)
	) name2434 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001 ,
		_w6482_
	);
	LUT3 #(
		.INIT('h01)
	) name2435 (
		_w6480_,
		_w6482_,
		_w6478_,
		_w6483_
	);
	LUT3 #(
		.INIT('h1b)
	) name2436 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001 ,
		_w6484_
	);
	LUT4 #(
		.INIT('ha820)
	) name2437 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001 ,
		_w6485_
	);
	LUT3 #(
		.INIT('h1b)
	) name2438 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001 ,
		_w6486_
	);
	LUT4 #(
		.INIT('ha820)
	) name2439 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001 ,
		_w6487_
	);
	LUT3 #(
		.INIT('h1b)
	) name2440 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001 ,
		_w6488_
	);
	LUT4 #(
		.INIT('ha820)
	) name2441 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001 ,
		_w6489_
	);
	LUT3 #(
		.INIT('h1b)
	) name2442 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001 ,
		_w6490_
	);
	LUT4 #(
		.INIT('ha820)
	) name2443 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001 ,
		_w6491_
	);
	LUT4 #(
		.INIT('h0001)
	) name2444 (
		_w6485_,
		_w6487_,
		_w6489_,
		_w6491_,
		_w6492_
	);
	LUT3 #(
		.INIT('h2a)
	) name2445 (
		_w5712_,
		_w6483_,
		_w6492_,
		_w6493_
	);
	LUT3 #(
		.INIT('h01)
	) name2446 (
		_w6476_,
		_w6493_,
		_w6463_,
		_w6494_
	);
	LUT2 #(
		.INIT('h8)
	) name2447 (
		_w6451_,
		_w6494_,
		_w6495_
	);
	LUT2 #(
		.INIT('h4)
	) name2448 (
		_w6429_,
		_w6495_,
		_w6496_
	);
	LUT3 #(
		.INIT('h10)
	) name2449 (
		_w6379_,
		_w6419_,
		_w6496_,
		_w6497_
	);
	LUT4 #(
		.INIT('h5455)
	) name2450 (
		\emc_DMDoe_reg/NET0131 ,
		_w6379_,
		_w6419_,
		_w6496_,
		_w6498_
	);
	LUT2 #(
		.INIT('h8)
	) name2451 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[2]/P0001 ,
		_w6499_
	);
	LUT3 #(
		.INIT('h08)
	) name2452 (
		_w5588_,
		_w5598_,
		_w6499_,
		_w6500_
	);
	LUT3 #(
		.INIT('h45)
	) name2453 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w6501_
	);
	LUT4 #(
		.INIT('h0200)
	) name2454 (
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w6502_
	);
	LUT4 #(
		.INIT('h0200)
	) name2455 (
		\core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w6503_
	);
	LUT4 #(
		.INIT('h0200)
	) name2456 (
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w6504_
	);
	LUT4 #(
		.INIT('h0200)
	) name2457 (
		\core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w6505_
	);
	LUT4 #(
		.INIT('h0001)
	) name2458 (
		_w6502_,
		_w6503_,
		_w6504_,
		_w6505_,
		_w6506_
	);
	LUT4 #(
		.INIT('h0200)
	) name2459 (
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w6507_
	);
	LUT4 #(
		.INIT('h0200)
	) name2460 (
		\core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w6508_
	);
	LUT4 #(
		.INIT('h0200)
	) name2461 (
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w6509_
	);
	LUT4 #(
		.INIT('h0200)
	) name2462 (
		\core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w6510_
	);
	LUT4 #(
		.INIT('h0001)
	) name2463 (
		_w6507_,
		_w6508_,
		_w6509_,
		_w6510_,
		_w6511_
	);
	LUT3 #(
		.INIT('hd0)
	) name2464 (
		_w4063_,
		_w6506_,
		_w6511_,
		_w6512_
	);
	LUT4 #(
		.INIT('h0200)
	) name2465 (
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w6513_
	);
	LUT4 #(
		.INIT('h0200)
	) name2466 (
		\core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w6514_
	);
	LUT4 #(
		.INIT('h0200)
	) name2467 (
		\core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w6515_
	);
	LUT4 #(
		.INIT('h0200)
	) name2468 (
		\core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w6516_
	);
	LUT3 #(
		.INIT('h01)
	) name2469 (
		_w6515_,
		_w6516_,
		_w6514_,
		_w6517_
	);
	LUT4 #(
		.INIT('h0200)
	) name2470 (
		\core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w6518_
	);
	LUT4 #(
		.INIT('h0200)
	) name2471 (
		\core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w6519_
	);
	LUT4 #(
		.INIT('h0200)
	) name2472 (
		\core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w6520_
	);
	LUT4 #(
		.INIT('h0200)
	) name2473 (
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w6521_
	);
	LUT4 #(
		.INIT('h0001)
	) name2474 (
		_w6518_,
		_w6519_,
		_w6520_,
		_w6521_,
		_w6522_
	);
	LUT4 #(
		.INIT('h45ef)
	) name2475 (
		_w4063_,
		_w6513_,
		_w6517_,
		_w6522_,
		_w6523_
	);
	LUT2 #(
		.INIT('h2)
	) name2476 (
		_w6512_,
		_w6523_,
		_w6524_
	);
	LUT4 #(
		.INIT('hefcd)
	) name2477 (
		_w5117_,
		_w5337_,
		_w6501_,
		_w6524_,
		_w6525_
	);
	LUT3 #(
		.INIT('h8a)
	) name2478 (
		_w5586_,
		_w6365_,
		_w6525_,
		_w6526_
	);
	LUT2 #(
		.INIT('h9)
	) name2479 (
		_w5503_,
		_w5506_,
		_w6527_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2480 (
		_w5502_,
		_w5512_,
		_w6212_,
		_w6527_,
		_w6528_
	);
	LUT3 #(
		.INIT('h10)
	) name2481 (
		_w5434_,
		_w6210_,
		_w6528_,
		_w6529_
	);
	LUT4 #(
		.INIT('h08a8)
	) name2482 (
		\core_dag_ilm2reg_I_reg[11]/NET0131 ,
		_w5353_,
		_w5370_,
		_w5381_,
		_w6530_
	);
	LUT4 #(
		.INIT('heee8)
	) name2483 (
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w5387_,
		_w5428_,
		_w5431_,
		_w6531_
	);
	LUT2 #(
		.INIT('h6)
	) name2484 (
		_w5504_,
		_w6531_,
		_w6532_
	);
	LUT4 #(
		.INIT('h010f)
	) name2485 (
		_w5434_,
		_w6210_,
		_w6530_,
		_w6532_,
		_w6533_
	);
	LUT4 #(
		.INIT('h0233)
	) name2486 (
		_w4063_,
		_w5049_,
		_w6506_,
		_w6511_,
		_w6534_
	);
	LUT4 #(
		.INIT('h0080)
	) name2487 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w6535_
	);
	LUT4 #(
		.INIT('h000b)
	) name2488 (
		_w4970_,
		_w6523_,
		_w6535_,
		_w6534_,
		_w6536_
	);
	LUT4 #(
		.INIT('ha222)
	) name2489 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w6537_
	);
	LUT4 #(
		.INIT('h4000)
	) name2490 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w6538_
	);
	LUT4 #(
		.INIT('h2a00)
	) name2491 (
		\idma_DCTL_reg[11]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w6539_
	);
	LUT2 #(
		.INIT('h1)
	) name2492 (
		_w6538_,
		_w6539_,
		_w6540_
	);
	LUT3 #(
		.INIT('h20)
	) name2493 (
		_w5539_,
		_w6537_,
		_w6540_,
		_w6541_
	);
	LUT3 #(
		.INIT('hd0)
	) name2494 (
		_w5059_,
		_w6536_,
		_w6541_,
		_w6542_
	);
	LUT4 #(
		.INIT('h5540)
	) name2495 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w6543_
	);
	LUT4 #(
		.INIT('h3332)
	) name2496 (
		_w5117_,
		_w5337_,
		_w6543_,
		_w6542_,
		_w6544_
	);
	LUT4 #(
		.INIT('h7500)
	) name2497 (
		_w5117_,
		_w6529_,
		_w6533_,
		_w6544_,
		_w6545_
	);
	LUT2 #(
		.INIT('h9)
	) name2498 (
		_w5178_,
		_w5296_,
		_w6546_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2499 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w6546_,
		_w6547_
	);
	LUT3 #(
		.INIT('h96)
	) name2500 (
		_w5169_,
		_w5177_,
		_w5178_,
		_w6548_
	);
	LUT4 #(
		.INIT('hab54)
	) name2501 (
		_w5187_,
		_w5188_,
		_w5191_,
		_w6548_,
		_w6549_
	);
	LUT4 #(
		.INIT('h0065)
	) name2502 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w6549_,
		_w6550_
	);
	LUT3 #(
		.INIT('h01)
	) name2503 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6550_,
		_w6547_,
		_w6551_
	);
	LUT3 #(
		.INIT('ha8)
	) name2504 (
		\core_dag_ilm1reg_I_reg[2]/NET0131 ,
		_w5165_,
		_w5167_,
		_w6552_
	);
	LUT3 #(
		.INIT('h10)
	) name2505 (
		_w5767_,
		_w5768_,
		_w6546_,
		_w6553_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2506 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5155_,
		_w5310_,
		_w6549_,
		_w6554_
	);
	LUT4 #(
		.INIT('h1011)
	) name2507 (
		_w6552_,
		_w6551_,
		_w6553_,
		_w6554_,
		_w6555_
	);
	LUT4 #(
		.INIT('h0200)
	) name2508 (
		\core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w6556_
	);
	LUT4 #(
		.INIT('h0200)
	) name2509 (
		\core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w6557_
	);
	LUT4 #(
		.INIT('h0200)
	) name2510 (
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w6558_
	);
	LUT4 #(
		.INIT('h0200)
	) name2511 (
		\core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w6559_
	);
	LUT3 #(
		.INIT('h01)
	) name2512 (
		_w6558_,
		_w6559_,
		_w6557_,
		_w6560_
	);
	LUT3 #(
		.INIT('h02)
	) name2513 (
		\core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 ,
		_w5070_,
		_w5073_,
		_w6561_
	);
	LUT4 #(
		.INIT('h0200)
	) name2514 (
		\core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w6562_
	);
	LUT4 #(
		.INIT('h0200)
	) name2515 (
		\core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w6563_
	);
	LUT4 #(
		.INIT('h0200)
	) name2516 (
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w6564_
	);
	LUT4 #(
		.INIT('h0200)
	) name2517 (
		\core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w6565_
	);
	LUT4 #(
		.INIT('h0001)
	) name2518 (
		_w6562_,
		_w6563_,
		_w6564_,
		_w6565_,
		_w6566_
	);
	LUT4 #(
		.INIT('h45ef)
	) name2519 (
		_w4063_,
		_w6556_,
		_w6560_,
		_w6566_,
		_w6567_
	);
	LUT3 #(
		.INIT('h8c)
	) name2520 (
		_w5117_,
		_w5337_,
		_w6567_,
		_w6568_
	);
	LUT4 #(
		.INIT('h0233)
	) name2521 (
		_w5117_,
		_w5586_,
		_w6555_,
		_w6568_,
		_w6569_
	);
	LUT3 #(
		.INIT('h45)
	) name2522 (
		_w6526_,
		_w6545_,
		_w6569_,
		_w6570_
	);
	LUT3 #(
		.INIT('hba)
	) name2523 (
		_w6526_,
		_w6545_,
		_w6569_,
		_w6571_
	);
	LUT4 #(
		.INIT('h708f)
	) name2524 (
		_w5391_,
		_w5428_,
		_w5432_,
		_w5519_,
		_w6572_
	);
	LUT2 #(
		.INIT('h9)
	) name2525 (
		_w5518_,
		_w5520_,
		_w6573_
	);
	LUT3 #(
		.INIT('hb4)
	) name2526 (
		_w5509_,
		_w5514_,
		_w6573_,
		_w6574_
	);
	LUT4 #(
		.INIT('h0100)
	) name2527 (
		_w5379_,
		_w5383_,
		_w5433_,
		_w6574_,
		_w6575_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2528 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5435_,
		_w6572_,
		_w6575_,
		_w6576_
	);
	LUT2 #(
		.INIT('h2)
	) name2529 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		_w5382_,
		_w6577_
	);
	LUT3 #(
		.INIT('h06)
	) name2530 (
		_w5443_,
		_w5525_,
		_w6572_,
		_w6578_
	);
	LUT4 #(
		.INIT('h1455)
	) name2531 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5443_,
		_w5525_,
		_w6574_,
		_w6579_
	);
	LUT3 #(
		.INIT('h45)
	) name2532 (
		_w6577_,
		_w6578_,
		_w6579_,
		_w6580_
	);
	LUT3 #(
		.INIT('h45)
	) name2533 (
		_w5337_,
		_w6576_,
		_w6580_,
		_w6581_
	);
	LUT3 #(
		.INIT('h87)
	) name2534 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w5182_,
		_w5185_,
		_w6582_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2535 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w6582_,
		_w6583_
	);
	LUT4 #(
		.INIT('h718e)
	) name2536 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w5182_,
		_w5183_,
		_w5186_,
		_w6584_
	);
	LUT4 #(
		.INIT('he718)
	) name2537 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w5182_,
		_w5183_,
		_w5186_,
		_w6585_
	);
	LUT4 #(
		.INIT('h6500)
	) name2538 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w6585_,
		_w6586_
	);
	LUT3 #(
		.INIT('h01)
	) name2539 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6586_,
		_w6583_,
		_w6587_
	);
	LUT2 #(
		.INIT('h8)
	) name2540 (
		\core_dag_ilm1reg_I_reg[1]/NET0131 ,
		_w5173_,
		_w6588_
	);
	LUT3 #(
		.INIT('h0e)
	) name2541 (
		_w5767_,
		_w5768_,
		_w6584_,
		_w6589_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2542 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5155_,
		_w5310_,
		_w6582_,
		_w6590_
	);
	LUT4 #(
		.INIT('h0045)
	) name2543 (
		_w6588_,
		_w6589_,
		_w6590_,
		_w6587_,
		_w6591_
	);
	LUT3 #(
		.INIT('ha2)
	) name2544 (
		_w5117_,
		_w5337_,
		_w6591_,
		_w6592_
	);
	LUT4 #(
		.INIT('h0200)
	) name2545 (
		\core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w6593_
	);
	LUT4 #(
		.INIT('h0200)
	) name2546 (
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w6594_
	);
	LUT4 #(
		.INIT('h0200)
	) name2547 (
		\core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w6595_
	);
	LUT4 #(
		.INIT('h0200)
	) name2548 (
		\core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w6596_
	);
	LUT3 #(
		.INIT('h01)
	) name2549 (
		_w6595_,
		_w6596_,
		_w6594_,
		_w6597_
	);
	LUT4 #(
		.INIT('h0200)
	) name2550 (
		\core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w6598_
	);
	LUT4 #(
		.INIT('h0200)
	) name2551 (
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w6599_
	);
	LUT4 #(
		.INIT('h0200)
	) name2552 (
		\core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w6600_
	);
	LUT4 #(
		.INIT('h0200)
	) name2553 (
		\core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w6601_
	);
	LUT4 #(
		.INIT('h0001)
	) name2554 (
		_w6598_,
		_w6599_,
		_w6600_,
		_w6601_,
		_w6602_
	);
	LUT4 #(
		.INIT('h45ef)
	) name2555 (
		_w4063_,
		_w6593_,
		_w6597_,
		_w6602_,
		_w6603_
	);
	LUT4 #(
		.INIT('h0200)
	) name2556 (
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w6604_
	);
	LUT4 #(
		.INIT('h0200)
	) name2557 (
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w6605_
	);
	LUT4 #(
		.INIT('h0200)
	) name2558 (
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w6606_
	);
	LUT4 #(
		.INIT('h0200)
	) name2559 (
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w6607_
	);
	LUT4 #(
		.INIT('h0001)
	) name2560 (
		_w6604_,
		_w6605_,
		_w6606_,
		_w6607_,
		_w6608_
	);
	LUT4 #(
		.INIT('h0200)
	) name2561 (
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w6609_
	);
	LUT4 #(
		.INIT('h0200)
	) name2562 (
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w6610_
	);
	LUT4 #(
		.INIT('h0200)
	) name2563 (
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w6611_
	);
	LUT4 #(
		.INIT('h0200)
	) name2564 (
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w6612_
	);
	LUT4 #(
		.INIT('h0001)
	) name2565 (
		_w6609_,
		_w6610_,
		_w6611_,
		_w6612_,
		_w6613_
	);
	LUT3 #(
		.INIT('hd0)
	) name2566 (
		_w4063_,
		_w6608_,
		_w6613_,
		_w6614_
	);
	LUT4 #(
		.INIT('h0233)
	) name2567 (
		_w4063_,
		_w5049_,
		_w6608_,
		_w6613_,
		_w6615_
	);
	LUT4 #(
		.INIT('h0080)
	) name2568 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w6616_
	);
	LUT4 #(
		.INIT('h0203)
	) name2569 (
		_w4970_,
		_w6615_,
		_w6616_,
		_w6603_,
		_w6617_
	);
	LUT4 #(
		.INIT('ha222)
	) name2570 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w6618_
	);
	LUT4 #(
		.INIT('h2a00)
	) name2571 (
		\idma_DCTL_reg[12]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w6619_
	);
	LUT4 #(
		.INIT('h4000)
	) name2572 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w6620_
	);
	LUT2 #(
		.INIT('h1)
	) name2573 (
		_w6619_,
		_w6620_,
		_w6621_
	);
	LUT3 #(
		.INIT('h20)
	) name2574 (
		_w5539_,
		_w6618_,
		_w6621_,
		_w6622_
	);
	LUT3 #(
		.INIT('hd0)
	) name2575 (
		_w5059_,
		_w6617_,
		_w6622_,
		_w6623_
	);
	LUT4 #(
		.INIT('h5540)
	) name2576 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w6624_
	);
	LUT3 #(
		.INIT('h01)
	) name2577 (
		_w5337_,
		_w6624_,
		_w6623_,
		_w6625_
	);
	LUT4 #(
		.INIT('h0200)
	) name2578 (
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w6626_
	);
	LUT3 #(
		.INIT('h02)
	) name2579 (
		\core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 ,
		_w5079_,
		_w5082_,
		_w6627_
	);
	LUT4 #(
		.INIT('h0200)
	) name2580 (
		\core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w6628_
	);
	LUT3 #(
		.INIT('h02)
	) name2581 (
		\core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 ,
		_w5061_,
		_w5065_,
		_w6629_
	);
	LUT4 #(
		.INIT('h0200)
	) name2582 (
		\core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w6630_
	);
	LUT4 #(
		.INIT('h0200)
	) name2583 (
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w6631_
	);
	LUT3 #(
		.INIT('h01)
	) name2584 (
		_w6630_,
		_w6631_,
		_w6628_,
		_w6632_
	);
	LUT4 #(
		.INIT('h0200)
	) name2585 (
		\core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w6633_
	);
	LUT4 #(
		.INIT('h0200)
	) name2586 (
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w6634_
	);
	LUT4 #(
		.INIT('h0200)
	) name2587 (
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w6635_
	);
	LUT4 #(
		.INIT('h0200)
	) name2588 (
		\core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w6636_
	);
	LUT4 #(
		.INIT('h0001)
	) name2589 (
		_w6633_,
		_w6634_,
		_w6635_,
		_w6636_,
		_w6637_
	);
	LUT4 #(
		.INIT('h45ef)
	) name2590 (
		_w4063_,
		_w6626_,
		_w6632_,
		_w6637_,
		_w6638_
	);
	LUT3 #(
		.INIT('h15)
	) name2591 (
		_w5117_,
		_w5337_,
		_w6638_,
		_w6639_
	);
	LUT3 #(
		.INIT('h45)
	) name2592 (
		_w5586_,
		_w6625_,
		_w6639_,
		_w6640_
	);
	LUT2 #(
		.INIT('h9)
	) name2593 (
		_w5281_,
		_w5283_,
		_w6641_
	);
	LUT4 #(
		.INIT('h708f)
	) name2594 (
		_w5251_,
		_w5270_,
		_w5275_,
		_w6641_,
		_w6642_
	);
	LUT3 #(
		.INIT('he0)
	) name2595 (
		_w5767_,
		_w5918_,
		_w6642_,
		_w6643_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2596 (
		\core_dag_ilm1reg_I_reg[12]/NET0131 ,
		_w5264_,
		_w5265_,
		_w5277_,
		_w6644_
	);
	LUT2 #(
		.INIT('h6)
	) name2597 (
		_w5282_,
		_w5309_,
		_w6645_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name2598 (
		_w5767_,
		_w5918_,
		_w6644_,
		_w6645_,
		_w6646_
	);
	LUT3 #(
		.INIT('ha8)
	) name2599 (
		\DM_rd0[12]_pad ,
		_w5610_,
		_w5612_,
		_w6647_
	);
	LUT4 #(
		.INIT('h135f)
	) name2600 (
		\DM_rdm[12]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w6648_
	);
	LUT4 #(
		.INIT('h135f)
	) name2601 (
		\DM_rd6[12]_pad ,
		\DM_rd7[12]_pad ,
		_w5596_,
		_w5591_,
		_w6649_
	);
	LUT2 #(
		.INIT('h8)
	) name2602 (
		_w6648_,
		_w6649_,
		_w6650_
	);
	LUT3 #(
		.INIT('h80)
	) name2603 (
		\DM_rd5[12]_pad ,
		_w5598_,
		_w5599_,
		_w6651_
	);
	LUT3 #(
		.INIT('h80)
	) name2604 (
		\DM_rd4[12]_pad ,
		_w5598_,
		_w5601_,
		_w6652_
	);
	LUT4 #(
		.INIT('h8000)
	) name2605 (
		\DM_rd2[12]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w6653_
	);
	LUT4 #(
		.INIT('h8000)
	) name2606 (
		\DM_rd1[12]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w6654_
	);
	LUT4 #(
		.INIT('h8000)
	) name2607 (
		\DM_rd3[12]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w6655_
	);
	LUT3 #(
		.INIT('h01)
	) name2608 (
		_w6654_,
		_w6655_,
		_w6653_,
		_w6656_
	);
	LUT3 #(
		.INIT('h10)
	) name2609 (
		_w6652_,
		_w6651_,
		_w6656_,
		_w6657_
	);
	LUT2 #(
		.INIT('h8)
	) name2610 (
		_w6650_,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h4)
	) name2611 (
		_w6647_,
		_w6658_,
		_w6659_
	);
	LUT4 #(
		.INIT('h4000)
	) name2612 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[12]/P0001 ,
		_w6660_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2613 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4210_,
		_w4207_,
		_w4215_,
		_w6661_
	);
	LUT3 #(
		.INIT('ha8)
	) name2614 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w6662_
	);
	LUT4 #(
		.INIT('h135f)
	) name2615 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w6663_
	);
	LUT2 #(
		.INIT('h4)
	) name2616 (
		_w6662_,
		_w6663_,
		_w6664_
	);
	LUT3 #(
		.INIT('h8a)
	) name2617 (
		_w5681_,
		_w6661_,
		_w6664_,
		_w6665_
	);
	LUT3 #(
		.INIT('h80)
	) name2618 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w5629_,
		_w5648_,
		_w6666_
	);
	LUT4 #(
		.INIT('h8000)
	) name2619 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_rxctl_SLOT1_EXT_reg[2]/NET0131 ,
		_w5634_,
		_w5660_,
		_w6667_
	);
	LUT4 #(
		.INIT('h8000)
	) name2620 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_rxctl_SLOT1_EXT_reg[2]/NET0131 ,
		_w5631_,
		_w5639_,
		_w6668_
	);
	LUT3 #(
		.INIT('h80)
	) name2621 (
		\memc_usysr_DO_reg[12]/NET0131 ,
		_w5631_,
		_w5660_,
		_w6669_
	);
	LUT3 #(
		.INIT('h80)
	) name2622 (
		\sport0_regs_AUTO_a_reg[12]/NET0131 ,
		_w5627_,
		_w5634_,
		_w6670_
	);
	LUT4 #(
		.INIT('h0001)
	) name2623 (
		_w6669_,
		_w6670_,
		_w6668_,
		_w6667_,
		_w6671_
	);
	LUT3 #(
		.INIT('h80)
	) name2624 (
		\bdma_BCTL_reg[12]/NET0131 ,
		_w5627_,
		_w5629_,
		_w6672_
	);
	LUT3 #(
		.INIT('h80)
	) name2625 (
		\bdma_BEAD_reg[12]/NET0131 ,
		_w5629_,
		_w5644_,
		_w6673_
	);
	LUT4 #(
		.INIT('h0100)
	) name2626 (
		_w6666_,
		_w6672_,
		_w6673_,
		_w6671_,
		_w6674_
	);
	LUT4 #(
		.INIT('h8000)
	) name2627 (
		\bdma_BWCOUNT_reg[12]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w6675_
	);
	LUT3 #(
		.INIT('h80)
	) name2628 (
		\PIO_out[8]_pad ,
		_w5628_,
		_w5635_,
		_w6676_
	);
	LUT3 #(
		.INIT('h80)
	) name2629 (
		\PIO_oe[8]_pad ,
		_w5628_,
		_w5632_,
		_w6677_
	);
	LUT3 #(
		.INIT('h80)
	) name2630 (
		\tm_tpr_reg_DO_reg[12]/NET0131 ,
		_w5631_,
		_w5635_,
		_w6678_
	);
	LUT3 #(
		.INIT('h80)
	) name2631 (
		\pio_PINT_reg[8]/NET0131 ,
		_w5670_,
		_w5672_,
		_w6679_
	);
	LUT4 #(
		.INIT('h0001)
	) name2632 (
		_w6676_,
		_w6677_,
		_w6678_,
		_w6679_,
		_w6680_
	);
	LUT3 #(
		.INIT('h80)
	) name2633 (
		\emc_WSCRreg_DO_reg[12]/NET0131 ,
		_w5631_,
		_w5632_,
		_w6681_
	);
	LUT3 #(
		.INIT('h80)
	) name2634 (
		\clkc_ckr_reg_DO_reg[12]/NET0131 ,
		_w5631_,
		_w5644_,
		_w6682_
	);
	LUT3 #(
		.INIT('h80)
	) name2635 (
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w5632_,
		_w5634_,
		_w6683_
	);
	LUT3 #(
		.INIT('h80)
	) name2636 (
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w5634_,
		_w5639_,
		_w6684_
	);
	LUT4 #(
		.INIT('h0001)
	) name2637 (
		_w6681_,
		_w6682_,
		_w6683_,
		_w6684_,
		_w6685_
	);
	LUT3 #(
		.INIT('h80)
	) name2638 (
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w5644_,
		_w5634_,
		_w6686_
	);
	LUT3 #(
		.INIT('h80)
	) name2639 (
		\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w5634_,
		_w5635_,
		_w6687_
	);
	LUT3 #(
		.INIT('h80)
	) name2640 (
		\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w5648_,
		_w5634_,
		_w6688_
	);
	LUT3 #(
		.INIT('h01)
	) name2641 (
		_w6687_,
		_w6688_,
		_w6686_,
		_w6689_
	);
	LUT3 #(
		.INIT('h80)
	) name2642 (
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w5634_,
		_w5637_,
		_w6690_
	);
	LUT3 #(
		.INIT('h80)
	) name2643 (
		\pio_pmask_reg_DO_reg[8]/NET0131 ,
		_w5628_,
		_w5660_,
		_w6691_
	);
	LUT3 #(
		.INIT('h80)
	) name2644 (
		\tm_TCR_TMP_reg[12]/NET0131 ,
		_w5631_,
		_w5637_,
		_w6692_
	);
	LUT3 #(
		.INIT('h80)
	) name2645 (
		\idma_DCTL_reg[12]/NET0131 ,
		_w5628_,
		_w5639_,
		_w6693_
	);
	LUT4 #(
		.INIT('h0001)
	) name2646 (
		_w6690_,
		_w6691_,
		_w6692_,
		_w6693_,
		_w6694_
	);
	LUT4 #(
		.INIT('h8000)
	) name2647 (
		_w6689_,
		_w6694_,
		_w6680_,
		_w6685_,
		_w6695_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2648 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w6675_,
		_w6695_,
		_w6674_,
		_w6696_
	);
	LUT4 #(
		.INIT('h135f)
	) name2649 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131 ,
		_w6697_
	);
	LUT4 #(
		.INIT('h135f)
	) name2650 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w6698_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		_w6697_,
		_w6698_,
		_w6699_
	);
	LUT4 #(
		.INIT('h135f)
	) name2652 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131 ,
		_w6700_
	);
	LUT4 #(
		.INIT('h135f)
	) name2653 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131 ,
		_w6701_
	);
	LUT4 #(
		.INIT('h135f)
	) name2654 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131 ,
		_w6702_
	);
	LUT4 #(
		.INIT('h135f)
	) name2655 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131 ,
		_w6703_
	);
	LUT4 #(
		.INIT('h8000)
	) name2656 (
		_w6702_,
		_w6703_,
		_w6700_,
		_w6701_,
		_w6704_
	);
	LUT3 #(
		.INIT('h2a)
	) name2657 (
		_w5687_,
		_w6699_,
		_w6704_,
		_w6705_
	);
	LUT4 #(
		.INIT('h135f)
	) name2658 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131 ,
		_w6706_
	);
	LUT4 #(
		.INIT('h135f)
	) name2659 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131 ,
		_w6707_
	);
	LUT2 #(
		.INIT('h8)
	) name2660 (
		_w6706_,
		_w6707_,
		_w6708_
	);
	LUT4 #(
		.INIT('h135f)
	) name2661 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131 ,
		_w6709_
	);
	LUT4 #(
		.INIT('h135f)
	) name2662 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131 ,
		_w6710_
	);
	LUT4 #(
		.INIT('h135f)
	) name2663 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131 ,
		_w6711_
	);
	LUT4 #(
		.INIT('h135f)
	) name2664 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131 ,
		_w6712_
	);
	LUT4 #(
		.INIT('h8000)
	) name2665 (
		_w6711_,
		_w6712_,
		_w6709_,
		_w6710_,
		_w6713_
	);
	LUT4 #(
		.INIT('h135f)
	) name2666 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[12]/P0001 ,
		\sport1_txctl_TX_reg[12]/P0001 ,
		_w6714_
	);
	LUT4 #(
		.INIT('h135f)
	) name2667 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[12]/P0001 ,
		\sport1_rxctl_RX_reg[12]/P0001 ,
		_w6715_
	);
	LUT3 #(
		.INIT('h2a)
	) name2668 (
		_w5706_,
		_w6714_,
		_w6715_,
		_w6716_
	);
	LUT4 #(
		.INIT('h00d5)
	) name2669 (
		_w5697_,
		_w6708_,
		_w6713_,
		_w6716_,
		_w6717_
	);
	LUT2 #(
		.INIT('h4)
	) name2670 (
		_w6705_,
		_w6717_,
		_w6718_
	);
	LUT3 #(
		.INIT('h1b)
	) name2671 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001 ,
		_w6719_
	);
	LUT4 #(
		.INIT('ha820)
	) name2672 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001 ,
		_w6720_
	);
	LUT3 #(
		.INIT('h1b)
	) name2673 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001 ,
		_w6721_
	);
	LUT4 #(
		.INIT('ha820)
	) name2674 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001 ,
		_w6722_
	);
	LUT3 #(
		.INIT('h1b)
	) name2675 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001 ,
		_w6723_
	);
	LUT4 #(
		.INIT('ha820)
	) name2676 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001 ,
		_w6724_
	);
	LUT3 #(
		.INIT('h01)
	) name2677 (
		_w6722_,
		_w6724_,
		_w6720_,
		_w6725_
	);
	LUT3 #(
		.INIT('h2a)
	) name2678 (
		_w5741_,
		_w5746_,
		_w6725_,
		_w6726_
	);
	LUT3 #(
		.INIT('h1b)
	) name2679 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001 ,
		_w6727_
	);
	LUT4 #(
		.INIT('ha820)
	) name2680 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001 ,
		_w6728_
	);
	LUT3 #(
		.INIT('h1b)
	) name2681 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001 ,
		_w6729_
	);
	LUT4 #(
		.INIT('ha820)
	) name2682 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001 ,
		_w6730_
	);
	LUT3 #(
		.INIT('h1b)
	) name2683 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001 ,
		_w6731_
	);
	LUT4 #(
		.INIT('ha820)
	) name2684 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001 ,
		_w6732_
	);
	LUT3 #(
		.INIT('h01)
	) name2685 (
		_w6730_,
		_w6732_,
		_w6728_,
		_w6733_
	);
	LUT3 #(
		.INIT('h1b)
	) name2686 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 ,
		_w6734_
	);
	LUT4 #(
		.INIT('ha820)
	) name2687 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 ,
		_w6735_
	);
	LUT3 #(
		.INIT('h1b)
	) name2688 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001 ,
		_w6736_
	);
	LUT4 #(
		.INIT('ha820)
	) name2689 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001 ,
		_w6737_
	);
	LUT3 #(
		.INIT('h1b)
	) name2690 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001 ,
		_w6738_
	);
	LUT4 #(
		.INIT('ha820)
	) name2691 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001 ,
		_w6739_
	);
	LUT4 #(
		.INIT('h0001)
	) name2692 (
		_w5714_,
		_w6735_,
		_w6737_,
		_w6739_,
		_w6740_
	);
	LUT3 #(
		.INIT('h2a)
	) name2693 (
		_w5712_,
		_w6733_,
		_w6740_,
		_w6741_
	);
	LUT3 #(
		.INIT('h1b)
	) name2694 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001 ,
		_w6742_
	);
	LUT4 #(
		.INIT('ha820)
	) name2695 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001 ,
		_w6743_
	);
	LUT4 #(
		.INIT('ha820)
	) name2696 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001 ,
		_w6744_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		_w6743_,
		_w6744_,
		_w6745_
	);
	LUT3 #(
		.INIT('h1b)
	) name2698 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001 ,
		_w6746_
	);
	LUT4 #(
		.INIT('ha820)
	) name2699 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001 ,
		_w6747_
	);
	LUT3 #(
		.INIT('h1b)
	) name2700 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001 ,
		_w6748_
	);
	LUT4 #(
		.INIT('ha820)
	) name2701 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001 ,
		_w6749_
	);
	LUT4 #(
		.INIT('ha820)
	) name2702 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001 ,
		_w6750_
	);
	LUT3 #(
		.INIT('h01)
	) name2703 (
		_w6749_,
		_w6750_,
		_w6747_,
		_w6751_
	);
	LUT3 #(
		.INIT('h2a)
	) name2704 (
		_w5730_,
		_w6745_,
		_w6751_,
		_w6752_
	);
	LUT3 #(
		.INIT('h01)
	) name2705 (
		_w6741_,
		_w6752_,
		_w6726_,
		_w6753_
	);
	LUT2 #(
		.INIT('h8)
	) name2706 (
		_w6718_,
		_w6753_,
		_w6754_
	);
	LUT4 #(
		.INIT('h0100)
	) name2707 (
		_w6660_,
		_w6696_,
		_w6665_,
		_w6754_,
		_w6755_
	);
	LUT2 #(
		.INIT('h8)
	) name2708 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[12]/P0001 ,
		_w6756_
	);
	LUT3 #(
		.INIT('h08)
	) name2709 (
		_w5588_,
		_w5598_,
		_w6756_,
		_w6757_
	);
	LUT4 #(
		.INIT('h0133)
	) name2710 (
		\emc_DMDoe_reg/NET0131 ,
		_w6659_,
		_w6755_,
		_w6757_,
		_w6758_
	);
	LUT4 #(
		.INIT('hc040)
	) name2711 (
		_w5117_,
		_w5337_,
		_w5586_,
		_w6758_,
		_w6759_
	);
	LUT4 #(
		.INIT('hef00)
	) name2712 (
		_w5117_,
		_w6643_,
		_w6646_,
		_w6759_,
		_w6760_
	);
	LUT2 #(
		.INIT('h2)
	) name2713 (
		_w6614_,
		_w6603_,
		_w6761_
	);
	LUT3 #(
		.INIT('ha8)
	) name2714 (
		\DM_rd0[1]_pad ,
		_w5610_,
		_w5612_,
		_w6762_
	);
	LUT4 #(
		.INIT('h135f)
	) name2715 (
		\DM_rdm[1]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w6763_
	);
	LUT4 #(
		.INIT('h135f)
	) name2716 (
		\DM_rd6[1]_pad ,
		\DM_rd7[1]_pad ,
		_w5596_,
		_w5591_,
		_w6764_
	);
	LUT2 #(
		.INIT('h8)
	) name2717 (
		_w6763_,
		_w6764_,
		_w6765_
	);
	LUT3 #(
		.INIT('h80)
	) name2718 (
		\DM_rd5[1]_pad ,
		_w5598_,
		_w5599_,
		_w6766_
	);
	LUT3 #(
		.INIT('h80)
	) name2719 (
		\DM_rd4[1]_pad ,
		_w5598_,
		_w5601_,
		_w6767_
	);
	LUT4 #(
		.INIT('h8000)
	) name2720 (
		\DM_rd2[1]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w6768_
	);
	LUT4 #(
		.INIT('h8000)
	) name2721 (
		\DM_rd1[1]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w6769_
	);
	LUT4 #(
		.INIT('h8000)
	) name2722 (
		\DM_rd3[1]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w6770_
	);
	LUT3 #(
		.INIT('h01)
	) name2723 (
		_w6769_,
		_w6770_,
		_w6768_,
		_w6771_
	);
	LUT3 #(
		.INIT('h10)
	) name2724 (
		_w6767_,
		_w6766_,
		_w6771_,
		_w6772_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		_w6765_,
		_w6772_,
		_w6773_
	);
	LUT2 #(
		.INIT('h4)
	) name2726 (
		_w6762_,
		_w6773_,
		_w6774_
	);
	LUT4 #(
		.INIT('h4000)
	) name2727 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[1]/P0001 ,
		_w6775_
	);
	LUT3 #(
		.INIT('h80)
	) name2728 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w5629_,
		_w5648_,
		_w6776_
	);
	LUT3 #(
		.INIT('h80)
	) name2729 (
		\emc_WSCRreg_DO_reg[1]/NET0131 ,
		_w5631_,
		_w5632_,
		_w6777_
	);
	LUT3 #(
		.INIT('h80)
	) name2730 (
		\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w5648_,
		_w5634_,
		_w6778_
	);
	LUT3 #(
		.INIT('h80)
	) name2731 (
		\idma_DOVL_reg[1]/NET0131 ,
		_w5804_,
		_w5824_,
		_w6779_
	);
	LUT3 #(
		.INIT('h80)
	) name2732 (
		\sport0_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w5627_,
		_w5634_,
		_w6780_
	);
	LUT4 #(
		.INIT('h0001)
	) name2733 (
		_w6777_,
		_w6778_,
		_w6779_,
		_w6780_,
		_w6781_
	);
	LUT3 #(
		.INIT('h80)
	) name2734 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w5632_,
		_w5634_,
		_w6782_
	);
	LUT3 #(
		.INIT('h80)
	) name2735 (
		\tm_tsr_reg_DO_reg[1]/NET0131 ,
		_w5627_,
		_w5631_,
		_w6783_
	);
	LUT3 #(
		.INIT('h80)
	) name2736 (
		\sport1_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w5631_,
		_w5639_,
		_w6784_
	);
	LUT4 #(
		.INIT('h0001)
	) name2737 (
		_w5795_,
		_w6782_,
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT3 #(
		.INIT('h40)
	) name2738 (
		_w6776_,
		_w6781_,
		_w6785_,
		_w6786_
	);
	LUT3 #(
		.INIT('h80)
	) name2739 (
		\bdma_BEAD_reg[1]/NET0131 ,
		_w5629_,
		_w5644_,
		_w6787_
	);
	LUT3 #(
		.INIT('h80)
	) name2740 (
		\bdma_BCTL_reg[1]/NET0131 ,
		_w5627_,
		_w5629_,
		_w6788_
	);
	LUT2 #(
		.INIT('h1)
	) name2741 (
		_w6787_,
		_w6788_,
		_w6789_
	);
	LUT2 #(
		.INIT('h8)
	) name2742 (
		_w6786_,
		_w6789_,
		_w6790_
	);
	LUT4 #(
		.INIT('h8000)
	) name2743 (
		\bdma_BOVL_reg[1]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w6791_
	);
	LUT4 #(
		.INIT('h8000)
	) name2744 (
		\bdma_BWCOUNT_reg[1]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w6792_
	);
	LUT3 #(
		.INIT('h80)
	) name2745 (
		\PIO_oe[1]_pad ,
		_w5628_,
		_w5632_,
		_w6793_
	);
	LUT3 #(
		.INIT('h80)
	) name2746 (
		\sport0_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w5634_,
		_w5660_,
		_w6794_
	);
	LUT3 #(
		.INIT('h80)
	) name2747 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w5628_,
		_w5639_,
		_w6795_
	);
	LUT3 #(
		.INIT('h80)
	) name2748 (
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w5634_,
		_w5639_,
		_w6796_
	);
	LUT4 #(
		.INIT('h0001)
	) name2749 (
		_w6793_,
		_w6794_,
		_w6795_,
		_w6796_,
		_w6797_
	);
	LUT3 #(
		.INIT('h80)
	) name2750 (
		\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w5634_,
		_w5635_,
		_w6798_
	);
	LUT3 #(
		.INIT('h80)
	) name2751 (
		\emc_WSCRext_reg_DO_reg[1]/NET0131 ,
		_w5670_,
		_w5790_,
		_w6799_
	);
	LUT3 #(
		.INIT('h80)
	) name2752 (
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w5634_,
		_w5637_,
		_w6800_
	);
	LUT3 #(
		.INIT('h80)
	) name2753 (
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w5670_,
		_w5810_,
		_w6801_
	);
	LUT4 #(
		.INIT('h0001)
	) name2754 (
		_w6798_,
		_w6799_,
		_w6800_,
		_w6801_,
		_w6802_
	);
	LUT3 #(
		.INIT('h80)
	) name2755 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w5644_,
		_w5634_,
		_w6803_
	);
	LUT3 #(
		.INIT('h80)
	) name2756 (
		\pio_pmask_reg_DO_reg[1]/NET0131 ,
		_w5628_,
		_w5660_,
		_w6804_
	);
	LUT3 #(
		.INIT('h80)
	) name2757 (
		\PIO_out[1]_pad ,
		_w5628_,
		_w5635_,
		_w6805_
	);
	LUT3 #(
		.INIT('h80)
	) name2758 (
		\tm_TCR_TMP_reg[1]/NET0131 ,
		_w5631_,
		_w5637_,
		_w6806_
	);
	LUT4 #(
		.INIT('h0001)
	) name2759 (
		_w6803_,
		_w6804_,
		_w6805_,
		_w6806_,
		_w6807_
	);
	LUT3 #(
		.INIT('h80)
	) name2760 (
		\memc_usysr_DO_reg[1]/NET0131 ,
		_w5631_,
		_w5660_,
		_w6808_
	);
	LUT3 #(
		.INIT('h80)
	) name2761 (
		\tm_tpr_reg_DO_reg[1]/NET0131 ,
		_w5631_,
		_w5635_,
		_w6809_
	);
	LUT3 #(
		.INIT('h80)
	) name2762 (
		\clkc_ckr_reg_DO_reg[1]/NET0131 ,
		_w5631_,
		_w5644_,
		_w6810_
	);
	LUT3 #(
		.INIT('h80)
	) name2763 (
		\pio_PINT_reg[1]/NET0131 ,
		_w5670_,
		_w5672_,
		_w6811_
	);
	LUT4 #(
		.INIT('h0001)
	) name2764 (
		_w6808_,
		_w6809_,
		_w6810_,
		_w6811_,
		_w6812_
	);
	LUT4 #(
		.INIT('h8000)
	) name2765 (
		_w6807_,
		_w6812_,
		_w6797_,
		_w6802_,
		_w6813_
	);
	LUT3 #(
		.INIT('h10)
	) name2766 (
		_w6792_,
		_w6791_,
		_w6813_,
		_w6814_
	);
	LUT3 #(
		.INIT('h2a)
	) name2767 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w6790_,
		_w6814_,
		_w6815_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2768 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4352_,
		_w4349_,
		_w4357_,
		_w6816_
	);
	LUT4 #(
		.INIT('h135f)
	) name2769 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_SSTAT_reg[1]/NET0131 ,
		_w6817_
	);
	LUT4 #(
		.INIT('h135f)
	) name2770 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_ICNTL_reg_DO_reg[1]/NET0131 ,
		_w6818_
	);
	LUT2 #(
		.INIT('h8)
	) name2771 (
		_w6817_,
		_w6818_,
		_w6819_
	);
	LUT3 #(
		.INIT('ha8)
	) name2772 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w6820_
	);
	LUT4 #(
		.INIT('h135f)
	) name2773 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w6821_
	);
	LUT4 #(
		.INIT('h153f)
	) name2774 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w6822_
	);
	LUT3 #(
		.INIT('h40)
	) name2775 (
		_w6820_,
		_w6821_,
		_w6822_,
		_w6823_
	);
	LUT2 #(
		.INIT('h8)
	) name2776 (
		_w6819_,
		_w6823_,
		_w6824_
	);
	LUT3 #(
		.INIT('h8a)
	) name2777 (
		_w5681_,
		_w6816_,
		_w6824_,
		_w6825_
	);
	LUT4 #(
		.INIT('h135f)
	) name2778 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131 ,
		_w6826_
	);
	LUT4 #(
		.INIT('h135f)
	) name2779 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131 ,
		_w6827_
	);
	LUT2 #(
		.INIT('h8)
	) name2780 (
		_w6826_,
		_w6827_,
		_w6828_
	);
	LUT4 #(
		.INIT('h135f)
	) name2781 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131 ,
		_w6829_
	);
	LUT4 #(
		.INIT('h135f)
	) name2782 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131 ,
		_w6830_
	);
	LUT4 #(
		.INIT('h135f)
	) name2783 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w6831_
	);
	LUT4 #(
		.INIT('h135f)
	) name2784 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w6832_
	);
	LUT4 #(
		.INIT('h8000)
	) name2785 (
		_w6831_,
		_w6832_,
		_w6829_,
		_w6830_,
		_w6833_
	);
	LUT3 #(
		.INIT('h2a)
	) name2786 (
		_w5687_,
		_w6828_,
		_w6833_,
		_w6834_
	);
	LUT4 #(
		.INIT('h135f)
	) name2787 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w6835_
	);
	LUT4 #(
		.INIT('h135f)
	) name2788 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131 ,
		_w6836_
	);
	LUT2 #(
		.INIT('h8)
	) name2789 (
		_w6835_,
		_w6836_,
		_w6837_
	);
	LUT4 #(
		.INIT('h135f)
	) name2790 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w6838_
	);
	LUT4 #(
		.INIT('h135f)
	) name2791 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131 ,
		_w6839_
	);
	LUT4 #(
		.INIT('h135f)
	) name2792 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131 ,
		_w6840_
	);
	LUT4 #(
		.INIT('h135f)
	) name2793 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131 ,
		_w6841_
	);
	LUT4 #(
		.INIT('h8000)
	) name2794 (
		_w6840_,
		_w6841_,
		_w6838_,
		_w6839_,
		_w6842_
	);
	LUT4 #(
		.INIT('h135f)
	) name2795 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		\sport1_txctl_TX_reg[1]/P0001 ,
		_w6843_
	);
	LUT4 #(
		.INIT('h135f)
	) name2796 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		\sport1_rxctl_RX_reg[1]/P0001 ,
		_w6844_
	);
	LUT3 #(
		.INIT('h2a)
	) name2797 (
		_w5706_,
		_w6843_,
		_w6844_,
		_w6845_
	);
	LUT4 #(
		.INIT('h00d5)
	) name2798 (
		_w5697_,
		_w6837_,
		_w6842_,
		_w6845_,
		_w6846_
	);
	LUT2 #(
		.INIT('h4)
	) name2799 (
		_w6834_,
		_w6846_,
		_w6847_
	);
	LUT3 #(
		.INIT('h1b)
	) name2800 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001 ,
		_w6848_
	);
	LUT4 #(
		.INIT('ha820)
	) name2801 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001 ,
		_w6849_
	);
	LUT2 #(
		.INIT('h8)
	) name2802 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w6850_
	);
	LUT2 #(
		.INIT('h1)
	) name2803 (
		_w6849_,
		_w6850_,
		_w6851_
	);
	LUT3 #(
		.INIT('h1b)
	) name2804 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001 ,
		_w6852_
	);
	LUT4 #(
		.INIT('ha820)
	) name2805 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001 ,
		_w6853_
	);
	LUT3 #(
		.INIT('h1b)
	) name2806 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001 ,
		_w6854_
	);
	LUT4 #(
		.INIT('ha820)
	) name2807 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001 ,
		_w6855_
	);
	LUT4 #(
		.INIT('ha820)
	) name2808 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001 ,
		_w6856_
	);
	LUT4 #(
		.INIT('ha820)
	) name2809 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001 ,
		_w6857_
	);
	LUT4 #(
		.INIT('h0001)
	) name2810 (
		_w6853_,
		_w6855_,
		_w6856_,
		_w6857_,
		_w6858_
	);
	LUT3 #(
		.INIT('h2a)
	) name2811 (
		_w5730_,
		_w6851_,
		_w6858_,
		_w6859_
	);
	LUT3 #(
		.INIT('h1b)
	) name2812 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 ,
		_w6860_
	);
	LUT4 #(
		.INIT('ha820)
	) name2813 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 ,
		_w6861_
	);
	LUT3 #(
		.INIT('h1b)
	) name2814 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001 ,
		_w6862_
	);
	LUT4 #(
		.INIT('ha820)
	) name2815 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001 ,
		_w6863_
	);
	LUT3 #(
		.INIT('h1b)
	) name2816 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001 ,
		_w6864_
	);
	LUT4 #(
		.INIT('ha820)
	) name2817 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001 ,
		_w6865_
	);
	LUT3 #(
		.INIT('h01)
	) name2818 (
		_w6863_,
		_w6865_,
		_w6861_,
		_w6866_
	);
	LUT3 #(
		.INIT('h1b)
	) name2819 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 ,
		_w6867_
	);
	LUT4 #(
		.INIT('ha820)
	) name2820 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 ,
		_w6868_
	);
	LUT3 #(
		.INIT('h1b)
	) name2821 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001 ,
		_w6869_
	);
	LUT4 #(
		.INIT('ha820)
	) name2822 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001 ,
		_w6870_
	);
	LUT3 #(
		.INIT('h1b)
	) name2823 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001 ,
		_w6871_
	);
	LUT4 #(
		.INIT('ha820)
	) name2824 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001 ,
		_w6872_
	);
	LUT3 #(
		.INIT('h1b)
	) name2825 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001 ,
		_w6873_
	);
	LUT4 #(
		.INIT('ha820)
	) name2826 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001 ,
		_w6874_
	);
	LUT4 #(
		.INIT('h0001)
	) name2827 (
		_w6868_,
		_w6870_,
		_w6872_,
		_w6874_,
		_w6875_
	);
	LUT3 #(
		.INIT('h2a)
	) name2828 (
		_w5712_,
		_w6866_,
		_w6875_,
		_w6876_
	);
	LUT3 #(
		.INIT('h1b)
	) name2829 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001 ,
		_w6877_
	);
	LUT4 #(
		.INIT('ha820)
	) name2830 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001 ,
		_w6878_
	);
	LUT3 #(
		.INIT('h1b)
	) name2831 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[1]/P0001 ,
		_w6879_
	);
	LUT4 #(
		.INIT('ha820)
	) name2832 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_SBs_reg[1]/P0001 ,
		_w6880_
	);
	LUT2 #(
		.INIT('h1)
	) name2833 (
		_w6878_,
		_w6880_,
		_w6881_
	);
	LUT3 #(
		.INIT('h1b)
	) name2834 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001 ,
		_w6882_
	);
	LUT4 #(
		.INIT('ha820)
	) name2835 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001 ,
		_w6883_
	);
	LUT3 #(
		.INIT('h1b)
	) name2836 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001 ,
		_w6884_
	);
	LUT4 #(
		.INIT('ha820)
	) name2837 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001 ,
		_w6885_
	);
	LUT3 #(
		.INIT('h1b)
	) name2838 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001 ,
		_w6886_
	);
	LUT4 #(
		.INIT('ha820)
	) name2839 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001 ,
		_w6887_
	);
	LUT3 #(
		.INIT('h01)
	) name2840 (
		_w6885_,
		_w6887_,
		_w6883_,
		_w6888_
	);
	LUT3 #(
		.INIT('h2a)
	) name2841 (
		_w5741_,
		_w6881_,
		_w6888_,
		_w6889_
	);
	LUT3 #(
		.INIT('h01)
	) name2842 (
		_w6876_,
		_w6889_,
		_w6859_,
		_w6890_
	);
	LUT2 #(
		.INIT('h8)
	) name2843 (
		_w6847_,
		_w6890_,
		_w6891_
	);
	LUT2 #(
		.INIT('h4)
	) name2844 (
		_w6825_,
		_w6891_,
		_w6892_
	);
	LUT3 #(
		.INIT('h10)
	) name2845 (
		_w6775_,
		_w6815_,
		_w6892_,
		_w6893_
	);
	LUT4 #(
		.INIT('h5455)
	) name2846 (
		\emc_DMDoe_reg/NET0131 ,
		_w6775_,
		_w6815_,
		_w6892_,
		_w6894_
	);
	LUT2 #(
		.INIT('h8)
	) name2847 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[1]/P0001 ,
		_w6895_
	);
	LUT3 #(
		.INIT('h08)
	) name2848 (
		_w5588_,
		_w5598_,
		_w6895_,
		_w6896_
	);
	LUT3 #(
		.INIT('h45)
	) name2849 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w6897_
	);
	LUT4 #(
		.INIT('hecfd)
	) name2850 (
		_w5117_,
		_w5337_,
		_w6761_,
		_w6897_,
		_w6898_
	);
	LUT2 #(
		.INIT('h2)
	) name2851 (
		_w5586_,
		_w6898_,
		_w6899_
	);
	LUT2 #(
		.INIT('h1)
	) name2852 (
		_w6760_,
		_w6899_,
		_w6900_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2853 (
		_w6581_,
		_w6592_,
		_w6640_,
		_w6900_,
		_w6901_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name2854 (
		_w6581_,
		_w6592_,
		_w6640_,
		_w6900_,
		_w6902_
	);
	LUT2 #(
		.INIT('h9)
	) name2855 (
		_w5515_,
		_w5517_,
		_w6903_
	);
	LUT4 #(
		.INIT('h00f4)
	) name2856 (
		_w5509_,
		_w5514_,
		_w5521_,
		_w5523_,
		_w6904_
	);
	LUT2 #(
		.INIT('h9)
	) name2857 (
		_w6903_,
		_w6904_,
		_w6905_
	);
	LUT2 #(
		.INIT('h6)
	) name2858 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5378_,
		_w6906_
	);
	LUT3 #(
		.INIT('h1e)
	) name2859 (
		_w5383_,
		_w5433_,
		_w6906_,
		_w6907_
	);
	LUT4 #(
		.INIT('h8882)
	) name2860 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5378_,
		_w5383_,
		_w5433_,
		_w6908_
	);
	LUT3 #(
		.INIT('hd0)
	) name2861 (
		_w5435_,
		_w6905_,
		_w6908_,
		_w6909_
	);
	LUT4 #(
		.INIT('h5140)
	) name2862 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5526_,
		_w6905_,
		_w6907_,
		_w6910_
	);
	LUT4 #(
		.INIT('h02a2)
	) name2863 (
		\core_dag_ilm2reg_I_reg[13]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w5370_,
		_w5377_,
		_w6911_
	);
	LUT4 #(
		.INIT('h5554)
	) name2864 (
		_w5337_,
		_w6909_,
		_w6910_,
		_w6911_,
		_w6912_
	);
	LUT3 #(
		.INIT('ha2)
	) name2865 (
		_w5117_,
		_w5337_,
		_w5771_,
		_w6913_
	);
	LUT4 #(
		.INIT('h0200)
	) name2866 (
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w6914_
	);
	LUT4 #(
		.INIT('h0200)
	) name2867 (
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w6915_
	);
	LUT4 #(
		.INIT('h0200)
	) name2868 (
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w6916_
	);
	LUT4 #(
		.INIT('h0200)
	) name2869 (
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w6917_
	);
	LUT4 #(
		.INIT('h0001)
	) name2870 (
		_w6914_,
		_w6915_,
		_w6916_,
		_w6917_,
		_w6918_
	);
	LUT4 #(
		.INIT('h0200)
	) name2871 (
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w6919_
	);
	LUT4 #(
		.INIT('h0200)
	) name2872 (
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w6920_
	);
	LUT4 #(
		.INIT('h0200)
	) name2873 (
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w6921_
	);
	LUT4 #(
		.INIT('h0200)
	) name2874 (
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w6922_
	);
	LUT4 #(
		.INIT('h0001)
	) name2875 (
		_w6919_,
		_w6920_,
		_w6921_,
		_w6922_,
		_w6923_
	);
	LUT3 #(
		.INIT('hd0)
	) name2876 (
		_w4063_,
		_w6918_,
		_w6923_,
		_w6924_
	);
	LUT4 #(
		.INIT('h0233)
	) name2877 (
		_w4063_,
		_w5049_,
		_w6918_,
		_w6923_,
		_w6925_
	);
	LUT4 #(
		.INIT('h0080)
	) name2878 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w6926_
	);
	LUT4 #(
		.INIT('h000b)
	) name2879 (
		_w4970_,
		_w5326_,
		_w6926_,
		_w6925_,
		_w6927_
	);
	LUT4 #(
		.INIT('ha222)
	) name2880 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w6928_
	);
	LUT4 #(
		.INIT('h4000)
	) name2881 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w6929_
	);
	LUT4 #(
		.INIT('h2a00)
	) name2882 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w6930_
	);
	LUT2 #(
		.INIT('h1)
	) name2883 (
		_w6929_,
		_w6930_,
		_w6931_
	);
	LUT3 #(
		.INIT('h20)
	) name2884 (
		_w5539_,
		_w6928_,
		_w6931_,
		_w6932_
	);
	LUT3 #(
		.INIT('hd0)
	) name2885 (
		_w5059_,
		_w6927_,
		_w6932_,
		_w6933_
	);
	LUT4 #(
		.INIT('h5540)
	) name2886 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w6934_
	);
	LUT3 #(
		.INIT('h01)
	) name2887 (
		_w5337_,
		_w6934_,
		_w6933_,
		_w6935_
	);
	LUT3 #(
		.INIT('h15)
	) name2888 (
		_w5117_,
		_w5337_,
		_w5563_,
		_w6936_
	);
	LUT3 #(
		.INIT('h45)
	) name2889 (
		_w5586_,
		_w6935_,
		_w6936_,
		_w6937_
	);
	LUT2 #(
		.INIT('h4)
	) name2890 (
		_w5326_,
		_w6924_,
		_w6938_
	);
	LUT4 #(
		.INIT('hefcd)
	) name2891 (
		_w5117_,
		_w5337_,
		_w5914_,
		_w6938_,
		_w6939_
	);
	LUT2 #(
		.INIT('h2)
	) name2892 (
		_w5586_,
		_w6939_,
		_w6940_
	);
	LUT4 #(
		.INIT('hc040)
	) name2893 (
		_w5117_,
		_w5337_,
		_w5586_,
		_w5760_,
		_w6941_
	);
	LUT4 #(
		.INIT('hef00)
	) name2894 (
		_w5117_,
		_w5312_,
		_w5315_,
		_w6941_,
		_w6942_
	);
	LUT2 #(
		.INIT('h1)
	) name2895 (
		_w6940_,
		_w6942_,
		_w6943_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2896 (
		_w6912_,
		_w6913_,
		_w6937_,
		_w6943_,
		_w6944_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name2897 (
		_w6912_,
		_w6913_,
		_w6937_,
		_w6943_,
		_w6945_
	);
	LUT4 #(
		.INIT('h0200)
	) name2898 (
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w6946_
	);
	LUT4 #(
		.INIT('h0200)
	) name2899 (
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w6947_
	);
	LUT4 #(
		.INIT('h0200)
	) name2900 (
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w6948_
	);
	LUT4 #(
		.INIT('h0200)
	) name2901 (
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w6949_
	);
	LUT4 #(
		.INIT('h0001)
	) name2902 (
		_w6946_,
		_w6947_,
		_w6948_,
		_w6949_,
		_w6950_
	);
	LUT4 #(
		.INIT('h0200)
	) name2903 (
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w6951_
	);
	LUT4 #(
		.INIT('h0200)
	) name2904 (
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w6952_
	);
	LUT4 #(
		.INIT('h0200)
	) name2905 (
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w6953_
	);
	LUT4 #(
		.INIT('h0200)
	) name2906 (
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w6954_
	);
	LUT4 #(
		.INIT('h0001)
	) name2907 (
		_w6951_,
		_w6952_,
		_w6953_,
		_w6954_,
		_w6955_
	);
	LUT3 #(
		.INIT('h1b)
	) name2908 (
		_w4063_,
		_w6950_,
		_w6955_,
		_w6956_
	);
	LUT2 #(
		.INIT('h1)
	) name2909 (
		_w6638_,
		_w6956_,
		_w6957_
	);
	LUT4 #(
		.INIT('h1032)
	) name2910 (
		_w5117_,
		_w5337_,
		_w6758_,
		_w6957_,
		_w6958_
	);
	LUT3 #(
		.INIT('hc4)
	) name2911 (
		_w5117_,
		_w5337_,
		_w6897_,
		_w6959_
	);
	LUT4 #(
		.INIT('h040f)
	) name2912 (
		_w5117_,
		_w6591_,
		_w6958_,
		_w6959_,
		_w6960_
	);
	LUT2 #(
		.INIT('h2)
	) name2913 (
		_w5586_,
		_w6960_,
		_w6961_
	);
	LUT3 #(
		.INIT('h69)
	) name2914 (
		\core_dag_ilm2reg_M_reg[1]/NET0131 ,
		_w5372_,
		_w5414_,
		_w6962_
	);
	LUT2 #(
		.INIT('h6)
	) name2915 (
		_w5480_,
		_w5481_,
		_w6963_
	);
	LUT4 #(
		.INIT('h0001)
	) name2916 (
		_w5379_,
		_w5383_,
		_w5433_,
		_w6963_,
		_w6964_
	);
	LUT4 #(
		.INIT('h080a)
	) name2917 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5435_,
		_w6964_,
		_w6962_,
		_w6965_
	);
	LUT3 #(
		.INIT('h20)
	) name2918 (
		\core_dag_ilm2reg_I_reg[1]/NET0131 ,
		_w5340_,
		_w5370_,
		_w6966_
	);
	LUT3 #(
		.INIT('h60)
	) name2919 (
		_w5443_,
		_w5525_,
		_w6962_,
		_w6967_
	);
	LUT3 #(
		.INIT('h69)
	) name2920 (
		_w5437_,
		_w5480_,
		_w5481_,
		_w6968_
	);
	LUT4 #(
		.INIT('h1455)
	) name2921 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w5443_,
		_w5525_,
		_w6968_,
		_w6969_
	);
	LUT3 #(
		.INIT('h45)
	) name2922 (
		_w6966_,
		_w6967_,
		_w6969_,
		_w6970_
	);
	LUT4 #(
		.INIT('h0123)
	) name2923 (
		_w4063_,
		_w5049_,
		_w6950_,
		_w6955_,
		_w6971_
	);
	LUT4 #(
		.INIT('h0800)
	) name2924 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w6972_
	);
	LUT4 #(
		.INIT('h000b)
	) name2925 (
		_w4970_,
		_w6638_,
		_w6971_,
		_w6972_,
		_w6973_
	);
	LUT4 #(
		.INIT('ha222)
	) name2926 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w6974_
	);
	LUT4 #(
		.INIT('h2a00)
	) name2927 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w6975_
	);
	LUT4 #(
		.INIT('h4000)
	) name2928 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[1]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w6976_
	);
	LUT2 #(
		.INIT('h1)
	) name2929 (
		_w6975_,
		_w6976_,
		_w6977_
	);
	LUT3 #(
		.INIT('h20)
	) name2930 (
		_w5539_,
		_w6974_,
		_w6977_,
		_w6978_
	);
	LUT3 #(
		.INIT('hd0)
	) name2931 (
		_w5059_,
		_w6973_,
		_w6978_,
		_w6979_
	);
	LUT4 #(
		.INIT('h5540)
	) name2932 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w6980_
	);
	LUT3 #(
		.INIT('h01)
	) name2933 (
		_w5117_,
		_w6980_,
		_w6979_,
		_w6981_
	);
	LUT4 #(
		.INIT('h0075)
	) name2934 (
		_w5117_,
		_w6965_,
		_w6970_,
		_w6981_,
		_w6982_
	);
	LUT3 #(
		.INIT('hc8)
	) name2935 (
		_w5117_,
		_w5337_,
		_w6603_,
		_w6983_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2936 (
		_w5117_,
		_w6643_,
		_w6646_,
		_w6983_,
		_w6984_
	);
	LUT4 #(
		.INIT('h3301)
	) name2937 (
		_w5337_,
		_w5586_,
		_w6982_,
		_w6984_,
		_w6985_
	);
	LUT2 #(
		.INIT('he)
	) name2938 (
		_w6961_,
		_w6985_,
		_w6986_
	);
	LUT4 #(
		.INIT('h0200)
	) name2939 (
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w6987_
	);
	LUT4 #(
		.INIT('h0200)
	) name2940 (
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w6988_
	);
	LUT4 #(
		.INIT('h0200)
	) name2941 (
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w6989_
	);
	LUT4 #(
		.INIT('h0200)
	) name2942 (
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w6990_
	);
	LUT4 #(
		.INIT('h0001)
	) name2943 (
		_w6987_,
		_w6988_,
		_w6989_,
		_w6990_,
		_w6991_
	);
	LUT4 #(
		.INIT('h0200)
	) name2944 (
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w6992_
	);
	LUT4 #(
		.INIT('h0200)
	) name2945 (
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w6993_
	);
	LUT4 #(
		.INIT('h0200)
	) name2946 (
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w6994_
	);
	LUT4 #(
		.INIT('h0200)
	) name2947 (
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w6995_
	);
	LUT4 #(
		.INIT('h0001)
	) name2948 (
		_w6992_,
		_w6993_,
		_w6994_,
		_w6995_,
		_w6996_
	);
	LUT3 #(
		.INIT('h1b)
	) name2949 (
		_w4063_,
		_w6991_,
		_w6996_,
		_w6997_
	);
	LUT2 #(
		.INIT('h1)
	) name2950 (
		_w6567_,
		_w6997_,
		_w6998_
	);
	LUT4 #(
		.INIT('h1032)
	) name2951 (
		_w5117_,
		_w5337_,
		_w6363_,
		_w6998_,
		_w6999_
	);
	LUT3 #(
		.INIT('hc4)
	) name2952 (
		_w5117_,
		_w5337_,
		_w6501_,
		_w7000_
	);
	LUT4 #(
		.INIT('h040f)
	) name2953 (
		_w5117_,
		_w6555_,
		_w6999_,
		_w7000_,
		_w7001_
	);
	LUT2 #(
		.INIT('h2)
	) name2954 (
		_w5586_,
		_w7001_,
		_w7002_
	);
	LUT2 #(
		.INIT('h6)
	) name2955 (
		_w5415_,
		_w5476_,
		_w7003_
	);
	LUT3 #(
		.INIT('he0)
	) name2956 (
		_w5434_,
		_w6210_,
		_w7003_,
		_w7004_
	);
	LUT4 #(
		.INIT('haa20)
	) name2957 (
		\core_dag_ilm2reg_I_reg[2]/NET0131 ,
		_w5341_,
		_w5370_,
		_w5411_,
		_w7005_
	);
	LUT2 #(
		.INIT('h9)
	) name2958 (
		_w5475_,
		_w5477_,
		_w7006_
	);
	LUT2 #(
		.INIT('h6)
	) name2959 (
		_w5483_,
		_w7006_,
		_w7007_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2960 (
		_w5434_,
		_w6210_,
		_w7005_,
		_w7007_,
		_w7008_
	);
	LUT4 #(
		.INIT('h0123)
	) name2961 (
		_w4063_,
		_w5049_,
		_w6991_,
		_w6996_,
		_w7009_
	);
	LUT4 #(
		.INIT('h0800)
	) name2962 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w7010_
	);
	LUT4 #(
		.INIT('h000b)
	) name2963 (
		_w4970_,
		_w6567_,
		_w7009_,
		_w7010_,
		_w7011_
	);
	LUT4 #(
		.INIT('ha222)
	) name2964 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w7012_
	);
	LUT4 #(
		.INIT('h2a00)
	) name2965 (
		\idma_DCTL_reg[2]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w7013_
	);
	LUT4 #(
		.INIT('h4000)
	) name2966 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[2]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w7014_
	);
	LUT2 #(
		.INIT('h1)
	) name2967 (
		_w7013_,
		_w7014_,
		_w7015_
	);
	LUT3 #(
		.INIT('h20)
	) name2968 (
		_w5539_,
		_w7012_,
		_w7015_,
		_w7016_
	);
	LUT3 #(
		.INIT('hd0)
	) name2969 (
		_w5059_,
		_w7011_,
		_w7016_,
		_w7017_
	);
	LUT4 #(
		.INIT('h5540)
	) name2970 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w7018_
	);
	LUT3 #(
		.INIT('h01)
	) name2971 (
		_w5117_,
		_w7018_,
		_w7017_,
		_w7019_
	);
	LUT4 #(
		.INIT('h0075)
	) name2972 (
		_w5117_,
		_w7004_,
		_w7008_,
		_w7019_,
		_w7020_
	);
	LUT3 #(
		.INIT('hc8)
	) name2973 (
		_w5117_,
		_w5337_,
		_w6523_,
		_w7021_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2974 (
		_w5117_,
		_w6245_,
		_w6250_,
		_w7021_,
		_w7022_
	);
	LUT4 #(
		.INIT('h3301)
	) name2975 (
		_w5337_,
		_w5586_,
		_w7020_,
		_w7022_,
		_w7023_
	);
	LUT2 #(
		.INIT('he)
	) name2976 (
		_w7002_,
		_w7023_,
		_w7024_
	);
	LUT4 #(
		.INIT('h0200)
	) name2977 (
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w7025_
	);
	LUT4 #(
		.INIT('h0200)
	) name2978 (
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w7026_
	);
	LUT4 #(
		.INIT('h0200)
	) name2979 (
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w7027_
	);
	LUT4 #(
		.INIT('h0200)
	) name2980 (
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w7028_
	);
	LUT4 #(
		.INIT('h0001)
	) name2981 (
		_w7025_,
		_w7026_,
		_w7027_,
		_w7028_,
		_w7029_
	);
	LUT4 #(
		.INIT('h0200)
	) name2982 (
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w7030_
	);
	LUT4 #(
		.INIT('h0200)
	) name2983 (
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w7031_
	);
	LUT4 #(
		.INIT('h0200)
	) name2984 (
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w7032_
	);
	LUT4 #(
		.INIT('h0200)
	) name2985 (
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w7033_
	);
	LUT4 #(
		.INIT('h0001)
	) name2986 (
		_w7030_,
		_w7031_,
		_w7032_,
		_w7033_,
		_w7034_
	);
	LUT3 #(
		.INIT('h1b)
	) name2987 (
		_w4063_,
		_w7029_,
		_w7034_,
		_w7035_
	);
	LUT2 #(
		.INIT('h1)
	) name2988 (
		_w6238_,
		_w7035_,
		_w7036_
	);
	LUT4 #(
		.INIT('h2301)
	) name2989 (
		_w5117_,
		_w5337_,
		_w6039_,
		_w7036_,
		_w7037_
	);
	LUT3 #(
		.INIT('h4c)
	) name2990 (
		_w5117_,
		_w5337_,
		_w6176_,
		_w7038_
	);
	LUT4 #(
		.INIT('hba00)
	) name2991 (
		_w5117_,
		_w6204_,
		_w6207_,
		_w7038_,
		_w7039_
	);
	LUT3 #(
		.INIT('ha8)
	) name2992 (
		_w5586_,
		_w7037_,
		_w7039_,
		_w7040_
	);
	LUT3 #(
		.INIT('h8c)
	) name2993 (
		_w5117_,
		_w5337_,
		_w6198_,
		_w7041_
	);
	LUT4 #(
		.INIT('h7500)
	) name2994 (
		_w5117_,
		_w5920_,
		_w5924_,
		_w7041_,
		_w7042_
	);
	LUT4 #(
		.INIT('h17e8)
	) name2995 (
		\core_dag_ilm2reg_M_reg[2]/NET0131 ,
		_w5412_,
		_w5415_,
		_w5470_,
		_w7043_
	);
	LUT3 #(
		.INIT('he0)
	) name2996 (
		_w5434_,
		_w6210_,
		_w7043_,
		_w7044_
	);
	LUT4 #(
		.INIT('haa08)
	) name2997 (
		\core_dag_ilm2reg_I_reg[3]/NET0131 ,
		_w5370_,
		_w5374_,
		_w5406_,
		_w7045_
	);
	LUT2 #(
		.INIT('h9)
	) name2998 (
		_w5469_,
		_w5471_,
		_w7046_
	);
	LUT4 #(
		.INIT('hab54)
	) name2999 (
		_w5478_,
		_w5479_,
		_w5483_,
		_w7046_,
		_w7047_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3000 (
		_w5434_,
		_w6210_,
		_w7045_,
		_w7047_,
		_w7048_
	);
	LUT4 #(
		.INIT('h0123)
	) name3001 (
		_w4063_,
		_w5049_,
		_w7029_,
		_w7034_,
		_w7049_
	);
	LUT4 #(
		.INIT('h0800)
	) name3002 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w7050_
	);
	LUT4 #(
		.INIT('h000b)
	) name3003 (
		_w4970_,
		_w6238_,
		_w7050_,
		_w7049_,
		_w7051_
	);
	LUT4 #(
		.INIT('ha222)
	) name3004 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w7052_
	);
	LUT4 #(
		.INIT('h2a00)
	) name3005 (
		\idma_DCTL_reg[3]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w7053_
	);
	LUT4 #(
		.INIT('h4000)
	) name3006 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[3]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w7054_
	);
	LUT2 #(
		.INIT('h1)
	) name3007 (
		_w7053_,
		_w7054_,
		_w7055_
	);
	LUT2 #(
		.INIT('h4)
	) name3008 (
		_w7052_,
		_w7055_,
		_w7056_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3009 (
		_w5059_,
		_w5539_,
		_w7051_,
		_w7056_,
		_w7057_
	);
	LUT4 #(
		.INIT('haa80)
	) name3010 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w7058_
	);
	LUT4 #(
		.INIT('h2223)
	) name3011 (
		_w5117_,
		_w5337_,
		_w7057_,
		_w7058_,
		_w7059_
	);
	LUT4 #(
		.INIT('h7500)
	) name3012 (
		_w5117_,
		_w7044_,
		_w7048_,
		_w7059_,
		_w7060_
	);
	LUT4 #(
		.INIT('h2223)
	) name3013 (
		_w5586_,
		_w7040_,
		_w7042_,
		_w7060_,
		_w7061_
	);
	LUT2 #(
		.INIT('h8)
	) name3014 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		_w5234_,
		_w7062_
	);
	LUT2 #(
		.INIT('h9)
	) name3015 (
		_w5239_,
		_w5245_,
		_w7063_
	);
	LUT4 #(
		.INIT('h004f)
	) name3016 (
		_w5193_,
		_w5227_,
		_w5232_,
		_w5249_,
		_w7064_
	);
	LUT3 #(
		.INIT('h36)
	) name3017 (
		_w5273_,
		_w7063_,
		_w7064_,
		_w7065_
	);
	LUT4 #(
		.INIT('hc993)
	) name3018 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w5237_,
		_w5241_,
		_w5302_,
		_w7066_
	);
	LUT4 #(
		.INIT('he0f1)
	) name3019 (
		_w5767_,
		_w5918_,
		_w7065_,
		_w7066_,
		_w7067_
	);
	LUT4 #(
		.INIT('h0200)
	) name3020 (
		\core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w7068_
	);
	LUT4 #(
		.INIT('h0200)
	) name3021 (
		\core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w7069_
	);
	LUT4 #(
		.INIT('h0200)
	) name3022 (
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w7070_
	);
	LUT4 #(
		.INIT('h0200)
	) name3023 (
		\core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w7071_
	);
	LUT3 #(
		.INIT('h01)
	) name3024 (
		_w7070_,
		_w7071_,
		_w7069_,
		_w7072_
	);
	LUT4 #(
		.INIT('h0200)
	) name3025 (
		\core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w7073_
	);
	LUT4 #(
		.INIT('h0200)
	) name3026 (
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w7074_
	);
	LUT4 #(
		.INIT('h0200)
	) name3027 (
		\core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w7075_
	);
	LUT4 #(
		.INIT('h0200)
	) name3028 (
		\core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w7076_
	);
	LUT4 #(
		.INIT('h0001)
	) name3029 (
		_w7073_,
		_w7074_,
		_w7075_,
		_w7076_,
		_w7077_
	);
	LUT4 #(
		.INIT('h45ef)
	) name3030 (
		_w4063_,
		_w7068_,
		_w7072_,
		_w7077_,
		_w7078_
	);
	LUT3 #(
		.INIT('h8c)
	) name3031 (
		_w5117_,
		_w5337_,
		_w7078_,
		_w7079_
	);
	LUT4 #(
		.INIT('h5700)
	) name3032 (
		_w5117_,
		_w7062_,
		_w7067_,
		_w7079_,
		_w7080_
	);
	LUT2 #(
		.INIT('h9)
	) name3033 (
		_w5459_,
		_w5461_,
		_w7081_
	);
	LUT3 #(
		.INIT('he1)
	) name3034 (
		_w5472_,
		_w5484_,
		_w7081_,
		_w7082_
	);
	LUT3 #(
		.INIT('h10)
	) name3035 (
		_w5434_,
		_w6210_,
		_w7082_,
		_w7083_
	);
	LUT4 #(
		.INIT('h08a8)
	) name3036 (
		\core_dag_ilm2reg_I_reg[4]/NET0131 ,
		_w5349_,
		_w5370_,
		_w5417_,
		_w7084_
	);
	LUT3 #(
		.INIT('he1)
	) name3037 (
		_w5408_,
		_w5416_,
		_w5460_,
		_w7085_
	);
	LUT4 #(
		.INIT('h010f)
	) name3038 (
		_w5434_,
		_w6210_,
		_w7084_,
		_w7085_,
		_w7086_
	);
	LUT4 #(
		.INIT('h0200)
	) name3039 (
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w7087_
	);
	LUT4 #(
		.INIT('h0200)
	) name3040 (
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w7088_
	);
	LUT4 #(
		.INIT('h0200)
	) name3041 (
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w7089_
	);
	LUT4 #(
		.INIT('h0200)
	) name3042 (
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w7090_
	);
	LUT4 #(
		.INIT('h0001)
	) name3043 (
		_w7087_,
		_w7088_,
		_w7089_,
		_w7090_,
		_w7091_
	);
	LUT4 #(
		.INIT('h0200)
	) name3044 (
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w7092_
	);
	LUT4 #(
		.INIT('h0200)
	) name3045 (
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w7093_
	);
	LUT4 #(
		.INIT('h0200)
	) name3046 (
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w7094_
	);
	LUT4 #(
		.INIT('h0200)
	) name3047 (
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w7095_
	);
	LUT4 #(
		.INIT('h0001)
	) name3048 (
		_w7092_,
		_w7093_,
		_w7094_,
		_w7095_,
		_w7096_
	);
	LUT3 #(
		.INIT('h1b)
	) name3049 (
		_w4063_,
		_w7091_,
		_w7096_,
		_w7097_
	);
	LUT4 #(
		.INIT('h0123)
	) name3050 (
		_w4063_,
		_w5049_,
		_w7091_,
		_w7096_,
		_w7098_
	);
	LUT4 #(
		.INIT('h0200)
	) name3051 (
		\core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w7099_
	);
	LUT4 #(
		.INIT('h0200)
	) name3052 (
		\core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w7100_
	);
	LUT4 #(
		.INIT('h0200)
	) name3053 (
		\core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w7101_
	);
	LUT4 #(
		.INIT('h0200)
	) name3054 (
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w7102_
	);
	LUT3 #(
		.INIT('h01)
	) name3055 (
		_w7101_,
		_w7102_,
		_w7100_,
		_w7103_
	);
	LUT4 #(
		.INIT('h0200)
	) name3056 (
		\core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w7104_
	);
	LUT4 #(
		.INIT('h0200)
	) name3057 (
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w7105_
	);
	LUT4 #(
		.INIT('h0200)
	) name3058 (
		\core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w7106_
	);
	LUT4 #(
		.INIT('h0200)
	) name3059 (
		\core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w7107_
	);
	LUT4 #(
		.INIT('h0001)
	) name3060 (
		_w7104_,
		_w7105_,
		_w7106_,
		_w7107_,
		_w7108_
	);
	LUT4 #(
		.INIT('h45ef)
	) name3061 (
		_w4063_,
		_w7099_,
		_w7103_,
		_w7108_,
		_w7109_
	);
	LUT4 #(
		.INIT('h0800)
	) name3062 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7110_
	);
	LUT4 #(
		.INIT('h000b)
	) name3063 (
		_w4970_,
		_w7109_,
		_w7110_,
		_w7098_,
		_w7111_
	);
	LUT4 #(
		.INIT('ha222)
	) name3064 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w7112_
	);
	LUT4 #(
		.INIT('h2a00)
	) name3065 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w7113_
	);
	LUT4 #(
		.INIT('h4000)
	) name3066 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[4]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w7114_
	);
	LUT2 #(
		.INIT('h1)
	) name3067 (
		_w7113_,
		_w7114_,
		_w7115_
	);
	LUT2 #(
		.INIT('h4)
	) name3068 (
		_w7112_,
		_w7115_,
		_w7116_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3069 (
		_w5059_,
		_w5539_,
		_w7111_,
		_w7116_,
		_w7117_
	);
	LUT4 #(
		.INIT('haa80)
	) name3070 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w7118_
	);
	LUT4 #(
		.INIT('h2223)
	) name3071 (
		_w5117_,
		_w5337_,
		_w7117_,
		_w7118_,
		_w7119_
	);
	LUT4 #(
		.INIT('h7500)
	) name3072 (
		_w5117_,
		_w7083_,
		_w7086_,
		_w7119_,
		_w7120_
	);
	LUT3 #(
		.INIT('hc9)
	) name3073 (
		_w5162_,
		_w5223_,
		_w5297_,
		_w7121_
	);
	LUT3 #(
		.INIT('h10)
	) name3074 (
		_w5767_,
		_w5918_,
		_w7121_,
		_w7122_
	);
	LUT4 #(
		.INIT('haa80)
	) name3075 (
		\core_dag_ilm1reg_I_reg[4]/NET0131 ,
		_w5125_,
		_w5195_,
		_w5216_,
		_w7123_
	);
	LUT2 #(
		.INIT('h9)
	) name3076 (
		_w5222_,
		_w5224_,
		_w7124_
	);
	LUT2 #(
		.INIT('h9)
	) name3077 (
		_w5193_,
		_w7124_,
		_w7125_
	);
	LUT4 #(
		.INIT('h010f)
	) name3078 (
		_w5767_,
		_w5918_,
		_w7123_,
		_w7125_,
		_w7126_
	);
	LUT3 #(
		.INIT('h20)
	) name3079 (
		_w5337_,
		_w7122_,
		_w7126_,
		_w7127_
	);
	LUT3 #(
		.INIT('ha8)
	) name3080 (
		\DM_rd0[9]_pad ,
		_w5610_,
		_w5612_,
		_w7128_
	);
	LUT4 #(
		.INIT('h135f)
	) name3081 (
		\DM_rdm[9]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w7129_
	);
	LUT4 #(
		.INIT('h135f)
	) name3082 (
		\DM_rd6[9]_pad ,
		\DM_rd7[9]_pad ,
		_w5596_,
		_w5591_,
		_w7130_
	);
	LUT2 #(
		.INIT('h8)
	) name3083 (
		_w7129_,
		_w7130_,
		_w7131_
	);
	LUT3 #(
		.INIT('h80)
	) name3084 (
		\DM_rd4[9]_pad ,
		_w5598_,
		_w5601_,
		_w7132_
	);
	LUT3 #(
		.INIT('h80)
	) name3085 (
		\DM_rd5[9]_pad ,
		_w5598_,
		_w5599_,
		_w7133_
	);
	LUT4 #(
		.INIT('h8000)
	) name3086 (
		\DM_rd2[9]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w7134_
	);
	LUT4 #(
		.INIT('h8000)
	) name3087 (
		\DM_rd1[9]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w7135_
	);
	LUT4 #(
		.INIT('h8000)
	) name3088 (
		\DM_rd3[9]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w7136_
	);
	LUT3 #(
		.INIT('h01)
	) name3089 (
		_w7135_,
		_w7136_,
		_w7134_,
		_w7137_
	);
	LUT3 #(
		.INIT('h10)
	) name3090 (
		_w7133_,
		_w7132_,
		_w7137_,
		_w7138_
	);
	LUT2 #(
		.INIT('h8)
	) name3091 (
		_w7131_,
		_w7138_,
		_w7139_
	);
	LUT2 #(
		.INIT('h4)
	) name3092 (
		_w7128_,
		_w7139_,
		_w7140_
	);
	LUT4 #(
		.INIT('h4000)
	) name3093 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[9]/P0001 ,
		_w7141_
	);
	LUT3 #(
		.INIT('h80)
	) name3094 (
		\bdma_BCTL_reg[9]/NET0131 ,
		_w5627_,
		_w5629_,
		_w7142_
	);
	LUT3 #(
		.INIT('h80)
	) name3095 (
		\tm_tpr_reg_DO_reg[9]/NET0131 ,
		_w5631_,
		_w5635_,
		_w7143_
	);
	LUT3 #(
		.INIT('h80)
	) name3096 (
		\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w5634_,
		_w5635_,
		_w7144_
	);
	LUT3 #(
		.INIT('h80)
	) name3097 (
		\idma_DOVL_reg[9]/NET0131 ,
		_w5804_,
		_w5824_,
		_w7145_
	);
	LUT4 #(
		.INIT('h0001)
	) name3098 (
		_w5795_,
		_w7143_,
		_w7144_,
		_w7145_,
		_w7146_
	);
	LUT4 #(
		.INIT('h8000)
	) name3099 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_txctl_Wcnt_reg[1]/NET0131 ,
		_w5634_,
		_w5660_,
		_w7147_
	);
	LUT4 #(
		.INIT('h8000)
	) name3100 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_txctl_Wcnt_reg[1]/NET0131 ,
		_w5631_,
		_w5639_,
		_w7148_
	);
	LUT2 #(
		.INIT('h1)
	) name3101 (
		_w7147_,
		_w7148_,
		_w7149_
	);
	LUT3 #(
		.INIT('h40)
	) name3102 (
		_w7142_,
		_w7146_,
		_w7149_,
		_w7150_
	);
	LUT3 #(
		.INIT('h80)
	) name3103 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w5629_,
		_w5648_,
		_w7151_
	);
	LUT3 #(
		.INIT('h80)
	) name3104 (
		\bdma_BEAD_reg[9]/NET0131 ,
		_w5629_,
		_w5644_,
		_w7152_
	);
	LUT2 #(
		.INIT('h1)
	) name3105 (
		_w7151_,
		_w7152_,
		_w7153_
	);
	LUT4 #(
		.INIT('h8000)
	) name3106 (
		\bdma_BWCOUNT_reg[9]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w7154_
	);
	LUT4 #(
		.INIT('h8000)
	) name3107 (
		\bdma_BOVL_reg[9]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w7155_
	);
	LUT3 #(
		.INIT('h80)
	) name3108 (
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w5634_,
		_w5637_,
		_w7156_
	);
	LUT3 #(
		.INIT('h80)
	) name3109 (
		\memc_usysr_DO_reg[9]/NET0131 ,
		_w5631_,
		_w5660_,
		_w7157_
	);
	LUT3 #(
		.INIT('h80)
	) name3110 (
		\clkc_ckr_reg_DO_reg[9]/NET0131 ,
		_w5631_,
		_w5644_,
		_w7158_
	);
	LUT3 #(
		.INIT('h80)
	) name3111 (
		\sport1_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w5670_,
		_w5810_,
		_w7159_
	);
	LUT4 #(
		.INIT('h0001)
	) name3112 (
		_w7156_,
		_w7157_,
		_w7158_,
		_w7159_,
		_w7160_
	);
	LUT3 #(
		.INIT('h80)
	) name3113 (
		\sport0_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w5627_,
		_w5634_,
		_w7161_
	);
	LUT3 #(
		.INIT('h80)
	) name3114 (
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w5634_,
		_w5639_,
		_w7162_
	);
	LUT3 #(
		.INIT('h80)
	) name3115 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w5628_,
		_w5639_,
		_w7163_
	);
	LUT3 #(
		.INIT('h80)
	) name3116 (
		\ITFS0_pad ,
		_w5632_,
		_w5634_,
		_w7164_
	);
	LUT4 #(
		.INIT('h0001)
	) name3117 (
		_w7161_,
		_w7162_,
		_w7163_,
		_w7164_,
		_w7165_
	);
	LUT3 #(
		.INIT('h80)
	) name3118 (
		\emc_WSCRreg_DO_reg[9]/NET0131 ,
		_w5631_,
		_w5632_,
		_w7166_
	);
	LUT3 #(
		.INIT('h80)
	) name3119 (
		\ITFS1_pad ,
		_w5644_,
		_w5634_,
		_w7167_
	);
	LUT3 #(
		.INIT('h80)
	) name3120 (
		\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w5648_,
		_w5634_,
		_w7168_
	);
	LUT3 #(
		.INIT('h80)
	) name3121 (
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w5631_,
		_w5637_,
		_w7169_
	);
	LUT4 #(
		.INIT('h0001)
	) name3122 (
		_w7166_,
		_w7167_,
		_w7168_,
		_w7169_,
		_w7170_
	);
	LUT4 #(
		.INIT('h4000)
	) name3123 (
		_w7155_,
		_w7160_,
		_w7165_,
		_w7170_,
		_w7171_
	);
	LUT4 #(
		.INIT('h4000)
	) name3124 (
		_w7154_,
		_w7150_,
		_w7153_,
		_w7171_,
		_w7172_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3125 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4224_,
		_w4221_,
		_w4229_,
		_w7173_
	);
	LUT3 #(
		.INIT('ha8)
	) name3126 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w7174_
	);
	LUT2 #(
		.INIT('h8)
	) name3127 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w7175_
	);
	LUT4 #(
		.INIT('h153f)
	) name3128 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w7176_
	);
	LUT3 #(
		.INIT('h10)
	) name3129 (
		_w7174_,
		_w7175_,
		_w7176_,
		_w7177_
	);
	LUT3 #(
		.INIT('h8a)
	) name3130 (
		_w5681_,
		_w7173_,
		_w7177_,
		_w7178_
	);
	LUT4 #(
		.INIT('h135f)
	) name3131 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131 ,
		_w7179_
	);
	LUT4 #(
		.INIT('h135f)
	) name3132 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131 ,
		_w7180_
	);
	LUT2 #(
		.INIT('h8)
	) name3133 (
		_w7179_,
		_w7180_,
		_w7181_
	);
	LUT4 #(
		.INIT('h135f)
	) name3134 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		_w7182_
	);
	LUT4 #(
		.INIT('h135f)
	) name3135 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131 ,
		_w7183_
	);
	LUT4 #(
		.INIT('h135f)
	) name3136 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131 ,
		_w7184_
	);
	LUT4 #(
		.INIT('h135f)
	) name3137 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131 ,
		_w7185_
	);
	LUT4 #(
		.INIT('h8000)
	) name3138 (
		_w7184_,
		_w7185_,
		_w7182_,
		_w7183_,
		_w7186_
	);
	LUT3 #(
		.INIT('h2a)
	) name3139 (
		_w5687_,
		_w7181_,
		_w7186_,
		_w7187_
	);
	LUT4 #(
		.INIT('h135f)
	) name3140 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 ,
		_w7188_
	);
	LUT4 #(
		.INIT('h135f)
	) name3141 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131 ,
		_w7189_
	);
	LUT2 #(
		.INIT('h8)
	) name3142 (
		_w7188_,
		_w7189_,
		_w7190_
	);
	LUT4 #(
		.INIT('h135f)
	) name3143 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131 ,
		_w7191_
	);
	LUT4 #(
		.INIT('h135f)
	) name3144 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131 ,
		_w7192_
	);
	LUT4 #(
		.INIT('h135f)
	) name3145 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131 ,
		_w7193_
	);
	LUT4 #(
		.INIT('h135f)
	) name3146 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131 ,
		_w7194_
	);
	LUT4 #(
		.INIT('h8000)
	) name3147 (
		_w7193_,
		_w7194_,
		_w7191_,
		_w7192_,
		_w7195_
	);
	LUT4 #(
		.INIT('h135f)
	) name3148 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[9]/P0001 ,
		\sport1_txctl_TX_reg[9]/P0001 ,
		_w7196_
	);
	LUT4 #(
		.INIT('h135f)
	) name3149 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[9]/P0001 ,
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w7197_
	);
	LUT3 #(
		.INIT('h2a)
	) name3150 (
		_w5706_,
		_w7196_,
		_w7197_,
		_w7198_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3151 (
		_w5697_,
		_w7190_,
		_w7195_,
		_w7198_,
		_w7199_
	);
	LUT2 #(
		.INIT('h4)
	) name3152 (
		_w7187_,
		_w7199_,
		_w7200_
	);
	LUT3 #(
		.INIT('h1b)
	) name3153 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001 ,
		_w7201_
	);
	LUT4 #(
		.INIT('ha820)
	) name3154 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001 ,
		_w7202_
	);
	LUT3 #(
		.INIT('h1b)
	) name3155 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001 ,
		_w7203_
	);
	LUT4 #(
		.INIT('ha820)
	) name3156 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001 ,
		_w7204_
	);
	LUT3 #(
		.INIT('h1b)
	) name3157 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001 ,
		_w7205_
	);
	LUT4 #(
		.INIT('ha820)
	) name3158 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001 ,
		_w7206_
	);
	LUT3 #(
		.INIT('h01)
	) name3159 (
		_w7204_,
		_w7206_,
		_w7202_,
		_w7207_
	);
	LUT3 #(
		.INIT('h2a)
	) name3160 (
		_w5741_,
		_w5746_,
		_w7207_,
		_w7208_
	);
	LUT3 #(
		.INIT('h1b)
	) name3161 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001 ,
		_w7209_
	);
	LUT4 #(
		.INIT('ha820)
	) name3162 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001 ,
		_w7210_
	);
	LUT3 #(
		.INIT('h1b)
	) name3163 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001 ,
		_w7211_
	);
	LUT4 #(
		.INIT('ha820)
	) name3164 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001 ,
		_w7212_
	);
	LUT3 #(
		.INIT('h1b)
	) name3165 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001 ,
		_w7213_
	);
	LUT4 #(
		.INIT('ha820)
	) name3166 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001 ,
		_w7214_
	);
	LUT3 #(
		.INIT('h01)
	) name3167 (
		_w7212_,
		_w7214_,
		_w7210_,
		_w7215_
	);
	LUT3 #(
		.INIT('h1b)
	) name3168 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 ,
		_w7216_
	);
	LUT4 #(
		.INIT('ha820)
	) name3169 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 ,
		_w7217_
	);
	LUT3 #(
		.INIT('h1b)
	) name3170 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001 ,
		_w7218_
	);
	LUT4 #(
		.INIT('ha820)
	) name3171 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001 ,
		_w7219_
	);
	LUT3 #(
		.INIT('h1b)
	) name3172 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001 ,
		_w7220_
	);
	LUT4 #(
		.INIT('ha820)
	) name3173 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001 ,
		_w7221_
	);
	LUT4 #(
		.INIT('h0001)
	) name3174 (
		_w5714_,
		_w7217_,
		_w7219_,
		_w7221_,
		_w7222_
	);
	LUT3 #(
		.INIT('h2a)
	) name3175 (
		_w5712_,
		_w7215_,
		_w7222_,
		_w7223_
	);
	LUT3 #(
		.INIT('h1b)
	) name3176 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001 ,
		_w7224_
	);
	LUT4 #(
		.INIT('ha820)
	) name3177 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001 ,
		_w7225_
	);
	LUT4 #(
		.INIT('ha820)
	) name3178 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001 ,
		_w7226_
	);
	LUT2 #(
		.INIT('h1)
	) name3179 (
		_w7225_,
		_w7226_,
		_w7227_
	);
	LUT3 #(
		.INIT('h1b)
	) name3180 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001 ,
		_w7228_
	);
	LUT4 #(
		.INIT('ha820)
	) name3181 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001 ,
		_w7229_
	);
	LUT3 #(
		.INIT('h1b)
	) name3182 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001 ,
		_w7230_
	);
	LUT4 #(
		.INIT('ha820)
	) name3183 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001 ,
		_w7231_
	);
	LUT4 #(
		.INIT('ha820)
	) name3184 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001 ,
		_w7232_
	);
	LUT3 #(
		.INIT('h01)
	) name3185 (
		_w7231_,
		_w7232_,
		_w7229_,
		_w7233_
	);
	LUT3 #(
		.INIT('h2a)
	) name3186 (
		_w5730_,
		_w7227_,
		_w7233_,
		_w7234_
	);
	LUT3 #(
		.INIT('h01)
	) name3187 (
		_w7223_,
		_w7234_,
		_w7208_,
		_w7235_
	);
	LUT2 #(
		.INIT('h8)
	) name3188 (
		_w7200_,
		_w7235_,
		_w7236_
	);
	LUT4 #(
		.INIT('h3100)
	) name3189 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w7178_,
		_w7172_,
		_w7236_,
		_w7237_
	);
	LUT2 #(
		.INIT('h8)
	) name3190 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[9]/P0001 ,
		_w7238_
	);
	LUT3 #(
		.INIT('h08)
	) name3191 (
		_w5588_,
		_w5598_,
		_w7238_,
		_w7239_
	);
	LUT4 #(
		.INIT('hba00)
	) name3192 (
		\emc_DMDoe_reg/NET0131 ,
		_w7141_,
		_w7237_,
		_w7239_,
		_w7240_
	);
	LUT2 #(
		.INIT('h1)
	) name3193 (
		_w7140_,
		_w7240_,
		_w7241_
	);
	LUT3 #(
		.INIT('h54)
	) name3194 (
		_w5117_,
		_w5337_,
		_w7241_,
		_w7242_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3195 (
		_w5337_,
		_w7122_,
		_w7126_,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('h1)
	) name3196 (
		_w7109_,
		_w7097_,
		_w7244_
	);
	LUT3 #(
		.INIT('ha8)
	) name3197 (
		\DM_rd0[4]_pad ,
		_w5610_,
		_w5612_,
		_w7245_
	);
	LUT4 #(
		.INIT('h135f)
	) name3198 (
		\DM_rdm[4]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w7246_
	);
	LUT4 #(
		.INIT('h135f)
	) name3199 (
		\DM_rd6[4]_pad ,
		\DM_rd7[4]_pad ,
		_w5596_,
		_w5591_,
		_w7247_
	);
	LUT2 #(
		.INIT('h8)
	) name3200 (
		_w7246_,
		_w7247_,
		_w7248_
	);
	LUT3 #(
		.INIT('h80)
	) name3201 (
		\DM_rd5[4]_pad ,
		_w5598_,
		_w5599_,
		_w7249_
	);
	LUT3 #(
		.INIT('h80)
	) name3202 (
		\DM_rd4[4]_pad ,
		_w5598_,
		_w5601_,
		_w7250_
	);
	LUT4 #(
		.INIT('h8000)
	) name3203 (
		\DM_rd2[4]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w7251_
	);
	LUT4 #(
		.INIT('h8000)
	) name3204 (
		\DM_rd1[4]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w7252_
	);
	LUT4 #(
		.INIT('h8000)
	) name3205 (
		\DM_rd3[4]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w7253_
	);
	LUT3 #(
		.INIT('h01)
	) name3206 (
		_w7252_,
		_w7253_,
		_w7251_,
		_w7254_
	);
	LUT3 #(
		.INIT('h10)
	) name3207 (
		_w7250_,
		_w7249_,
		_w7254_,
		_w7255_
	);
	LUT2 #(
		.INIT('h8)
	) name3208 (
		_w7248_,
		_w7255_,
		_w7256_
	);
	LUT2 #(
		.INIT('h4)
	) name3209 (
		_w7245_,
		_w7256_,
		_w7257_
	);
	LUT4 #(
		.INIT('h4000)
	) name3210 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[4]/P0001 ,
		_w7258_
	);
	LUT3 #(
		.INIT('h80)
	) name3211 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w5629_,
		_w5648_,
		_w7259_
	);
	LUT3 #(
		.INIT('h80)
	) name3212 (
		\emc_WSCRreg_DO_reg[4]/NET0131 ,
		_w5631_,
		_w5632_,
		_w7260_
	);
	LUT3 #(
		.INIT('h80)
	) name3213 (
		\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w5634_,
		_w5635_,
		_w7261_
	);
	LUT3 #(
		.INIT('h80)
	) name3214 (
		\sport1_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w5631_,
		_w5639_,
		_w7262_
	);
	LUT3 #(
		.INIT('h80)
	) name3215 (
		\tm_tsr_reg_DO_reg[4]/NET0131 ,
		_w5627_,
		_w5631_,
		_w7263_
	);
	LUT4 #(
		.INIT('h0001)
	) name3216 (
		_w7260_,
		_w7261_,
		_w7262_,
		_w7263_,
		_w7264_
	);
	LUT3 #(
		.INIT('h80)
	) name3217 (
		\idma_DOVL_reg[4]/NET0131 ,
		_w5804_,
		_w5824_,
		_w7265_
	);
	LUT3 #(
		.INIT('h80)
	) name3218 (
		\sport0_regs_AUTOreg_DO_reg[4]/NET0131 ,
		_w5627_,
		_w5634_,
		_w7266_
	);
	LUT3 #(
		.INIT('h80)
	) name3219 (
		\tm_tpr_reg_DO_reg[4]/NET0131 ,
		_w5631_,
		_w5635_,
		_w7267_
	);
	LUT4 #(
		.INIT('h0001)
	) name3220 (
		_w5795_,
		_w7265_,
		_w7266_,
		_w7267_,
		_w7268_
	);
	LUT3 #(
		.INIT('h40)
	) name3221 (
		_w7259_,
		_w7264_,
		_w7268_,
		_w7269_
	);
	LUT3 #(
		.INIT('h80)
	) name3222 (
		\bdma_BEAD_reg[4]/NET0131 ,
		_w5629_,
		_w5644_,
		_w7270_
	);
	LUT3 #(
		.INIT('h80)
	) name3223 (
		\bdma_BCTL_reg[4]/NET0131 ,
		_w5627_,
		_w5629_,
		_w7271_
	);
	LUT2 #(
		.INIT('h1)
	) name3224 (
		_w7270_,
		_w7271_,
		_w7272_
	);
	LUT2 #(
		.INIT('h8)
	) name3225 (
		_w7269_,
		_w7272_,
		_w7273_
	);
	LUT4 #(
		.INIT('h8000)
	) name3226 (
		\bdma_BOVL_reg[4]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w7274_
	);
	LUT4 #(
		.INIT('h8000)
	) name3227 (
		\bdma_BWCOUNT_reg[4]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w7275_
	);
	LUT3 #(
		.INIT('h80)
	) name3228 (
		\pio_pmask_reg_DO_reg[4]/NET0131 ,
		_w5628_,
		_w5660_,
		_w7276_
	);
	LUT3 #(
		.INIT('h80)
	) name3229 (
		\sport0_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w5634_,
		_w5660_,
		_w7277_
	);
	LUT3 #(
		.INIT('h80)
	) name3230 (
		\sport1_regs_AUTOreg_DO_reg[4]/NET0131 ,
		_w5670_,
		_w5810_,
		_w7278_
	);
	LUT3 #(
		.INIT('h80)
	) name3231 (
		\tm_TCR_TMP_reg[4]/NET0131 ,
		_w5631_,
		_w5637_,
		_w7279_
	);
	LUT4 #(
		.INIT('h0001)
	) name3232 (
		_w7276_,
		_w7277_,
		_w7278_,
		_w7279_,
		_w7280_
	);
	LUT3 #(
		.INIT('h80)
	) name3233 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w5632_,
		_w5634_,
		_w7281_
	);
	LUT3 #(
		.INIT('h80)
	) name3234 (
		\emc_WSCRext_reg_DO_reg[4]/NET0131 ,
		_w5670_,
		_w5790_,
		_w7282_
	);
	LUT3 #(
		.INIT('h80)
	) name3235 (
		\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w5648_,
		_w5634_,
		_w7283_
	);
	LUT3 #(
		.INIT('h80)
	) name3236 (
		\sport1_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w5644_,
		_w5634_,
		_w7284_
	);
	LUT4 #(
		.INIT('h0001)
	) name3237 (
		_w7281_,
		_w7282_,
		_w7283_,
		_w7284_,
		_w7285_
	);
	LUT3 #(
		.INIT('h80)
	) name3238 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w5628_,
		_w5639_,
		_w7286_
	);
	LUT3 #(
		.INIT('h80)
	) name3239 (
		\PIO_out[4]_pad ,
		_w5628_,
		_w5635_,
		_w7287_
	);
	LUT3 #(
		.INIT('h80)
	) name3240 (
		\PIO_oe[4]_pad ,
		_w5628_,
		_w5632_,
		_w7288_
	);
	LUT3 #(
		.INIT('h80)
	) name3241 (
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w5634_,
		_w5639_,
		_w7289_
	);
	LUT4 #(
		.INIT('h0001)
	) name3242 (
		_w7286_,
		_w7287_,
		_w7288_,
		_w7289_,
		_w7290_
	);
	LUT3 #(
		.INIT('h80)
	) name3243 (
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w5634_,
		_w5637_,
		_w7291_
	);
	LUT3 #(
		.INIT('h80)
	) name3244 (
		\clkc_ckr_reg_DO_reg[4]/NET0131 ,
		_w5631_,
		_w5644_,
		_w7292_
	);
	LUT3 #(
		.INIT('h80)
	) name3245 (
		\memc_usysr_DO_reg[4]/NET0131 ,
		_w5631_,
		_w5660_,
		_w7293_
	);
	LUT3 #(
		.INIT('h80)
	) name3246 (
		\pio_PINT_reg[4]/NET0131 ,
		_w5670_,
		_w5672_,
		_w7294_
	);
	LUT4 #(
		.INIT('h0001)
	) name3247 (
		_w7291_,
		_w7292_,
		_w7293_,
		_w7294_,
		_w7295_
	);
	LUT4 #(
		.INIT('h8000)
	) name3248 (
		_w7290_,
		_w7295_,
		_w7280_,
		_w7285_,
		_w7296_
	);
	LUT3 #(
		.INIT('h10)
	) name3249 (
		_w7275_,
		_w7274_,
		_w7296_,
		_w7297_
	);
	LUT3 #(
		.INIT('h2a)
	) name3250 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w7273_,
		_w7297_,
		_w7298_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3251 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4197_,
		_w4194_,
		_w4202_,
		_w7299_
	);
	LUT2 #(
		.INIT('h8)
	) name3252 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[4]/NET0131 ,
		_w7300_
	);
	LUT4 #(
		.INIT('h135f)
	) name3253 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		_w7301_
	);
	LUT2 #(
		.INIT('h4)
	) name3254 (
		_w7300_,
		_w7301_,
		_w7302_
	);
	LUT3 #(
		.INIT('ha8)
	) name3255 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w7303_
	);
	LUT4 #(
		.INIT('h135f)
	) name3256 (
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w7304_
	);
	LUT4 #(
		.INIT('h135f)
	) name3257 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w7305_
	);
	LUT3 #(
		.INIT('h40)
	) name3258 (
		_w7303_,
		_w7304_,
		_w7305_,
		_w7306_
	);
	LUT2 #(
		.INIT('h8)
	) name3259 (
		_w7302_,
		_w7306_,
		_w7307_
	);
	LUT3 #(
		.INIT('h8a)
	) name3260 (
		_w5681_,
		_w7299_,
		_w7307_,
		_w7308_
	);
	LUT4 #(
		.INIT('h135f)
	) name3261 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131 ,
		_w7309_
	);
	LUT4 #(
		.INIT('h135f)
	) name3262 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131 ,
		_w7310_
	);
	LUT2 #(
		.INIT('h8)
	) name3263 (
		_w7309_,
		_w7310_,
		_w7311_
	);
	LUT4 #(
		.INIT('h135f)
	) name3264 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131 ,
		_w7312_
	);
	LUT4 #(
		.INIT('h135f)
	) name3265 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w7313_
	);
	LUT4 #(
		.INIT('h135f)
	) name3266 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w7314_
	);
	LUT4 #(
		.INIT('h135f)
	) name3267 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131 ,
		_w7315_
	);
	LUT4 #(
		.INIT('h8000)
	) name3268 (
		_w7314_,
		_w7315_,
		_w7312_,
		_w7313_,
		_w7316_
	);
	LUT3 #(
		.INIT('h2a)
	) name3269 (
		_w5687_,
		_w7311_,
		_w7316_,
		_w7317_
	);
	LUT4 #(
		.INIT('h135f)
	) name3270 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 ,
		_w7318_
	);
	LUT4 #(
		.INIT('h135f)
	) name3271 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w7319_
	);
	LUT2 #(
		.INIT('h8)
	) name3272 (
		_w7318_,
		_w7319_,
		_w7320_
	);
	LUT4 #(
		.INIT('h135f)
	) name3273 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131 ,
		_w7321_
	);
	LUT4 #(
		.INIT('h135f)
	) name3274 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131 ,
		_w7322_
	);
	LUT4 #(
		.INIT('h135f)
	) name3275 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131 ,
		_w7323_
	);
	LUT4 #(
		.INIT('h135f)
	) name3276 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131 ,
		_w7324_
	);
	LUT4 #(
		.INIT('h8000)
	) name3277 (
		_w7323_,
		_w7324_,
		_w7321_,
		_w7322_,
		_w7325_
	);
	LUT4 #(
		.INIT('h135f)
	) name3278 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[4]/P0001 ,
		\sport1_txctl_TX_reg[4]/P0001 ,
		_w7326_
	);
	LUT4 #(
		.INIT('h135f)
	) name3279 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport1_rxctl_RX_reg[4]/P0001 ,
		_w7327_
	);
	LUT3 #(
		.INIT('h2a)
	) name3280 (
		_w5706_,
		_w7326_,
		_w7327_,
		_w7328_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3281 (
		_w5697_,
		_w7320_,
		_w7325_,
		_w7328_,
		_w7329_
	);
	LUT2 #(
		.INIT('h4)
	) name3282 (
		_w7317_,
		_w7329_,
		_w7330_
	);
	LUT3 #(
		.INIT('h1b)
	) name3283 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001 ,
		_w7331_
	);
	LUT4 #(
		.INIT('ha820)
	) name3284 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001 ,
		_w7332_
	);
	LUT2 #(
		.INIT('h1)
	) name3285 (
		_w5743_,
		_w7332_,
		_w7333_
	);
	LUT3 #(
		.INIT('h1b)
	) name3286 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001 ,
		_w7334_
	);
	LUT4 #(
		.INIT('ha820)
	) name3287 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001 ,
		_w7335_
	);
	LUT3 #(
		.INIT('h1b)
	) name3288 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001 ,
		_w7336_
	);
	LUT4 #(
		.INIT('ha820)
	) name3289 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001 ,
		_w7337_
	);
	LUT3 #(
		.INIT('h1b)
	) name3290 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001 ,
		_w7338_
	);
	LUT4 #(
		.INIT('ha820)
	) name3291 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001 ,
		_w7339_
	);
	LUT3 #(
		.INIT('h01)
	) name3292 (
		_w7337_,
		_w7339_,
		_w7335_,
		_w7340_
	);
	LUT3 #(
		.INIT('h2a)
	) name3293 (
		_w5741_,
		_w7333_,
		_w7340_,
		_w7341_
	);
	LUT3 #(
		.INIT('h1b)
	) name3294 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001 ,
		_w7342_
	);
	LUT4 #(
		.INIT('ha820)
	) name3295 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001 ,
		_w7343_
	);
	LUT3 #(
		.INIT('h1b)
	) name3296 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001 ,
		_w7344_
	);
	LUT4 #(
		.INIT('ha820)
	) name3297 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001 ,
		_w7345_
	);
	LUT3 #(
		.INIT('h1b)
	) name3298 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001 ,
		_w7346_
	);
	LUT4 #(
		.INIT('ha820)
	) name3299 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001 ,
		_w7347_
	);
	LUT3 #(
		.INIT('h01)
	) name3300 (
		_w7345_,
		_w7347_,
		_w7343_,
		_w7348_
	);
	LUT3 #(
		.INIT('h1b)
	) name3301 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 ,
		_w7349_
	);
	LUT4 #(
		.INIT('ha820)
	) name3302 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 ,
		_w7350_
	);
	LUT3 #(
		.INIT('h1b)
	) name3303 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001 ,
		_w7351_
	);
	LUT4 #(
		.INIT('ha820)
	) name3304 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001 ,
		_w7352_
	);
	LUT3 #(
		.INIT('h1b)
	) name3305 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001 ,
		_w7353_
	);
	LUT4 #(
		.INIT('ha820)
	) name3306 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001 ,
		_w7354_
	);
	LUT3 #(
		.INIT('h1b)
	) name3307 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001 ,
		_w7355_
	);
	LUT4 #(
		.INIT('ha820)
	) name3308 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001 ,
		_w7356_
	);
	LUT4 #(
		.INIT('h0001)
	) name3309 (
		_w7350_,
		_w7352_,
		_w7354_,
		_w7356_,
		_w7357_
	);
	LUT3 #(
		.INIT('h2a)
	) name3310 (
		_w5712_,
		_w7348_,
		_w7357_,
		_w7358_
	);
	LUT3 #(
		.INIT('h1b)
	) name3311 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001 ,
		_w7359_
	);
	LUT4 #(
		.INIT('ha820)
	) name3312 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001 ,
		_w7360_
	);
	LUT2 #(
		.INIT('h8)
	) name3313 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w7361_
	);
	LUT2 #(
		.INIT('h1)
	) name3314 (
		_w7360_,
		_w7361_,
		_w7362_
	);
	LUT3 #(
		.INIT('h1b)
	) name3315 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001 ,
		_w7363_
	);
	LUT4 #(
		.INIT('ha820)
	) name3316 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001 ,
		_w7364_
	);
	LUT3 #(
		.INIT('h1b)
	) name3317 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001 ,
		_w7365_
	);
	LUT4 #(
		.INIT('ha820)
	) name3318 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001 ,
		_w7366_
	);
	LUT4 #(
		.INIT('ha820)
	) name3319 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001 ,
		_w7367_
	);
	LUT4 #(
		.INIT('ha820)
	) name3320 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001 ,
		_w7368_
	);
	LUT4 #(
		.INIT('h0001)
	) name3321 (
		_w7364_,
		_w7366_,
		_w7367_,
		_w7368_,
		_w7369_
	);
	LUT3 #(
		.INIT('h2a)
	) name3322 (
		_w5730_,
		_w7362_,
		_w7369_,
		_w7370_
	);
	LUT3 #(
		.INIT('h01)
	) name3323 (
		_w7358_,
		_w7370_,
		_w7341_,
		_w7371_
	);
	LUT2 #(
		.INIT('h8)
	) name3324 (
		_w7330_,
		_w7371_,
		_w7372_
	);
	LUT2 #(
		.INIT('h4)
	) name3325 (
		_w7308_,
		_w7372_,
		_w7373_
	);
	LUT3 #(
		.INIT('h10)
	) name3326 (
		_w7258_,
		_w7298_,
		_w7373_,
		_w7374_
	);
	LUT4 #(
		.INIT('h5455)
	) name3327 (
		\emc_DMDoe_reg/NET0131 ,
		_w7258_,
		_w7298_,
		_w7373_,
		_w7375_
	);
	LUT2 #(
		.INIT('h8)
	) name3328 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[4]/P0001 ,
		_w7376_
	);
	LUT3 #(
		.INIT('h08)
	) name3329 (
		_w5588_,
		_w5598_,
		_w7376_,
		_w7377_
	);
	LUT3 #(
		.INIT('h45)
	) name3330 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w7378_
	);
	LUT4 #(
		.INIT('h80a2)
	) name3331 (
		_w5117_,
		_w5337_,
		_w7378_,
		_w7244_,
		_w7379_
	);
	LUT2 #(
		.INIT('h2)
	) name3332 (
		_w5586_,
		_w7379_,
		_w7380_
	);
	LUT2 #(
		.INIT('h4)
	) name3333 (
		_w7243_,
		_w7380_,
		_w7381_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3334 (
		_w5586_,
		_w7080_,
		_w7120_,
		_w7381_,
		_w7382_
	);
	LUT2 #(
		.INIT('h9)
	) name3335 (
		_w5455_,
		_w5457_,
		_w7383_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3336 (
		_w5462_,
		_w5472_,
		_w5484_,
		_w5485_,
		_w7384_
	);
	LUT2 #(
		.INIT('h6)
	) name3337 (
		_w7383_,
		_w7384_,
		_w7385_
	);
	LUT3 #(
		.INIT('h10)
	) name3338 (
		_w5434_,
		_w6210_,
		_w7385_,
		_w7386_
	);
	LUT2 #(
		.INIT('h8)
	) name3339 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		_w5418_,
		_w7387_
	);
	LUT4 #(
		.INIT('hab02)
	) name3340 (
		\core_dag_ilm2reg_M_reg[4]/NET0131 ,
		_w5408_,
		_w5416_,
		_w5421_,
		_w7388_
	);
	LUT2 #(
		.INIT('h6)
	) name3341 (
		_w5456_,
		_w7388_,
		_w7389_
	);
	LUT4 #(
		.INIT('h010f)
	) name3342 (
		_w5434_,
		_w6210_,
		_w7387_,
		_w7389_,
		_w7390_
	);
	LUT2 #(
		.INIT('h9)
	) name3343 (
		_w5246_,
		_w5248_,
		_w7391_
	);
	LUT4 #(
		.INIT('hb04f)
	) name3344 (
		_w5193_,
		_w5227_,
		_w5232_,
		_w7391_,
		_w7392_
	);
	LUT4 #(
		.INIT('h0065)
	) name3345 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w7392_,
		_w7393_
	);
	LUT2 #(
		.INIT('h9)
	) name3346 (
		_w5247_,
		_w5302_,
		_w7394_
	);
	LUT4 #(
		.INIT('h9a00)
	) name3347 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w7394_,
		_w7395_
	);
	LUT3 #(
		.INIT('h01)
	) name3348 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w7395_,
		_w7393_,
		_w7396_
	);
	LUT4 #(
		.INIT('h008a)
	) name3349 (
		\core_dag_ilm1reg_I_reg[8]/NET0131 ,
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		_w5153_,
		_w5240_,
		_w7397_
	);
	LUT3 #(
		.INIT('h0e)
	) name3350 (
		_w5767_,
		_w5768_,
		_w7392_,
		_w7398_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3351 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5155_,
		_w5310_,
		_w7394_,
		_w7399_
	);
	LUT4 #(
		.INIT('h0045)
	) name3352 (
		_w7397_,
		_w7398_,
		_w7399_,
		_w7396_,
		_w7400_
	);
	LUT4 #(
		.INIT('h45ef)
	) name3353 (
		_w5337_,
		_w7386_,
		_w7390_,
		_w7400_,
		_w7401_
	);
	LUT4 #(
		.INIT('h0200)
	) name3354 (
		\core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w7402_
	);
	LUT4 #(
		.INIT('h0200)
	) name3355 (
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w7403_
	);
	LUT3 #(
		.INIT('h02)
	) name3356 (
		\core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 ,
		_w5061_,
		_w5065_,
		_w7404_
	);
	LUT4 #(
		.INIT('h0200)
	) name3357 (
		\core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w7405_
	);
	LUT3 #(
		.INIT('h02)
	) name3358 (
		\core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 ,
		_w5070_,
		_w5073_,
		_w7406_
	);
	LUT4 #(
		.INIT('h0200)
	) name3359 (
		\core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w7407_
	);
	LUT3 #(
		.INIT('h01)
	) name3360 (
		_w7405_,
		_w7407_,
		_w7403_,
		_w7408_
	);
	LUT4 #(
		.INIT('h0200)
	) name3361 (
		\core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w7409_
	);
	LUT4 #(
		.INIT('h0200)
	) name3362 (
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w7410_
	);
	LUT4 #(
		.INIT('h0200)
	) name3363 (
		\core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w7411_
	);
	LUT4 #(
		.INIT('h0200)
	) name3364 (
		\core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w7412_
	);
	LUT4 #(
		.INIT('h0001)
	) name3365 (
		_w7409_,
		_w7410_,
		_w7411_,
		_w7412_,
		_w7413_
	);
	LUT4 #(
		.INIT('h45ef)
	) name3366 (
		_w4063_,
		_w7402_,
		_w7408_,
		_w7413_,
		_w7414_
	);
	LUT4 #(
		.INIT('h0200)
	) name3367 (
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w7415_
	);
	LUT4 #(
		.INIT('h0200)
	) name3368 (
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w7416_
	);
	LUT4 #(
		.INIT('h0200)
	) name3369 (
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w7417_
	);
	LUT4 #(
		.INIT('h0200)
	) name3370 (
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w7418_
	);
	LUT4 #(
		.INIT('h0001)
	) name3371 (
		_w7415_,
		_w7416_,
		_w7417_,
		_w7418_,
		_w7419_
	);
	LUT4 #(
		.INIT('h0200)
	) name3372 (
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w7420_
	);
	LUT4 #(
		.INIT('h0200)
	) name3373 (
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w7421_
	);
	LUT4 #(
		.INIT('h0200)
	) name3374 (
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w7422_
	);
	LUT4 #(
		.INIT('h0200)
	) name3375 (
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w7423_
	);
	LUT4 #(
		.INIT('h0001)
	) name3376 (
		_w7420_,
		_w7421_,
		_w7422_,
		_w7423_,
		_w7424_
	);
	LUT3 #(
		.INIT('hd0)
	) name3377 (
		_w4063_,
		_w7419_,
		_w7424_,
		_w7425_
	);
	LUT4 #(
		.INIT('h0233)
	) name3378 (
		_w4063_,
		_w5049_,
		_w7419_,
		_w7424_,
		_w7426_
	);
	LUT4 #(
		.INIT('h0800)
	) name3379 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w7427_
	);
	LUT4 #(
		.INIT('h0203)
	) name3380 (
		_w4970_,
		_w7426_,
		_w7427_,
		_w7414_,
		_w7428_
	);
	LUT4 #(
		.INIT('ha222)
	) name3381 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w7429_
	);
	LUT4 #(
		.INIT('h2a00)
	) name3382 (
		\idma_DCTL_reg[5]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w7430_
	);
	LUT4 #(
		.INIT('h4000)
	) name3383 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w7431_
	);
	LUT2 #(
		.INIT('h1)
	) name3384 (
		_w7430_,
		_w7431_,
		_w7432_
	);
	LUT3 #(
		.INIT('h20)
	) name3385 (
		_w5539_,
		_w7429_,
		_w7432_,
		_w7433_
	);
	LUT3 #(
		.INIT('hd0)
	) name3386 (
		_w5059_,
		_w7428_,
		_w7433_,
		_w7434_
	);
	LUT4 #(
		.INIT('h5540)
	) name3387 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w7435_
	);
	LUT3 #(
		.INIT('h01)
	) name3388 (
		_w5337_,
		_w7435_,
		_w7434_,
		_w7436_
	);
	LUT3 #(
		.INIT('h02)
	) name3389 (
		\core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 ,
		_w5070_,
		_w5073_,
		_w7437_
	);
	LUT4 #(
		.INIT('h0200)
	) name3390 (
		\core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w7438_
	);
	LUT3 #(
		.INIT('h02)
	) name3391 (
		\core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131 ,
		_w5079_,
		_w5082_,
		_w7439_
	);
	LUT4 #(
		.INIT('h0200)
	) name3392 (
		\core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w7440_
	);
	LUT4 #(
		.INIT('h0200)
	) name3393 (
		\core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w7441_
	);
	LUT4 #(
		.INIT('h0200)
	) name3394 (
		\core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w7442_
	);
	LUT3 #(
		.INIT('h01)
	) name3395 (
		_w7441_,
		_w7442_,
		_w7440_,
		_w7443_
	);
	LUT4 #(
		.INIT('h0200)
	) name3396 (
		\core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w7444_
	);
	LUT4 #(
		.INIT('h0200)
	) name3397 (
		\core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w7445_
	);
	LUT4 #(
		.INIT('h0200)
	) name3398 (
		\core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w7446_
	);
	LUT4 #(
		.INIT('h0200)
	) name3399 (
		\core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w7447_
	);
	LUT4 #(
		.INIT('h0001)
	) name3400 (
		_w7444_,
		_w7445_,
		_w7446_,
		_w7447_,
		_w7448_
	);
	LUT4 #(
		.INIT('h45ef)
	) name3401 (
		_w4063_,
		_w7438_,
		_w7443_,
		_w7448_,
		_w7449_
	);
	LUT3 #(
		.INIT('h15)
	) name3402 (
		_w5117_,
		_w5337_,
		_w7449_,
		_w7450_
	);
	LUT3 #(
		.INIT('h45)
	) name3403 (
		_w5586_,
		_w7436_,
		_w7450_,
		_w7451_
	);
	LUT2 #(
		.INIT('h2)
	) name3404 (
		_w7425_,
		_w7414_,
		_w7452_
	);
	LUT3 #(
		.INIT('ha8)
	) name3405 (
		\DM_rd0[8]_pad ,
		_w5610_,
		_w5612_,
		_w7453_
	);
	LUT4 #(
		.INIT('h135f)
	) name3406 (
		\DM_rdm[8]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w7454_
	);
	LUT4 #(
		.INIT('h135f)
	) name3407 (
		\DM_rd6[8]_pad ,
		\DM_rd7[8]_pad ,
		_w5596_,
		_w5591_,
		_w7455_
	);
	LUT2 #(
		.INIT('h8)
	) name3408 (
		_w7454_,
		_w7455_,
		_w7456_
	);
	LUT3 #(
		.INIT('h80)
	) name3409 (
		\DM_rd5[8]_pad ,
		_w5598_,
		_w5599_,
		_w7457_
	);
	LUT3 #(
		.INIT('h80)
	) name3410 (
		\DM_rd4[8]_pad ,
		_w5598_,
		_w5601_,
		_w7458_
	);
	LUT4 #(
		.INIT('h8000)
	) name3411 (
		\DM_rd2[8]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w7459_
	);
	LUT4 #(
		.INIT('h8000)
	) name3412 (
		\DM_rd1[8]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w7460_
	);
	LUT4 #(
		.INIT('h8000)
	) name3413 (
		\DM_rd3[8]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w7461_
	);
	LUT3 #(
		.INIT('h01)
	) name3414 (
		_w7460_,
		_w7461_,
		_w7459_,
		_w7462_
	);
	LUT3 #(
		.INIT('h10)
	) name3415 (
		_w7458_,
		_w7457_,
		_w7462_,
		_w7463_
	);
	LUT2 #(
		.INIT('h8)
	) name3416 (
		_w7456_,
		_w7463_,
		_w7464_
	);
	LUT2 #(
		.INIT('h4)
	) name3417 (
		_w7453_,
		_w7464_,
		_w7465_
	);
	LUT4 #(
		.INIT('h4000)
	) name3418 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[8]/P0001 ,
		_w7466_
	);
	LUT3 #(
		.INIT('h80)
	) name3419 (
		\bdma_BCTL_reg[8]/NET0131 ,
		_w5627_,
		_w5629_,
		_w7467_
	);
	LUT3 #(
		.INIT('h80)
	) name3420 (
		\tm_tpr_reg_DO_reg[8]/NET0131 ,
		_w5631_,
		_w5635_,
		_w7468_
	);
	LUT3 #(
		.INIT('h80)
	) name3421 (
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w5634_,
		_w5639_,
		_w7469_
	);
	LUT3 #(
		.INIT('h80)
	) name3422 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w5628_,
		_w5639_,
		_w7470_
	);
	LUT4 #(
		.INIT('h0001)
	) name3423 (
		_w5795_,
		_w7468_,
		_w7469_,
		_w7470_,
		_w7471_
	);
	LUT4 #(
		.INIT('h8000)
	) name3424 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_txctl_Wcnt_reg[0]/NET0131 ,
		_w5631_,
		_w5639_,
		_w7472_
	);
	LUT4 #(
		.INIT('h8000)
	) name3425 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_txctl_Wcnt_reg[0]/NET0131 ,
		_w5634_,
		_w5660_,
		_w7473_
	);
	LUT2 #(
		.INIT('h1)
	) name3426 (
		_w7472_,
		_w7473_,
		_w7474_
	);
	LUT3 #(
		.INIT('h40)
	) name3427 (
		_w7467_,
		_w7471_,
		_w7474_,
		_w7475_
	);
	LUT3 #(
		.INIT('h80)
	) name3428 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w5629_,
		_w5648_,
		_w7476_
	);
	LUT3 #(
		.INIT('h80)
	) name3429 (
		\bdma_BEAD_reg[8]/NET0131 ,
		_w5629_,
		_w5644_,
		_w7477_
	);
	LUT2 #(
		.INIT('h1)
	) name3430 (
		_w7476_,
		_w7477_,
		_w7478_
	);
	LUT4 #(
		.INIT('h8000)
	) name3431 (
		\bdma_BWCOUNT_reg[8]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w7479_
	);
	LUT4 #(
		.INIT('h8000)
	) name3432 (
		\bdma_BOVL_reg[8]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w7480_
	);
	LUT3 #(
		.INIT('h80)
	) name3433 (
		\IRFS1_pad ,
		_w5644_,
		_w5634_,
		_w7481_
	);
	LUT3 #(
		.INIT('h80)
	) name3434 (
		\memc_usysr_DO_reg[8]/NET0131 ,
		_w5631_,
		_w5660_,
		_w7482_
	);
	LUT3 #(
		.INIT('h80)
	) name3435 (
		\clkc_ckr_reg_DO_reg[8]/NET0131 ,
		_w5631_,
		_w5644_,
		_w7483_
	);
	LUT3 #(
		.INIT('h80)
	) name3436 (
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w5634_,
		_w5637_,
		_w7484_
	);
	LUT4 #(
		.INIT('h0001)
	) name3437 (
		_w7481_,
		_w7482_,
		_w7483_,
		_w7484_,
		_w7485_
	);
	LUT3 #(
		.INIT('h80)
	) name3438 (
		\sport0_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w5627_,
		_w5634_,
		_w7486_
	);
	LUT3 #(
		.INIT('h80)
	) name3439 (
		\emc_WSCRreg_DO_reg[8]/NET0131 ,
		_w5631_,
		_w5632_,
		_w7487_
	);
	LUT3 #(
		.INIT('h80)
	) name3440 (
		\sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w5648_,
		_w5634_,
		_w7488_
	);
	LUT3 #(
		.INIT('h80)
	) name3441 (
		\sport1_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w5670_,
		_w5810_,
		_w7489_
	);
	LUT4 #(
		.INIT('h0001)
	) name3442 (
		_w7486_,
		_w7487_,
		_w7488_,
		_w7489_,
		_w7490_
	);
	LUT3 #(
		.INIT('h80)
	) name3443 (
		\idma_DOVL_reg[8]/NET0131 ,
		_w5804_,
		_w5824_,
		_w7491_
	);
	LUT3 #(
		.INIT('h80)
	) name3444 (
		\IRFS0_pad ,
		_w5632_,
		_w5634_,
		_w7492_
	);
	LUT3 #(
		.INIT('h80)
	) name3445 (
		\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w5634_,
		_w5635_,
		_w7493_
	);
	LUT3 #(
		.INIT('h80)
	) name3446 (
		\tm_TCR_TMP_reg[8]/NET0131 ,
		_w5631_,
		_w5637_,
		_w7494_
	);
	LUT4 #(
		.INIT('h0001)
	) name3447 (
		_w7491_,
		_w7492_,
		_w7493_,
		_w7494_,
		_w7495_
	);
	LUT4 #(
		.INIT('h4000)
	) name3448 (
		_w7480_,
		_w7485_,
		_w7490_,
		_w7495_,
		_w7496_
	);
	LUT4 #(
		.INIT('h4000)
	) name3449 (
		_w7479_,
		_w7475_,
		_w7478_,
		_w7496_,
		_w7497_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3450 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4184_,
		_w4181_,
		_w4189_,
		_w7498_
	);
	LUT3 #(
		.INIT('ha8)
	) name3451 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w7499_
	);
	LUT2 #(
		.INIT('h8)
	) name3452 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w7500_
	);
	LUT4 #(
		.INIT('h135f)
	) name3453 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w7501_
	);
	LUT3 #(
		.INIT('h10)
	) name3454 (
		_w7499_,
		_w7500_,
		_w7501_,
		_w7502_
	);
	LUT3 #(
		.INIT('h8a)
	) name3455 (
		_w5681_,
		_w7498_,
		_w7502_,
		_w7503_
	);
	LUT4 #(
		.INIT('h135f)
	) name3456 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131 ,
		_w7504_
	);
	LUT4 #(
		.INIT('h135f)
	) name3457 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131 ,
		_w7505_
	);
	LUT2 #(
		.INIT('h8)
	) name3458 (
		_w7504_,
		_w7505_,
		_w7506_
	);
	LUT4 #(
		.INIT('h135f)
	) name3459 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131 ,
		_w7507_
	);
	LUT4 #(
		.INIT('h135f)
	) name3460 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131 ,
		_w7508_
	);
	LUT4 #(
		.INIT('h135f)
	) name3461 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131 ,
		_w7509_
	);
	LUT4 #(
		.INIT('h135f)
	) name3462 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131 ,
		_w7510_
	);
	LUT4 #(
		.INIT('h8000)
	) name3463 (
		_w7509_,
		_w7510_,
		_w7507_,
		_w7508_,
		_w7511_
	);
	LUT3 #(
		.INIT('h2a)
	) name3464 (
		_w5697_,
		_w7506_,
		_w7511_,
		_w7512_
	);
	LUT4 #(
		.INIT('h135f)
	) name3465 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131 ,
		_w7513_
	);
	LUT4 #(
		.INIT('h135f)
	) name3466 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131 ,
		_w7514_
	);
	LUT2 #(
		.INIT('h8)
	) name3467 (
		_w7513_,
		_w7514_,
		_w7515_
	);
	LUT4 #(
		.INIT('h135f)
	) name3468 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131 ,
		_w7516_
	);
	LUT4 #(
		.INIT('h135f)
	) name3469 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131 ,
		_w7517_
	);
	LUT4 #(
		.INIT('h135f)
	) name3470 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131 ,
		_w7518_
	);
	LUT4 #(
		.INIT('h135f)
	) name3471 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 ,
		_w7519_
	);
	LUT4 #(
		.INIT('h8000)
	) name3472 (
		_w7518_,
		_w7519_,
		_w7516_,
		_w7517_,
		_w7520_
	);
	LUT4 #(
		.INIT('h135f)
	) name3473 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[8]/P0001 ,
		\sport1_txctl_TX_reg[8]/P0001 ,
		_w7521_
	);
	LUT4 #(
		.INIT('h135f)
	) name3474 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[8]/P0001 ,
		\sport1_rxctl_RX_reg[8]/P0001 ,
		_w7522_
	);
	LUT3 #(
		.INIT('h2a)
	) name3475 (
		_w5706_,
		_w7521_,
		_w7522_,
		_w7523_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3476 (
		_w5687_,
		_w7515_,
		_w7520_,
		_w7523_,
		_w7524_
	);
	LUT2 #(
		.INIT('h4)
	) name3477 (
		_w7512_,
		_w7524_,
		_w7525_
	);
	LUT3 #(
		.INIT('h1b)
	) name3478 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001 ,
		_w7526_
	);
	LUT4 #(
		.INIT('ha820)
	) name3479 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001 ,
		_w7527_
	);
	LUT3 #(
		.INIT('h1b)
	) name3480 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001 ,
		_w7528_
	);
	LUT4 #(
		.INIT('ha820)
	) name3481 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001 ,
		_w7529_
	);
	LUT3 #(
		.INIT('h1b)
	) name3482 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001 ,
		_w7530_
	);
	LUT4 #(
		.INIT('ha820)
	) name3483 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001 ,
		_w7531_
	);
	LUT3 #(
		.INIT('h01)
	) name3484 (
		_w7529_,
		_w7531_,
		_w7527_,
		_w7532_
	);
	LUT3 #(
		.INIT('h2a)
	) name3485 (
		_w5741_,
		_w5746_,
		_w7532_,
		_w7533_
	);
	LUT3 #(
		.INIT('h1b)
	) name3486 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001 ,
		_w7534_
	);
	LUT4 #(
		.INIT('ha820)
	) name3487 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001 ,
		_w7535_
	);
	LUT4 #(
		.INIT('ha820)
	) name3488 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001 ,
		_w7536_
	);
	LUT2 #(
		.INIT('h1)
	) name3489 (
		_w7535_,
		_w7536_,
		_w7537_
	);
	LUT3 #(
		.INIT('h1b)
	) name3490 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001 ,
		_w7538_
	);
	LUT4 #(
		.INIT('ha820)
	) name3491 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001 ,
		_w7539_
	);
	LUT3 #(
		.INIT('h1b)
	) name3492 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001 ,
		_w7540_
	);
	LUT4 #(
		.INIT('ha820)
	) name3493 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001 ,
		_w7541_
	);
	LUT4 #(
		.INIT('ha820)
	) name3494 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001 ,
		_w7542_
	);
	LUT3 #(
		.INIT('h01)
	) name3495 (
		_w7541_,
		_w7542_,
		_w7539_,
		_w7543_
	);
	LUT3 #(
		.INIT('h2a)
	) name3496 (
		_w5730_,
		_w7537_,
		_w7543_,
		_w7544_
	);
	LUT3 #(
		.INIT('h1b)
	) name3497 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 ,
		_w7545_
	);
	LUT4 #(
		.INIT('ha820)
	) name3498 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 ,
		_w7546_
	);
	LUT3 #(
		.INIT('h1b)
	) name3499 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001 ,
		_w7547_
	);
	LUT4 #(
		.INIT('ha820)
	) name3500 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001 ,
		_w7548_
	);
	LUT3 #(
		.INIT('h1b)
	) name3501 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001 ,
		_w7549_
	);
	LUT4 #(
		.INIT('ha820)
	) name3502 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001 ,
		_w7550_
	);
	LUT3 #(
		.INIT('h01)
	) name3503 (
		_w7548_,
		_w7550_,
		_w7546_,
		_w7551_
	);
	LUT3 #(
		.INIT('h1b)
	) name3504 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001 ,
		_w7552_
	);
	LUT4 #(
		.INIT('ha820)
	) name3505 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001 ,
		_w7553_
	);
	LUT3 #(
		.INIT('h1b)
	) name3506 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001 ,
		_w7554_
	);
	LUT4 #(
		.INIT('ha820)
	) name3507 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001 ,
		_w7555_
	);
	LUT3 #(
		.INIT('h1b)
	) name3508 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001 ,
		_w7556_
	);
	LUT4 #(
		.INIT('ha820)
	) name3509 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001 ,
		_w7557_
	);
	LUT4 #(
		.INIT('h0001)
	) name3510 (
		_w5714_,
		_w7553_,
		_w7555_,
		_w7557_,
		_w7558_
	);
	LUT3 #(
		.INIT('h2a)
	) name3511 (
		_w5712_,
		_w7551_,
		_w7558_,
		_w7559_
	);
	LUT3 #(
		.INIT('h01)
	) name3512 (
		_w7544_,
		_w7559_,
		_w7533_,
		_w7560_
	);
	LUT2 #(
		.INIT('h8)
	) name3513 (
		_w7525_,
		_w7560_,
		_w7561_
	);
	LUT4 #(
		.INIT('h3100)
	) name3514 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w7503_,
		_w7497_,
		_w7561_,
		_w7562_
	);
	LUT2 #(
		.INIT('h8)
	) name3515 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[8]/P0001 ,
		_w7563_
	);
	LUT3 #(
		.INIT('h08)
	) name3516 (
		_w5588_,
		_w5598_,
		_w7563_,
		_w7564_
	);
	LUT4 #(
		.INIT('hba00)
	) name3517 (
		\emc_DMDoe_reg/NET0131 ,
		_w7466_,
		_w7562_,
		_w7564_,
		_w7565_
	);
	LUT2 #(
		.INIT('h1)
	) name3518 (
		_w7465_,
		_w7565_,
		_w7566_
	);
	LUT4 #(
		.INIT('hecfd)
	) name3519 (
		_w5117_,
		_w5337_,
		_w7452_,
		_w7566_,
		_w7567_
	);
	LUT2 #(
		.INIT('h2)
	) name3520 (
		_w5586_,
		_w7567_,
		_w7568_
	);
	LUT4 #(
		.INIT('h888e)
	) name3521 (
		\core_dag_ilm1reg_M_reg[4]/NET0131 ,
		_w5217_,
		_w5162_,
		_w5297_,
		_w7569_
	);
	LUT2 #(
		.INIT('h9)
	) name3522 (
		_w5220_,
		_w7569_,
		_w7570_
	);
	LUT4 #(
		.INIT('h9a00)
	) name3523 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w7570_,
		_w7571_
	);
	LUT2 #(
		.INIT('h9)
	) name3524 (
		_w5219_,
		_w5221_,
		_w7572_
	);
	LUT4 #(
		.INIT('hf10e)
	) name3525 (
		_w5225_,
		_w5193_,
		_w5228_,
		_w7572_,
		_w7573_
	);
	LUT4 #(
		.INIT('h6500)
	) name3526 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w7573_,
		_w7574_
	);
	LUT3 #(
		.INIT('h01)
	) name3527 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w7574_,
		_w7571_,
		_w7575_
	);
	LUT4 #(
		.INIT('haa20)
	) name3528 (
		\core_dag_ilm1reg_I_reg[5]/NET0131 ,
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w5195_,
		_w5201_,
		_w7576_
	);
	LUT3 #(
		.INIT('h10)
	) name3529 (
		_w5767_,
		_w5768_,
		_w7570_,
		_w7577_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3530 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5155_,
		_w5310_,
		_w7573_,
		_w7578_
	);
	LUT4 #(
		.INIT('h0045)
	) name3531 (
		_w7576_,
		_w7577_,
		_w7578_,
		_w7575_,
		_w7579_
	);
	LUT3 #(
		.INIT('ha8)
	) name3532 (
		\DM_rd0[5]_pad ,
		_w5610_,
		_w5612_,
		_w7580_
	);
	LUT4 #(
		.INIT('h135f)
	) name3533 (
		\DM_rdm[5]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w7581_
	);
	LUT4 #(
		.INIT('h135f)
	) name3534 (
		\DM_rd6[5]_pad ,
		\DM_rd7[5]_pad ,
		_w5596_,
		_w5591_,
		_w7582_
	);
	LUT2 #(
		.INIT('h8)
	) name3535 (
		_w7581_,
		_w7582_,
		_w7583_
	);
	LUT3 #(
		.INIT('h80)
	) name3536 (
		\DM_rd5[5]_pad ,
		_w5598_,
		_w5599_,
		_w7584_
	);
	LUT3 #(
		.INIT('h80)
	) name3537 (
		\DM_rd4[5]_pad ,
		_w5598_,
		_w5601_,
		_w7585_
	);
	LUT4 #(
		.INIT('h8000)
	) name3538 (
		\DM_rd2[5]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w7586_
	);
	LUT4 #(
		.INIT('h8000)
	) name3539 (
		\DM_rd1[5]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w7587_
	);
	LUT4 #(
		.INIT('h8000)
	) name3540 (
		\DM_rd3[5]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w7588_
	);
	LUT3 #(
		.INIT('h01)
	) name3541 (
		_w7587_,
		_w7588_,
		_w7586_,
		_w7589_
	);
	LUT3 #(
		.INIT('h10)
	) name3542 (
		_w7585_,
		_w7584_,
		_w7589_,
		_w7590_
	);
	LUT2 #(
		.INIT('h8)
	) name3543 (
		_w7583_,
		_w7590_,
		_w7591_
	);
	LUT2 #(
		.INIT('h4)
	) name3544 (
		_w7580_,
		_w7591_,
		_w7592_
	);
	LUT4 #(
		.INIT('h4000)
	) name3545 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[5]/P0001 ,
		_w7593_
	);
	LUT3 #(
		.INIT('h80)
	) name3546 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w5629_,
		_w5648_,
		_w7594_
	);
	LUT3 #(
		.INIT('h80)
	) name3547 (
		\emc_WSCRreg_DO_reg[5]/NET0131 ,
		_w5631_,
		_w5632_,
		_w7595_
	);
	LUT3 #(
		.INIT('h80)
	) name3548 (
		\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w5634_,
		_w5635_,
		_w7596_
	);
	LUT3 #(
		.INIT('h80)
	) name3549 (
		\sport1_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w5631_,
		_w5639_,
		_w7597_
	);
	LUT3 #(
		.INIT('h80)
	) name3550 (
		\tm_tsr_reg_DO_reg[5]/NET0131 ,
		_w5627_,
		_w5631_,
		_w7598_
	);
	LUT4 #(
		.INIT('h0001)
	) name3551 (
		_w7595_,
		_w7596_,
		_w7597_,
		_w7598_,
		_w7599_
	);
	LUT3 #(
		.INIT('h80)
	) name3552 (
		\idma_DOVL_reg[5]/NET0131 ,
		_w5804_,
		_w5824_,
		_w7600_
	);
	LUT3 #(
		.INIT('h80)
	) name3553 (
		\sport0_regs_AUTOreg_DO_reg[5]/NET0131 ,
		_w5627_,
		_w5634_,
		_w7601_
	);
	LUT3 #(
		.INIT('h80)
	) name3554 (
		\tm_tpr_reg_DO_reg[5]/NET0131 ,
		_w5631_,
		_w5635_,
		_w7602_
	);
	LUT4 #(
		.INIT('h0001)
	) name3555 (
		_w5795_,
		_w7600_,
		_w7601_,
		_w7602_,
		_w7603_
	);
	LUT3 #(
		.INIT('h40)
	) name3556 (
		_w7594_,
		_w7599_,
		_w7603_,
		_w7604_
	);
	LUT3 #(
		.INIT('h80)
	) name3557 (
		\bdma_BEAD_reg[5]/NET0131 ,
		_w5629_,
		_w5644_,
		_w7605_
	);
	LUT3 #(
		.INIT('h80)
	) name3558 (
		\bdma_BCTL_reg[5]/NET0131 ,
		_w5627_,
		_w5629_,
		_w7606_
	);
	LUT2 #(
		.INIT('h1)
	) name3559 (
		_w7605_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h8)
	) name3560 (
		_w7604_,
		_w7607_,
		_w7608_
	);
	LUT4 #(
		.INIT('h8000)
	) name3561 (
		\bdma_BOVL_reg[5]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w7609_
	);
	LUT3 #(
		.INIT('h1b)
	) name3562 (
		\bdma_BDMA_boot_reg/NET0131_reg_syn_10 ,
		\bdma_BWCOUNT_reg[5]/NET0131_reg_syn_2 ,
		\bdma_BWCOUNT_reg[5]/NET0131_reg_syn_8 ,
		_w7610_
	);
	LUT4 #(
		.INIT('h0080)
	) name3563 (
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w7610_,
		_w7611_
	);
	LUT3 #(
		.INIT('h80)
	) name3564 (
		\pio_pmask_reg_DO_reg[5]/NET0131 ,
		_w5628_,
		_w5660_,
		_w7612_
	);
	LUT3 #(
		.INIT('h80)
	) name3565 (
		\sport0_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w5634_,
		_w5660_,
		_w7613_
	);
	LUT3 #(
		.INIT('h80)
	) name3566 (
		\sport1_regs_AUTOreg_DO_reg[5]/NET0131 ,
		_w5670_,
		_w5810_,
		_w7614_
	);
	LUT3 #(
		.INIT('h80)
	) name3567 (
		\tm_TCR_TMP_reg[5]/NET0131 ,
		_w5631_,
		_w5637_,
		_w7615_
	);
	LUT4 #(
		.INIT('h0001)
	) name3568 (
		_w7612_,
		_w7613_,
		_w7614_,
		_w7615_,
		_w7616_
	);
	LUT3 #(
		.INIT('h80)
	) name3569 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w5632_,
		_w5634_,
		_w7617_
	);
	LUT3 #(
		.INIT('h80)
	) name3570 (
		\emc_WSCRext_reg_DO_reg[5]/NET0131 ,
		_w5670_,
		_w5790_,
		_w7618_
	);
	LUT3 #(
		.INIT('h80)
	) name3571 (
		\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w5648_,
		_w5634_,
		_w7619_
	);
	LUT3 #(
		.INIT('h80)
	) name3572 (
		\sport1_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w5644_,
		_w5634_,
		_w7620_
	);
	LUT4 #(
		.INIT('h0001)
	) name3573 (
		_w7617_,
		_w7618_,
		_w7619_,
		_w7620_,
		_w7621_
	);
	LUT3 #(
		.INIT('h80)
	) name3574 (
		\idma_DCTL_reg[5]/NET0131 ,
		_w5628_,
		_w5639_,
		_w7622_
	);
	LUT3 #(
		.INIT('h80)
	) name3575 (
		\PIO_out[5]_pad ,
		_w5628_,
		_w5635_,
		_w7623_
	);
	LUT3 #(
		.INIT('h80)
	) name3576 (
		\PIO_oe[5]_pad ,
		_w5628_,
		_w5632_,
		_w7624_
	);
	LUT3 #(
		.INIT('h80)
	) name3577 (
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w5634_,
		_w5639_,
		_w7625_
	);
	LUT4 #(
		.INIT('h0001)
	) name3578 (
		_w7622_,
		_w7623_,
		_w7624_,
		_w7625_,
		_w7626_
	);
	LUT3 #(
		.INIT('h80)
	) name3579 (
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w5634_,
		_w5637_,
		_w7627_
	);
	LUT3 #(
		.INIT('h80)
	) name3580 (
		\clkc_ckr_reg_DO_reg[5]/NET0131 ,
		_w5631_,
		_w5644_,
		_w7628_
	);
	LUT3 #(
		.INIT('h80)
	) name3581 (
		\memc_usysr_DO_reg[5]/NET0131 ,
		_w5631_,
		_w5660_,
		_w7629_
	);
	LUT3 #(
		.INIT('h80)
	) name3582 (
		\pio_PINT_reg[5]/NET0131 ,
		_w5670_,
		_w5672_,
		_w7630_
	);
	LUT4 #(
		.INIT('h0001)
	) name3583 (
		_w7627_,
		_w7628_,
		_w7629_,
		_w7630_,
		_w7631_
	);
	LUT4 #(
		.INIT('h8000)
	) name3584 (
		_w7626_,
		_w7631_,
		_w7616_,
		_w7621_,
		_w7632_
	);
	LUT3 #(
		.INIT('h10)
	) name3585 (
		_w7611_,
		_w7609_,
		_w7632_,
		_w7633_
	);
	LUT3 #(
		.INIT('h2a)
	) name3586 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w7608_,
		_w7633_,
		_w7634_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3587 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4322_,
		_w4319_,
		_w4327_,
		_w7635_
	);
	LUT4 #(
		.INIT('h135f)
	) name3588 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w7636_
	);
	LUT4 #(
		.INIT('h153f)
	) name3589 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[5]/NET0131 ,
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w7637_
	);
	LUT3 #(
		.INIT('ha8)
	) name3590 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w7638_
	);
	LUT4 #(
		.INIT('h135f)
	) name3591 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		_w7639_
	);
	LUT4 #(
		.INIT('h4000)
	) name3592 (
		_w7638_,
		_w7639_,
		_w7636_,
		_w7637_,
		_w7640_
	);
	LUT3 #(
		.INIT('h8a)
	) name3593 (
		_w5681_,
		_w7635_,
		_w7640_,
		_w7641_
	);
	LUT4 #(
		.INIT('h135f)
	) name3594 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131 ,
		_w7642_
	);
	LUT4 #(
		.INIT('h135f)
	) name3595 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131 ,
		_w7643_
	);
	LUT2 #(
		.INIT('h8)
	) name3596 (
		_w7642_,
		_w7643_,
		_w7644_
	);
	LUT4 #(
		.INIT('h135f)
	) name3597 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131 ,
		_w7645_
	);
	LUT4 #(
		.INIT('h135f)
	) name3598 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w7646_
	);
	LUT4 #(
		.INIT('h135f)
	) name3599 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131 ,
		_w7647_
	);
	LUT4 #(
		.INIT('h135f)
	) name3600 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131 ,
		_w7648_
	);
	LUT4 #(
		.INIT('h8000)
	) name3601 (
		_w7647_,
		_w7648_,
		_w7645_,
		_w7646_,
		_w7649_
	);
	LUT3 #(
		.INIT('h2a)
	) name3602 (
		_w5687_,
		_w7644_,
		_w7649_,
		_w7650_
	);
	LUT4 #(
		.INIT('h135f)
	) name3603 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w7651_
	);
	LUT4 #(
		.INIT('h135f)
	) name3604 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 ,
		_w7652_
	);
	LUT2 #(
		.INIT('h8)
	) name3605 (
		_w7651_,
		_w7652_,
		_w7653_
	);
	LUT4 #(
		.INIT('h135f)
	) name3606 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131 ,
		_w7654_
	);
	LUT4 #(
		.INIT('h135f)
	) name3607 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131 ,
		_w7655_
	);
	LUT4 #(
		.INIT('h135f)
	) name3608 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131 ,
		_w7656_
	);
	LUT4 #(
		.INIT('h135f)
	) name3609 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131 ,
		_w7657_
	);
	LUT4 #(
		.INIT('h8000)
	) name3610 (
		_w7656_,
		_w7657_,
		_w7654_,
		_w7655_,
		_w7658_
	);
	LUT4 #(
		.INIT('h135f)
	) name3611 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[5]/P0001 ,
		\sport1_txctl_TX_reg[5]/P0001 ,
		_w7659_
	);
	LUT4 #(
		.INIT('h135f)
	) name3612 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport1_rxctl_RX_reg[5]/P0001 ,
		_w7660_
	);
	LUT3 #(
		.INIT('h2a)
	) name3613 (
		_w5706_,
		_w7659_,
		_w7660_,
		_w7661_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3614 (
		_w5697_,
		_w7653_,
		_w7658_,
		_w7661_,
		_w7662_
	);
	LUT2 #(
		.INIT('h4)
	) name3615 (
		_w7650_,
		_w7662_,
		_w7663_
	);
	LUT3 #(
		.INIT('h1b)
	) name3616 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001 ,
		_w7664_
	);
	LUT4 #(
		.INIT('ha820)
	) name3617 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001 ,
		_w7665_
	);
	LUT3 #(
		.INIT('h1b)
	) name3618 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001 ,
		_w7666_
	);
	LUT4 #(
		.INIT('ha820)
	) name3619 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001 ,
		_w7667_
	);
	LUT3 #(
		.INIT('h1b)
	) name3620 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001 ,
		_w7668_
	);
	LUT4 #(
		.INIT('ha820)
	) name3621 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001 ,
		_w7669_
	);
	LUT3 #(
		.INIT('h01)
	) name3622 (
		_w7667_,
		_w7669_,
		_w7665_,
		_w7670_
	);
	LUT3 #(
		.INIT('h1b)
	) name3623 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 ,
		_w7671_
	);
	LUT4 #(
		.INIT('ha820)
	) name3624 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 ,
		_w7672_
	);
	LUT3 #(
		.INIT('h1b)
	) name3625 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001 ,
		_w7673_
	);
	LUT4 #(
		.INIT('ha820)
	) name3626 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001 ,
		_w7674_
	);
	LUT3 #(
		.INIT('h1b)
	) name3627 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001 ,
		_w7675_
	);
	LUT4 #(
		.INIT('ha820)
	) name3628 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001 ,
		_w7676_
	);
	LUT3 #(
		.INIT('h1b)
	) name3629 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001 ,
		_w7677_
	);
	LUT4 #(
		.INIT('ha820)
	) name3630 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001 ,
		_w7678_
	);
	LUT4 #(
		.INIT('h0001)
	) name3631 (
		_w7672_,
		_w7674_,
		_w7676_,
		_w7678_,
		_w7679_
	);
	LUT3 #(
		.INIT('h2a)
	) name3632 (
		_w5712_,
		_w7670_,
		_w7679_,
		_w7680_
	);
	LUT3 #(
		.INIT('h1b)
	) name3633 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001 ,
		_w7681_
	);
	LUT4 #(
		.INIT('ha820)
	) name3634 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001 ,
		_w7682_
	);
	LUT2 #(
		.INIT('h8)
	) name3635 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w7683_
	);
	LUT2 #(
		.INIT('h1)
	) name3636 (
		_w7682_,
		_w7683_,
		_w7684_
	);
	LUT4 #(
		.INIT('ha820)
	) name3637 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001 ,
		_w7685_
	);
	LUT3 #(
		.INIT('h1b)
	) name3638 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001 ,
		_w7686_
	);
	LUT4 #(
		.INIT('ha820)
	) name3639 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001 ,
		_w7687_
	);
	LUT4 #(
		.INIT('ha820)
	) name3640 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001 ,
		_w7688_
	);
	LUT4 #(
		.INIT('ha820)
	) name3641 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001 ,
		_w7689_
	);
	LUT4 #(
		.INIT('h0001)
	) name3642 (
		_w7685_,
		_w7687_,
		_w7688_,
		_w7689_,
		_w7690_
	);
	LUT3 #(
		.INIT('h2a)
	) name3643 (
		_w5730_,
		_w7684_,
		_w7690_,
		_w7691_
	);
	LUT3 #(
		.INIT('h1b)
	) name3644 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001 ,
		_w7692_
	);
	LUT4 #(
		.INIT('ha820)
	) name3645 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001 ,
		_w7693_
	);
	LUT2 #(
		.INIT('h1)
	) name3646 (
		_w5743_,
		_w7693_,
		_w7694_
	);
	LUT3 #(
		.INIT('h1b)
	) name3647 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001 ,
		_w7695_
	);
	LUT4 #(
		.INIT('ha820)
	) name3648 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001 ,
		_w7696_
	);
	LUT3 #(
		.INIT('h1b)
	) name3649 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001 ,
		_w7697_
	);
	LUT4 #(
		.INIT('ha820)
	) name3650 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001 ,
		_w7698_
	);
	LUT3 #(
		.INIT('h1b)
	) name3651 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001 ,
		_w7699_
	);
	LUT4 #(
		.INIT('ha820)
	) name3652 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001 ,
		_w7700_
	);
	LUT3 #(
		.INIT('h01)
	) name3653 (
		_w7698_,
		_w7700_,
		_w7696_,
		_w7701_
	);
	LUT3 #(
		.INIT('h2a)
	) name3654 (
		_w5741_,
		_w7694_,
		_w7701_,
		_w7702_
	);
	LUT3 #(
		.INIT('h01)
	) name3655 (
		_w7691_,
		_w7702_,
		_w7680_,
		_w7703_
	);
	LUT2 #(
		.INIT('h8)
	) name3656 (
		_w7663_,
		_w7703_,
		_w7704_
	);
	LUT2 #(
		.INIT('h4)
	) name3657 (
		_w7641_,
		_w7704_,
		_w7705_
	);
	LUT3 #(
		.INIT('h10)
	) name3658 (
		_w7593_,
		_w7634_,
		_w7705_,
		_w7706_
	);
	LUT4 #(
		.INIT('h5455)
	) name3659 (
		\emc_DMDoe_reg/NET0131 ,
		_w7593_,
		_w7634_,
		_w7705_,
		_w7707_
	);
	LUT2 #(
		.INIT('h8)
	) name3660 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[5]/P0001 ,
		_w7708_
	);
	LUT3 #(
		.INIT('h08)
	) name3661 (
		_w5588_,
		_w5598_,
		_w7708_,
		_w7709_
	);
	LUT3 #(
		.INIT('h45)
	) name3662 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w7710_
	);
	LUT4 #(
		.INIT('hc040)
	) name3663 (
		_w5117_,
		_w5337_,
		_w5586_,
		_w7710_,
		_w7711_
	);
	LUT4 #(
		.INIT('h1033)
	) name3664 (
		_w5117_,
		_w7568_,
		_w7579_,
		_w7711_,
		_w7712_
	);
	LUT4 #(
		.INIT('h2f00)
	) name3665 (
		_w5117_,
		_w7401_,
		_w7451_,
		_w7712_,
		_w7713_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name3666 (
		_w5117_,
		_w7401_,
		_w7451_,
		_w7712_,
		_w7714_
	);
	LUT4 #(
		.INIT('haa20)
	) name3667 (
		\core_dag_ilm2reg_I_reg[6]/NET0131 ,
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w5399_,
		_w5400_,
		_w7715_
	);
	LUT4 #(
		.INIT('h6996)
	) name3668 (
		\core_dag_ilm2reg_M_reg[6]/NET0131 ,
		_w5405_,
		_w5447_,
		_w5451_,
		_w7716_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3669 (
		_w5463_,
		_w5472_,
		_w5484_,
		_w5486_,
		_w7717_
	);
	LUT2 #(
		.INIT('h6)
	) name3670 (
		_w7716_,
		_w7717_,
		_w7718_
	);
	LUT2 #(
		.INIT('h6)
	) name3671 (
		_w5426_,
		_w5452_,
		_w7719_
	);
	LUT4 #(
		.INIT('h01ef)
	) name3672 (
		_w5434_,
		_w6210_,
		_w7718_,
		_w7719_,
		_w7720_
	);
	LUT4 #(
		.INIT('h781e)
	) name3673 (
		\core_dag_ilm1reg_M_reg[6]/NET0131 ,
		_w5196_,
		_w5210_,
		_w5300_,
		_w7721_
	);
	LUT4 #(
		.INIT('h009a)
	) name3674 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w7721_,
		_w7722_
	);
	LUT2 #(
		.INIT('h9)
	) name3675 (
		_w5212_,
		_w5213_,
		_w7723_
	);
	LUT4 #(
		.INIT('h0455)
	) name3676 (
		_w5205_,
		_w5226_,
		_w5193_,
		_w5229_,
		_w7724_
	);
	LUT3 #(
		.INIT('hc9)
	) name3677 (
		_w5230_,
		_w7723_,
		_w7724_,
		_w7725_
	);
	LUT4 #(
		.INIT('h6500)
	) name3678 (
		_w5156_,
		_w5286_,
		_w5288_,
		_w7725_,
		_w7726_
	);
	LUT3 #(
		.INIT('h01)
	) name3679 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w7726_,
		_w7722_,
		_w7727_
	);
	LUT3 #(
		.INIT('h02)
	) name3680 (
		\core_dag_ilm1reg_I_reg[7]/NET0131 ,
		_w5153_,
		_w5206_,
		_w7728_
	);
	LUT3 #(
		.INIT('h01)
	) name3681 (
		_w5767_,
		_w5768_,
		_w7721_,
		_w7729_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3682 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w5155_,
		_w5310_,
		_w7725_,
		_w7730_
	);
	LUT4 #(
		.INIT('h0045)
	) name3683 (
		_w7728_,
		_w7729_,
		_w7730_,
		_w7727_,
		_w7731_
	);
	LUT4 #(
		.INIT('h54fe)
	) name3684 (
		_w5337_,
		_w7715_,
		_w7720_,
		_w7731_,
		_w7732_
	);
	LUT4 #(
		.INIT('h0200)
	) name3685 (
		\core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w7733_
	);
	LUT4 #(
		.INIT('h0200)
	) name3686 (
		\core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w7734_
	);
	LUT4 #(
		.INIT('h0200)
	) name3687 (
		\core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w7735_
	);
	LUT4 #(
		.INIT('h0200)
	) name3688 (
		\core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w7736_
	);
	LUT3 #(
		.INIT('h01)
	) name3689 (
		_w7735_,
		_w7736_,
		_w7734_,
		_w7737_
	);
	LUT4 #(
		.INIT('h0200)
	) name3690 (
		\core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w7738_
	);
	LUT4 #(
		.INIT('h0200)
	) name3691 (
		\core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w7739_
	);
	LUT4 #(
		.INIT('h0200)
	) name3692 (
		\core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w7740_
	);
	LUT4 #(
		.INIT('h0200)
	) name3693 (
		\core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w7741_
	);
	LUT4 #(
		.INIT('h0001)
	) name3694 (
		_w7738_,
		_w7739_,
		_w7740_,
		_w7741_,
		_w7742_
	);
	LUT4 #(
		.INIT('h45ef)
	) name3695 (
		_w4063_,
		_w7733_,
		_w7737_,
		_w7742_,
		_w7743_
	);
	LUT4 #(
		.INIT('h0200)
	) name3696 (
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w7744_
	);
	LUT4 #(
		.INIT('h0200)
	) name3697 (
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w7745_
	);
	LUT4 #(
		.INIT('h0200)
	) name3698 (
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w7746_
	);
	LUT4 #(
		.INIT('h0200)
	) name3699 (
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w7747_
	);
	LUT4 #(
		.INIT('h0001)
	) name3700 (
		_w7744_,
		_w7745_,
		_w7746_,
		_w7747_,
		_w7748_
	);
	LUT4 #(
		.INIT('h0200)
	) name3701 (
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w7749_
	);
	LUT4 #(
		.INIT('h0200)
	) name3702 (
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w7750_
	);
	LUT4 #(
		.INIT('h0200)
	) name3703 (
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w7751_
	);
	LUT4 #(
		.INIT('h0200)
	) name3704 (
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w7752_
	);
	LUT4 #(
		.INIT('h0001)
	) name3705 (
		_w7749_,
		_w7750_,
		_w7751_,
		_w7752_,
		_w7753_
	);
	LUT3 #(
		.INIT('hd0)
	) name3706 (
		_w4063_,
		_w7748_,
		_w7753_,
		_w7754_
	);
	LUT4 #(
		.INIT('h0233)
	) name3707 (
		_w4063_,
		_w5049_,
		_w7748_,
		_w7753_,
		_w7755_
	);
	LUT4 #(
		.INIT('h0080)
	) name3708 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w7756_
	);
	LUT4 #(
		.INIT('h0203)
	) name3709 (
		_w4970_,
		_w7755_,
		_w7756_,
		_w7743_,
		_w7757_
	);
	LUT4 #(
		.INIT('ha222)
	) name3710 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w7758_
	);
	LUT4 #(
		.INIT('h2a00)
	) name3711 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w7759_
	);
	LUT4 #(
		.INIT('h4000)
	) name3712 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w7760_
	);
	LUT2 #(
		.INIT('h1)
	) name3713 (
		_w7759_,
		_w7760_,
		_w7761_
	);
	LUT3 #(
		.INIT('h20)
	) name3714 (
		_w5539_,
		_w7758_,
		_w7761_,
		_w7762_
	);
	LUT3 #(
		.INIT('hd0)
	) name3715 (
		_w5059_,
		_w7757_,
		_w7762_,
		_w7763_
	);
	LUT4 #(
		.INIT('h5540)
	) name3716 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w7764_
	);
	LUT3 #(
		.INIT('h01)
	) name3717 (
		_w5337_,
		_w7764_,
		_w7763_,
		_w7765_
	);
	LUT3 #(
		.INIT('h02)
	) name3718 (
		\core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 ,
		_w5070_,
		_w5073_,
		_w7766_
	);
	LUT4 #(
		.INIT('h0200)
	) name3719 (
		\core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5076_,
		_w7767_
	);
	LUT4 #(
		.INIT('h0200)
	) name3720 (
		\core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5068_,
		_w7768_
	);
	LUT4 #(
		.INIT('h0200)
	) name3721 (
		\core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5093_,
		_w7769_
	);
	LUT4 #(
		.INIT('h0200)
	) name3722 (
		\core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5085_,
		_w7770_
	);
	LUT3 #(
		.INIT('h01)
	) name3723 (
		_w7769_,
		_w7770_,
		_w7768_,
		_w7771_
	);
	LUT4 #(
		.INIT('h0200)
	) name3724 (
		\core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 ,
		_w5061_,
		_w5065_,
		_w5098_,
		_w7772_
	);
	LUT4 #(
		.INIT('h0200)
	) name3725 (
		\core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 ,
		_w5079_,
		_w5082_,
		_w5096_,
		_w7773_
	);
	LUT4 #(
		.INIT('h0200)
	) name3726 (
		\core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 ,
		_w5087_,
		_w5090_,
		_w5102_,
		_w7774_
	);
	LUT4 #(
		.INIT('h0200)
	) name3727 (
		\core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 ,
		_w5070_,
		_w5073_,
		_w5100_,
		_w7775_
	);
	LUT4 #(
		.INIT('h0001)
	) name3728 (
		_w7772_,
		_w7773_,
		_w7774_,
		_w7775_,
		_w7776_
	);
	LUT4 #(
		.INIT('h45ef)
	) name3729 (
		_w4063_,
		_w7767_,
		_w7771_,
		_w7776_,
		_w7777_
	);
	LUT3 #(
		.INIT('h15)
	) name3730 (
		_w5117_,
		_w5337_,
		_w7777_,
		_w7778_
	);
	LUT3 #(
		.INIT('h45)
	) name3731 (
		_w5586_,
		_w7765_,
		_w7778_,
		_w7779_
	);
	LUT2 #(
		.INIT('h2)
	) name3732 (
		_w7754_,
		_w7743_,
		_w7780_
	);
	LUT3 #(
		.INIT('ha8)
	) name3733 (
		\DM_rd0[7]_pad ,
		_w5610_,
		_w5612_,
		_w7781_
	);
	LUT4 #(
		.INIT('h135f)
	) name3734 (
		\DM_rdm[7]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w7782_
	);
	LUT4 #(
		.INIT('h135f)
	) name3735 (
		\DM_rd6[7]_pad ,
		\DM_rd7[7]_pad ,
		_w5596_,
		_w5591_,
		_w7783_
	);
	LUT2 #(
		.INIT('h8)
	) name3736 (
		_w7782_,
		_w7783_,
		_w7784_
	);
	LUT3 #(
		.INIT('h80)
	) name3737 (
		\DM_rd5[7]_pad ,
		_w5598_,
		_w5599_,
		_w7785_
	);
	LUT3 #(
		.INIT('h80)
	) name3738 (
		\DM_rd4[7]_pad ,
		_w5598_,
		_w5601_,
		_w7786_
	);
	LUT4 #(
		.INIT('h8000)
	) name3739 (
		\DM_rd2[7]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w7787_
	);
	LUT4 #(
		.INIT('h8000)
	) name3740 (
		\DM_rd1[7]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w7788_
	);
	LUT4 #(
		.INIT('h8000)
	) name3741 (
		\DM_rd3[7]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w7789_
	);
	LUT3 #(
		.INIT('h01)
	) name3742 (
		_w7788_,
		_w7789_,
		_w7787_,
		_w7790_
	);
	LUT3 #(
		.INIT('h10)
	) name3743 (
		_w7786_,
		_w7785_,
		_w7790_,
		_w7791_
	);
	LUT2 #(
		.INIT('h8)
	) name3744 (
		_w7784_,
		_w7791_,
		_w7792_
	);
	LUT2 #(
		.INIT('h4)
	) name3745 (
		_w7781_,
		_w7792_,
		_w7793_
	);
	LUT4 #(
		.INIT('h4000)
	) name3746 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[7]/P0001 ,
		_w7794_
	);
	LUT3 #(
		.INIT('h80)
	) name3747 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w5629_,
		_w5648_,
		_w7795_
	);
	LUT3 #(
		.INIT('h80)
	) name3748 (
		\emc_WSCRreg_DO_reg[7]/NET0131 ,
		_w5631_,
		_w5632_,
		_w7796_
	);
	LUT3 #(
		.INIT('h80)
	) name3749 (
		\tm_TCR_TMP_reg[7]/NET0131 ,
		_w5631_,
		_w5637_,
		_w7797_
	);
	LUT3 #(
		.INIT('h80)
	) name3750 (
		\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w5634_,
		_w5635_,
		_w7798_
	);
	LUT3 #(
		.INIT('h80)
	) name3751 (
		\sport0_regs_AUTOreg_DO_reg[7]/NET0131 ,
		_w5627_,
		_w5634_,
		_w7799_
	);
	LUT4 #(
		.INIT('h0001)
	) name3752 (
		_w7796_,
		_w7797_,
		_w7798_,
		_w7799_,
		_w7800_
	);
	LUT3 #(
		.INIT('h80)
	) name3753 (
		\sport1_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w5631_,
		_w5639_,
		_w7801_
	);
	LUT3 #(
		.INIT('h80)
	) name3754 (
		\emc_WSCRext_reg_DO_reg[7]/NET0131 ,
		_w5670_,
		_w5790_,
		_w7802_
	);
	LUT3 #(
		.INIT('h80)
	) name3755 (
		\tm_tpr_reg_DO_reg[7]/NET0131 ,
		_w5631_,
		_w5635_,
		_w7803_
	);
	LUT4 #(
		.INIT('h0001)
	) name3756 (
		_w5795_,
		_w7801_,
		_w7802_,
		_w7803_,
		_w7804_
	);
	LUT3 #(
		.INIT('h40)
	) name3757 (
		_w7795_,
		_w7800_,
		_w7804_,
		_w7805_
	);
	LUT3 #(
		.INIT('h80)
	) name3758 (
		\bdma_BEAD_reg[7]/NET0131 ,
		_w5629_,
		_w5644_,
		_w7806_
	);
	LUT3 #(
		.INIT('h80)
	) name3759 (
		\bdma_BCTL_reg[7]/NET0131 ,
		_w5627_,
		_w5629_,
		_w7807_
	);
	LUT2 #(
		.INIT('h1)
	) name3760 (
		_w7806_,
		_w7807_,
		_w7808_
	);
	LUT2 #(
		.INIT('h8)
	) name3761 (
		_w7805_,
		_w7808_,
		_w7809_
	);
	LUT4 #(
		.INIT('h8000)
	) name3762 (
		\bdma_BOVL_reg[7]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w7810_
	);
	LUT4 #(
		.INIT('h8000)
	) name3763 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w7811_
	);
	LUT3 #(
		.INIT('h80)
	) name3764 (
		\pio_pmask_reg_DO_reg[7]/NET0131 ,
		_w5628_,
		_w5660_,
		_w7812_
	);
	LUT3 #(
		.INIT('h80)
	) name3765 (
		\sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w5648_,
		_w5634_,
		_w7813_
	);
	LUT3 #(
		.INIT('h80)
	) name3766 (
		\sport0_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w5634_,
		_w5660_,
		_w7814_
	);
	LUT3 #(
		.INIT('h80)
	) name3767 (
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w5632_,
		_w5634_,
		_w7815_
	);
	LUT4 #(
		.INIT('h0001)
	) name3768 (
		_w7812_,
		_w7813_,
		_w7814_,
		_w7815_,
		_w7816_
	);
	LUT3 #(
		.INIT('h80)
	) name3769 (
		\idma_DOVL_reg[7]/NET0131 ,
		_w5804_,
		_w5824_,
		_w7817_
	);
	LUT3 #(
		.INIT('h80)
	) name3770 (
		\tm_tsr_reg_DO_reg[7]/NET0131 ,
		_w5627_,
		_w5631_,
		_w7818_
	);
	LUT3 #(
		.INIT('h80)
	) name3771 (
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w5634_,
		_w5639_,
		_w7819_
	);
	LUT3 #(
		.INIT('h80)
	) name3772 (
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w5634_,
		_w5637_,
		_w7820_
	);
	LUT4 #(
		.INIT('h0001)
	) name3773 (
		_w7817_,
		_w7818_,
		_w7819_,
		_w7820_,
		_w7821_
	);
	LUT3 #(
		.INIT('h80)
	) name3774 (
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w5644_,
		_w5634_,
		_w7822_
	);
	LUT3 #(
		.INIT('h80)
	) name3775 (
		\PIO_out[7]_pad ,
		_w5628_,
		_w5635_,
		_w7823_
	);
	LUT3 #(
		.INIT('h80)
	) name3776 (
		\PIO_oe[7]_pad ,
		_w5628_,
		_w5632_,
		_w7824_
	);
	LUT3 #(
		.INIT('h80)
	) name3777 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w5628_,
		_w5639_,
		_w7825_
	);
	LUT4 #(
		.INIT('h0001)
	) name3778 (
		_w7822_,
		_w7823_,
		_w7824_,
		_w7825_,
		_w7826_
	);
	LUT3 #(
		.INIT('h80)
	) name3779 (
		\sport1_regs_AUTOreg_DO_reg[7]/NET0131 ,
		_w5670_,
		_w5810_,
		_w7827_
	);
	LUT3 #(
		.INIT('h80)
	) name3780 (
		\clkc_ckr_reg_DO_reg[7]/NET0131 ,
		_w5631_,
		_w5644_,
		_w7828_
	);
	LUT3 #(
		.INIT('h80)
	) name3781 (
		\memc_usysr_DO_reg[7]/NET0131 ,
		_w5631_,
		_w5660_,
		_w7829_
	);
	LUT3 #(
		.INIT('h80)
	) name3782 (
		\pio_PINT_reg[7]/NET0131 ,
		_w5670_,
		_w5672_,
		_w7830_
	);
	LUT4 #(
		.INIT('h0001)
	) name3783 (
		_w7827_,
		_w7828_,
		_w7829_,
		_w7830_,
		_w7831_
	);
	LUT4 #(
		.INIT('h8000)
	) name3784 (
		_w7826_,
		_w7831_,
		_w7816_,
		_w7821_,
		_w7832_
	);
	LUT3 #(
		.INIT('h10)
	) name3785 (
		_w7811_,
		_w7810_,
		_w7832_,
		_w7833_
	);
	LUT3 #(
		.INIT('h2a)
	) name3786 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w7809_,
		_w7833_,
		_w7834_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3787 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4263_,
		_w4260_,
		_w4268_,
		_w7835_
	);
	LUT2 #(
		.INIT('h8)
	) name3788 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w7836_
	);
	LUT4 #(
		.INIT('h153f)
	) name3789 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[7]/NET0131 ,
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w7837_
	);
	LUT3 #(
		.INIT('ha8)
	) name3790 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w7838_
	);
	LUT4 #(
		.INIT('h135f)
	) name3791 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w7839_
	);
	LUT4 #(
		.INIT('h1000)
	) name3792 (
		_w7838_,
		_w7836_,
		_w7839_,
		_w7837_,
		_w7840_
	);
	LUT3 #(
		.INIT('h8a)
	) name3793 (
		_w5681_,
		_w7835_,
		_w7840_,
		_w7841_
	);
	LUT4 #(
		.INIT('h135f)
	) name3794 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131 ,
		_w7842_
	);
	LUT4 #(
		.INIT('h135f)
	) name3795 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131 ,
		_w7843_
	);
	LUT2 #(
		.INIT('h8)
	) name3796 (
		_w7842_,
		_w7843_,
		_w7844_
	);
	LUT4 #(
		.INIT('h135f)
	) name3797 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131 ,
		_w7845_
	);
	LUT4 #(
		.INIT('h135f)
	) name3798 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131 ,
		_w7846_
	);
	LUT4 #(
		.INIT('h135f)
	) name3799 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131 ,
		_w7847_
	);
	LUT4 #(
		.INIT('h135f)
	) name3800 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131 ,
		_w7848_
	);
	LUT4 #(
		.INIT('h8000)
	) name3801 (
		_w7847_,
		_w7848_,
		_w7845_,
		_w7846_,
		_w7849_
	);
	LUT3 #(
		.INIT('h2a)
	) name3802 (
		_w5687_,
		_w7844_,
		_w7849_,
		_w7850_
	);
	LUT4 #(
		.INIT('h135f)
	) name3803 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 ,
		_w7851_
	);
	LUT4 #(
		.INIT('h135f)
	) name3804 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131 ,
		_w7852_
	);
	LUT2 #(
		.INIT('h8)
	) name3805 (
		_w7851_,
		_w7852_,
		_w7853_
	);
	LUT4 #(
		.INIT('h135f)
	) name3806 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131 ,
		_w7854_
	);
	LUT4 #(
		.INIT('h135f)
	) name3807 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131 ,
		_w7855_
	);
	LUT4 #(
		.INIT('h135f)
	) name3808 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131 ,
		_w7856_
	);
	LUT4 #(
		.INIT('h135f)
	) name3809 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131 ,
		_w7857_
	);
	LUT4 #(
		.INIT('h8000)
	) name3810 (
		_w7856_,
		_w7857_,
		_w7854_,
		_w7855_,
		_w7858_
	);
	LUT4 #(
		.INIT('h135f)
	) name3811 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[7]/P0001 ,
		\sport1_txctl_TX_reg[7]/P0001 ,
		_w7859_
	);
	LUT4 #(
		.INIT('h135f)
	) name3812 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[7]/P0001 ,
		\sport1_rxctl_RX_reg[7]/P0001 ,
		_w7860_
	);
	LUT3 #(
		.INIT('h2a)
	) name3813 (
		_w5706_,
		_w7859_,
		_w7860_,
		_w7861_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3814 (
		_w5697_,
		_w7853_,
		_w7858_,
		_w7861_,
		_w7862_
	);
	LUT2 #(
		.INIT('h4)
	) name3815 (
		_w7850_,
		_w7862_,
		_w7863_
	);
	LUT3 #(
		.INIT('h1b)
	) name3816 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001 ,
		_w7864_
	);
	LUT4 #(
		.INIT('ha820)
	) name3817 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001 ,
		_w7865_
	);
	LUT3 #(
		.INIT('h1b)
	) name3818 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001 ,
		_w7866_
	);
	LUT4 #(
		.INIT('ha820)
	) name3819 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001 ,
		_w7867_
	);
	LUT3 #(
		.INIT('h1b)
	) name3820 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001 ,
		_w7868_
	);
	LUT4 #(
		.INIT('ha820)
	) name3821 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001 ,
		_w7869_
	);
	LUT3 #(
		.INIT('h01)
	) name3822 (
		_w7867_,
		_w7869_,
		_w7865_,
		_w7870_
	);
	LUT3 #(
		.INIT('h2a)
	) name3823 (
		_w5741_,
		_w5746_,
		_w7870_,
		_w7871_
	);
	LUT3 #(
		.INIT('h1b)
	) name3824 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001 ,
		_w7872_
	);
	LUT4 #(
		.INIT('ha820)
	) name3825 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001 ,
		_w7873_
	);
	LUT2 #(
		.INIT('h8)
	) name3826 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w7874_
	);
	LUT2 #(
		.INIT('h1)
	) name3827 (
		_w7873_,
		_w7874_,
		_w7875_
	);
	LUT3 #(
		.INIT('h1b)
	) name3828 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001 ,
		_w7876_
	);
	LUT4 #(
		.INIT('ha820)
	) name3829 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001 ,
		_w7877_
	);
	LUT3 #(
		.INIT('h1b)
	) name3830 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001 ,
		_w7878_
	);
	LUT4 #(
		.INIT('ha820)
	) name3831 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001 ,
		_w7879_
	);
	LUT4 #(
		.INIT('ha820)
	) name3832 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001 ,
		_w7880_
	);
	LUT4 #(
		.INIT('ha820)
	) name3833 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001 ,
		_w7881_
	);
	LUT4 #(
		.INIT('h0001)
	) name3834 (
		_w7877_,
		_w7879_,
		_w7880_,
		_w7881_,
		_w7882_
	);
	LUT3 #(
		.INIT('h2a)
	) name3835 (
		_w5730_,
		_w7875_,
		_w7882_,
		_w7883_
	);
	LUT3 #(
		.INIT('h1b)
	) name3836 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 ,
		_w7884_
	);
	LUT4 #(
		.INIT('ha820)
	) name3837 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 ,
		_w7885_
	);
	LUT3 #(
		.INIT('h1b)
	) name3838 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001 ,
		_w7886_
	);
	LUT4 #(
		.INIT('ha820)
	) name3839 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001 ,
		_w7887_
	);
	LUT3 #(
		.INIT('h1b)
	) name3840 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001 ,
		_w7888_
	);
	LUT4 #(
		.INIT('ha820)
	) name3841 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001 ,
		_w7889_
	);
	LUT3 #(
		.INIT('h01)
	) name3842 (
		_w7887_,
		_w7889_,
		_w7885_,
		_w7890_
	);
	LUT3 #(
		.INIT('h1b)
	) name3843 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001 ,
		_w7891_
	);
	LUT4 #(
		.INIT('ha820)
	) name3844 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001 ,
		_w7892_
	);
	LUT3 #(
		.INIT('h1b)
	) name3845 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001 ,
		_w7893_
	);
	LUT4 #(
		.INIT('ha820)
	) name3846 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001 ,
		_w7894_
	);
	LUT3 #(
		.INIT('h1b)
	) name3847 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001 ,
		_w7895_
	);
	LUT4 #(
		.INIT('ha820)
	) name3848 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001 ,
		_w7896_
	);
	LUT4 #(
		.INIT('h0001)
	) name3849 (
		_w5714_,
		_w7892_,
		_w7894_,
		_w7896_,
		_w7897_
	);
	LUT3 #(
		.INIT('h2a)
	) name3850 (
		_w5712_,
		_w7890_,
		_w7897_,
		_w7898_
	);
	LUT3 #(
		.INIT('h01)
	) name3851 (
		_w7883_,
		_w7898_,
		_w7871_,
		_w7899_
	);
	LUT2 #(
		.INIT('h8)
	) name3852 (
		_w7863_,
		_w7899_,
		_w7900_
	);
	LUT2 #(
		.INIT('h4)
	) name3853 (
		_w7841_,
		_w7900_,
		_w7901_
	);
	LUT3 #(
		.INIT('h10)
	) name3854 (
		_w7794_,
		_w7834_,
		_w7901_,
		_w7902_
	);
	LUT4 #(
		.INIT('h5455)
	) name3855 (
		\emc_DMDoe_reg/NET0131 ,
		_w7794_,
		_w7834_,
		_w7901_,
		_w7903_
	);
	LUT2 #(
		.INIT('h8)
	) name3856 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[7]/P0001 ,
		_w7904_
	);
	LUT3 #(
		.INIT('h08)
	) name3857 (
		_w5588_,
		_w5598_,
		_w7904_,
		_w7905_
	);
	LUT3 #(
		.INIT('h45)
	) name3858 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w7906_
	);
	LUT4 #(
		.INIT('hecfd)
	) name3859 (
		_w5117_,
		_w5337_,
		_w7780_,
		_w7906_,
		_w7907_
	);
	LUT2 #(
		.INIT('h2)
	) name3860 (
		_w5586_,
		_w7907_,
		_w7908_
	);
	LUT2 #(
		.INIT('h9)
	) name3861 (
		_w5200_,
		_w5204_,
		_w7909_
	);
	LUT4 #(
		.INIT('hd02f)
	) name3862 (
		_w5226_,
		_w5193_,
		_w5229_,
		_w7909_,
		_w7910_
	);
	LUT3 #(
		.INIT('he0)
	) name3863 (
		_w5767_,
		_w5918_,
		_w7910_,
		_w7911_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3864 (
		\core_dag_ilm1reg_I_reg[6]/NET0131 ,
		_w5195_,
		_w5158_,
		_w5194_,
		_w7912_
	);
	LUT2 #(
		.INIT('h6)
	) name3865 (
		_w5198_,
		_w5300_,
		_w7913_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name3866 (
		_w5767_,
		_w5918_,
		_w7912_,
		_w7913_,
		_w7914_
	);
	LUT3 #(
		.INIT('ha8)
	) name3867 (
		\DM_rd0[6]_pad ,
		_w5610_,
		_w5612_,
		_w7915_
	);
	LUT4 #(
		.INIT('h135f)
	) name3868 (
		\DM_rdm[6]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w7916_
	);
	LUT4 #(
		.INIT('h135f)
	) name3869 (
		\DM_rd6[6]_pad ,
		\DM_rd7[6]_pad ,
		_w5596_,
		_w5591_,
		_w7917_
	);
	LUT2 #(
		.INIT('h8)
	) name3870 (
		_w7916_,
		_w7917_,
		_w7918_
	);
	LUT3 #(
		.INIT('h80)
	) name3871 (
		\DM_rd5[6]_pad ,
		_w5598_,
		_w5599_,
		_w7919_
	);
	LUT3 #(
		.INIT('h80)
	) name3872 (
		\DM_rd4[6]_pad ,
		_w5598_,
		_w5601_,
		_w7920_
	);
	LUT4 #(
		.INIT('h8000)
	) name3873 (
		\DM_rd2[6]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w7921_
	);
	LUT4 #(
		.INIT('h8000)
	) name3874 (
		\DM_rd1[6]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w7922_
	);
	LUT4 #(
		.INIT('h8000)
	) name3875 (
		\DM_rd3[6]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w7923_
	);
	LUT3 #(
		.INIT('h01)
	) name3876 (
		_w7922_,
		_w7923_,
		_w7921_,
		_w7924_
	);
	LUT3 #(
		.INIT('h10)
	) name3877 (
		_w7920_,
		_w7919_,
		_w7924_,
		_w7925_
	);
	LUT2 #(
		.INIT('h8)
	) name3878 (
		_w7918_,
		_w7925_,
		_w7926_
	);
	LUT2 #(
		.INIT('h4)
	) name3879 (
		_w7915_,
		_w7926_,
		_w7927_
	);
	LUT4 #(
		.INIT('h4000)
	) name3880 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[6]/P0001 ,
		_w7928_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3881 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4145_,
		_w4154_,
		_w7929_
	);
	LUT4 #(
		.INIT('ha820)
	) name3882 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001 ,
		_w7930_
	);
	LUT3 #(
		.INIT('h1b)
	) name3883 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001 ,
		_w7931_
	);
	LUT4 #(
		.INIT('ha820)
	) name3884 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001 ,
		_w7932_
	);
	LUT2 #(
		.INIT('h1)
	) name3885 (
		_w7930_,
		_w7932_,
		_w7933_
	);
	LUT3 #(
		.INIT('h1b)
	) name3886 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001 ,
		_w7934_
	);
	LUT4 #(
		.INIT('ha820)
	) name3887 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001 ,
		_w7935_
	);
	LUT3 #(
		.INIT('h1b)
	) name3888 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001 ,
		_w7936_
	);
	LUT4 #(
		.INIT('ha820)
	) name3889 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001 ,
		_w7937_
	);
	LUT4 #(
		.INIT('ha820)
	) name3890 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001 ,
		_w7938_
	);
	LUT3 #(
		.INIT('h01)
	) name3891 (
		_w7937_,
		_w7938_,
		_w7935_,
		_w7939_
	);
	LUT2 #(
		.INIT('h8)
	) name3892 (
		_w7933_,
		_w7939_,
		_w7940_
	);
	LUT3 #(
		.INIT('h8a)
	) name3893 (
		_w5730_,
		_w7929_,
		_w7940_,
		_w7941_
	);
	LUT3 #(
		.INIT('h80)
	) name3894 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w5629_,
		_w5648_,
		_w7942_
	);
	LUT3 #(
		.INIT('h80)
	) name3895 (
		\emc_WSCRreg_DO_reg[6]/NET0131 ,
		_w5631_,
		_w5632_,
		_w7943_
	);
	LUT3 #(
		.INIT('h80)
	) name3896 (
		\tm_TCR_TMP_reg[6]/NET0131 ,
		_w5631_,
		_w5637_,
		_w7944_
	);
	LUT3 #(
		.INIT('h80)
	) name3897 (
		\sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w5634_,
		_w5635_,
		_w7945_
	);
	LUT3 #(
		.INIT('h80)
	) name3898 (
		\sport0_regs_AUTOreg_DO_reg[6]/NET0131 ,
		_w5627_,
		_w5634_,
		_w7946_
	);
	LUT4 #(
		.INIT('h0001)
	) name3899 (
		_w7943_,
		_w7944_,
		_w7945_,
		_w7946_,
		_w7947_
	);
	LUT3 #(
		.INIT('h80)
	) name3900 (
		\sport1_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w5631_,
		_w5639_,
		_w7948_
	);
	LUT3 #(
		.INIT('h80)
	) name3901 (
		\emc_WSCRext_reg_DO_reg[6]/NET0131 ,
		_w5670_,
		_w5790_,
		_w7949_
	);
	LUT3 #(
		.INIT('h80)
	) name3902 (
		\tm_tpr_reg_DO_reg[6]/NET0131 ,
		_w5631_,
		_w5635_,
		_w7950_
	);
	LUT4 #(
		.INIT('h0001)
	) name3903 (
		_w5795_,
		_w7948_,
		_w7949_,
		_w7950_,
		_w7951_
	);
	LUT3 #(
		.INIT('h40)
	) name3904 (
		_w7942_,
		_w7947_,
		_w7951_,
		_w7952_
	);
	LUT3 #(
		.INIT('h80)
	) name3905 (
		\bdma_BEAD_reg[6]/NET0131 ,
		_w5629_,
		_w5644_,
		_w7953_
	);
	LUT3 #(
		.INIT('h80)
	) name3906 (
		\bdma_BCTL_reg[6]/NET0131 ,
		_w5627_,
		_w5629_,
		_w7954_
	);
	LUT2 #(
		.INIT('h1)
	) name3907 (
		_w7953_,
		_w7954_,
		_w7955_
	);
	LUT2 #(
		.INIT('h8)
	) name3908 (
		_w7952_,
		_w7955_,
		_w7956_
	);
	LUT4 #(
		.INIT('h8000)
	) name3909 (
		\bdma_BOVL_reg[6]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5658_,
		_w5804_,
		_w7957_
	);
	LUT4 #(
		.INIT('h8000)
	) name3910 (
		\bdma_BWCOUNT_reg[6]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w5657_,
		_w5658_,
		_w7958_
	);
	LUT3 #(
		.INIT('h80)
	) name3911 (
		\pio_pmask_reg_DO_reg[6]/NET0131 ,
		_w5628_,
		_w5660_,
		_w7959_
	);
	LUT3 #(
		.INIT('h80)
	) name3912 (
		\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w5648_,
		_w5634_,
		_w7960_
	);
	LUT3 #(
		.INIT('h80)
	) name3913 (
		\sport0_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w5634_,
		_w5660_,
		_w7961_
	);
	LUT3 #(
		.INIT('h80)
	) name3914 (
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w5632_,
		_w5634_,
		_w7962_
	);
	LUT4 #(
		.INIT('h0001)
	) name3915 (
		_w7959_,
		_w7960_,
		_w7961_,
		_w7962_,
		_w7963_
	);
	LUT3 #(
		.INIT('h80)
	) name3916 (
		\idma_DOVL_reg[6]/NET0131 ,
		_w5804_,
		_w5824_,
		_w7964_
	);
	LUT3 #(
		.INIT('h80)
	) name3917 (
		\tm_tsr_reg_DO_reg[6]/NET0131 ,
		_w5627_,
		_w5631_,
		_w7965_
	);
	LUT3 #(
		.INIT('h80)
	) name3918 (
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w5634_,
		_w5639_,
		_w7966_
	);
	LUT3 #(
		.INIT('h80)
	) name3919 (
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w5634_,
		_w5637_,
		_w7967_
	);
	LUT4 #(
		.INIT('h0001)
	) name3920 (
		_w7964_,
		_w7965_,
		_w7966_,
		_w7967_,
		_w7968_
	);
	LUT3 #(
		.INIT('h80)
	) name3921 (
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w5644_,
		_w5634_,
		_w7969_
	);
	LUT3 #(
		.INIT('h80)
	) name3922 (
		\PIO_out[6]_pad ,
		_w5628_,
		_w5635_,
		_w7970_
	);
	LUT3 #(
		.INIT('h80)
	) name3923 (
		\PIO_oe[6]_pad ,
		_w5628_,
		_w5632_,
		_w7971_
	);
	LUT3 #(
		.INIT('h80)
	) name3924 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w5628_,
		_w5639_,
		_w7972_
	);
	LUT4 #(
		.INIT('h0001)
	) name3925 (
		_w7969_,
		_w7970_,
		_w7971_,
		_w7972_,
		_w7973_
	);
	LUT3 #(
		.INIT('h80)
	) name3926 (
		\sport1_regs_AUTOreg_DO_reg[6]/NET0131 ,
		_w5670_,
		_w5810_,
		_w7974_
	);
	LUT3 #(
		.INIT('h80)
	) name3927 (
		\clkc_ckr_reg_DO_reg[6]/NET0131 ,
		_w5631_,
		_w5644_,
		_w7975_
	);
	LUT3 #(
		.INIT('h80)
	) name3928 (
		\memc_usysr_DO_reg[6]/NET0131 ,
		_w5631_,
		_w5660_,
		_w7976_
	);
	LUT3 #(
		.INIT('h80)
	) name3929 (
		\pio_PINT_reg[6]/NET0131 ,
		_w5670_,
		_w5672_,
		_w7977_
	);
	LUT4 #(
		.INIT('h0001)
	) name3930 (
		_w7974_,
		_w7975_,
		_w7976_,
		_w7977_,
		_w7978_
	);
	LUT4 #(
		.INIT('h8000)
	) name3931 (
		_w7973_,
		_w7978_,
		_w7963_,
		_w7968_,
		_w7979_
	);
	LUT3 #(
		.INIT('h10)
	) name3932 (
		_w7958_,
		_w7957_,
		_w7979_,
		_w7980_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3933 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4295_,
		_w4292_,
		_w4300_,
		_w7981_
	);
	LUT4 #(
		.INIT('h153f)
	) name3934 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w7982_
	);
	LUT4 #(
		.INIT('h135f)
	) name3935 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		\core_c_psq_SSTAT_reg[6]/NET0131 ,
		_w7983_
	);
	LUT3 #(
		.INIT('ha8)
	) name3936 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w7984_
	);
	LUT4 #(
		.INIT('h135f)
	) name3937 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w7985_
	);
	LUT4 #(
		.INIT('h4000)
	) name3938 (
		_w7984_,
		_w7985_,
		_w7982_,
		_w7983_,
		_w7986_
	);
	LUT4 #(
		.INIT('h135f)
	) name3939 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w7987_
	);
	LUT4 #(
		.INIT('h135f)
	) name3940 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w7988_
	);
	LUT2 #(
		.INIT('h8)
	) name3941 (
		_w7987_,
		_w7988_,
		_w7989_
	);
	LUT4 #(
		.INIT('h135f)
	) name3942 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131 ,
		_w7990_
	);
	LUT4 #(
		.INIT('h135f)
	) name3943 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131 ,
		_w7991_
	);
	LUT4 #(
		.INIT('h135f)
	) name3944 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131 ,
		_w7992_
	);
	LUT4 #(
		.INIT('h135f)
	) name3945 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131 ,
		_w7993_
	);
	LUT4 #(
		.INIT('h8000)
	) name3946 (
		_w7992_,
		_w7993_,
		_w7990_,
		_w7991_,
		_w7994_
	);
	LUT3 #(
		.INIT('h2a)
	) name3947 (
		_w5687_,
		_w7989_,
		_w7994_,
		_w7995_
	);
	LUT4 #(
		.INIT('h135f)
	) name3948 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131 ,
		_w7996_
	);
	LUT4 #(
		.INIT('h135f)
	) name3949 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131 ,
		_w7997_
	);
	LUT2 #(
		.INIT('h8)
	) name3950 (
		_w7996_,
		_w7997_,
		_w7998_
	);
	LUT4 #(
		.INIT('h135f)
	) name3951 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131 ,
		_w7999_
	);
	LUT4 #(
		.INIT('h135f)
	) name3952 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131 ,
		_w8000_
	);
	LUT4 #(
		.INIT('h135f)
	) name3953 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 ,
		_w8001_
	);
	LUT4 #(
		.INIT('h135f)
	) name3954 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 ,
		_w8002_
	);
	LUT4 #(
		.INIT('h8000)
	) name3955 (
		_w8001_,
		_w8002_,
		_w7999_,
		_w8000_,
		_w8003_
	);
	LUT4 #(
		.INIT('h135f)
	) name3956 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[6]/P0001 ,
		\sport1_txctl_TX_reg[6]/P0001 ,
		_w8004_
	);
	LUT4 #(
		.INIT('h135f)
	) name3957 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		\sport1_rxctl_RX_reg[6]/P0001 ,
		_w8005_
	);
	LUT3 #(
		.INIT('h2a)
	) name3958 (
		_w5706_,
		_w8004_,
		_w8005_,
		_w8006_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3959 (
		_w5697_,
		_w7998_,
		_w8003_,
		_w8006_,
		_w8007_
	);
	LUT3 #(
		.INIT('h1b)
	) name3960 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001 ,
		_w8008_
	);
	LUT4 #(
		.INIT('ha820)
	) name3961 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001 ,
		_w8009_
	);
	LUT2 #(
		.INIT('h1)
	) name3962 (
		_w5743_,
		_w8009_,
		_w8010_
	);
	LUT3 #(
		.INIT('h1b)
	) name3963 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001 ,
		_w8011_
	);
	LUT4 #(
		.INIT('ha820)
	) name3964 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001 ,
		_w8012_
	);
	LUT3 #(
		.INIT('h1b)
	) name3965 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001 ,
		_w8013_
	);
	LUT4 #(
		.INIT('ha820)
	) name3966 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001 ,
		_w8014_
	);
	LUT3 #(
		.INIT('h1b)
	) name3967 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001 ,
		_w8015_
	);
	LUT4 #(
		.INIT('ha820)
	) name3968 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001 ,
		_w8016_
	);
	LUT3 #(
		.INIT('h01)
	) name3969 (
		_w8014_,
		_w8016_,
		_w8012_,
		_w8017_
	);
	LUT3 #(
		.INIT('h2a)
	) name3970 (
		_w5741_,
		_w8010_,
		_w8017_,
		_w8018_
	);
	LUT3 #(
		.INIT('h1b)
	) name3971 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 ,
		_w8019_
	);
	LUT4 #(
		.INIT('ha820)
	) name3972 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 ,
		_w8020_
	);
	LUT3 #(
		.INIT('h1b)
	) name3973 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001 ,
		_w8021_
	);
	LUT4 #(
		.INIT('ha820)
	) name3974 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001 ,
		_w8022_
	);
	LUT3 #(
		.INIT('h1b)
	) name3975 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001 ,
		_w8023_
	);
	LUT4 #(
		.INIT('ha820)
	) name3976 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001 ,
		_w8024_
	);
	LUT3 #(
		.INIT('h01)
	) name3977 (
		_w8022_,
		_w8024_,
		_w8020_,
		_w8025_
	);
	LUT3 #(
		.INIT('h1b)
	) name3978 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001 ,
		_w8026_
	);
	LUT4 #(
		.INIT('ha820)
	) name3979 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001 ,
		_w8027_
	);
	LUT3 #(
		.INIT('h1b)
	) name3980 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001 ,
		_w8028_
	);
	LUT4 #(
		.INIT('ha820)
	) name3981 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001 ,
		_w8029_
	);
	LUT3 #(
		.INIT('h1b)
	) name3982 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001 ,
		_w8030_
	);
	LUT4 #(
		.INIT('ha820)
	) name3983 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001 ,
		_w8031_
	);
	LUT3 #(
		.INIT('h1b)
	) name3984 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001 ,
		_w8032_
	);
	LUT4 #(
		.INIT('ha820)
	) name3985 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001 ,
		_w8033_
	);
	LUT4 #(
		.INIT('h0001)
	) name3986 (
		_w8027_,
		_w8029_,
		_w8031_,
		_w8033_,
		_w8034_
	);
	LUT3 #(
		.INIT('h2a)
	) name3987 (
		_w5712_,
		_w8025_,
		_w8034_,
		_w8035_
	);
	LUT4 #(
		.INIT('h0100)
	) name3988 (
		_w8018_,
		_w8035_,
		_w7995_,
		_w8007_,
		_w8036_
	);
	LUT4 #(
		.INIT('h7500)
	) name3989 (
		_w5681_,
		_w7981_,
		_w7986_,
		_w8036_,
		_w8037_
	);
	LUT4 #(
		.INIT('hd500)
	) name3990 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w7956_,
		_w7980_,
		_w8037_,
		_w8038_
	);
	LUT3 #(
		.INIT('h10)
	) name3991 (
		_w7928_,
		_w7941_,
		_w8038_,
		_w8039_
	);
	LUT4 #(
		.INIT('h5455)
	) name3992 (
		\emc_DMDoe_reg/NET0131 ,
		_w7928_,
		_w7941_,
		_w8038_,
		_w8040_
	);
	LUT2 #(
		.INIT('h8)
	) name3993 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[6]/P0001 ,
		_w8041_
	);
	LUT3 #(
		.INIT('h08)
	) name3994 (
		_w5588_,
		_w5598_,
		_w8041_,
		_w8042_
	);
	LUT3 #(
		.INIT('h45)
	) name3995 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w8043_
	);
	LUT4 #(
		.INIT('hc040)
	) name3996 (
		_w5117_,
		_w5337_,
		_w5586_,
		_w8043_,
		_w8044_
	);
	LUT4 #(
		.INIT('hef00)
	) name3997 (
		_w5117_,
		_w7911_,
		_w7914_,
		_w8044_,
		_w8045_
	);
	LUT2 #(
		.INIT('h1)
	) name3998 (
		_w7908_,
		_w8045_,
		_w8046_
	);
	LUT4 #(
		.INIT('h2f00)
	) name3999 (
		_w5117_,
		_w7732_,
		_w7779_,
		_w8046_,
		_w8047_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name4000 (
		_w5117_,
		_w7732_,
		_w7779_,
		_w8046_,
		_w8048_
	);
	LUT3 #(
		.INIT('h8a)
	) name4001 (
		_w5337_,
		_w7911_,
		_w7914_,
		_w8049_
	);
	LUT2 #(
		.INIT('h9)
	) name4002 (
		_w5446_,
		_w5448_,
		_w8050_
	);
	LUT4 #(
		.INIT('hba45)
	) name4003 (
		_w5453_,
		_w5465_,
		_w7717_,
		_w8050_,
		_w8051_
	);
	LUT3 #(
		.INIT('h10)
	) name4004 (
		_w5434_,
		_w6210_,
		_w8051_,
		_w8052_
	);
	LUT3 #(
		.INIT('h8a)
	) name4005 (
		\core_dag_ilm2reg_I_reg[7]/NET0131 ,
		_w5399_,
		_w5401_,
		_w8053_
	);
	LUT4 #(
		.INIT('h718e)
	) name4006 (
		\core_dag_ilm2reg_M_reg[6]/NET0131 ,
		_w5405_,
		_w5426_,
		_w5444_,
		_w8054_
	);
	LUT4 #(
		.INIT('h010f)
	) name4007 (
		_w5434_,
		_w6210_,
		_w8053_,
		_w8054_,
		_w8055_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4008 (
		_w5117_,
		_w5337_,
		_w8052_,
		_w8055_,
		_w8056_
	);
	LUT4 #(
		.INIT('h0200)
	) name4009 (
		\core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w8057_
	);
	LUT4 #(
		.INIT('h0200)
	) name4010 (
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w8058_
	);
	LUT4 #(
		.INIT('h0200)
	) name4011 (
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w8059_
	);
	LUT4 #(
		.INIT('h0200)
	) name4012 (
		\core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w8060_
	);
	LUT4 #(
		.INIT('h0001)
	) name4013 (
		_w8057_,
		_w8058_,
		_w8059_,
		_w8060_,
		_w8061_
	);
	LUT4 #(
		.INIT('h0200)
	) name4014 (
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w8062_
	);
	LUT4 #(
		.INIT('h0200)
	) name4015 (
		\core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w8063_
	);
	LUT4 #(
		.INIT('h0200)
	) name4016 (
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w8064_
	);
	LUT4 #(
		.INIT('h0200)
	) name4017 (
		\core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w8065_
	);
	LUT4 #(
		.INIT('h0001)
	) name4018 (
		_w8062_,
		_w8063_,
		_w8064_,
		_w8065_,
		_w8066_
	);
	LUT3 #(
		.INIT('hd0)
	) name4019 (
		_w4063_,
		_w8061_,
		_w8066_,
		_w8067_
	);
	LUT4 #(
		.INIT('h0233)
	) name4020 (
		_w4063_,
		_w5049_,
		_w8061_,
		_w8066_,
		_w8068_
	);
	LUT4 #(
		.INIT('h0080)
	) name4021 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w8069_
	);
	LUT4 #(
		.INIT('h000b)
	) name4022 (
		_w4970_,
		_w7777_,
		_w8068_,
		_w8069_,
		_w8070_
	);
	LUT4 #(
		.INIT('ha222)
	) name4023 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w8071_
	);
	LUT4 #(
		.INIT('h4000)
	) name4024 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w8072_
	);
	LUT4 #(
		.INIT('h2a00)
	) name4025 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w8073_
	);
	LUT2 #(
		.INIT('h1)
	) name4026 (
		_w8072_,
		_w8073_,
		_w8074_
	);
	LUT3 #(
		.INIT('h20)
	) name4027 (
		_w5539_,
		_w8071_,
		_w8074_,
		_w8075_
	);
	LUT3 #(
		.INIT('hd0)
	) name4028 (
		_w5059_,
		_w8070_,
		_w8075_,
		_w8076_
	);
	LUT4 #(
		.INIT('h5540)
	) name4029 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w8077_
	);
	LUT3 #(
		.INIT('h01)
	) name4030 (
		_w5337_,
		_w8077_,
		_w8076_,
		_w8078_
	);
	LUT3 #(
		.INIT('h15)
	) name4031 (
		_w5117_,
		_w5337_,
		_w7743_,
		_w8079_
	);
	LUT3 #(
		.INIT('h45)
	) name4032 (
		_w5586_,
		_w8078_,
		_w8079_,
		_w8080_
	);
	LUT3 #(
		.INIT('hb0)
	) name4033 (
		_w8049_,
		_w8056_,
		_w8080_,
		_w8081_
	);
	LUT4 #(
		.INIT('h4051)
	) name4034 (
		_w5117_,
		_w5337_,
		_w7731_,
		_w8043_,
		_w8082_
	);
	LUT2 #(
		.INIT('h4)
	) name4035 (
		_w7777_,
		_w8067_,
		_w8083_
	);
	LUT4 #(
		.INIT('h2a08)
	) name4036 (
		_w5117_,
		_w5337_,
		_w7906_,
		_w8083_,
		_w8084_
	);
	LUT2 #(
		.INIT('h2)
	) name4037 (
		_w5586_,
		_w8084_,
		_w8085_
	);
	LUT2 #(
		.INIT('h4)
	) name4038 (
		_w8082_,
		_w8085_,
		_w8086_
	);
	LUT2 #(
		.INIT('he)
	) name4039 (
		_w8081_,
		_w8086_,
		_w8087_
	);
	LUT4 #(
		.INIT('h80c4)
	) name4040 (
		_w5337_,
		_w5586_,
		_w7400_,
		_w7710_,
		_w8088_
	);
	LUT4 #(
		.INIT('h0200)
	) name4041 (
		\core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w8089_
	);
	LUT4 #(
		.INIT('h0200)
	) name4042 (
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w8090_
	);
	LUT4 #(
		.INIT('h0200)
	) name4043 (
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w8091_
	);
	LUT4 #(
		.INIT('h0200)
	) name4044 (
		\core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w8092_
	);
	LUT4 #(
		.INIT('h0001)
	) name4045 (
		_w8089_,
		_w8090_,
		_w8091_,
		_w8092_,
		_w8093_
	);
	LUT4 #(
		.INIT('h0200)
	) name4046 (
		\core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w8094_
	);
	LUT4 #(
		.INIT('h0200)
	) name4047 (
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w8095_
	);
	LUT4 #(
		.INIT('h0200)
	) name4048 (
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w8096_
	);
	LUT4 #(
		.INIT('h0200)
	) name4049 (
		\core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w8097_
	);
	LUT4 #(
		.INIT('h0001)
	) name4050 (
		_w8094_,
		_w8095_,
		_w8096_,
		_w8097_,
		_w8098_
	);
	LUT3 #(
		.INIT('hd0)
	) name4051 (
		_w4063_,
		_w8093_,
		_w8098_,
		_w8099_
	);
	LUT4 #(
		.INIT('h0233)
	) name4052 (
		_w4063_,
		_w5049_,
		_w8093_,
		_w8098_,
		_w8100_
	);
	LUT4 #(
		.INIT('h0080)
	) name4053 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w8101_
	);
	LUT4 #(
		.INIT('h000b)
	) name4054 (
		_w4970_,
		_w7449_,
		_w8100_,
		_w8101_,
		_w8102_
	);
	LUT4 #(
		.INIT('ha222)
	) name4055 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w8103_
	);
	LUT4 #(
		.INIT('h2a00)
	) name4056 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w8104_
	);
	LUT4 #(
		.INIT('h4000)
	) name4057 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w8105_
	);
	LUT2 #(
		.INIT('h1)
	) name4058 (
		_w8104_,
		_w8105_,
		_w8106_
	);
	LUT2 #(
		.INIT('h4)
	) name4059 (
		_w8103_,
		_w8106_,
		_w8107_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4060 (
		_w5059_,
		_w5539_,
		_w8102_,
		_w8107_,
		_w8108_
	);
	LUT4 #(
		.INIT('haa80)
	) name4061 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w8109_
	);
	LUT3 #(
		.INIT('h54)
	) name4062 (
		_w5337_,
		_w8108_,
		_w8109_,
		_w8110_
	);
	LUT3 #(
		.INIT('h13)
	) name4063 (
		_w5337_,
		_w5586_,
		_w7414_,
		_w8111_
	);
	LUT2 #(
		.INIT('h4)
	) name4064 (
		_w8110_,
		_w8111_,
		_w8112_
	);
	LUT3 #(
		.INIT('h54)
	) name4065 (
		_w5117_,
		_w8088_,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('h4)
	) name4066 (
		_w7449_,
		_w8099_,
		_w8114_
	);
	LUT4 #(
		.INIT('h4c08)
	) name4067 (
		_w5337_,
		_w5586_,
		_w7566_,
		_w8114_,
		_w8115_
	);
	LUT2 #(
		.INIT('h9)
	) name4068 (
		_w5494_,
		_w5496_,
		_w8116_
	);
	LUT3 #(
		.INIT('h1e)
	) name4069 (
		_w5467_,
		_w5488_,
		_w8116_,
		_w8117_
	);
	LUT3 #(
		.INIT('h10)
	) name4070 (
		_w5434_,
		_w6210_,
		_w8117_,
		_w8118_
	);
	LUT4 #(
		.INIT('haa20)
	) name4071 (
		\core_dag_ilm2reg_I_reg[8]/NET0131 ,
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		_w5393_,
		_w5396_,
		_w8119_
	);
	LUT3 #(
		.INIT('he1)
	) name4072 (
		_w5403_,
		_w5427_,
		_w5495_,
		_w8120_
	);
	LUT4 #(
		.INIT('h010f)
	) name4073 (
		_w5434_,
		_w6210_,
		_w8119_,
		_w8120_,
		_w8121_
	);
	LUT3 #(
		.INIT('h45)
	) name4074 (
		_w5337_,
		_w8118_,
		_w8121_,
		_w8122_
	);
	LUT3 #(
		.INIT('h31)
	) name4075 (
		_w5337_,
		_w5586_,
		_w7579_,
		_w8123_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4076 (
		_w5117_,
		_w8115_,
		_w8122_,
		_w8123_,
		_w8124_
	);
	LUT2 #(
		.INIT('h1)
	) name4077 (
		_w8113_,
		_w8124_,
		_w8125_
	);
	LUT3 #(
		.INIT('hc4)
	) name4078 (
		_w5117_,
		_w5337_,
		_w7241_,
		_w8126_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4079 (
		_w5117_,
		_w7062_,
		_w7067_,
		_w8126_,
		_w8127_
	);
	LUT4 #(
		.INIT('h0200)
	) name4080 (
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5039_,
		_w8128_
	);
	LUT4 #(
		.INIT('h0200)
	) name4081 (
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5035_,
		_w8129_
	);
	LUT4 #(
		.INIT('h0200)
	) name4082 (
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5037_,
		_w8130_
	);
	LUT4 #(
		.INIT('h0200)
	) name4083 (
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		_w4976_,
		_w4978_,
		_w5033_,
		_w8131_
	);
	LUT4 #(
		.INIT('h0001)
	) name4084 (
		_w8128_,
		_w8129_,
		_w8130_,
		_w8131_,
		_w8132_
	);
	LUT4 #(
		.INIT('h0200)
	) name4085 (
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		_w4976_,
		_w4978_,
		_w4999_,
		_w8133_
	);
	LUT4 #(
		.INIT('h0200)
	) name4086 (
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		_w5004_,
		_w5006_,
		_w5009_,
		_w8134_
	);
	LUT4 #(
		.INIT('h0200)
	) name4087 (
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		_w5013_,
		_w5014_,
		_w5016_,
		_w8135_
	);
	LUT4 #(
		.INIT('h0200)
	) name4088 (
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		_w5020_,
		_w5021_,
		_w5023_,
		_w8136_
	);
	LUT4 #(
		.INIT('h0001)
	) name4089 (
		_w8133_,
		_w8134_,
		_w8135_,
		_w8136_,
		_w8137_
	);
	LUT3 #(
		.INIT('hd0)
	) name4090 (
		_w4063_,
		_w8132_,
		_w8137_,
		_w8138_
	);
	LUT2 #(
		.INIT('h4)
	) name4091 (
		_w7078_,
		_w8138_,
		_w8139_
	);
	LUT4 #(
		.INIT('hefcd)
	) name4092 (
		_w5117_,
		_w5337_,
		_w7378_,
		_w8139_,
		_w8140_
	);
	LUT3 #(
		.INIT('h8a)
	) name4093 (
		_w5586_,
		_w8127_,
		_w8140_,
		_w8141_
	);
	LUT4 #(
		.INIT('h0233)
	) name4094 (
		_w4063_,
		_w5049_,
		_w8132_,
		_w8137_,
		_w8142_
	);
	LUT4 #(
		.INIT('h0080)
	) name4095 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w8143_
	);
	LUT4 #(
		.INIT('h000b)
	) name4096 (
		_w4970_,
		_w7078_,
		_w8142_,
		_w8143_,
		_w8144_
	);
	LUT4 #(
		.INIT('ha222)
	) name4097 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		_w5569_,
		_w5570_,
		_w5571_,
		_w8145_
	);
	LUT4 #(
		.INIT('h4000)
	) name4098 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w8146_
	);
	LUT4 #(
		.INIT('h2a00)
	) name4099 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w4067_,
		_w4845_,
		_w5573_,
		_w8147_
	);
	LUT2 #(
		.INIT('h1)
	) name4100 (
		_w8146_,
		_w8147_,
		_w8148_
	);
	LUT2 #(
		.INIT('h4)
	) name4101 (
		_w8145_,
		_w8148_,
		_w8149_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4102 (
		_w5059_,
		_w5539_,
		_w8144_,
		_w8149_,
		_w8150_
	);
	LUT4 #(
		.INIT('haa80)
	) name4103 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w5530_,
		_w5534_,
		_w5538_,
		_w8151_
	);
	LUT3 #(
		.INIT('h01)
	) name4104 (
		_w5337_,
		_w8150_,
		_w8151_,
		_w8152_
	);
	LUT3 #(
		.INIT('h51)
	) name4105 (
		_w5117_,
		_w5337_,
		_w7109_,
		_w8153_
	);
	LUT2 #(
		.INIT('h4)
	) name4106 (
		_w8152_,
		_w8153_,
		_w8154_
	);
	LUT4 #(
		.INIT('h7771)
	) name4107 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		_w5397_,
		_w5403_,
		_w5427_,
		_w8155_
	);
	LUT2 #(
		.INIT('h9)
	) name4108 (
		_w5489_,
		_w8155_,
		_w8156_
	);
	LUT3 #(
		.INIT('he0)
	) name4109 (
		_w5434_,
		_w6210_,
		_w8156_,
		_w8157_
	);
	LUT3 #(
		.INIT('ha8)
	) name4110 (
		\core_dag_ilm2reg_I_reg[9]/NET0131 ,
		_w5392_,
		_w5393_,
		_w8158_
	);
	LUT2 #(
		.INIT('h9)
	) name4111 (
		_w5491_,
		_w5493_,
		_w8159_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4112 (
		_w5467_,
		_w5488_,
		_w5497_,
		_w5510_,
		_w8160_
	);
	LUT2 #(
		.INIT('h9)
	) name4113 (
		_w8159_,
		_w8160_,
		_w8161_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name4114 (
		_w5434_,
		_w6210_,
		_w8158_,
		_w8161_,
		_w8162_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4115 (
		_w5117_,
		_w5337_,
		_w8157_,
		_w8162_,
		_w8163_
	);
	LUT4 #(
		.INIT('h5150)
	) name4116 (
		_w5586_,
		_w7127_,
		_w8154_,
		_w8163_,
		_w8164_
	);
	LUT2 #(
		.INIT('h1)
	) name4117 (
		_w8141_,
		_w8164_,
		_w8165_
	);
	LUT2 #(
		.INIT('he)
	) name4118 (
		_w8141_,
		_w8164_,
		_w8166_
	);
	LUT3 #(
		.INIT('h01)
	) name4119 (
		_w6570_,
		_w8113_,
		_w8124_,
		_w8167_
	);
	LUT4 #(
		.INIT('h1110)
	) name4120 (
		_w7713_,
		_w8047_,
		_w8081_,
		_w8086_,
		_w8168_
	);
	LUT3 #(
		.INIT('h01)
	) name4121 (
		_w6241_,
		_w6901_,
		_w6944_,
		_w8169_
	);
	LUT4 #(
		.INIT('h4000)
	) name4122 (
		_w8165_,
		_w8168_,
		_w8169_,
		_w8167_,
		_w8170_
	);
	LUT4 #(
		.INIT('h2000)
	) name4123 (
		\memc_Dread_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w8171_
	);
	LUT2 #(
		.INIT('h1)
	) name4124 (
		\core_c_dec_Long_Cg_reg/P0001 ,
		\core_c_dec_Prderr_Cg_reg/NET0131 ,
		_w8172_
	);
	LUT3 #(
		.INIT('h10)
	) name4125 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4428_,
		_w8172_,
		_w8173_
	);
	LUT4 #(
		.INIT('h0100)
	) name4126 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4104_,
		_w4428_,
		_w8172_,
		_w8174_
	);
	LUT4 #(
		.INIT('h4000)
	) name4127 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w5044_,
		_w5045_,
		_w5046_,
		_w8175_
	);
	LUT3 #(
		.INIT('h04)
	) name4128 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w4090_,
		_w4091_,
		_w8176_
	);
	LUT4 #(
		.INIT('h0040)
	) name4129 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w8177_
	);
	LUT4 #(
		.INIT('hf3bf)
	) name4130 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w8178_
	);
	LUT4 #(
		.INIT('hfb00)
	) name4131 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w4090_,
		_w4091_,
		_w8178_,
		_w8179_
	);
	LUT2 #(
		.INIT('h4)
	) name4132 (
		_w8175_,
		_w8179_,
		_w8180_
	);
	LUT4 #(
		.INIT('h3313)
	) name4133 (
		_w5058_,
		_w8171_,
		_w8174_,
		_w8180_,
		_w8181_
	);
	LUT2 #(
		.INIT('h8)
	) name4134 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_RDcyc_reg/NET0131 ,
		_w8182_
	);
	LUT4 #(
		.INIT('h2000)
	) name4135 (
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w8182_,
		_w8183_
	);
	LUT4 #(
		.INIT('haeaf)
	) name4136 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		\sport1_txctl_TSreq_reg/NET0131 ,
		_w8184_
	);
	LUT4 #(
		.INIT('h0700)
	) name4137 (
		_w4519_,
		_w5536_,
		_w8183_,
		_w8184_,
		_w8185_
	);
	LUT4 #(
		.INIT('h00df)
	) name4138 (
		_w4067_,
		_w4068_,
		_w4845_,
		_w8185_,
		_w8186_
	);
	LUT2 #(
		.INIT('h2)
	) name4139 (
		_w8181_,
		_w8186_,
		_w8187_
	);
	LUT3 #(
		.INIT('h47)
	) name4140 (
		\memc_Dwrite_C_reg/NET0131 ,
		_w4971_,
		_w5571_,
		_w8188_
	);
	LUT3 #(
		.INIT('h07)
	) name4141 (
		_w4061_,
		_w4062_,
		_w4984_,
		_w8189_
	);
	LUT4 #(
		.INIT('h00df)
	) name4142 (
		_w4067_,
		_w4068_,
		_w4845_,
		_w8189_,
		_w8190_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4143 (
		\idma_WRcyc_reg/NET0131 ,
		_w4067_,
		_w4068_,
		_w4845_,
		_w8191_
	);
	LUT4 #(
		.INIT('h0777)
	) name4144 (
		_w5530_,
		_w5534_,
		_w5573_,
		_w8191_,
		_w8192_
	);
	LUT3 #(
		.INIT('h20)
	) name4145 (
		_w8188_,
		_w8190_,
		_w8192_,
		_w8193_
	);
	LUT3 #(
		.INIT('h20)
	) name4146 (
		_w8181_,
		_w8186_,
		_w8193_,
		_w8194_
	);
	LUT3 #(
		.INIT('h01)
	) name4147 (
		_w6944_,
		_w8170_,
		_w8194_,
		_w8195_
	);
	LUT2 #(
		.INIT('h1)
	) name4148 (
		_w4088_,
		_w8189_,
		_w8196_
	);
	LUT2 #(
		.INIT('h2)
	) name4149 (
		_w8192_,
		_w8196_,
		_w8197_
	);
	LUT3 #(
		.INIT('h80)
	) name4150 (
		\bdma_BRdataBUF_reg[0]/P0001 ,
		_w5530_,
		_w5534_,
		_w8198_
	);
	LUT3 #(
		.INIT('h80)
	) name4151 (
		\idma_DTMP_H_reg[0]/P0001 ,
		_w5573_,
		_w8191_,
		_w8199_
	);
	LUT3 #(
		.INIT('h20)
	) name4152 (
		\sport1_rxctl_RX_reg[0]/P0001 ,
		_w4088_,
		_w4980_,
		_w8200_
	);
	LUT3 #(
		.INIT('h20)
	) name4153 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		_w4088_,
		_w4984_,
		_w8201_
	);
	LUT2 #(
		.INIT('h1)
	) name4154 (
		_w8200_,
		_w8201_,
		_w8202_
	);
	LUT3 #(
		.INIT('h10)
	) name4155 (
		_w8199_,
		_w8198_,
		_w8202_,
		_w8203_
	);
	LUT3 #(
		.INIT('h4f)
	) name4156 (
		_w5910_,
		_w8197_,
		_w8203_,
		_w8204_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4157 (
		_w5938_,
		_w6035_,
		_w8192_,
		_w8196_,
		_w8205_
	);
	LUT3 #(
		.INIT('h80)
	) name4158 (
		\bdma_BRdataBUF_reg[10]/P0001 ,
		_w5530_,
		_w5534_,
		_w8206_
	);
	LUT3 #(
		.INIT('h80)
	) name4159 (
		\idma_DTMP_H_reg[10]/P0001 ,
		_w5573_,
		_w8191_,
		_w8207_
	);
	LUT3 #(
		.INIT('h20)
	) name4160 (
		\sport0_rxctl_RX_reg[10]/P0001 ,
		_w4088_,
		_w4984_,
		_w8208_
	);
	LUT3 #(
		.INIT('h20)
	) name4161 (
		\sport1_rxctl_RX_reg[10]/P0001 ,
		_w4088_,
		_w4980_,
		_w8209_
	);
	LUT2 #(
		.INIT('h1)
	) name4162 (
		_w8208_,
		_w8209_,
		_w8210_
	);
	LUT3 #(
		.INIT('h10)
	) name4163 (
		_w8207_,
		_w8206_,
		_w8210_,
		_w8211_
	);
	LUT2 #(
		.INIT('hb)
	) name4164 (
		_w8205_,
		_w8211_,
		_w8212_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4165 (
		_w6264_,
		_w6359_,
		_w8192_,
		_w8196_,
		_w8213_
	);
	LUT3 #(
		.INIT('h80)
	) name4166 (
		\bdma_BRdataBUF_reg[11]/P0001 ,
		_w5530_,
		_w5534_,
		_w8214_
	);
	LUT3 #(
		.INIT('h80)
	) name4167 (
		\idma_DTMP_H_reg[11]/P0001 ,
		_w5573_,
		_w8191_,
		_w8215_
	);
	LUT3 #(
		.INIT('h20)
	) name4168 (
		\sport1_rxctl_RX_reg[11]/P0001 ,
		_w4088_,
		_w4980_,
		_w8216_
	);
	LUT3 #(
		.INIT('h20)
	) name4169 (
		\sport0_rxctl_RX_reg[11]/P0001 ,
		_w4088_,
		_w4984_,
		_w8217_
	);
	LUT2 #(
		.INIT('h1)
	) name4170 (
		_w8216_,
		_w8217_,
		_w8218_
	);
	LUT3 #(
		.INIT('h10)
	) name4171 (
		_w8215_,
		_w8214_,
		_w8218_,
		_w8219_
	);
	LUT2 #(
		.INIT('hb)
	) name4172 (
		_w8213_,
		_w8219_,
		_w8220_
	);
	LUT3 #(
		.INIT('h04)
	) name4173 (
		_w6755_,
		_w8192_,
		_w8196_,
		_w8221_
	);
	LUT3 #(
		.INIT('h80)
	) name4174 (
		\bdma_BRdataBUF_reg[12]/P0001 ,
		_w5530_,
		_w5534_,
		_w8222_
	);
	LUT3 #(
		.INIT('h80)
	) name4175 (
		\idma_DTMP_H_reg[12]/P0001 ,
		_w5573_,
		_w8191_,
		_w8223_
	);
	LUT3 #(
		.INIT('h20)
	) name4176 (
		\sport0_rxctl_RX_reg[12]/P0001 ,
		_w4088_,
		_w4984_,
		_w8224_
	);
	LUT3 #(
		.INIT('h20)
	) name4177 (
		\sport1_rxctl_RX_reg[12]/P0001 ,
		_w4088_,
		_w4980_,
		_w8225_
	);
	LUT2 #(
		.INIT('h1)
	) name4178 (
		_w8224_,
		_w8225_,
		_w8226_
	);
	LUT3 #(
		.INIT('h10)
	) name4179 (
		_w8223_,
		_w8222_,
		_w8226_,
		_w8227_
	);
	LUT2 #(
		.INIT('hb)
	) name4180 (
		_w8221_,
		_w8227_,
		_w8228_
	);
	LUT3 #(
		.INIT('h04)
	) name4181 (
		_w5757_,
		_w8192_,
		_w8196_,
		_w8229_
	);
	LUT3 #(
		.INIT('h80)
	) name4182 (
		\bdma_BRdataBUF_reg[13]/P0001 ,
		_w5530_,
		_w5534_,
		_w8230_
	);
	LUT3 #(
		.INIT('h80)
	) name4183 (
		\idma_DTMP_H_reg[13]/P0001 ,
		_w5573_,
		_w8191_,
		_w8231_
	);
	LUT3 #(
		.INIT('h20)
	) name4184 (
		\sport0_rxctl_RX_reg[13]/P0001 ,
		_w4088_,
		_w4984_,
		_w8232_
	);
	LUT3 #(
		.INIT('h20)
	) name4185 (
		\sport1_rxctl_RX_reg[13]/P0001 ,
		_w4088_,
		_w4980_,
		_w8233_
	);
	LUT2 #(
		.INIT('h1)
	) name4186 (
		_w8232_,
		_w8233_,
		_w8234_
	);
	LUT3 #(
		.INIT('h10)
	) name4187 (
		_w8231_,
		_w8230_,
		_w8234_,
		_w8235_
	);
	LUT2 #(
		.INIT('hb)
	) name4188 (
		_w8229_,
		_w8235_,
		_w8236_
	);
	LUT4 #(
		.INIT('h4000)
	) name4189 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[14]/P0001 ,
		_w8237_
	);
	LUT3 #(
		.INIT('h80)
	) name4190 (
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w5634_,
		_w5637_,
		_w8238_
	);
	LUT3 #(
		.INIT('h80)
	) name4191 (
		PM_bdry_sel_pad,
		_w5671_,
		_w5794_,
		_w8239_
	);
	LUT3 #(
		.INIT('h80)
	) name4192 (
		\memc_usysr_DO_reg[14]/NET0131 ,
		_w5631_,
		_w5660_,
		_w8240_
	);
	LUT3 #(
		.INIT('h80)
	) name4193 (
		\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w5634_,
		_w5635_,
		_w8241_
	);
	LUT4 #(
		.INIT('h0001)
	) name4194 (
		_w8238_,
		_w8239_,
		_w8240_,
		_w8241_,
		_w8242_
	);
	LUT3 #(
		.INIT('h80)
	) name4195 (
		\tm_tpr_reg_DO_reg[14]/NET0131 ,
		_w5631_,
		_w5635_,
		_w8243_
	);
	LUT3 #(
		.INIT('h80)
	) name4196 (
		\pio_pmask_reg_DO_reg[10]/NET0131 ,
		_w5628_,
		_w5660_,
		_w8244_
	);
	LUT3 #(
		.INIT('h80)
	) name4197 (
		\sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w5648_,
		_w5634_,
		_w8245_
	);
	LUT3 #(
		.INIT('h80)
	) name4198 (
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w5634_,
		_w5639_,
		_w8246_
	);
	LUT4 #(
		.INIT('h0001)
	) name4199 (
		_w8243_,
		_w8244_,
		_w8245_,
		_w8246_,
		_w8247_
	);
	LUT3 #(
		.INIT('h80)
	) name4200 (
		\PIO_oe[10]_pad ,
		_w5628_,
		_w5632_,
		_w8248_
	);
	LUT3 #(
		.INIT('h80)
	) name4201 (
		\tm_TCR_TMP_reg[14]/NET0131 ,
		_w5631_,
		_w5637_,
		_w8249_
	);
	LUT3 #(
		.INIT('h80)
	) name4202 (
		\sport0_regs_AUTO_a_reg[14]/NET0131 ,
		_w5627_,
		_w5634_,
		_w8250_
	);
	LUT3 #(
		.INIT('h80)
	) name4203 (
		\ISCLK1_pad ,
		_w5644_,
		_w5634_,
		_w8251_
	);
	LUT4 #(
		.INIT('h0001)
	) name4204 (
		_w8248_,
		_w8249_,
		_w8250_,
		_w8251_,
		_w8252_
	);
	LUT3 #(
		.INIT('h80)
	) name4205 (
		_w8242_,
		_w8247_,
		_w8252_,
		_w8253_
	);
	LUT3 #(
		.INIT('h80)
	) name4206 (
		\bdma_BCTL_reg[14]/NET0131 ,
		_w5627_,
		_w5629_,
		_w8254_
	);
	LUT3 #(
		.INIT('h80)
	) name4207 (
		\ISCLK0_pad ,
		_w5632_,
		_w5634_,
		_w8255_
	);
	LUT3 #(
		.INIT('h80)
	) name4208 (
		\clkc_ckr_reg_DO_reg[14]/NET0131 ,
		_w5631_,
		_w5644_,
		_w8256_
	);
	LUT3 #(
		.INIT('h80)
	) name4209 (
		\idma_DCTL_reg[14]/NET0131 ,
		_w5628_,
		_w5639_,
		_w8257_
	);
	LUT3 #(
		.INIT('h80)
	) name4210 (
		\emc_WSCRreg_DO_reg[14]/NET0131 ,
		_w5631_,
		_w5632_,
		_w8258_
	);
	LUT4 #(
		.INIT('h0001)
	) name4211 (
		_w8255_,
		_w8256_,
		_w8257_,
		_w8258_,
		_w8259_
	);
	LUT3 #(
		.INIT('h80)
	) name4212 (
		\PIO_out[10]_pad ,
		_w5628_,
		_w5635_,
		_w8260_
	);
	LUT3 #(
		.INIT('h80)
	) name4213 (
		\pio_PINT_reg[10]/NET0131 ,
		_w5670_,
		_w5672_,
		_w8261_
	);
	LUT4 #(
		.INIT('h0001)
	) name4214 (
		_w5945_,
		_w5947_,
		_w8260_,
		_w8261_,
		_w8262_
	);
	LUT3 #(
		.INIT('h40)
	) name4215 (
		_w8254_,
		_w8259_,
		_w8262_,
		_w8263_
	);
	LUT4 #(
		.INIT('ha820)
	) name4216 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001 ,
		_w8264_
	);
	LUT4 #(
		.INIT('ha820)
	) name4217 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001 ,
		_w8265_
	);
	LUT2 #(
		.INIT('h1)
	) name4218 (
		_w8264_,
		_w8265_,
		_w8266_
	);
	LUT3 #(
		.INIT('h1b)
	) name4219 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001 ,
		_w8267_
	);
	LUT4 #(
		.INIT('ha820)
	) name4220 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001 ,
		_w8268_
	);
	LUT3 #(
		.INIT('h1b)
	) name4221 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001 ,
		_w8269_
	);
	LUT4 #(
		.INIT('ha820)
	) name4222 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001 ,
		_w8270_
	);
	LUT3 #(
		.INIT('h1b)
	) name4223 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001 ,
		_w8271_
	);
	LUT4 #(
		.INIT('ha820)
	) name4224 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001 ,
		_w8272_
	);
	LUT3 #(
		.INIT('h01)
	) name4225 (
		_w8270_,
		_w8272_,
		_w8268_,
		_w8273_
	);
	LUT3 #(
		.INIT('h2a)
	) name4226 (
		_w5730_,
		_w8266_,
		_w8273_,
		_w8274_
	);
	LUT3 #(
		.INIT('h2a)
	) name4227 (
		_w5697_,
		_w5698_,
		_w5699_,
		_w8275_
	);
	LUT3 #(
		.INIT('h2a)
	) name4228 (
		_w5687_,
		_w5688_,
		_w5689_,
		_w8276_
	);
	LUT4 #(
		.INIT('h135f)
	) name4229 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport0_txctl_TX_reg[14]/P0001 ,
		\sport1_txctl_TX_reg[14]/P0001 ,
		_w8277_
	);
	LUT4 #(
		.INIT('h135f)
	) name4230 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[14]/P0001 ,
		\sport1_rxctl_RX_reg[14]/P0001 ,
		_w8278_
	);
	LUT3 #(
		.INIT('h2a)
	) name4231 (
		_w5706_,
		_w8277_,
		_w8278_,
		_w8279_
	);
	LUT2 #(
		.INIT('h8)
	) name4232 (
		\core_c_dec_IRE_reg[18]/NET0131 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w8280_
	);
	LUT4 #(
		.INIT('h135f)
	) name4233 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w8281_
	);
	LUT3 #(
		.INIT('h8a)
	) name4234 (
		_w5681_,
		_w8280_,
		_w8281_,
		_w8282_
	);
	LUT4 #(
		.INIT('h0001)
	) name4235 (
		_w8279_,
		_w8282_,
		_w8275_,
		_w8276_,
		_w8283_
	);
	LUT3 #(
		.INIT('h1b)
	) name4236 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001 ,
		_w8284_
	);
	LUT4 #(
		.INIT('ha820)
	) name4237 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001 ,
		_w8285_
	);
	LUT3 #(
		.INIT('h1b)
	) name4238 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001 ,
		_w8286_
	);
	LUT4 #(
		.INIT('ha820)
	) name4239 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001 ,
		_w8287_
	);
	LUT3 #(
		.INIT('h1b)
	) name4240 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001 ,
		_w8288_
	);
	LUT4 #(
		.INIT('ha820)
	) name4241 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001 ,
		_w8289_
	);
	LUT3 #(
		.INIT('h01)
	) name4242 (
		_w8287_,
		_w8289_,
		_w8285_,
		_w8290_
	);
	LUT3 #(
		.INIT('h2a)
	) name4243 (
		_w5741_,
		_w5746_,
		_w8290_,
		_w8291_
	);
	LUT3 #(
		.INIT('h1b)
	) name4244 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 ,
		_w8292_
	);
	LUT4 #(
		.INIT('ha820)
	) name4245 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 ,
		_w8293_
	);
	LUT3 #(
		.INIT('h1b)
	) name4246 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001 ,
		_w8294_
	);
	LUT4 #(
		.INIT('ha820)
	) name4247 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001 ,
		_w8295_
	);
	LUT3 #(
		.INIT('h1b)
	) name4248 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001 ,
		_w8296_
	);
	LUT4 #(
		.INIT('ha820)
	) name4249 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001 ,
		_w8297_
	);
	LUT3 #(
		.INIT('h01)
	) name4250 (
		_w8295_,
		_w8297_,
		_w8293_,
		_w8298_
	);
	LUT3 #(
		.INIT('h1b)
	) name4251 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001 ,
		_w8299_
	);
	LUT4 #(
		.INIT('ha820)
	) name4252 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001 ,
		_w8300_
	);
	LUT3 #(
		.INIT('h1b)
	) name4253 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001 ,
		_w8301_
	);
	LUT4 #(
		.INIT('ha820)
	) name4254 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001 ,
		_w8302_
	);
	LUT3 #(
		.INIT('h1b)
	) name4255 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001 ,
		_w8303_
	);
	LUT4 #(
		.INIT('ha820)
	) name4256 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001 ,
		_w8304_
	);
	LUT4 #(
		.INIT('h0001)
	) name4257 (
		_w5714_,
		_w8300_,
		_w8302_,
		_w8304_,
		_w8305_
	);
	LUT3 #(
		.INIT('h2a)
	) name4258 (
		_w5712_,
		_w8298_,
		_w8305_,
		_w8306_
	);
	LUT4 #(
		.INIT('h0100)
	) name4259 (
		_w8274_,
		_w8291_,
		_w8306_,
		_w8283_,
		_w8307_
	);
	LUT4 #(
		.INIT('hd500)
	) name4260 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w8253_,
		_w8263_,
		_w8307_,
		_w8308_
	);
	LUT2 #(
		.INIT('h4)
	) name4261 (
		_w8237_,
		_w8308_,
		_w8309_
	);
	LUT3 #(
		.INIT('h02)
	) name4262 (
		_w8192_,
		_w8196_,
		_w8309_,
		_w8310_
	);
	LUT3 #(
		.INIT('h80)
	) name4263 (
		\bdma_BRdataBUF_reg[14]/P0001 ,
		_w5530_,
		_w5534_,
		_w8311_
	);
	LUT3 #(
		.INIT('h80)
	) name4264 (
		\idma_DTMP_H_reg[14]/P0001 ,
		_w5573_,
		_w8191_,
		_w8312_
	);
	LUT3 #(
		.INIT('h20)
	) name4265 (
		\sport0_rxctl_RX_reg[14]/P0001 ,
		_w4088_,
		_w4984_,
		_w8313_
	);
	LUT3 #(
		.INIT('h20)
	) name4266 (
		\sport1_rxctl_RX_reg[14]/P0001 ,
		_w4088_,
		_w4980_,
		_w8314_
	);
	LUT2 #(
		.INIT('h1)
	) name4267 (
		_w8313_,
		_w8314_,
		_w8315_
	);
	LUT3 #(
		.INIT('h10)
	) name4268 (
		_w8312_,
		_w8311_,
		_w8315_,
		_w8316_
	);
	LUT2 #(
		.INIT('hb)
	) name4269 (
		_w8310_,
		_w8316_,
		_w8317_
	);
	LUT4 #(
		.INIT('h4000)
	) name4270 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		\regout_STD_C_reg[15]/P0001 ,
		_w8318_
	);
	LUT3 #(
		.INIT('h80)
	) name4271 (
		\PIO_out[11]_pad ,
		_w5628_,
		_w5635_,
		_w8319_
	);
	LUT3 #(
		.INIT('h80)
	) name4272 (
		\tm_TCR_TMP_reg[15]/NET0131 ,
		_w5631_,
		_w5637_,
		_w8320_
	);
	LUT3 #(
		.INIT('h80)
	) name4273 (
		\clkc_ckr_reg_DO_reg[15]/NET0131 ,
		_w5631_,
		_w5644_,
		_w8321_
	);
	LUT3 #(
		.INIT('h01)
	) name4274 (
		_w8320_,
		_w8321_,
		_w8319_,
		_w8322_
	);
	LUT3 #(
		.INIT('h80)
	) name4275 (
		\pio_pmask_reg_DO_reg[11]/NET0131 ,
		_w5628_,
		_w5660_,
		_w8323_
	);
	LUT3 #(
		.INIT('h80)
	) name4276 (
		\sice_ICYC_en_reg/NET0131 ,
		_w5671_,
		_w5794_,
		_w8324_
	);
	LUT3 #(
		.INIT('h80)
	) name4277 (
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w5634_,
		_w5639_,
		_w8325_
	);
	LUT3 #(
		.INIT('h80)
	) name4278 (
		\memc_usysr_DO_reg[15]/NET0131 ,
		_w5631_,
		_w5660_,
		_w8326_
	);
	LUT4 #(
		.INIT('h0001)
	) name4279 (
		_w8323_,
		_w8324_,
		_w8325_,
		_w8326_,
		_w8327_
	);
	LUT3 #(
		.INIT('h80)
	) name4280 (
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w5632_,
		_w5634_,
		_w8328_
	);
	LUT3 #(
		.INIT('h80)
	) name4281 (
		\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w5648_,
		_w5634_,
		_w8329_
	);
	LUT3 #(
		.INIT('h80)
	) name4282 (
		\pio_PINT_reg[11]/NET0131 ,
		_w5670_,
		_w5672_,
		_w8330_
	);
	LUT3 #(
		.INIT('h80)
	) name4283 (
		\sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w5634_,
		_w5635_,
		_w8331_
	);
	LUT4 #(
		.INIT('h0001)
	) name4284 (
		_w8328_,
		_w8329_,
		_w8330_,
		_w8331_,
		_w8332_
	);
	LUT3 #(
		.INIT('h80)
	) name4285 (
		_w8322_,
		_w8327_,
		_w8332_,
		_w8333_
	);
	LUT3 #(
		.INIT('h80)
	) name4286 (
		\bdma_BCTL_reg[15]/NET0131 ,
		_w5627_,
		_w5629_,
		_w8334_
	);
	LUT3 #(
		.INIT('h80)
	) name4287 (
		\tm_tpr_reg_DO_reg[15]/NET0131 ,
		_w5631_,
		_w5635_,
		_w8335_
	);
	LUT3 #(
		.INIT('h80)
	) name4288 (
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w5627_,
		_w5634_,
		_w8336_
	);
	LUT3 #(
		.INIT('h80)
	) name4289 (
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w5634_,
		_w5637_,
		_w8337_
	);
	LUT3 #(
		.INIT('h80)
	) name4290 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w5634_,
		_w5660_,
		_w8338_
	);
	LUT4 #(
		.INIT('h0001)
	) name4291 (
		_w8335_,
		_w8336_,
		_w8337_,
		_w8338_,
		_w8339_
	);
	LUT3 #(
		.INIT('h80)
	) name4292 (
		\tm_tsr_reg_DO_reg[8]/NET0131 ,
		_w5627_,
		_w5631_,
		_w8340_
	);
	LUT3 #(
		.INIT('h80)
	) name4293 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w5631_,
		_w5639_,
		_w8341_
	);
	LUT3 #(
		.INIT('h80)
	) name4294 (
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w5644_,
		_w5634_,
		_w8342_
	);
	LUT3 #(
		.INIT('h80)
	) name4295 (
		\PIO_oe[11]_pad ,
		_w5628_,
		_w5632_,
		_w8343_
	);
	LUT4 #(
		.INIT('h0001)
	) name4296 (
		_w8340_,
		_w8341_,
		_w8342_,
		_w8343_,
		_w8344_
	);
	LUT3 #(
		.INIT('h40)
	) name4297 (
		_w8334_,
		_w8339_,
		_w8344_,
		_w8345_
	);
	LUT4 #(
		.INIT('ha820)
	) name4298 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001 ,
		_w8346_
	);
	LUT4 #(
		.INIT('ha820)
	) name4299 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001 ,
		_w8347_
	);
	LUT2 #(
		.INIT('h1)
	) name4300 (
		_w8346_,
		_w8347_,
		_w8348_
	);
	LUT3 #(
		.INIT('h1b)
	) name4301 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001 ,
		_w8349_
	);
	LUT4 #(
		.INIT('ha820)
	) name4302 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001 ,
		_w8350_
	);
	LUT3 #(
		.INIT('h1b)
	) name4303 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001 ,
		_w8351_
	);
	LUT4 #(
		.INIT('ha820)
	) name4304 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001 ,
		_w8352_
	);
	LUT4 #(
		.INIT('ha820)
	) name4305 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001 ,
		_w8353_
	);
	LUT3 #(
		.INIT('h01)
	) name4306 (
		_w8352_,
		_w8353_,
		_w8350_,
		_w8354_
	);
	LUT3 #(
		.INIT('h2a)
	) name4307 (
		_w5730_,
		_w8348_,
		_w8354_,
		_w8355_
	);
	LUT4 #(
		.INIT('h135f)
	) name4308 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[15]/P0001 ,
		\sport1_txctl_TX_reg[15]/P0001 ,
		_w8356_
	);
	LUT4 #(
		.INIT('h135f)
	) name4309 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w8357_
	);
	LUT3 #(
		.INIT('h2a)
	) name4310 (
		_w5706_,
		_w8356_,
		_w8357_,
		_w8358_
	);
	LUT2 #(
		.INIT('h8)
	) name4311 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w8359_
	);
	LUT4 #(
		.INIT('h135f)
	) name4312 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		\core_c_dec_IRE_reg[19]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w8360_
	);
	LUT3 #(
		.INIT('h8a)
	) name4313 (
		_w5681_,
		_w8359_,
		_w8360_,
		_w8361_
	);
	LUT4 #(
		.INIT('h0001)
	) name4314 (
		_w8275_,
		_w8276_,
		_w8358_,
		_w8361_,
		_w8362_
	);
	LUT3 #(
		.INIT('h1b)
	) name4315 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001 ,
		_w8363_
	);
	LUT4 #(
		.INIT('ha820)
	) name4316 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001 ,
		_w8364_
	);
	LUT3 #(
		.INIT('h1b)
	) name4317 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001 ,
		_w8365_
	);
	LUT4 #(
		.INIT('ha820)
	) name4318 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001 ,
		_w8366_
	);
	LUT3 #(
		.INIT('h1b)
	) name4319 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001 ,
		_w8367_
	);
	LUT4 #(
		.INIT('ha820)
	) name4320 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001 ,
		_w8368_
	);
	LUT3 #(
		.INIT('h01)
	) name4321 (
		_w8366_,
		_w8368_,
		_w8364_,
		_w8369_
	);
	LUT3 #(
		.INIT('h2a)
	) name4322 (
		_w5741_,
		_w5746_,
		_w8369_,
		_w8370_
	);
	LUT3 #(
		.INIT('h1b)
	) name4323 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 ,
		_w8371_
	);
	LUT4 #(
		.INIT('ha820)
	) name4324 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 ,
		_w8372_
	);
	LUT3 #(
		.INIT('h1b)
	) name4325 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001 ,
		_w8373_
	);
	LUT4 #(
		.INIT('ha820)
	) name4326 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001 ,
		_w8374_
	);
	LUT3 #(
		.INIT('h1b)
	) name4327 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001 ,
		_w8375_
	);
	LUT4 #(
		.INIT('ha820)
	) name4328 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001 ,
		_w8376_
	);
	LUT3 #(
		.INIT('h01)
	) name4329 (
		_w8374_,
		_w8376_,
		_w8372_,
		_w8377_
	);
	LUT3 #(
		.INIT('h1b)
	) name4330 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001 ,
		_w8378_
	);
	LUT4 #(
		.INIT('ha820)
	) name4331 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001 ,
		_w8379_
	);
	LUT3 #(
		.INIT('h1b)
	) name4332 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001 ,
		_w8380_
	);
	LUT4 #(
		.INIT('ha820)
	) name4333 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001 ,
		_w8381_
	);
	LUT3 #(
		.INIT('h1b)
	) name4334 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001 ,
		_w8382_
	);
	LUT4 #(
		.INIT('ha820)
	) name4335 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001 ,
		_w8383_
	);
	LUT4 #(
		.INIT('h0001)
	) name4336 (
		_w5714_,
		_w8379_,
		_w8381_,
		_w8383_,
		_w8384_
	);
	LUT3 #(
		.INIT('h2a)
	) name4337 (
		_w5712_,
		_w8377_,
		_w8384_,
		_w8385_
	);
	LUT4 #(
		.INIT('h0100)
	) name4338 (
		_w8355_,
		_w8370_,
		_w8385_,
		_w8362_,
		_w8386_
	);
	LUT4 #(
		.INIT('hd500)
	) name4339 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w8333_,
		_w8345_,
		_w8386_,
		_w8387_
	);
	LUT2 #(
		.INIT('h4)
	) name4340 (
		_w8318_,
		_w8387_,
		_w8388_
	);
	LUT3 #(
		.INIT('h02)
	) name4341 (
		_w8192_,
		_w8196_,
		_w8388_,
		_w8389_
	);
	LUT3 #(
		.INIT('h80)
	) name4342 (
		\bdma_BRdataBUF_reg[15]/P0001 ,
		_w5530_,
		_w5534_,
		_w8390_
	);
	LUT3 #(
		.INIT('h80)
	) name4343 (
		\idma_DTMP_H_reg[15]/P0001 ,
		_w5573_,
		_w8191_,
		_w8391_
	);
	LUT3 #(
		.INIT('h20)
	) name4344 (
		\sport0_rxctl_RX_reg[15]/P0001 ,
		_w4088_,
		_w4984_,
		_w8392_
	);
	LUT3 #(
		.INIT('h20)
	) name4345 (
		\sport1_rxctl_RX_reg[15]/P0001 ,
		_w4088_,
		_w4980_,
		_w8393_
	);
	LUT2 #(
		.INIT('h1)
	) name4346 (
		_w8392_,
		_w8393_,
		_w8394_
	);
	LUT3 #(
		.INIT('h10)
	) name4347 (
		_w8391_,
		_w8390_,
		_w8394_,
		_w8395_
	);
	LUT2 #(
		.INIT('hb)
	) name4348 (
		_w8389_,
		_w8395_,
		_w8396_
	);
	LUT3 #(
		.INIT('h80)
	) name4349 (
		\bdma_BRdataBUF_reg[1]/P0001 ,
		_w5530_,
		_w5534_,
		_w8397_
	);
	LUT3 #(
		.INIT('h80)
	) name4350 (
		\idma_DTMP_H_reg[1]/P0001 ,
		_w5573_,
		_w8191_,
		_w8398_
	);
	LUT3 #(
		.INIT('h20)
	) name4351 (
		\sport1_rxctl_RX_reg[1]/P0001 ,
		_w4088_,
		_w4980_,
		_w8399_
	);
	LUT3 #(
		.INIT('h20)
	) name4352 (
		\sport0_rxctl_RX_reg[1]/P0001 ,
		_w4088_,
		_w4984_,
		_w8400_
	);
	LUT2 #(
		.INIT('h1)
	) name4353 (
		_w8399_,
		_w8400_,
		_w8401_
	);
	LUT3 #(
		.INIT('h10)
	) name4354 (
		_w8398_,
		_w8397_,
		_w8401_,
		_w8402_
	);
	LUT3 #(
		.INIT('h4f)
	) name4355 (
		_w6893_,
		_w8197_,
		_w8402_,
		_w8403_
	);
	LUT3 #(
		.INIT('h80)
	) name4356 (
		\bdma_BRdataBUF_reg[2]/P0001 ,
		_w5530_,
		_w5534_,
		_w8404_
	);
	LUT3 #(
		.INIT('h80)
	) name4357 (
		\idma_DTMP_H_reg[2]/P0001 ,
		_w5573_,
		_w8191_,
		_w8405_
	);
	LUT3 #(
		.INIT('h20)
	) name4358 (
		\sport1_rxctl_RX_reg[2]/P0001 ,
		_w4088_,
		_w4980_,
		_w8406_
	);
	LUT3 #(
		.INIT('h20)
	) name4359 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		_w4088_,
		_w4984_,
		_w8407_
	);
	LUT2 #(
		.INIT('h1)
	) name4360 (
		_w8406_,
		_w8407_,
		_w8408_
	);
	LUT3 #(
		.INIT('h10)
	) name4361 (
		_w8405_,
		_w8404_,
		_w8408_,
		_w8409_
	);
	LUT3 #(
		.INIT('h4f)
	) name4362 (
		_w6497_,
		_w8197_,
		_w8409_,
		_w8410_
	);
	LUT3 #(
		.INIT('h80)
	) name4363 (
		\bdma_BRdataBUF_reg[3]/P0001 ,
		_w5530_,
		_w5534_,
		_w8411_
	);
	LUT3 #(
		.INIT('h80)
	) name4364 (
		\idma_DTMP_H_reg[3]/P0001 ,
		_w5573_,
		_w8191_,
		_w8412_
	);
	LUT3 #(
		.INIT('h20)
	) name4365 (
		\sport1_rxctl_RX_reg[3]/P0001 ,
		_w4088_,
		_w4980_,
		_w8413_
	);
	LUT3 #(
		.INIT('h20)
	) name4366 (
		\sport0_rxctl_RX_reg[3]/P0001 ,
		_w4088_,
		_w4984_,
		_w8414_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		_w8413_,
		_w8414_,
		_w8415_
	);
	LUT3 #(
		.INIT('h10)
	) name4368 (
		_w8412_,
		_w8411_,
		_w8415_,
		_w8416_
	);
	LUT3 #(
		.INIT('h4f)
	) name4369 (
		_w6172_,
		_w8197_,
		_w8416_,
		_w8417_
	);
	LUT3 #(
		.INIT('h80)
	) name4370 (
		\bdma_BRdataBUF_reg[4]/P0001 ,
		_w5530_,
		_w5534_,
		_w8418_
	);
	LUT3 #(
		.INIT('h80)
	) name4371 (
		\idma_DTMP_H_reg[4]/P0001 ,
		_w5573_,
		_w8191_,
		_w8419_
	);
	LUT3 #(
		.INIT('h20)
	) name4372 (
		\sport1_rxctl_RX_reg[4]/P0001 ,
		_w4088_,
		_w4980_,
		_w8420_
	);
	LUT3 #(
		.INIT('h20)
	) name4373 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w4088_,
		_w4984_,
		_w8421_
	);
	LUT2 #(
		.INIT('h1)
	) name4374 (
		_w8420_,
		_w8421_,
		_w8422_
	);
	LUT3 #(
		.INIT('h10)
	) name4375 (
		_w8419_,
		_w8418_,
		_w8422_,
		_w8423_
	);
	LUT3 #(
		.INIT('h4f)
	) name4376 (
		_w7374_,
		_w8197_,
		_w8423_,
		_w8424_
	);
	LUT3 #(
		.INIT('h80)
	) name4377 (
		\bdma_BRdataBUF_reg[5]/P0001 ,
		_w5530_,
		_w5534_,
		_w8425_
	);
	LUT3 #(
		.INIT('h80)
	) name4378 (
		\idma_DTMP_H_reg[5]/P0001 ,
		_w5573_,
		_w8191_,
		_w8426_
	);
	LUT3 #(
		.INIT('h20)
	) name4379 (
		\sport1_rxctl_RX_reg[5]/P0001 ,
		_w4088_,
		_w4980_,
		_w8427_
	);
	LUT3 #(
		.INIT('h20)
	) name4380 (
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w4088_,
		_w4984_,
		_w8428_
	);
	LUT2 #(
		.INIT('h1)
	) name4381 (
		_w8427_,
		_w8428_,
		_w8429_
	);
	LUT3 #(
		.INIT('h10)
	) name4382 (
		_w8426_,
		_w8425_,
		_w8429_,
		_w8430_
	);
	LUT3 #(
		.INIT('h4f)
	) name4383 (
		_w7706_,
		_w8197_,
		_w8430_,
		_w8431_
	);
	LUT3 #(
		.INIT('h80)
	) name4384 (
		\bdma_BRdataBUF_reg[6]/P0001 ,
		_w5530_,
		_w5534_,
		_w8432_
	);
	LUT3 #(
		.INIT('h80)
	) name4385 (
		\idma_DTMP_H_reg[6]/P0001 ,
		_w5573_,
		_w8191_,
		_w8433_
	);
	LUT3 #(
		.INIT('h20)
	) name4386 (
		\sport1_rxctl_RX_reg[6]/P0001 ,
		_w4088_,
		_w4980_,
		_w8434_
	);
	LUT3 #(
		.INIT('h20)
	) name4387 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w4088_,
		_w4984_,
		_w8435_
	);
	LUT2 #(
		.INIT('h1)
	) name4388 (
		_w8434_,
		_w8435_,
		_w8436_
	);
	LUT3 #(
		.INIT('h10)
	) name4389 (
		_w8433_,
		_w8432_,
		_w8436_,
		_w8437_
	);
	LUT3 #(
		.INIT('h4f)
	) name4390 (
		_w8039_,
		_w8197_,
		_w8437_,
		_w8438_
	);
	LUT3 #(
		.INIT('h80)
	) name4391 (
		\idma_DTMP_H_reg[7]/P0001 ,
		_w5573_,
		_w8191_,
		_w8439_
	);
	LUT3 #(
		.INIT('h80)
	) name4392 (
		\bdma_BRdataBUF_reg[7]/P0001 ,
		_w5530_,
		_w5534_,
		_w8440_
	);
	LUT3 #(
		.INIT('h20)
	) name4393 (
		\sport1_rxctl_RX_reg[7]/P0001 ,
		_w4088_,
		_w4980_,
		_w8441_
	);
	LUT3 #(
		.INIT('h20)
	) name4394 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w4088_,
		_w4984_,
		_w8442_
	);
	LUT2 #(
		.INIT('h1)
	) name4395 (
		_w8441_,
		_w8442_,
		_w8443_
	);
	LUT3 #(
		.INIT('h10)
	) name4396 (
		_w8440_,
		_w8439_,
		_w8443_,
		_w8444_
	);
	LUT3 #(
		.INIT('h4f)
	) name4397 (
		_w7902_,
		_w8197_,
		_w8444_,
		_w8445_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4398 (
		_w7466_,
		_w7562_,
		_w8192_,
		_w8196_,
		_w8446_
	);
	LUT3 #(
		.INIT('h80)
	) name4399 (
		\bdma_BRdataBUF_reg[8]/P0001 ,
		_w5530_,
		_w5534_,
		_w8447_
	);
	LUT3 #(
		.INIT('h80)
	) name4400 (
		\idma_DTMP_H_reg[8]/P0001 ,
		_w5573_,
		_w8191_,
		_w8448_
	);
	LUT3 #(
		.INIT('h20)
	) name4401 (
		\sport1_rxctl_RX_reg[8]/P0001 ,
		_w4088_,
		_w4980_,
		_w8449_
	);
	LUT3 #(
		.INIT('h20)
	) name4402 (
		\sport0_rxctl_RX_reg[8]/P0001 ,
		_w4088_,
		_w4984_,
		_w8450_
	);
	LUT2 #(
		.INIT('h1)
	) name4403 (
		_w8449_,
		_w8450_,
		_w8451_
	);
	LUT3 #(
		.INIT('h10)
	) name4404 (
		_w8448_,
		_w8447_,
		_w8451_,
		_w8452_
	);
	LUT2 #(
		.INIT('hb)
	) name4405 (
		_w8446_,
		_w8452_,
		_w8453_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4406 (
		_w7141_,
		_w7237_,
		_w8192_,
		_w8196_,
		_w8454_
	);
	LUT3 #(
		.INIT('h80)
	) name4407 (
		\bdma_BRdataBUF_reg[9]/P0001 ,
		_w5530_,
		_w5534_,
		_w8455_
	);
	LUT3 #(
		.INIT('h80)
	) name4408 (
		\idma_DTMP_H_reg[9]/P0001 ,
		_w5573_,
		_w8191_,
		_w8456_
	);
	LUT3 #(
		.INIT('h20)
	) name4409 (
		\sport0_rxctl_RX_reg[9]/P0001 ,
		_w4088_,
		_w4984_,
		_w8457_
	);
	LUT3 #(
		.INIT('h20)
	) name4410 (
		\sport1_rxctl_RX_reg[9]/P0001 ,
		_w4088_,
		_w4980_,
		_w8458_
	);
	LUT2 #(
		.INIT('h1)
	) name4411 (
		_w8457_,
		_w8458_,
		_w8459_
	);
	LUT3 #(
		.INIT('h10)
	) name4412 (
		_w8456_,
		_w8455_,
		_w8459_,
		_w8460_
	);
	LUT2 #(
		.INIT('hb)
	) name4413 (
		_w8454_,
		_w8460_,
		_w8461_
	);
	LUT3 #(
		.INIT('h53)
	) name4414 (
		\bdma_BOVL_reg[6]/NET0131 ,
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		_w4519_,
		_w8462_
	);
	LUT3 #(
		.INIT('h74)
	) name4415 (
		\idma_DOVL_reg[6]/NET0131 ,
		_w4946_,
		_w8462_,
		_w8463_
	);
	LUT3 #(
		.INIT('h53)
	) name4416 (
		\bdma_BOVL_reg[7]/NET0131 ,
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		_w4519_,
		_w8464_
	);
	LUT3 #(
		.INIT('h74)
	) name4417 (
		\idma_DOVL_reg[7]/NET0131 ,
		_w4946_,
		_w8464_,
		_w8465_
	);
	LUT3 #(
		.INIT('h53)
	) name4418 (
		\bdma_BOVL_reg[4]/NET0131 ,
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		_w4519_,
		_w8466_
	);
	LUT3 #(
		.INIT('h74)
	) name4419 (
		\idma_DOVL_reg[4]/NET0131 ,
		_w4946_,
		_w8466_,
		_w8467_
	);
	LUT3 #(
		.INIT('h80)
	) name4420 (
		_w8463_,
		_w8465_,
		_w8467_,
		_w8468_
	);
	LUT3 #(
		.INIT('h53)
	) name4421 (
		\bdma_BOVL_reg[5]/NET0131 ,
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		_w4519_,
		_w8469_
	);
	LUT3 #(
		.INIT('h74)
	) name4422 (
		\idma_DOVL_reg[5]/NET0131 ,
		_w4946_,
		_w8469_,
		_w8470_
	);
	LUT4 #(
		.INIT('h2000)
	) name4423 (
		_w6944_,
		_w8194_,
		_w8468_,
		_w8470_,
		_w8471_
	);
	LUT3 #(
		.INIT('h08)
	) name4424 (
		_w8463_,
		_w8465_,
		_w8467_,
		_w8472_
	);
	LUT4 #(
		.INIT('h2000)
	) name4425 (
		_w6944_,
		_w8194_,
		_w8470_,
		_w8472_,
		_w8473_
	);
	LUT4 #(
		.INIT('h0020)
	) name4426 (
		_w6944_,
		_w8194_,
		_w8468_,
		_w8470_,
		_w8474_
	);
	LUT4 #(
		.INIT('h0200)
	) name4427 (
		_w6944_,
		_w8194_,
		_w8470_,
		_w8472_,
		_w8475_
	);
	LUT3 #(
		.INIT('h40)
	) name4428 (
		_w8463_,
		_w8465_,
		_w8467_,
		_w8476_
	);
	LUT4 #(
		.INIT('h2000)
	) name4429 (
		_w6944_,
		_w8194_,
		_w8470_,
		_w8476_,
		_w8477_
	);
	LUT3 #(
		.INIT('h04)
	) name4430 (
		_w8463_,
		_w8465_,
		_w8467_,
		_w8478_
	);
	LUT4 #(
		.INIT('h2000)
	) name4431 (
		_w6944_,
		_w8194_,
		_w8470_,
		_w8478_,
		_w8479_
	);
	LUT4 #(
		.INIT('h0200)
	) name4432 (
		_w6944_,
		_w8194_,
		_w8470_,
		_w8476_,
		_w8480_
	);
	LUT4 #(
		.INIT('h0200)
	) name4433 (
		_w6944_,
		_w8194_,
		_w8470_,
		_w8478_,
		_w8481_
	);
	LUT2 #(
		.INIT('h8)
	) name4434 (
		T_ICE_RSTn_pad,
		T_RSTn_pad,
		_w8482_
	);
	LUT2 #(
		.INIT('h7)
	) name4435 (
		T_ICE_RSTn_pad,
		T_RSTn_pad,
		_w8483_
	);
	LUT3 #(
		.INIT('h80)
	) name4436 (
		T_ICE_RSTn_pad,
		T_RSTn_pad,
		\clkc_DSPoff_reg/NET0131 ,
		_w8484_
	);
	LUT3 #(
		.INIT('h80)
	) name4437 (
		T_ICE_RSTn_pad,
		T_RSTn_pad,
		\clkc_SlowDn_reg/NET0131 ,
		_w8485_
	);
	LUT3 #(
		.INIT('h80)
	) name4438 (
		T_ICE_RSTn_pad,
		T_RSTn_pad,
		\clkc_OSCoff_reg/NET0131 ,
		_w8486_
	);
	LUT3 #(
		.INIT('h7f)
	) name4439 (
		T_ICE_RSTn_pad,
		T_RSTn_pad,
		\clkc_OSCoff_reg/NET0131 ,
		_w8487_
	);
	LUT3 #(
		.INIT('hca)
	) name4440 (
		T_CLKI_OSC_pad,
		T_CLKI_PLL_pad,
		T_Sel_PLL_pad,
		_w8488_
	);
	LUT2 #(
		.INIT('h4)
	) name4441 (
		_w8486_,
		_w8488_,
		_w8489_
	);
	LUT4 #(
		.INIT('h7477)
	) name4442 (
		\clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131 ,
		_w8485_,
		_w8486_,
		_w8488_,
		_w8490_
	);
	LUT2 #(
		.INIT('h4)
	) name4443 (
		_w8484_,
		_w8490_,
		_w8491_
	);
	LUT2 #(
		.INIT('hb)
	) name4444 (
		_w8484_,
		_w8490_,
		_w8492_
	);
	LUT4 #(
		.INIT('h8088)
	) name4445 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8493_
	);
	LUT3 #(
		.INIT('h20)
	) name4446 (
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w8494_
	);
	LUT4 #(
		.INIT('h3f77)
	) name4447 (
		\emc_ECMA_reg[0]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[4]/P0001 ,
		_w8494_,
		_w8495_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4448 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8496_
	);
	LUT4 #(
		.INIT('h8088)
	) name4449 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8497_
	);
	LUT4 #(
		.INIT('h0100)
	) name4450 (
		_w8493_,
		_w8496_,
		_w8497_,
		_w8495_,
		_w8498_
	);
	LUT3 #(
		.INIT('h8b)
	) name4451 (
		\bdma_BEAD_reg[0]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8498_,
		_w8499_
	);
	LUT4 #(
		.INIT('h8088)
	) name4452 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8500_
	);
	LUT2 #(
		.INIT('h8)
	) name4453 (
		\emc_ECMA_reg[10]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w8501_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4454 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8502_
	);
	LUT4 #(
		.INIT('h8088)
	) name4455 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8503_
	);
	LUT4 #(
		.INIT('h0001)
	) name4456 (
		_w8500_,
		_w8502_,
		_w8501_,
		_w8503_,
		_w8504_
	);
	LUT3 #(
		.INIT('h8b)
	) name4457 (
		\bdma_BEAD_reg[10]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8504_,
		_w8505_
	);
	LUT2 #(
		.INIT('h8)
	) name4458 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w8506_
	);
	LUT4 #(
		.INIT('h0004)
	) name4459 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4825_,
		_w4843_,
		_w8506_,
		_w8507_
	);
	LUT4 #(
		.INIT('h4450)
	) name4460 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\emc_ECMA_reg[12]/P0001 ,
		_w8507_,
		_w8508_
	);
	LUT3 #(
		.INIT('h02)
	) name4461 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4825_,
		_w8509_
	);
	LUT3 #(
		.INIT('h01)
	) name4462 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\emc_ECMA_reg[12]/P0001 ,
		_w8510_
	);
	LUT3 #(
		.INIT('h04)
	) name4463 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w4843_,
		_w8510_,
		_w8511_
	);
	LUT2 #(
		.INIT('h8)
	) name4464 (
		_w8509_,
		_w8511_,
		_w8512_
	);
	LUT4 #(
		.INIT('h8088)
	) name4465 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8513_
	);
	LUT3 #(
		.INIT('he4)
	) name4466 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		_w8514_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4467 (
		_w4721_,
		_w4804_,
		_w4805_,
		_w8514_,
		_w8515_
	);
	LUT2 #(
		.INIT('h1)
	) name4468 (
		_w8513_,
		_w8515_,
		_w8516_
	);
	LUT4 #(
		.INIT('h5700)
	) name4469 (
		\emc_ECMcs_reg/NET0131 ,
		_w8508_,
		_w8512_,
		_w8516_,
		_w8517_
	);
	LUT3 #(
		.INIT('h8b)
	) name4470 (
		\bdma_BEAD_reg[12]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8517_,
		_w8518_
	);
	LUT3 #(
		.INIT('h9f)
	) name4471 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w4843_,
		_w8519_
	);
	LUT3 #(
		.INIT('h01)
	) name4472 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4843_,
		_w8520_
	);
	LUT2 #(
		.INIT('h4)
	) name4473 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w4825_,
		_w8521_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name4474 (
		_w8509_,
		_w8519_,
		_w8520_,
		_w8521_,
		_w8522_
	);
	LUT4 #(
		.INIT('h8088)
	) name4475 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8523_
	);
	LUT3 #(
		.INIT('hd8)
	) name4476 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		_w8524_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4477 (
		_w4721_,
		_w4804_,
		_w4805_,
		_w8524_,
		_w8525_
	);
	LUT2 #(
		.INIT('h1)
	) name4478 (
		_w8523_,
		_w8525_,
		_w8526_
	);
	LUT4 #(
		.INIT('h0455)
	) name4479 (
		\bdma_BM_cyc_reg/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w8522_,
		_w8526_,
		_w8527_
	);
	LUT2 #(
		.INIT('h8)
	) name4480 (
		\bdma_BEAD_reg[13]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8528_
	);
	LUT2 #(
		.INIT('he)
	) name4481 (
		_w8527_,
		_w8528_,
		_w8529_
	);
	LUT4 #(
		.INIT('h87ff)
	) name4482 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4843_,
		_w8530_
	);
	LUT3 #(
		.INIT('h60)
	) name4483 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4825_,
		_w8531_
	);
	LUT4 #(
		.INIT('h31f5)
	) name4484 (
		_w8509_,
		_w8520_,
		_w8530_,
		_w8531_,
		_w8532_
	);
	LUT4 #(
		.INIT('h8088)
	) name4485 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8533_
	);
	LUT3 #(
		.INIT('hd8)
	) name4486 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		_w8534_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4487 (
		_w4721_,
		_w4804_,
		_w4805_,
		_w8534_,
		_w8535_
	);
	LUT2 #(
		.INIT('h1)
	) name4488 (
		_w8533_,
		_w8535_,
		_w8536_
	);
	LUT4 #(
		.INIT('h0455)
	) name4489 (
		\bdma_BM_cyc_reg/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w8532_,
		_w8536_,
		_w8537_
	);
	LUT2 #(
		.INIT('h8)
	) name4490 (
		\bdma_BCTL_reg[8]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8538_
	);
	LUT2 #(
		.INIT('he)
	) name4491 (
		_w8537_,
		_w8538_,
		_w8539_
	);
	LUT4 #(
		.INIT('h8088)
	) name4492 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8540_
	);
	LUT4 #(
		.INIT('h3f77)
	) name4493 (
		\emc_ECMA_reg[1]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[5]/P0001 ,
		_w8494_,
		_w8541_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4494 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8542_
	);
	LUT4 #(
		.INIT('h8088)
	) name4495 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8543_
	);
	LUT4 #(
		.INIT('h0100)
	) name4496 (
		_w8540_,
		_w8542_,
		_w8543_,
		_w8541_,
		_w8544_
	);
	LUT3 #(
		.INIT('h8b)
	) name4497 (
		\bdma_BEAD_reg[1]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8544_,
		_w8545_
	);
	LUT4 #(
		.INIT('h8088)
	) name4498 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8546_
	);
	LUT4 #(
		.INIT('h3f77)
	) name4499 (
		\emc_ECMA_reg[2]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[6]/P0001 ,
		_w8494_,
		_w8547_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4500 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8548_
	);
	LUT4 #(
		.INIT('h8088)
	) name4501 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8549_
	);
	LUT4 #(
		.INIT('h0100)
	) name4502 (
		_w8546_,
		_w8548_,
		_w8549_,
		_w8547_,
		_w8550_
	);
	LUT3 #(
		.INIT('h8b)
	) name4503 (
		\bdma_BEAD_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8550_,
		_w8551_
	);
	LUT4 #(
		.INIT('h8088)
	) name4504 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8552_
	);
	LUT4 #(
		.INIT('h3f77)
	) name4505 (
		\emc_ECMA_reg[3]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[7]/P0001 ,
		_w8494_,
		_w8553_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4506 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8554_
	);
	LUT4 #(
		.INIT('h8088)
	) name4507 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8555_
	);
	LUT4 #(
		.INIT('h0100)
	) name4508 (
		_w8552_,
		_w8554_,
		_w8555_,
		_w8553_,
		_w8556_
	);
	LUT3 #(
		.INIT('h8b)
	) name4509 (
		\bdma_BEAD_reg[3]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8556_,
		_w8557_
	);
	LUT4 #(
		.INIT('h8088)
	) name4510 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8558_
	);
	LUT4 #(
		.INIT('h3f77)
	) name4511 (
		\emc_ECMA_reg[4]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[8]/P0001 ,
		_w8494_,
		_w8559_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4512 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8560_
	);
	LUT4 #(
		.INIT('h8088)
	) name4513 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8561_
	);
	LUT4 #(
		.INIT('h0100)
	) name4514 (
		_w8558_,
		_w8560_,
		_w8561_,
		_w8559_,
		_w8562_
	);
	LUT3 #(
		.INIT('h8b)
	) name4515 (
		\bdma_BEAD_reg[4]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8562_,
		_w8563_
	);
	LUT4 #(
		.INIT('h8088)
	) name4516 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8564_
	);
	LUT4 #(
		.INIT('h3f77)
	) name4517 (
		\emc_ECMA_reg[5]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[9]/P0001 ,
		_w8494_,
		_w8565_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4518 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8566_
	);
	LUT4 #(
		.INIT('h8088)
	) name4519 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8567_
	);
	LUT4 #(
		.INIT('h0100)
	) name4520 (
		_w8564_,
		_w8566_,
		_w8567_,
		_w8565_,
		_w8568_
	);
	LUT3 #(
		.INIT('h8b)
	) name4521 (
		\bdma_BEAD_reg[5]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8568_,
		_w8569_
	);
	LUT4 #(
		.INIT('h8088)
	) name4522 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8570_
	);
	LUT4 #(
		.INIT('h3f77)
	) name4523 (
		\emc_ECMA_reg[6]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[10]/P0001 ,
		_w8494_,
		_w8571_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4524 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8572_
	);
	LUT4 #(
		.INIT('h8088)
	) name4525 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8573_
	);
	LUT4 #(
		.INIT('h0100)
	) name4526 (
		_w8570_,
		_w8572_,
		_w8573_,
		_w8571_,
		_w8574_
	);
	LUT3 #(
		.INIT('h8b)
	) name4527 (
		\bdma_BEAD_reg[6]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8574_,
		_w8575_
	);
	LUT4 #(
		.INIT('h8088)
	) name4528 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8576_
	);
	LUT4 #(
		.INIT('h3f77)
	) name4529 (
		\emc_ECMA_reg[7]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[11]/P0001 ,
		_w8494_,
		_w8577_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4530 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8578_
	);
	LUT4 #(
		.INIT('h8088)
	) name4531 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8579_
	);
	LUT4 #(
		.INIT('h0100)
	) name4532 (
		_w8576_,
		_w8578_,
		_w8579_,
		_w8577_,
		_w8580_
	);
	LUT3 #(
		.INIT('h8b)
	) name4533 (
		\bdma_BEAD_reg[7]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8580_,
		_w8581_
	);
	LUT4 #(
		.INIT('h8088)
	) name4534 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8582_
	);
	LUT2 #(
		.INIT('h8)
	) name4535 (
		\emc_ECMA_reg[8]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w8583_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4536 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8584_
	);
	LUT4 #(
		.INIT('h8088)
	) name4537 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8585_
	);
	LUT4 #(
		.INIT('h0001)
	) name4538 (
		_w8582_,
		_w8584_,
		_w8583_,
		_w8585_,
		_w8586_
	);
	LUT3 #(
		.INIT('h8b)
	) name4539 (
		\bdma_BEAD_reg[8]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8586_,
		_w8587_
	);
	LUT4 #(
		.INIT('h8088)
	) name4540 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8588_
	);
	LUT2 #(
		.INIT('h8)
	) name4541 (
		\emc_ECMA_reg[9]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w8589_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4542 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8590_
	);
	LUT4 #(
		.INIT('h8088)
	) name4543 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8591_
	);
	LUT4 #(
		.INIT('h0001)
	) name4544 (
		_w8588_,
		_w8590_,
		_w8589_,
		_w8591_,
		_w8592_
	);
	LUT3 #(
		.INIT('h8b)
	) name4545 (
		\bdma_BEAD_reg[9]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8592_,
		_w8593_
	);
	LUT4 #(
		.INIT('h1f11)
	) name4546 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w8594_
	);
	LUT4 #(
		.INIT('h0100)
	) name4547 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w8595_
	);
	LUT2 #(
		.INIT('h2)
	) name4548 (
		\core_c_dec_accCM_E_reg/NET0131 ,
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w8596_
	);
	LUT4 #(
		.INIT('h0111)
	) name4549 (
		\bdma_BM_cyc_reg/P0001 ,
		_w4750_,
		_w8494_,
		_w8596_,
		_w8597_
	);
	LUT2 #(
		.INIT('h4)
	) name4550 (
		_w8595_,
		_w8597_,
		_w8598_
	);
	LUT4 #(
		.INIT('h0100)
	) name4551 (
		_w4721_,
		_w4804_,
		_w4805_,
		_w8598_,
		_w8599_
	);
	LUT3 #(
		.INIT('h15)
	) name4552 (
		\core_c_psq_MGNT_reg/NET0131 ,
		_w8594_,
		_w8599_,
		_w8600_
	);
	LUT2 #(
		.INIT('h4)
	) name4553 (
		\core_c_psq_MGNT_reg/NET0131 ,
		\emc_ED_oei_reg/P0001 ,
		_w8601_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4554 (
		\emc_selPMDi_reg/P0001 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w8602_
	);
	LUT3 #(
		.INIT('h02)
	) name4555 (
		\emc_selDMDi_reg/P0001 ,
		_w8594_,
		_w8602_,
		_w8603_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4556 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w8594_,
		_w8602_,
		_w8604_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name4557 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_pMFMAC_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w8605_
	);
	LUT3 #(
		.INIT('h70)
	) name4558 (
		_w5871_,
		_w5880_,
		_w8605_,
		_w8606_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name4559 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_pMFSHT_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w8607_
	);
	LUT3 #(
		.INIT('h70)
	) name4560 (
		_w5886_,
		_w5893_,
		_w8607_,
		_w8608_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name4561 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_pMFALU_Ei_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_STI_Cg_reg/NET0131 ,
		_w8609_
	);
	LUT3 #(
		.INIT('h70)
	) name4562 (
		_w5898_,
		_w5905_,
		_w8609_,
		_w8610_
	);
	LUT4 #(
		.INIT('h5554)
	) name4563 (
		\emc_PMDoe_reg/NET0131 ,
		_w8608_,
		_w8610_,
		_w8606_,
		_w8611_
	);
	LUT2 #(
		.INIT('h8)
	) name4564 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[0]/P0001 ,
		_w8612_
	);
	LUT2 #(
		.INIT('h1)
	) name4565 (
		\memc_PMo_oe2_reg/P0001 ,
		\memc_PMo_oe3_reg/P0001 ,
		_w8613_
	);
	LUT2 #(
		.INIT('h1)
	) name4566 (
		\memc_PMo_oe4_reg/P0001 ,
		\memc_PMo_oe5_reg/P0001 ,
		_w8614_
	);
	LUT4 #(
		.INIT('h0001)
	) name4567 (
		\memc_PMo_oe4_reg/P0001 ,
		\memc_PMo_oe5_reg/P0001 ,
		\memc_PMo_oe6_reg/P0001 ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8615_
	);
	LUT2 #(
		.INIT('h1)
	) name4568 (
		\memc_PMo_oe0_reg/P0001 ,
		\memc_PMo_oe1_reg/P0001 ,
		_w8616_
	);
	LUT3 #(
		.INIT('h80)
	) name4569 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8617_
	);
	LUT4 #(
		.INIT('h4000)
	) name4570 (
		_w8612_,
		_w8613_,
		_w8615_,
		_w8616_,
		_w8618_
	);
	LUT2 #(
		.INIT('h2)
	) name4571 (
		\memc_PMo_oe2_reg/P0001 ,
		\memc_PMo_oe3_reg/P0001 ,
		_w8619_
	);
	LUT3 #(
		.INIT('h80)
	) name4572 (
		_w8615_,
		_w8616_,
		_w8619_,
		_w8620_
	);
	LUT4 #(
		.INIT('h0001)
	) name4573 (
		\memc_PMo_oe0_reg/P0001 ,
		\memc_PMo_oe1_reg/P0001 ,
		\memc_PMo_oe2_reg/P0001 ,
		\memc_PMo_oe3_reg/P0001 ,
		_w8621_
	);
	LUT3 #(
		.INIT('h10)
	) name4574 (
		\memc_PMo_oe4_reg/P0001 ,
		\memc_PMo_oe5_reg/P0001 ,
		\memc_PMo_oe6_reg/P0001 ,
		_w8622_
	);
	LUT4 #(
		.INIT('h0100)
	) name4575 (
		\memc_PMo_oe4_reg/P0001 ,
		\memc_PMo_oe5_reg/P0001 ,
		\memc_PMo_oe6_reg/P0001 ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8623_
	);
	LUT4 #(
		.INIT('h9fff)
	) name4576 (
		\memc_PMo_oe6_reg/P0001 ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8614_,
		_w8621_,
		_w8624_
	);
	LUT2 #(
		.INIT('h4)
	) name4577 (
		_w8620_,
		_w8624_,
		_w8625_
	);
	LUT2 #(
		.INIT('h2)
	) name4578 (
		\memc_PMo_oe4_reg/P0001 ,
		\memc_PMo_oe5_reg/P0001 ,
		_w8626_
	);
	LUT4 #(
		.INIT('h1000)
	) name4579 (
		\memc_PMo_oe6_reg/P0001 ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8626_,
		_w8627_
	);
	LUT2 #(
		.INIT('h4)
	) name4580 (
		\memc_PMo_oe0_reg/P0001 ,
		\memc_PMo_oe1_reg/P0001 ,
		_w8628_
	);
	LUT3 #(
		.INIT('h80)
	) name4581 (
		_w8613_,
		_w8615_,
		_w8628_,
		_w8629_
	);
	LUT2 #(
		.INIT('h4)
	) name4582 (
		\memc_PMo_oe2_reg/P0001 ,
		\memc_PMo_oe3_reg/P0001 ,
		_w8630_
	);
	LUT3 #(
		.INIT('h80)
	) name4583 (
		_w8615_,
		_w8616_,
		_w8630_,
		_w8631_
	);
	LUT2 #(
		.INIT('h4)
	) name4584 (
		\memc_PMo_oe4_reg/P0001 ,
		\memc_PMo_oe5_reg/P0001 ,
		_w8632_
	);
	LUT4 #(
		.INIT('h1000)
	) name4585 (
		\memc_PMo_oe6_reg/P0001 ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8632_,
		_w8633_
	);
	LUT4 #(
		.INIT('h0001)
	) name4586 (
		_w8627_,
		_w8629_,
		_w8631_,
		_w8633_,
		_w8634_
	);
	LUT2 #(
		.INIT('h2)
	) name4587 (
		\memc_PMo_oe0_reg/P0001 ,
		\memc_PMo_oe1_reg/P0001 ,
		_w8635_
	);
	LUT3 #(
		.INIT('h80)
	) name4588 (
		_w8613_,
		_w8615_,
		_w8635_,
		_w8636_
	);
	LUT4 #(
		.INIT('haa80)
	) name4589 (
		\PM_rd0[0]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8637_
	);
	LUT4 #(
		.INIT('h8000)
	) name4590 (
		\PM_rd3[0]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8638_
	);
	LUT4 #(
		.INIT('h8000)
	) name4591 (
		\PM_rd1[0]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8639_
	);
	LUT4 #(
		.INIT('h0007)
	) name4592 (
		\PM_rd5[0]_pad ,
		_w8633_,
		_w8638_,
		_w8639_,
		_w8640_
	);
	LUT3 #(
		.INIT('h80)
	) name4593 (
		\PM_rd7[0]_pad ,
		_w8621_,
		_w8623_,
		_w8641_
	);
	LUT4 #(
		.INIT('h2000)
	) name4594 (
		\PM_rd6[0]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8642_
	);
	LUT3 #(
		.INIT('h01)
	) name4595 (
		_w8617_,
		_w8642_,
		_w8641_,
		_w8643_
	);
	LUT4 #(
		.INIT('h8000)
	) name4596 (
		\PM_rd2[0]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8644_
	);
	LUT3 #(
		.INIT('h13)
	) name4597 (
		\PM_rd4[0]_pad ,
		_w8644_,
		_w8627_,
		_w8645_
	);
	LUT3 #(
		.INIT('h80)
	) name4598 (
		_w8643_,
		_w8645_,
		_w8640_,
		_w8646_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4599 (
		_w8611_,
		_w8618_,
		_w8637_,
		_w8646_,
		_w8647_
	);
	LUT2 #(
		.INIT('h8)
	) name4600 (
		_w8602_,
		_w8647_,
		_w8648_
	);
	LUT4 #(
		.INIT('h0013)
	) name4601 (
		_w5914_,
		_w8604_,
		_w8603_,
		_w8648_,
		_w8649_
	);
	LUT3 #(
		.INIT('h80)
	) name4602 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWdataBUF_reg[0]/P0001 ,
		_w8650_
	);
	LUT3 #(
		.INIT('hf2)
	) name4603 (
		_w8601_,
		_w8649_,
		_w8650_,
		_w8651_
	);
	LUT2 #(
		.INIT('h8)
	) name4604 (
		\bdma_BCTL_reg[11]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8652_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4605 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w8594_,
		_w8602_,
		_w8653_
	);
	LUT3 #(
		.INIT('h70)
	) name4606 (
		_w6025_,
		_w6031_,
		_w8609_,
		_w8654_
	);
	LUT3 #(
		.INIT('h70)
	) name4607 (
		_w6013_,
		_w6020_,
		_w8605_,
		_w8655_
	);
	LUT3 #(
		.INIT('h70)
	) name4608 (
		_w5746_,
		_w6005_,
		_w8607_,
		_w8656_
	);
	LUT3 #(
		.INIT('h01)
	) name4609 (
		_w8655_,
		_w8656_,
		_w8654_,
		_w8657_
	);
	LUT4 #(
		.INIT('h5554)
	) name4610 (
		\emc_PMDoe_reg/NET0131 ,
		_w8655_,
		_w8656_,
		_w8654_,
		_w8658_
	);
	LUT2 #(
		.INIT('h8)
	) name4611 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[10]/P0001 ,
		_w8659_
	);
	LUT4 #(
		.INIT('h0080)
	) name4612 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8659_,
		_w8660_
	);
	LUT4 #(
		.INIT('haa80)
	) name4613 (
		\PM_rd0[10]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8661_
	);
	LUT4 #(
		.INIT('h8000)
	) name4614 (
		\PM_rd3[10]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8662_
	);
	LUT4 #(
		.INIT('h8000)
	) name4615 (
		\PM_rd1[10]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8663_
	);
	LUT4 #(
		.INIT('h0007)
	) name4616 (
		\PM_rd5[10]_pad ,
		_w8633_,
		_w8662_,
		_w8663_,
		_w8664_
	);
	LUT3 #(
		.INIT('h80)
	) name4617 (
		\PM_rd7[10]_pad ,
		_w8621_,
		_w8623_,
		_w8665_
	);
	LUT4 #(
		.INIT('h2000)
	) name4618 (
		\PM_rd6[10]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8666_
	);
	LUT3 #(
		.INIT('h01)
	) name4619 (
		_w8617_,
		_w8666_,
		_w8665_,
		_w8667_
	);
	LUT4 #(
		.INIT('h8000)
	) name4620 (
		\PM_rd2[10]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8668_
	);
	LUT3 #(
		.INIT('h07)
	) name4621 (
		\PM_rd4[10]_pad ,
		_w8627_,
		_w8668_,
		_w8669_
	);
	LUT3 #(
		.INIT('h80)
	) name4622 (
		_w8667_,
		_w8669_,
		_w8664_,
		_w8670_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4623 (
		_w8658_,
		_w8660_,
		_w8661_,
		_w8670_,
		_w8671_
	);
	LUT2 #(
		.INIT('h8)
	) name4624 (
		_w8602_,
		_w8671_,
		_w8672_
	);
	LUT4 #(
		.INIT('h0007)
	) name4625 (
		_w6039_,
		_w8603_,
		_w8653_,
		_w8672_,
		_w8673_
	);
	LUT3 #(
		.INIT('hce)
	) name4626 (
		_w8601_,
		_w8652_,
		_w8673_,
		_w8674_
	);
	LUT2 #(
		.INIT('h8)
	) name4627 (
		\bdma_BCTL_reg[12]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8675_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4628 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w8594_,
		_w8602_,
		_w8676_
	);
	LUT3 #(
		.INIT('h70)
	) name4629 (
		_w6348_,
		_w6355_,
		_w8609_,
		_w8677_
	);
	LUT3 #(
		.INIT('h70)
	) name4630 (
		_w6337_,
		_w6344_,
		_w8605_,
		_w8678_
	);
	LUT3 #(
		.INIT('h70)
	) name4631 (
		_w5746_,
		_w6329_,
		_w8607_,
		_w8679_
	);
	LUT3 #(
		.INIT('h01)
	) name4632 (
		_w8678_,
		_w8679_,
		_w8677_,
		_w8680_
	);
	LUT4 #(
		.INIT('h5554)
	) name4633 (
		\emc_PMDoe_reg/NET0131 ,
		_w8678_,
		_w8679_,
		_w8677_,
		_w8681_
	);
	LUT2 #(
		.INIT('h8)
	) name4634 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[11]/P0001 ,
		_w8682_
	);
	LUT4 #(
		.INIT('h0080)
	) name4635 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8682_,
		_w8683_
	);
	LUT4 #(
		.INIT('haa80)
	) name4636 (
		\PM_rd0[11]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8684_
	);
	LUT4 #(
		.INIT('h8000)
	) name4637 (
		\PM_rd3[11]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8685_
	);
	LUT4 #(
		.INIT('h8000)
	) name4638 (
		\PM_rd1[11]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8686_
	);
	LUT4 #(
		.INIT('h0007)
	) name4639 (
		\PM_rd5[11]_pad ,
		_w8633_,
		_w8685_,
		_w8686_,
		_w8687_
	);
	LUT3 #(
		.INIT('h80)
	) name4640 (
		\PM_rd7[11]_pad ,
		_w8621_,
		_w8623_,
		_w8688_
	);
	LUT4 #(
		.INIT('h2000)
	) name4641 (
		\PM_rd6[11]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8689_
	);
	LUT3 #(
		.INIT('h01)
	) name4642 (
		_w8617_,
		_w8689_,
		_w8688_,
		_w8690_
	);
	LUT4 #(
		.INIT('h8000)
	) name4643 (
		\PM_rd2[11]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8691_
	);
	LUT3 #(
		.INIT('h07)
	) name4644 (
		\PM_rd4[11]_pad ,
		_w8627_,
		_w8691_,
		_w8692_
	);
	LUT3 #(
		.INIT('h80)
	) name4645 (
		_w8690_,
		_w8692_,
		_w8687_,
		_w8693_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4646 (
		_w8681_,
		_w8683_,
		_w8684_,
		_w8693_,
		_w8694_
	);
	LUT2 #(
		.INIT('h8)
	) name4647 (
		_w8602_,
		_w8694_,
		_w8695_
	);
	LUT4 #(
		.INIT('h0007)
	) name4648 (
		_w6363_,
		_w8603_,
		_w8676_,
		_w8695_,
		_w8696_
	);
	LUT3 #(
		.INIT('hce)
	) name4649 (
		_w8601_,
		_w8675_,
		_w8696_,
		_w8697_
	);
	LUT2 #(
		.INIT('h8)
	) name4650 (
		\bdma_BCTL_reg[13]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8698_
	);
	LUT4 #(
		.INIT('h0008)
	) name4651 (
		\emc_selDMDi_reg/P0001 ,
		_w6758_,
		_w8594_,
		_w8602_,
		_w8699_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4652 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w8594_,
		_w8602_,
		_w8700_
	);
	LUT3 #(
		.INIT('h70)
	) name4653 (
		_w6745_,
		_w6751_,
		_w8609_,
		_w8701_
	);
	LUT3 #(
		.INIT('h70)
	) name4654 (
		_w6733_,
		_w6740_,
		_w8605_,
		_w8702_
	);
	LUT3 #(
		.INIT('h70)
	) name4655 (
		_w5746_,
		_w6725_,
		_w8607_,
		_w8703_
	);
	LUT4 #(
		.INIT('h5554)
	) name4656 (
		\emc_PMDoe_reg/NET0131 ,
		_w8702_,
		_w8703_,
		_w8701_,
		_w8704_
	);
	LUT2 #(
		.INIT('h8)
	) name4657 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[12]/P0001 ,
		_w8705_
	);
	LUT4 #(
		.INIT('h0080)
	) name4658 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8705_,
		_w8706_
	);
	LUT4 #(
		.INIT('haa80)
	) name4659 (
		\PM_rd0[12]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8707_
	);
	LUT4 #(
		.INIT('h8000)
	) name4660 (
		\PM_rd3[12]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8708_
	);
	LUT4 #(
		.INIT('h8000)
	) name4661 (
		\PM_rd1[12]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8709_
	);
	LUT4 #(
		.INIT('h0007)
	) name4662 (
		\PM_rd5[12]_pad ,
		_w8633_,
		_w8708_,
		_w8709_,
		_w8710_
	);
	LUT3 #(
		.INIT('h80)
	) name4663 (
		\PM_rd7[12]_pad ,
		_w8621_,
		_w8623_,
		_w8711_
	);
	LUT4 #(
		.INIT('h2000)
	) name4664 (
		\PM_rd6[12]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8712_
	);
	LUT3 #(
		.INIT('h01)
	) name4665 (
		_w8617_,
		_w8712_,
		_w8711_,
		_w8713_
	);
	LUT4 #(
		.INIT('h8000)
	) name4666 (
		\PM_rd2[12]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8714_
	);
	LUT3 #(
		.INIT('h07)
	) name4667 (
		\PM_rd4[12]_pad ,
		_w8627_,
		_w8714_,
		_w8715_
	);
	LUT3 #(
		.INIT('h80)
	) name4668 (
		_w8713_,
		_w8715_,
		_w8710_,
		_w8716_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4669 (
		_w8704_,
		_w8706_,
		_w8707_,
		_w8716_,
		_w8717_
	);
	LUT2 #(
		.INIT('h8)
	) name4670 (
		_w8602_,
		_w8717_,
		_w8718_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4671 (
		_w8601_,
		_w8700_,
		_w8699_,
		_w8718_,
		_w8719_
	);
	LUT2 #(
		.INIT('he)
	) name4672 (
		_w8698_,
		_w8719_,
		_w8720_
	);
	LUT2 #(
		.INIT('h8)
	) name4673 (
		\bdma_BCTL_reg[14]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8721_
	);
	LUT4 #(
		.INIT('h0008)
	) name4674 (
		\emc_selDMDi_reg/P0001 ,
		_w5760_,
		_w8594_,
		_w8602_,
		_w8722_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4675 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w8594_,
		_w8602_,
		_w8723_
	);
	LUT3 #(
		.INIT('h70)
	) name4676 (
		_w5733_,
		_w5739_,
		_w8609_,
		_w8724_
	);
	LUT3 #(
		.INIT('h70)
	) name4677 (
		_w5719_,
		_w5728_,
		_w8605_,
		_w8725_
	);
	LUT3 #(
		.INIT('h70)
	) name4678 (
		_w5746_,
		_w5753_,
		_w8607_,
		_w8726_
	);
	LUT4 #(
		.INIT('h5554)
	) name4679 (
		\emc_PMDoe_reg/NET0131 ,
		_w8725_,
		_w8726_,
		_w8724_,
		_w8727_
	);
	LUT2 #(
		.INIT('h8)
	) name4680 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[13]/P0001 ,
		_w8728_
	);
	LUT4 #(
		.INIT('h0080)
	) name4681 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8728_,
		_w8729_
	);
	LUT4 #(
		.INIT('haa80)
	) name4682 (
		\PM_rd0[13]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8730_
	);
	LUT4 #(
		.INIT('h8000)
	) name4683 (
		\PM_rd3[13]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8731_
	);
	LUT4 #(
		.INIT('h8000)
	) name4684 (
		\PM_rd1[13]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8732_
	);
	LUT4 #(
		.INIT('h0007)
	) name4685 (
		\PM_rd5[13]_pad ,
		_w8633_,
		_w8731_,
		_w8732_,
		_w8733_
	);
	LUT3 #(
		.INIT('h80)
	) name4686 (
		\PM_rd7[13]_pad ,
		_w8621_,
		_w8623_,
		_w8734_
	);
	LUT4 #(
		.INIT('h2000)
	) name4687 (
		\PM_rd6[13]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8735_
	);
	LUT3 #(
		.INIT('h01)
	) name4688 (
		_w8617_,
		_w8735_,
		_w8734_,
		_w8736_
	);
	LUT4 #(
		.INIT('h8000)
	) name4689 (
		\PM_rd2[13]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8737_
	);
	LUT3 #(
		.INIT('h07)
	) name4690 (
		\PM_rd4[13]_pad ,
		_w8627_,
		_w8737_,
		_w8738_
	);
	LUT3 #(
		.INIT('h80)
	) name4691 (
		_w8736_,
		_w8738_,
		_w8733_,
		_w8739_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4692 (
		_w8727_,
		_w8729_,
		_w8730_,
		_w8739_,
		_w8740_
	);
	LUT2 #(
		.INIT('h8)
	) name4693 (
		_w8602_,
		_w8740_,
		_w8741_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4694 (
		_w8601_,
		_w8723_,
		_w8722_,
		_w8741_,
		_w8742_
	);
	LUT2 #(
		.INIT('he)
	) name4695 (
		_w8721_,
		_w8742_,
		_w8743_
	);
	LUT2 #(
		.INIT('h8)
	) name4696 (
		\bdma_BCTL_reg[15]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8744_
	);
	LUT3 #(
		.INIT('ha8)
	) name4697 (
		\DM_rd0[14]_pad ,
		_w5610_,
		_w5612_,
		_w8745_
	);
	LUT4 #(
		.INIT('h135f)
	) name4698 (
		\DM_rdm[14]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w8746_
	);
	LUT4 #(
		.INIT('h135f)
	) name4699 (
		\DM_rd6[14]_pad ,
		\DM_rd7[14]_pad ,
		_w5596_,
		_w5591_,
		_w8747_
	);
	LUT2 #(
		.INIT('h8)
	) name4700 (
		_w8746_,
		_w8747_,
		_w8748_
	);
	LUT3 #(
		.INIT('h80)
	) name4701 (
		\DM_rd5[14]_pad ,
		_w5598_,
		_w5599_,
		_w8749_
	);
	LUT3 #(
		.INIT('h80)
	) name4702 (
		\DM_rd4[14]_pad ,
		_w5598_,
		_w5601_,
		_w8750_
	);
	LUT4 #(
		.INIT('h8000)
	) name4703 (
		\DM_rd2[14]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w8751_
	);
	LUT4 #(
		.INIT('h8000)
	) name4704 (
		\DM_rd1[14]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w8752_
	);
	LUT4 #(
		.INIT('h8000)
	) name4705 (
		\DM_rd3[14]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w8753_
	);
	LUT3 #(
		.INIT('h01)
	) name4706 (
		_w8752_,
		_w8753_,
		_w8751_,
		_w8754_
	);
	LUT3 #(
		.INIT('h10)
	) name4707 (
		_w8750_,
		_w8749_,
		_w8754_,
		_w8755_
	);
	LUT2 #(
		.INIT('h8)
	) name4708 (
		_w8748_,
		_w8755_,
		_w8756_
	);
	LUT2 #(
		.INIT('h4)
	) name4709 (
		_w8745_,
		_w8756_,
		_w8757_
	);
	LUT2 #(
		.INIT('h8)
	) name4710 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[14]/P0001 ,
		_w8758_
	);
	LUT3 #(
		.INIT('h08)
	) name4711 (
		_w5588_,
		_w5598_,
		_w8758_,
		_w8759_
	);
	LUT4 #(
		.INIT('hba00)
	) name4712 (
		\emc_DMDoe_reg/NET0131 ,
		_w8237_,
		_w8308_,
		_w8759_,
		_w8760_
	);
	LUT2 #(
		.INIT('h1)
	) name4713 (
		_w8757_,
		_w8760_,
		_w8761_
	);
	LUT4 #(
		.INIT('h0200)
	) name4714 (
		\emc_selDMDi_reg/P0001 ,
		_w8594_,
		_w8602_,
		_w8761_,
		_w8762_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4715 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w8594_,
		_w8602_,
		_w8763_
	);
	LUT3 #(
		.INIT('h70)
	) name4716 (
		_w8298_,
		_w8305_,
		_w8605_,
		_w8764_
	);
	LUT3 #(
		.INIT('h70)
	) name4717 (
		_w8266_,
		_w8273_,
		_w8609_,
		_w8765_
	);
	LUT3 #(
		.INIT('h70)
	) name4718 (
		_w5746_,
		_w8290_,
		_w8607_,
		_w8766_
	);
	LUT3 #(
		.INIT('h01)
	) name4719 (
		_w8765_,
		_w8766_,
		_w8764_,
		_w8767_
	);
	LUT4 #(
		.INIT('h5554)
	) name4720 (
		\emc_PMDoe_reg/NET0131 ,
		_w8765_,
		_w8766_,
		_w8764_,
		_w8768_
	);
	LUT2 #(
		.INIT('h8)
	) name4721 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[14]/P0001 ,
		_w8769_
	);
	LUT4 #(
		.INIT('h0080)
	) name4722 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8769_,
		_w8770_
	);
	LUT4 #(
		.INIT('haa80)
	) name4723 (
		\PM_rd0[14]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8771_
	);
	LUT4 #(
		.INIT('h8000)
	) name4724 (
		\PM_rd3[14]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8772_
	);
	LUT4 #(
		.INIT('h8000)
	) name4725 (
		\PM_rd1[14]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8773_
	);
	LUT4 #(
		.INIT('h0007)
	) name4726 (
		\PM_rd5[14]_pad ,
		_w8633_,
		_w8772_,
		_w8773_,
		_w8774_
	);
	LUT3 #(
		.INIT('h80)
	) name4727 (
		\PM_rd7[14]_pad ,
		_w8621_,
		_w8623_,
		_w8775_
	);
	LUT4 #(
		.INIT('h2000)
	) name4728 (
		\PM_rd6[14]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8776_
	);
	LUT3 #(
		.INIT('h01)
	) name4729 (
		_w8617_,
		_w8776_,
		_w8775_,
		_w8777_
	);
	LUT4 #(
		.INIT('h8000)
	) name4730 (
		\PM_rd2[14]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8778_
	);
	LUT3 #(
		.INIT('h07)
	) name4731 (
		\PM_rd4[14]_pad ,
		_w8627_,
		_w8778_,
		_w8779_
	);
	LUT3 #(
		.INIT('h80)
	) name4732 (
		_w8777_,
		_w8779_,
		_w8774_,
		_w8780_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4733 (
		_w8768_,
		_w8770_,
		_w8771_,
		_w8780_,
		_w8781_
	);
	LUT2 #(
		.INIT('h8)
	) name4734 (
		_w8602_,
		_w8781_,
		_w8782_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4735 (
		_w8601_,
		_w8763_,
		_w8762_,
		_w8782_,
		_w8783_
	);
	LUT2 #(
		.INIT('he)
	) name4736 (
		_w8744_,
		_w8783_,
		_w8784_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4737 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w8594_,
		_w8602_,
		_w8785_
	);
	LUT3 #(
		.INIT('ha8)
	) name4738 (
		\DM_rd0[15]_pad ,
		_w5610_,
		_w5612_,
		_w8786_
	);
	LUT4 #(
		.INIT('h135f)
	) name4739 (
		\DM_rdm[15]_pad ,
		_w5588_,
		_w5593_,
		_w5598_,
		_w8787_
	);
	LUT4 #(
		.INIT('h135f)
	) name4740 (
		\DM_rd6[15]_pad ,
		\DM_rd7[15]_pad ,
		_w5596_,
		_w5591_,
		_w8788_
	);
	LUT2 #(
		.INIT('h8)
	) name4741 (
		_w8787_,
		_w8788_,
		_w8789_
	);
	LUT3 #(
		.INIT('h80)
	) name4742 (
		\DM_rd5[15]_pad ,
		_w5598_,
		_w5599_,
		_w8790_
	);
	LUT3 #(
		.INIT('h80)
	) name4743 (
		\DM_rd4[15]_pad ,
		_w5598_,
		_w5601_,
		_w8791_
	);
	LUT4 #(
		.INIT('h8000)
	) name4744 (
		\DM_rd2[15]_pad ,
		_w5589_,
		_w5594_,
		_w5603_,
		_w8792_
	);
	LUT4 #(
		.INIT('h8000)
	) name4745 (
		\DM_rd1[15]_pad ,
		_w5589_,
		_w5594_,
		_w5605_,
		_w8793_
	);
	LUT4 #(
		.INIT('h8000)
	) name4746 (
		\DM_rd3[15]_pad ,
		_w5587_,
		_w5594_,
		_w5607_,
		_w8794_
	);
	LUT3 #(
		.INIT('h01)
	) name4747 (
		_w8793_,
		_w8794_,
		_w8792_,
		_w8795_
	);
	LUT3 #(
		.INIT('h10)
	) name4748 (
		_w8791_,
		_w8790_,
		_w8795_,
		_w8796_
	);
	LUT2 #(
		.INIT('h8)
	) name4749 (
		_w8789_,
		_w8796_,
		_w8797_
	);
	LUT2 #(
		.INIT('h4)
	) name4750 (
		_w8786_,
		_w8797_,
		_w8798_
	);
	LUT2 #(
		.INIT('h8)
	) name4751 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[15]/P0001 ,
		_w8799_
	);
	LUT3 #(
		.INIT('h08)
	) name4752 (
		_w5588_,
		_w5598_,
		_w8799_,
		_w8800_
	);
	LUT4 #(
		.INIT('hba00)
	) name4753 (
		\emc_DMDoe_reg/NET0131 ,
		_w8318_,
		_w8387_,
		_w8800_,
		_w8801_
	);
	LUT2 #(
		.INIT('h1)
	) name4754 (
		_w8798_,
		_w8801_,
		_w8802_
	);
	LUT4 #(
		.INIT('h0200)
	) name4755 (
		\emc_selDMDi_reg/P0001 ,
		_w8594_,
		_w8602_,
		_w8802_,
		_w8803_
	);
	LUT3 #(
		.INIT('h70)
	) name4756 (
		_w8377_,
		_w8384_,
		_w8605_,
		_w8804_
	);
	LUT3 #(
		.INIT('h70)
	) name4757 (
		_w8348_,
		_w8354_,
		_w8609_,
		_w8805_
	);
	LUT3 #(
		.INIT('h70)
	) name4758 (
		_w5746_,
		_w8369_,
		_w8607_,
		_w8806_
	);
	LUT3 #(
		.INIT('h01)
	) name4759 (
		_w8805_,
		_w8806_,
		_w8804_,
		_w8807_
	);
	LUT4 #(
		.INIT('h5554)
	) name4760 (
		\emc_PMDoe_reg/NET0131 ,
		_w8805_,
		_w8806_,
		_w8804_,
		_w8808_
	);
	LUT2 #(
		.INIT('h8)
	) name4761 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[15]/P0001 ,
		_w8809_
	);
	LUT4 #(
		.INIT('h0080)
	) name4762 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8809_,
		_w8810_
	);
	LUT4 #(
		.INIT('haa80)
	) name4763 (
		\PM_rd0[15]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8811_
	);
	LUT4 #(
		.INIT('h8000)
	) name4764 (
		\PM_rd3[15]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8812_
	);
	LUT4 #(
		.INIT('h8000)
	) name4765 (
		\PM_rd1[15]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8813_
	);
	LUT4 #(
		.INIT('h0007)
	) name4766 (
		\PM_rd5[15]_pad ,
		_w8633_,
		_w8812_,
		_w8813_,
		_w8814_
	);
	LUT3 #(
		.INIT('h80)
	) name4767 (
		\PM_rd7[15]_pad ,
		_w8621_,
		_w8623_,
		_w8815_
	);
	LUT4 #(
		.INIT('h2000)
	) name4768 (
		\PM_rd6[15]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8816_
	);
	LUT3 #(
		.INIT('h01)
	) name4769 (
		_w8617_,
		_w8816_,
		_w8815_,
		_w8817_
	);
	LUT4 #(
		.INIT('h8000)
	) name4770 (
		\PM_rd2[15]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8818_
	);
	LUT3 #(
		.INIT('h07)
	) name4771 (
		\PM_rd4[15]_pad ,
		_w8627_,
		_w8818_,
		_w8819_
	);
	LUT3 #(
		.INIT('h80)
	) name4772 (
		_w8817_,
		_w8819_,
		_w8814_,
		_w8820_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4773 (
		_w8808_,
		_w8810_,
		_w8811_,
		_w8820_,
		_w8821_
	);
	LUT2 #(
		.INIT('h8)
	) name4774 (
		_w8602_,
		_w8821_,
		_w8822_
	);
	LUT3 #(
		.INIT('hfe)
	) name4775 (
		_w8803_,
		_w8785_,
		_w8822_,
		_w8823_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4776 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w8594_,
		_w8602_,
		_w8824_
	);
	LUT3 #(
		.INIT('h70)
	) name4777 (
		_w6866_,
		_w6875_,
		_w8605_,
		_w8825_
	);
	LUT3 #(
		.INIT('h70)
	) name4778 (
		_w6881_,
		_w6888_,
		_w8607_,
		_w8826_
	);
	LUT3 #(
		.INIT('h70)
	) name4779 (
		_w6851_,
		_w6858_,
		_w8609_,
		_w8827_
	);
	LUT4 #(
		.INIT('h5554)
	) name4780 (
		\emc_PMDoe_reg/NET0131 ,
		_w8826_,
		_w8827_,
		_w8825_,
		_w8828_
	);
	LUT2 #(
		.INIT('h8)
	) name4781 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[1]/P0001 ,
		_w8829_
	);
	LUT4 #(
		.INIT('h0080)
	) name4782 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8829_,
		_w8830_
	);
	LUT4 #(
		.INIT('haa80)
	) name4783 (
		\PM_rd0[1]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8831_
	);
	LUT4 #(
		.INIT('h8000)
	) name4784 (
		\PM_rd3[1]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8832_
	);
	LUT4 #(
		.INIT('h8000)
	) name4785 (
		\PM_rd1[1]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8833_
	);
	LUT4 #(
		.INIT('h0007)
	) name4786 (
		\PM_rd5[1]_pad ,
		_w8633_,
		_w8832_,
		_w8833_,
		_w8834_
	);
	LUT3 #(
		.INIT('h80)
	) name4787 (
		\PM_rd7[1]_pad ,
		_w8621_,
		_w8623_,
		_w8835_
	);
	LUT4 #(
		.INIT('h2000)
	) name4788 (
		\PM_rd6[1]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8836_
	);
	LUT3 #(
		.INIT('h01)
	) name4789 (
		_w8617_,
		_w8836_,
		_w8835_,
		_w8837_
	);
	LUT4 #(
		.INIT('h8000)
	) name4790 (
		\PM_rd2[1]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8838_
	);
	LUT3 #(
		.INIT('h07)
	) name4791 (
		\PM_rd4[1]_pad ,
		_w8627_,
		_w8838_,
		_w8839_
	);
	LUT3 #(
		.INIT('h80)
	) name4792 (
		_w8837_,
		_w8839_,
		_w8834_,
		_w8840_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4793 (
		_w8828_,
		_w8830_,
		_w8831_,
		_w8840_,
		_w8841_
	);
	LUT2 #(
		.INIT('h8)
	) name4794 (
		_w8602_,
		_w8841_,
		_w8842_
	);
	LUT4 #(
		.INIT('h0007)
	) name4795 (
		_w6897_,
		_w8603_,
		_w8824_,
		_w8842_,
		_w8843_
	);
	LUT3 #(
		.INIT('h80)
	) name4796 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWdataBUF_reg[1]/P0001 ,
		_w8844_
	);
	LUT3 #(
		.INIT('hf2)
	) name4797 (
		_w8601_,
		_w8843_,
		_w8844_,
		_w8845_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4798 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w8594_,
		_w8602_,
		_w8846_
	);
	LUT3 #(
		.INIT('h70)
	) name4799 (
		_w6468_,
		_w6475_,
		_w8607_,
		_w8847_
	);
	LUT3 #(
		.INIT('h70)
	) name4800 (
		_w6483_,
		_w6492_,
		_w8605_,
		_w8848_
	);
	LUT3 #(
		.INIT('h70)
	) name4801 (
		_w6455_,
		_w6462_,
		_w8609_,
		_w8849_
	);
	LUT4 #(
		.INIT('h5554)
	) name4802 (
		\emc_PMDoe_reg/NET0131 ,
		_w8848_,
		_w8849_,
		_w8847_,
		_w8850_
	);
	LUT2 #(
		.INIT('h8)
	) name4803 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[2]/P0001 ,
		_w8851_
	);
	LUT4 #(
		.INIT('h0080)
	) name4804 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8851_,
		_w8852_
	);
	LUT4 #(
		.INIT('haa80)
	) name4805 (
		\PM_rd0[2]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8853_
	);
	LUT4 #(
		.INIT('h8000)
	) name4806 (
		\PM_rd3[2]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8854_
	);
	LUT4 #(
		.INIT('h8000)
	) name4807 (
		\PM_rd1[2]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8855_
	);
	LUT4 #(
		.INIT('h0007)
	) name4808 (
		\PM_rd5[2]_pad ,
		_w8633_,
		_w8854_,
		_w8855_,
		_w8856_
	);
	LUT3 #(
		.INIT('h80)
	) name4809 (
		\PM_rd7[2]_pad ,
		_w8621_,
		_w8623_,
		_w8857_
	);
	LUT4 #(
		.INIT('h2000)
	) name4810 (
		\PM_rd6[2]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8858_
	);
	LUT3 #(
		.INIT('h01)
	) name4811 (
		_w8617_,
		_w8858_,
		_w8857_,
		_w8859_
	);
	LUT4 #(
		.INIT('h8000)
	) name4812 (
		\PM_rd2[2]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8860_
	);
	LUT3 #(
		.INIT('h07)
	) name4813 (
		\PM_rd4[2]_pad ,
		_w8627_,
		_w8860_,
		_w8861_
	);
	LUT3 #(
		.INIT('h80)
	) name4814 (
		_w8859_,
		_w8861_,
		_w8856_,
		_w8862_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4815 (
		_w8850_,
		_w8852_,
		_w8853_,
		_w8862_,
		_w8863_
	);
	LUT2 #(
		.INIT('h8)
	) name4816 (
		_w8602_,
		_w8863_,
		_w8864_
	);
	LUT4 #(
		.INIT('h0007)
	) name4817 (
		_w6501_,
		_w8603_,
		_w8846_,
		_w8864_,
		_w8865_
	);
	LUT3 #(
		.INIT('h80)
	) name4818 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWdataBUF_reg[2]/P0001 ,
		_w8866_
	);
	LUT3 #(
		.INIT('hf2)
	) name4819 (
		_w8601_,
		_w8865_,
		_w8866_,
		_w8867_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4820 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w8594_,
		_w8602_,
		_w8868_
	);
	LUT3 #(
		.INIT('h70)
	) name4821 (
		_w6147_,
		_w6156_,
		_w8605_,
		_w8869_
	);
	LUT3 #(
		.INIT('h70)
	) name4822 (
		_w6132_,
		_w6139_,
		_w8607_,
		_w8870_
	);
	LUT3 #(
		.INIT('h70)
	) name4823 (
		_w6161_,
		_w6167_,
		_w8609_,
		_w8871_
	);
	LUT4 #(
		.INIT('h5554)
	) name4824 (
		\emc_PMDoe_reg/NET0131 ,
		_w8870_,
		_w8871_,
		_w8869_,
		_w8872_
	);
	LUT2 #(
		.INIT('h8)
	) name4825 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[3]/P0001 ,
		_w8873_
	);
	LUT4 #(
		.INIT('h0080)
	) name4826 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8873_,
		_w8874_
	);
	LUT4 #(
		.INIT('haa80)
	) name4827 (
		\PM_rd0[3]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8875_
	);
	LUT4 #(
		.INIT('h8000)
	) name4828 (
		\PM_rd3[3]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8876_
	);
	LUT4 #(
		.INIT('h8000)
	) name4829 (
		\PM_rd1[3]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8877_
	);
	LUT4 #(
		.INIT('h0007)
	) name4830 (
		\PM_rd5[3]_pad ,
		_w8633_,
		_w8876_,
		_w8877_,
		_w8878_
	);
	LUT3 #(
		.INIT('h80)
	) name4831 (
		\PM_rd7[3]_pad ,
		_w8621_,
		_w8623_,
		_w8879_
	);
	LUT4 #(
		.INIT('h2000)
	) name4832 (
		\PM_rd6[3]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8880_
	);
	LUT3 #(
		.INIT('h01)
	) name4833 (
		_w8617_,
		_w8880_,
		_w8879_,
		_w8881_
	);
	LUT4 #(
		.INIT('h8000)
	) name4834 (
		\PM_rd2[3]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8882_
	);
	LUT3 #(
		.INIT('h07)
	) name4835 (
		\PM_rd4[3]_pad ,
		_w8627_,
		_w8882_,
		_w8883_
	);
	LUT3 #(
		.INIT('h80)
	) name4836 (
		_w8881_,
		_w8883_,
		_w8878_,
		_w8884_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4837 (
		_w8872_,
		_w8874_,
		_w8875_,
		_w8884_,
		_w8885_
	);
	LUT2 #(
		.INIT('h8)
	) name4838 (
		_w8602_,
		_w8885_,
		_w8886_
	);
	LUT4 #(
		.INIT('h0007)
	) name4839 (
		_w6176_,
		_w8603_,
		_w8868_,
		_w8886_,
		_w8887_
	);
	LUT3 #(
		.INIT('h80)
	) name4840 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWdataBUF_reg[3]/P0001 ,
		_w8888_
	);
	LUT3 #(
		.INIT('hf2)
	) name4841 (
		_w8601_,
		_w8887_,
		_w8888_,
		_w8889_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4842 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w8594_,
		_w8602_,
		_w8890_
	);
	LUT3 #(
		.INIT('h70)
	) name4843 (
		_w7348_,
		_w7357_,
		_w8605_,
		_w8891_
	);
	LUT3 #(
		.INIT('h70)
	) name4844 (
		_w7362_,
		_w7369_,
		_w8609_,
		_w8892_
	);
	LUT3 #(
		.INIT('h70)
	) name4845 (
		_w7333_,
		_w7340_,
		_w8607_,
		_w8893_
	);
	LUT4 #(
		.INIT('h5554)
	) name4846 (
		\emc_PMDoe_reg/NET0131 ,
		_w8892_,
		_w8893_,
		_w8891_,
		_w8894_
	);
	LUT2 #(
		.INIT('h8)
	) name4847 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[4]/P0001 ,
		_w8895_
	);
	LUT4 #(
		.INIT('h0080)
	) name4848 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8895_,
		_w8896_
	);
	LUT4 #(
		.INIT('haa80)
	) name4849 (
		\PM_rd0[4]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8897_
	);
	LUT4 #(
		.INIT('h8000)
	) name4850 (
		\PM_rd3[4]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8898_
	);
	LUT4 #(
		.INIT('h8000)
	) name4851 (
		\PM_rd1[4]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8899_
	);
	LUT4 #(
		.INIT('h0007)
	) name4852 (
		\PM_rd5[4]_pad ,
		_w8633_,
		_w8898_,
		_w8899_,
		_w8900_
	);
	LUT3 #(
		.INIT('h80)
	) name4853 (
		\PM_rd7[4]_pad ,
		_w8621_,
		_w8623_,
		_w8901_
	);
	LUT4 #(
		.INIT('h2000)
	) name4854 (
		\PM_rd6[4]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8902_
	);
	LUT3 #(
		.INIT('h01)
	) name4855 (
		_w8617_,
		_w8902_,
		_w8901_,
		_w8903_
	);
	LUT4 #(
		.INIT('h8000)
	) name4856 (
		\PM_rd2[4]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8904_
	);
	LUT3 #(
		.INIT('h07)
	) name4857 (
		\PM_rd4[4]_pad ,
		_w8627_,
		_w8904_,
		_w8905_
	);
	LUT3 #(
		.INIT('h80)
	) name4858 (
		_w8903_,
		_w8905_,
		_w8900_,
		_w8906_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4859 (
		_w8894_,
		_w8896_,
		_w8897_,
		_w8906_,
		_w8907_
	);
	LUT2 #(
		.INIT('h8)
	) name4860 (
		_w8602_,
		_w8907_,
		_w8908_
	);
	LUT4 #(
		.INIT('h0007)
	) name4861 (
		_w7378_,
		_w8603_,
		_w8890_,
		_w8908_,
		_w8909_
	);
	LUT3 #(
		.INIT('h80)
	) name4862 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWdataBUF_reg[4]/P0001 ,
		_w8910_
	);
	LUT3 #(
		.INIT('hf2)
	) name4863 (
		_w8601_,
		_w8909_,
		_w8910_,
		_w8911_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4864 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w8594_,
		_w8602_,
		_w8912_
	);
	LUT3 #(
		.INIT('h70)
	) name4865 (
		_w7670_,
		_w7679_,
		_w8605_,
		_w8913_
	);
	LUT3 #(
		.INIT('h70)
	) name4866 (
		_w7684_,
		_w7690_,
		_w8609_,
		_w8914_
	);
	LUT3 #(
		.INIT('h70)
	) name4867 (
		_w7694_,
		_w7701_,
		_w8607_,
		_w8915_
	);
	LUT4 #(
		.INIT('h5554)
	) name4868 (
		\emc_PMDoe_reg/NET0131 ,
		_w8914_,
		_w8915_,
		_w8913_,
		_w8916_
	);
	LUT2 #(
		.INIT('h8)
	) name4869 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[5]/P0001 ,
		_w8917_
	);
	LUT4 #(
		.INIT('h0080)
	) name4870 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8917_,
		_w8918_
	);
	LUT4 #(
		.INIT('haa80)
	) name4871 (
		\PM_rd0[5]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8919_
	);
	LUT4 #(
		.INIT('h8000)
	) name4872 (
		\PM_rd3[5]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8920_
	);
	LUT4 #(
		.INIT('h8000)
	) name4873 (
		\PM_rd1[5]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8921_
	);
	LUT4 #(
		.INIT('h0007)
	) name4874 (
		\PM_rd5[5]_pad ,
		_w8633_,
		_w8920_,
		_w8921_,
		_w8922_
	);
	LUT3 #(
		.INIT('h80)
	) name4875 (
		\PM_rd7[5]_pad ,
		_w8621_,
		_w8623_,
		_w8923_
	);
	LUT4 #(
		.INIT('h2000)
	) name4876 (
		\PM_rd6[5]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8924_
	);
	LUT3 #(
		.INIT('h01)
	) name4877 (
		_w8617_,
		_w8924_,
		_w8923_,
		_w8925_
	);
	LUT4 #(
		.INIT('h8000)
	) name4878 (
		\PM_rd2[5]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8926_
	);
	LUT3 #(
		.INIT('h07)
	) name4879 (
		\PM_rd4[5]_pad ,
		_w8627_,
		_w8926_,
		_w8927_
	);
	LUT3 #(
		.INIT('h80)
	) name4880 (
		_w8925_,
		_w8927_,
		_w8922_,
		_w8928_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4881 (
		_w8916_,
		_w8918_,
		_w8919_,
		_w8928_,
		_w8929_
	);
	LUT2 #(
		.INIT('h8)
	) name4882 (
		_w8602_,
		_w8929_,
		_w8930_
	);
	LUT4 #(
		.INIT('h0007)
	) name4883 (
		_w7710_,
		_w8603_,
		_w8912_,
		_w8930_,
		_w8931_
	);
	LUT3 #(
		.INIT('h80)
	) name4884 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWdataBUF_reg[5]/P0001 ,
		_w8932_
	);
	LUT3 #(
		.INIT('hf2)
	) name4885 (
		_w8601_,
		_w8931_,
		_w8932_,
		_w8933_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4886 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w8594_,
		_w8602_,
		_w8934_
	);
	LUT4 #(
		.INIT('haa80)
	) name4887 (
		\PM_rd0[6]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8935_
	);
	LUT4 #(
		.INIT('h8000)
	) name4888 (
		\PM_rd1[6]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8936_
	);
	LUT4 #(
		.INIT('h8000)
	) name4889 (
		\PM_rd2[6]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8937_
	);
	LUT4 #(
		.INIT('h0007)
	) name4890 (
		\PM_rd5[6]_pad ,
		_w8633_,
		_w8937_,
		_w8936_,
		_w8938_
	);
	LUT3 #(
		.INIT('h80)
	) name4891 (
		\PM_rd7[6]_pad ,
		_w8621_,
		_w8623_,
		_w8939_
	);
	LUT4 #(
		.INIT('h2000)
	) name4892 (
		\PM_rd6[6]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8940_
	);
	LUT3 #(
		.INIT('h01)
	) name4893 (
		_w8617_,
		_w8940_,
		_w8939_,
		_w8941_
	);
	LUT4 #(
		.INIT('h8000)
	) name4894 (
		\PM_rd3[6]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8942_
	);
	LUT3 #(
		.INIT('h07)
	) name4895 (
		\PM_rd4[6]_pad ,
		_w8627_,
		_w8942_,
		_w8943_
	);
	LUT3 #(
		.INIT('h80)
	) name4896 (
		_w8941_,
		_w8943_,
		_w8938_,
		_w8944_
	);
	LUT2 #(
		.INIT('h4)
	) name4897 (
		_w8935_,
		_w8944_,
		_w8945_
	);
	LUT3 #(
		.INIT('h70)
	) name4898 (
		_w8025_,
		_w8034_,
		_w8605_,
		_w8946_
	);
	LUT3 #(
		.INIT('h70)
	) name4899 (
		_w8010_,
		_w8017_,
		_w8607_,
		_w8947_
	);
	LUT2 #(
		.INIT('h1)
	) name4900 (
		_w8946_,
		_w8947_,
		_w8948_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4901 (
		_w7929_,
		_w7940_,
		_w8609_,
		_w8948_,
		_w8949_
	);
	LUT2 #(
		.INIT('h8)
	) name4902 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[6]/P0001 ,
		_w8950_
	);
	LUT4 #(
		.INIT('h0080)
	) name4903 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8950_,
		_w8951_
	);
	LUT4 #(
		.INIT('h0133)
	) name4904 (
		\emc_PMDoe_reg/NET0131 ,
		_w8945_,
		_w8949_,
		_w8951_,
		_w8952_
	);
	LUT2 #(
		.INIT('h8)
	) name4905 (
		_w8602_,
		_w8952_,
		_w8953_
	);
	LUT4 #(
		.INIT('h0007)
	) name4906 (
		_w8043_,
		_w8603_,
		_w8934_,
		_w8953_,
		_w8954_
	);
	LUT3 #(
		.INIT('h80)
	) name4907 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWdataBUF_reg[6]/P0001 ,
		_w8955_
	);
	LUT3 #(
		.INIT('hf2)
	) name4908 (
		_w8601_,
		_w8954_,
		_w8955_,
		_w8956_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4909 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w8594_,
		_w8602_,
		_w8957_
	);
	LUT3 #(
		.INIT('h70)
	) name4910 (
		_w7890_,
		_w7897_,
		_w8605_,
		_w8958_
	);
	LUT3 #(
		.INIT('h70)
	) name4911 (
		_w7875_,
		_w7882_,
		_w8609_,
		_w8959_
	);
	LUT3 #(
		.INIT('h70)
	) name4912 (
		_w5746_,
		_w7870_,
		_w8607_,
		_w8960_
	);
	LUT4 #(
		.INIT('h5554)
	) name4913 (
		\emc_PMDoe_reg/NET0131 ,
		_w8959_,
		_w8960_,
		_w8958_,
		_w8961_
	);
	LUT2 #(
		.INIT('h8)
	) name4914 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[7]/P0001 ,
		_w8962_
	);
	LUT4 #(
		.INIT('h0080)
	) name4915 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8962_,
		_w8963_
	);
	LUT4 #(
		.INIT('haa80)
	) name4916 (
		\PM_rd0[7]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8964_
	);
	LUT4 #(
		.INIT('h8000)
	) name4917 (
		\PM_rd3[7]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8965_
	);
	LUT4 #(
		.INIT('h8000)
	) name4918 (
		\PM_rd1[7]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8966_
	);
	LUT4 #(
		.INIT('h0007)
	) name4919 (
		\PM_rd5[7]_pad ,
		_w8633_,
		_w8965_,
		_w8966_,
		_w8967_
	);
	LUT3 #(
		.INIT('h80)
	) name4920 (
		\PM_rd7[7]_pad ,
		_w8621_,
		_w8623_,
		_w8968_
	);
	LUT4 #(
		.INIT('h2000)
	) name4921 (
		\PM_rd6[7]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8969_
	);
	LUT3 #(
		.INIT('h01)
	) name4922 (
		_w8617_,
		_w8969_,
		_w8968_,
		_w8970_
	);
	LUT4 #(
		.INIT('h8000)
	) name4923 (
		\PM_rd2[7]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8971_
	);
	LUT3 #(
		.INIT('h07)
	) name4924 (
		\PM_rd4[7]_pad ,
		_w8627_,
		_w8971_,
		_w8972_
	);
	LUT3 #(
		.INIT('h80)
	) name4925 (
		_w8970_,
		_w8972_,
		_w8967_,
		_w8973_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4926 (
		_w8961_,
		_w8963_,
		_w8964_,
		_w8973_,
		_w8974_
	);
	LUT2 #(
		.INIT('h8)
	) name4927 (
		_w8602_,
		_w8974_,
		_w8975_
	);
	LUT4 #(
		.INIT('h0007)
	) name4928 (
		_w7906_,
		_w8603_,
		_w8957_,
		_w8975_,
		_w8976_
	);
	LUT3 #(
		.INIT('h80)
	) name4929 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWdataBUF_reg[7]/P0001 ,
		_w8977_
	);
	LUT3 #(
		.INIT('hf2)
	) name4930 (
		_w8601_,
		_w8976_,
		_w8977_,
		_w8978_
	);
	LUT2 #(
		.INIT('h8)
	) name4931 (
		\bdma_BCTL_reg[9]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w8979_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4932 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w8594_,
		_w8602_,
		_w8980_
	);
	LUT3 #(
		.INIT('h70)
	) name4933 (
		_w7537_,
		_w7543_,
		_w8609_,
		_w8981_
	);
	LUT3 #(
		.INIT('h70)
	) name4934 (
		_w7551_,
		_w7558_,
		_w8605_,
		_w8982_
	);
	LUT3 #(
		.INIT('h70)
	) name4935 (
		_w5746_,
		_w7532_,
		_w8607_,
		_w8983_
	);
	LUT3 #(
		.INIT('h01)
	) name4936 (
		_w8982_,
		_w8983_,
		_w8981_,
		_w8984_
	);
	LUT4 #(
		.INIT('h5554)
	) name4937 (
		\emc_PMDoe_reg/NET0131 ,
		_w8982_,
		_w8983_,
		_w8981_,
		_w8985_
	);
	LUT2 #(
		.INIT('h8)
	) name4938 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[8]/P0001 ,
		_w8986_
	);
	LUT4 #(
		.INIT('h0080)
	) name4939 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w8986_,
		_w8987_
	);
	LUT4 #(
		.INIT('haa80)
	) name4940 (
		\PM_rd0[8]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w8988_
	);
	LUT4 #(
		.INIT('h8000)
	) name4941 (
		\PM_rd3[8]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w8989_
	);
	LUT4 #(
		.INIT('h8000)
	) name4942 (
		\PM_rd1[8]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w8990_
	);
	LUT4 #(
		.INIT('h0007)
	) name4943 (
		\PM_rd5[8]_pad ,
		_w8633_,
		_w8989_,
		_w8990_,
		_w8991_
	);
	LUT3 #(
		.INIT('h80)
	) name4944 (
		\PM_rd7[8]_pad ,
		_w8621_,
		_w8623_,
		_w8992_
	);
	LUT4 #(
		.INIT('h2000)
	) name4945 (
		\PM_rd6[8]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w8993_
	);
	LUT3 #(
		.INIT('h01)
	) name4946 (
		_w8617_,
		_w8993_,
		_w8992_,
		_w8994_
	);
	LUT4 #(
		.INIT('h8000)
	) name4947 (
		\PM_rd2[8]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w8995_
	);
	LUT3 #(
		.INIT('h07)
	) name4948 (
		\PM_rd4[8]_pad ,
		_w8627_,
		_w8995_,
		_w8996_
	);
	LUT3 #(
		.INIT('h80)
	) name4949 (
		_w8994_,
		_w8996_,
		_w8991_,
		_w8997_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4950 (
		_w8985_,
		_w8987_,
		_w8988_,
		_w8997_,
		_w8998_
	);
	LUT2 #(
		.INIT('h8)
	) name4951 (
		_w8602_,
		_w8998_,
		_w8999_
	);
	LUT4 #(
		.INIT('h0007)
	) name4952 (
		_w7566_,
		_w8603_,
		_w8980_,
		_w8999_,
		_w9000_
	);
	LUT3 #(
		.INIT('hce)
	) name4953 (
		_w8601_,
		_w8979_,
		_w9000_,
		_w9001_
	);
	LUT2 #(
		.INIT('h8)
	) name4954 (
		\bdma_BCTL_reg[10]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w9002_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4955 (
		\emc_selDMDi_reg/P0001 ,
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w8594_,
		_w8602_,
		_w9003_
	);
	LUT3 #(
		.INIT('h70)
	) name4956 (
		_w7227_,
		_w7233_,
		_w8609_,
		_w9004_
	);
	LUT3 #(
		.INIT('h70)
	) name4957 (
		_w7215_,
		_w7222_,
		_w8605_,
		_w9005_
	);
	LUT3 #(
		.INIT('h70)
	) name4958 (
		_w5746_,
		_w7207_,
		_w8607_,
		_w9006_
	);
	LUT3 #(
		.INIT('h01)
	) name4959 (
		_w9005_,
		_w9006_,
		_w9004_,
		_w9007_
	);
	LUT4 #(
		.INIT('h5554)
	) name4960 (
		\emc_PMDoe_reg/NET0131 ,
		_w9005_,
		_w9006_,
		_w9004_,
		_w9008_
	);
	LUT2 #(
		.INIT('h8)
	) name4961 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[9]/P0001 ,
		_w9009_
	);
	LUT4 #(
		.INIT('h0080)
	) name4962 (
		_w8613_,
		_w8615_,
		_w8616_,
		_w9009_,
		_w9010_
	);
	LUT4 #(
		.INIT('haa80)
	) name4963 (
		\PM_rd0[9]_pad ,
		_w8625_,
		_w8634_,
		_w8636_,
		_w9011_
	);
	LUT4 #(
		.INIT('h8000)
	) name4964 (
		\PM_rd3[9]_pad ,
		_w8615_,
		_w8616_,
		_w8630_,
		_w9012_
	);
	LUT4 #(
		.INIT('h8000)
	) name4965 (
		\PM_rd1[9]_pad ,
		_w8613_,
		_w8615_,
		_w8628_,
		_w9013_
	);
	LUT4 #(
		.INIT('h0007)
	) name4966 (
		\PM_rd5[9]_pad ,
		_w8633_,
		_w9012_,
		_w9013_,
		_w9014_
	);
	LUT3 #(
		.INIT('h80)
	) name4967 (
		\PM_rd7[9]_pad ,
		_w8621_,
		_w8623_,
		_w9015_
	);
	LUT4 #(
		.INIT('h2000)
	) name4968 (
		\PM_rd6[9]_pad ,
		\memc_PMo_oe7_reg/P0001 ,
		_w8621_,
		_w8622_,
		_w9016_
	);
	LUT3 #(
		.INIT('h01)
	) name4969 (
		_w8617_,
		_w9016_,
		_w9015_,
		_w9017_
	);
	LUT4 #(
		.INIT('h8000)
	) name4970 (
		\PM_rd2[9]_pad ,
		_w8615_,
		_w8616_,
		_w8619_,
		_w9018_
	);
	LUT3 #(
		.INIT('h07)
	) name4971 (
		\PM_rd4[9]_pad ,
		_w8627_,
		_w9018_,
		_w9019_
	);
	LUT3 #(
		.INIT('h80)
	) name4972 (
		_w9017_,
		_w9019_,
		_w9014_,
		_w9020_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4973 (
		_w9008_,
		_w9010_,
		_w9011_,
		_w9020_,
		_w9021_
	);
	LUT2 #(
		.INIT('h8)
	) name4974 (
		_w8602_,
		_w9021_,
		_w9022_
	);
	LUT4 #(
		.INIT('h0007)
	) name4975 (
		_w7241_,
		_w8603_,
		_w9003_,
		_w9022_,
		_w9023_
	);
	LUT3 #(
		.INIT('hce)
	) name4976 (
		_w8601_,
		_w9002_,
		_w9023_,
		_w9024_
	);
	LUT3 #(
		.INIT('hba)
	) name4977 (
		\bdma_BM_cyc_reg/P0001 ,
		\core_c_psq_MGNT_reg/NET0131 ,
		\emc_ED_oei_reg/P0001 ,
		_w9025_
	);
	LUT4 #(
		.INIT('h8f88)
	) name4978 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\core_c_psq_MGNT_reg/NET0131 ,
		\emc_ED_oei_reg/P0001 ,
		_w9026_
	);
	LUT3 #(
		.INIT('h01)
	) name4979 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_L_reg[0]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9027_
	);
	LUT4 #(
		.INIT('h5051)
	) name4980 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[0]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9028_
	);
	LUT2 #(
		.INIT('h4)
	) name4981 (
		_w9027_,
		_w9028_,
		_w9029_
	);
	LUT4 #(
		.INIT('hfaea)
	) name4982 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[10]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9030_
	);
	LUT4 #(
		.INIT('h5040)
	) name4983 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[11]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9031_
	);
	LUT4 #(
		.INIT('h5040)
	) name4984 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[12]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9032_
	);
	LUT4 #(
		.INIT('hfaea)
	) name4985 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[13]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9033_
	);
	LUT4 #(
		.INIT('h5040)
	) name4986 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[14]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9034_
	);
	LUT4 #(
		.INIT('hfaea)
	) name4987 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[15]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9035_
	);
	LUT3 #(
		.INIT('h01)
	) name4988 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_L_reg[1]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9036_
	);
	LUT4 #(
		.INIT('h5051)
	) name4989 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[1]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9037_
	);
	LUT2 #(
		.INIT('h4)
	) name4990 (
		_w9036_,
		_w9037_,
		_w9038_
	);
	LUT3 #(
		.INIT('hc8)
	) name4991 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[2]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9039_
	);
	LUT4 #(
		.INIT('h5545)
	) name4992 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_L_reg[2]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9040_
	);
	LUT2 #(
		.INIT('hb)
	) name4993 (
		_w9039_,
		_w9040_,
		_w9041_
	);
	LUT3 #(
		.INIT('h01)
	) name4994 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_L_reg[3]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9042_
	);
	LUT4 #(
		.INIT('h5051)
	) name4995 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[3]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9043_
	);
	LUT2 #(
		.INIT('h4)
	) name4996 (
		_w9042_,
		_w9043_,
		_w9044_
	);
	LUT3 #(
		.INIT('h01)
	) name4997 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_L_reg[4]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9045_
	);
	LUT4 #(
		.INIT('h5051)
	) name4998 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[4]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9046_
	);
	LUT2 #(
		.INIT('h4)
	) name4999 (
		_w9045_,
		_w9046_,
		_w9047_
	);
	LUT3 #(
		.INIT('hc8)
	) name5000 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[5]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9048_
	);
	LUT4 #(
		.INIT('h5545)
	) name5001 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_L_reg[5]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9049_
	);
	LUT2 #(
		.INIT('hb)
	) name5002 (
		_w9048_,
		_w9049_,
		_w9050_
	);
	LUT3 #(
		.INIT('h01)
	) name5003 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_L_reg[6]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9051_
	);
	LUT4 #(
		.INIT('h5051)
	) name5004 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[6]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9052_
	);
	LUT2 #(
		.INIT('h4)
	) name5005 (
		_w9051_,
		_w9052_,
		_w9053_
	);
	LUT3 #(
		.INIT('hc8)
	) name5006 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[7]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9054_
	);
	LUT4 #(
		.INIT('h5545)
	) name5007 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_L_reg[7]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9055_
	);
	LUT2 #(
		.INIT('hb)
	) name5008 (
		_w9054_,
		_w9055_,
		_w9056_
	);
	LUT4 #(
		.INIT('h5040)
	) name5009 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[8]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9057_
	);
	LUT4 #(
		.INIT('h5040)
	) name5010 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_DTMP_H_reg[9]/P0001 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w9058_
	);
	LUT2 #(
		.INIT('he)
	) name5011 (
		\idma_RDCMD_reg/P0001 ,
		\idma_RDcyc_reg/NET0131 ,
		_w9059_
	);
	LUT2 #(
		.INIT('h4)
	) name5012 (
		T_IMS_pad,
		\sice_OE_reg/P0001 ,
		_w9060_
	);
	LUT2 #(
		.INIT('h4)
	) name5013 (
		\memc_EXTC_E_reg/NET0131 ,
		\memc_Pwrite_E_reg/NET0131 ,
		_w9061_
	);
	LUT3 #(
		.INIT('h10)
	) name5014 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\memc_EXTC_E_reg/NET0131 ,
		\memc_Pwrite_E_reg/NET0131 ,
		_w9062_
	);
	LUT4 #(
		.INIT('h00ea)
	) name5015 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w9062_,
		_w9063_
	);
	LUT2 #(
		.INIT('h4)
	) name5016 (
		_w4104_,
		_w9063_,
		_w9064_
	);
	LUT2 #(
		.INIT('h2)
	) name5017 (
		_w5025_,
		_w9064_,
		_w9065_
	);
	LUT2 #(
		.INIT('h8)
	) name5018 (
		_w5041_,
		_w9064_,
		_w9066_
	);
	LUT3 #(
		.INIT('h23)
	) name5019 (
		_w4104_,
		_w4966_,
		_w9063_,
		_w9067_
	);
	LUT3 #(
		.INIT('h07)
	) name5020 (
		_w5041_,
		_w9064_,
		_w9067_,
		_w9068_
	);
	LUT4 #(
		.INIT('h30a0)
	) name5021 (
		_w4966_,
		_w5041_,
		_w5327_,
		_w9064_,
		_w9069_
	);
	LUT2 #(
		.INIT('h4)
	) name5022 (
		_w9065_,
		_w9069_,
		_w9070_
	);
	LUT3 #(
		.INIT('h80)
	) name5023 (
		_w5041_,
		_w5549_,
		_w9064_,
		_w9071_
	);
	LUT3 #(
		.INIT('h0d)
	) name5024 (
		_w5025_,
		_w9064_,
		_w9067_,
		_w9072_
	);
	LUT2 #(
		.INIT('h4)
	) name5025 (
		_w9071_,
		_w9072_,
		_w9073_
	);
	LUT4 #(
		.INIT('hbf00)
	) name5026 (
		_w5439_,
		_w5529_,
		_w9068_,
		_w9073_,
		_w9074_
	);
	LUT2 #(
		.INIT('h2)
	) name5027 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		\bdma_CMcnt_reg[1]/NET0131 ,
		_w9075_
	);
	LUT2 #(
		.INIT('h8)
	) name5028 (
		_w4884_,
		_w9075_,
		_w9076_
	);
	LUT3 #(
		.INIT('h80)
	) name5029 (
		_w4885_,
		_w4884_,
		_w9075_,
		_w9077_
	);
	LUT4 #(
		.INIT('h4000)
	) name5030 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w4885_,
		_w4884_,
		_w9075_,
		_w9078_
	);
	LUT2 #(
		.INIT('h1)
	) name5031 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		\bdma_CMcnt_reg[1]/NET0131 ,
		_w9079_
	);
	LUT2 #(
		.INIT('h8)
	) name5032 (
		_w4884_,
		_w9079_,
		_w9080_
	);
	LUT3 #(
		.INIT('h80)
	) name5033 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w4884_,
		_w9079_,
		_w9081_
	);
	LUT4 #(
		.INIT('h8000)
	) name5034 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w4885_,
		_w4884_,
		_w9079_,
		_w9082_
	);
	LUT2 #(
		.INIT('h1)
	) name5035 (
		_w9078_,
		_w9082_,
		_w9083_
	);
	LUT2 #(
		.INIT('h2)
	) name5036 (
		_w5530_,
		_w9083_,
		_w9084_
	);
	LUT4 #(
		.INIT('hea00)
	) name5037 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w9061_,
		_w9085_
	);
	LUT4 #(
		.INIT('ha222)
	) name5038 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9086_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5039 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9087_
	);
	LUT2 #(
		.INIT('h1)
	) name5040 (
		_w5576_,
		_w9087_,
		_w9088_
	);
	LUT3 #(
		.INIT('h45)
	) name5041 (
		_w9084_,
		_w9086_,
		_w9088_,
		_w9089_
	);
	LUT3 #(
		.INIT('h08)
	) name5042 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9090_
	);
	LUT4 #(
		.INIT('h00c5)
	) name5043 (
		_w4966_,
		_w5041_,
		_w9064_,
		_w9090_,
		_w9091_
	);
	LUT4 #(
		.INIT('h30a0)
	) name5044 (
		_w4966_,
		_w5041_,
		_w5544_,
		_w9064_,
		_w9092_
	);
	LUT4 #(
		.INIT('h0045)
	) name5045 (
		_w9072_,
		_w9089_,
		_w9091_,
		_w9092_,
		_w9093_
	);
	LUT2 #(
		.INIT('h8)
	) name5046 (
		_w5914_,
		_w9070_,
		_w9094_
	);
	LUT4 #(
		.INIT('hff54)
	) name5047 (
		_w9070_,
		_w9074_,
		_w9093_,
		_w9094_,
		_w9095_
	);
	LUT3 #(
		.INIT('h80)
	) name5048 (
		_w5041_,
		_w6181_,
		_w9064_,
		_w9096_
	);
	LUT2 #(
		.INIT('h2)
	) name5049 (
		_w9072_,
		_w9096_,
		_w9097_
	);
	LUT4 #(
		.INIT('hef00)
	) name5050 (
		_w6209_,
		_w6215_,
		_w9068_,
		_w9097_,
		_w9098_
	);
	LUT4 #(
		.INIT('ha222)
	) name5051 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9099_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5052 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9100_
	);
	LUT2 #(
		.INIT('h1)
	) name5053 (
		_w6222_,
		_w9100_,
		_w9101_
	);
	LUT3 #(
		.INIT('h45)
	) name5054 (
		_w9084_,
		_w9099_,
		_w9101_,
		_w9102_
	);
	LUT3 #(
		.INIT('h08)
	) name5055 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9103_
	);
	LUT4 #(
		.INIT('h00c5)
	) name5056 (
		_w4966_,
		_w5041_,
		_w9064_,
		_w9103_,
		_w9104_
	);
	LUT4 #(
		.INIT('h30a0)
	) name5057 (
		_w4966_,
		_w5041_,
		_w6186_,
		_w9064_,
		_w9105_
	);
	LUT4 #(
		.INIT('h0045)
	) name5058 (
		_w9072_,
		_w9102_,
		_w9104_,
		_w9105_,
		_w9106_
	);
	LUT4 #(
		.INIT('h0100)
	) name5059 (
		_w5937_,
		_w6038_,
		_w9065_,
		_w9069_,
		_w9107_
	);
	LUT4 #(
		.INIT('hff54)
	) name5060 (
		_w9070_,
		_w9098_,
		_w9106_,
		_w9107_,
		_w9108_
	);
	LUT3 #(
		.INIT('h80)
	) name5061 (
		_w5041_,
		_w6506_,
		_w9064_,
		_w9109_
	);
	LUT2 #(
		.INIT('h2)
	) name5062 (
		_w9072_,
		_w9109_,
		_w9110_
	);
	LUT4 #(
		.INIT('hbf00)
	) name5063 (
		_w6529_,
		_w6533_,
		_w9068_,
		_w9110_,
		_w9111_
	);
	LUT4 #(
		.INIT('ha222)
	) name5064 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9112_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5065 (
		\idma_DCTL_reg[11]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9113_
	);
	LUT2 #(
		.INIT('h1)
	) name5066 (
		_w6538_,
		_w9113_,
		_w9114_
	);
	LUT3 #(
		.INIT('h45)
	) name5067 (
		_w9084_,
		_w9112_,
		_w9114_,
		_w9115_
	);
	LUT3 #(
		.INIT('h08)
	) name5068 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9116_
	);
	LUT4 #(
		.INIT('h00c5)
	) name5069 (
		_w4966_,
		_w5041_,
		_w9064_,
		_w9116_,
		_w9117_
	);
	LUT4 #(
		.INIT('h30a0)
	) name5070 (
		_w4966_,
		_w5041_,
		_w6511_,
		_w9064_,
		_w9118_
	);
	LUT4 #(
		.INIT('h0045)
	) name5071 (
		_w9072_,
		_w9115_,
		_w9117_,
		_w9118_,
		_w9119_
	);
	LUT4 #(
		.INIT('h0100)
	) name5072 (
		_w6263_,
		_w6362_,
		_w9065_,
		_w9069_,
		_w9120_
	);
	LUT4 #(
		.INIT('hff54)
	) name5073 (
		_w9070_,
		_w9111_,
		_w9119_,
		_w9120_,
		_w9121_
	);
	LUT3 #(
		.INIT('h80)
	) name5074 (
		_w5041_,
		_w6955_,
		_w9064_,
		_w9122_
	);
	LUT2 #(
		.INIT('h2)
	) name5075 (
		_w9072_,
		_w9122_,
		_w9123_
	);
	LUT4 #(
		.INIT('hbf00)
	) name5076 (
		_w6965_,
		_w6970_,
		_w9068_,
		_w9123_,
		_w9124_
	);
	LUT4 #(
		.INIT('ha222)
	) name5077 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9125_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5078 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9126_
	);
	LUT2 #(
		.INIT('h1)
	) name5079 (
		_w6976_,
		_w9126_,
		_w9127_
	);
	LUT3 #(
		.INIT('h45)
	) name5080 (
		_w9084_,
		_w9125_,
		_w9127_,
		_w9128_
	);
	LUT3 #(
		.INIT('h08)
	) name5081 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9129_
	);
	LUT4 #(
		.INIT('h00c5)
	) name5082 (
		_w4966_,
		_w5041_,
		_w9064_,
		_w9129_,
		_w9130_
	);
	LUT4 #(
		.INIT('h30a0)
	) name5083 (
		_w4966_,
		_w5041_,
		_w6950_,
		_w9064_,
		_w9131_
	);
	LUT4 #(
		.INIT('h0045)
	) name5084 (
		_w9072_,
		_w9128_,
		_w9130_,
		_w9131_,
		_w9132_
	);
	LUT2 #(
		.INIT('h8)
	) name5085 (
		_w6897_,
		_w9070_,
		_w9133_
	);
	LUT4 #(
		.INIT('hff54)
	) name5086 (
		_w9070_,
		_w9124_,
		_w9132_,
		_w9133_,
		_w9134_
	);
	LUT3 #(
		.INIT('h80)
	) name5087 (
		_w5041_,
		_w6996_,
		_w9064_,
		_w9135_
	);
	LUT2 #(
		.INIT('h2)
	) name5088 (
		_w9072_,
		_w9135_,
		_w9136_
	);
	LUT4 #(
		.INIT('hbf00)
	) name5089 (
		_w7004_,
		_w7008_,
		_w9068_,
		_w9136_,
		_w9137_
	);
	LUT4 #(
		.INIT('ha222)
	) name5090 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9138_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5091 (
		\idma_DCTL_reg[2]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9139_
	);
	LUT2 #(
		.INIT('h1)
	) name5092 (
		_w7014_,
		_w9139_,
		_w9140_
	);
	LUT3 #(
		.INIT('h45)
	) name5093 (
		_w9084_,
		_w9138_,
		_w9140_,
		_w9141_
	);
	LUT3 #(
		.INIT('h08)
	) name5094 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9142_
	);
	LUT4 #(
		.INIT('h00c5)
	) name5095 (
		_w4966_,
		_w5041_,
		_w9064_,
		_w9142_,
		_w9143_
	);
	LUT4 #(
		.INIT('h30a0)
	) name5096 (
		_w4966_,
		_w5041_,
		_w6991_,
		_w9064_,
		_w9144_
	);
	LUT4 #(
		.INIT('h0045)
	) name5097 (
		_w9072_,
		_w9141_,
		_w9143_,
		_w9144_,
		_w9145_
	);
	LUT2 #(
		.INIT('h8)
	) name5098 (
		_w6501_,
		_w9070_,
		_w9146_
	);
	LUT4 #(
		.INIT('hff54)
	) name5099 (
		_w9070_,
		_w9137_,
		_w9145_,
		_w9146_,
		_w9147_
	);
	LUT4 #(
		.INIT('ha222)
	) name5100 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9148_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5101 (
		\idma_DCTL_reg[3]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9149_
	);
	LUT2 #(
		.INIT('h1)
	) name5102 (
		_w7054_,
		_w9149_,
		_w9150_
	);
	LUT3 #(
		.INIT('h45)
	) name5103 (
		_w9084_,
		_w9148_,
		_w9150_,
		_w9151_
	);
	LUT3 #(
		.INIT('h08)
	) name5104 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9152_
	);
	LUT2 #(
		.INIT('h2)
	) name5105 (
		_w9067_,
		_w9152_,
		_w9153_
	);
	LUT2 #(
		.INIT('h4)
	) name5106 (
		_w9151_,
		_w9153_,
		_w9154_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5107 (
		_w5327_,
		_w6054_,
		_w6173_,
		_w6175_,
		_w9155_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5108 (
		_w5327_,
		_w7044_,
		_w7048_,
		_w9155_,
		_w9156_
	);
	LUT4 #(
		.INIT('h0704)
	) name5109 (
		_w7029_,
		_w9065_,
		_w9066_,
		_w9156_,
		_w9157_
	);
	LUT4 #(
		.INIT('h00df)
	) name5110 (
		_w5041_,
		_w7034_,
		_w9064_,
		_w9067_,
		_w9158_
	);
	LUT3 #(
		.INIT('h45)
	) name5111 (
		_w9154_,
		_w9157_,
		_w9158_,
		_w9159_
	);
	LUT4 #(
		.INIT('h0010)
	) name5112 (
		_w5327_,
		_w7083_,
		_w7086_,
		_w9065_,
		_w9160_
	);
	LUT4 #(
		.INIT('h335f)
	) name5113 (
		_w5025_,
		_w5041_,
		_w7091_,
		_w9064_,
		_w9161_
	);
	LUT4 #(
		.INIT('h00df)
	) name5114 (
		_w5041_,
		_w7096_,
		_w9064_,
		_w9067_,
		_w9162_
	);
	LUT4 #(
		.INIT('ha222)
	) name5115 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9163_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5116 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9164_
	);
	LUT2 #(
		.INIT('h1)
	) name5117 (
		_w7114_,
		_w9164_,
		_w9165_
	);
	LUT3 #(
		.INIT('h45)
	) name5118 (
		_w9084_,
		_w9163_,
		_w9165_,
		_w9166_
	);
	LUT3 #(
		.INIT('h08)
	) name5119 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9167_
	);
	LUT2 #(
		.INIT('h2)
	) name5120 (
		_w9067_,
		_w9167_,
		_w9168_
	);
	LUT2 #(
		.INIT('h4)
	) name5121 (
		_w9166_,
		_w9168_,
		_w9169_
	);
	LUT3 #(
		.INIT('h0b)
	) name5122 (
		_w7378_,
		_w9070_,
		_w9169_,
		_w9170_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5123 (
		_w9160_,
		_w9161_,
		_w9162_,
		_w9170_,
		_w9171_
	);
	LUT4 #(
		.INIT('h0010)
	) name5124 (
		_w5327_,
		_w7386_,
		_w7390_,
		_w9065_,
		_w9172_
	);
	LUT4 #(
		.INIT('h335f)
	) name5125 (
		_w5025_,
		_w5041_,
		_w7424_,
		_w9064_,
		_w9173_
	);
	LUT4 #(
		.INIT('h00df)
	) name5126 (
		_w5041_,
		_w7419_,
		_w9064_,
		_w9067_,
		_w9174_
	);
	LUT4 #(
		.INIT('ha222)
	) name5127 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9175_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5128 (
		\idma_DCTL_reg[5]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9176_
	);
	LUT2 #(
		.INIT('h1)
	) name5129 (
		_w7431_,
		_w9176_,
		_w9177_
	);
	LUT3 #(
		.INIT('h45)
	) name5130 (
		_w9084_,
		_w9175_,
		_w9177_,
		_w9178_
	);
	LUT3 #(
		.INIT('h08)
	) name5131 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9179_
	);
	LUT2 #(
		.INIT('h2)
	) name5132 (
		_w9067_,
		_w9179_,
		_w9180_
	);
	LUT2 #(
		.INIT('h4)
	) name5133 (
		_w9178_,
		_w9180_,
		_w9181_
	);
	LUT3 #(
		.INIT('h0b)
	) name5134 (
		_w7710_,
		_w9070_,
		_w9181_,
		_w9182_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5135 (
		_w9172_,
		_w9173_,
		_w9174_,
		_w9182_,
		_w9183_
	);
	LUT4 #(
		.INIT('h0001)
	) name5136 (
		_w5327_,
		_w7715_,
		_w7720_,
		_w9065_,
		_w9184_
	);
	LUT4 #(
		.INIT('h335f)
	) name5137 (
		_w5025_,
		_w5041_,
		_w7753_,
		_w9064_,
		_w9185_
	);
	LUT4 #(
		.INIT('h00df)
	) name5138 (
		_w5041_,
		_w7748_,
		_w9064_,
		_w9067_,
		_w9186_
	);
	LUT4 #(
		.INIT('ha222)
	) name5139 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9187_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5140 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9188_
	);
	LUT2 #(
		.INIT('h1)
	) name5141 (
		_w7760_,
		_w9188_,
		_w9189_
	);
	LUT3 #(
		.INIT('h45)
	) name5142 (
		_w9084_,
		_w9187_,
		_w9189_,
		_w9190_
	);
	LUT3 #(
		.INIT('h08)
	) name5143 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9191_
	);
	LUT2 #(
		.INIT('h2)
	) name5144 (
		_w9067_,
		_w9191_,
		_w9192_
	);
	LUT2 #(
		.INIT('h4)
	) name5145 (
		_w9190_,
		_w9192_,
		_w9193_
	);
	LUT3 #(
		.INIT('h0b)
	) name5146 (
		_w8043_,
		_w9070_,
		_w9193_,
		_w9194_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5147 (
		_w9184_,
		_w9185_,
		_w9186_,
		_w9194_,
		_w9195_
	);
	LUT4 #(
		.INIT('h0010)
	) name5148 (
		_w5327_,
		_w8052_,
		_w8055_,
		_w9065_,
		_w9196_
	);
	LUT4 #(
		.INIT('h335f)
	) name5149 (
		_w5025_,
		_w5041_,
		_w8066_,
		_w9064_,
		_w9197_
	);
	LUT4 #(
		.INIT('h00df)
	) name5150 (
		_w5041_,
		_w8061_,
		_w9064_,
		_w9067_,
		_w9198_
	);
	LUT4 #(
		.INIT('ha222)
	) name5151 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9199_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5152 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9200_
	);
	LUT2 #(
		.INIT('h1)
	) name5153 (
		_w8072_,
		_w9200_,
		_w9201_
	);
	LUT3 #(
		.INIT('h45)
	) name5154 (
		_w9084_,
		_w9199_,
		_w9201_,
		_w9202_
	);
	LUT3 #(
		.INIT('h08)
	) name5155 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9203_
	);
	LUT2 #(
		.INIT('h2)
	) name5156 (
		_w9067_,
		_w9203_,
		_w9204_
	);
	LUT2 #(
		.INIT('h4)
	) name5157 (
		_w9202_,
		_w9204_,
		_w9205_
	);
	LUT3 #(
		.INIT('h0b)
	) name5158 (
		_w7906_,
		_w9070_,
		_w9205_,
		_w9206_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5159 (
		_w9196_,
		_w9197_,
		_w9198_,
		_w9206_,
		_w9207_
	);
	LUT4 #(
		.INIT('h0010)
	) name5160 (
		_w5327_,
		_w8118_,
		_w8121_,
		_w9065_,
		_w9208_
	);
	LUT4 #(
		.INIT('h335f)
	) name5161 (
		_w5025_,
		_w5041_,
		_w8098_,
		_w9064_,
		_w9209_
	);
	LUT4 #(
		.INIT('h00df)
	) name5162 (
		_w5041_,
		_w8093_,
		_w9064_,
		_w9067_,
		_w9210_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5163 (
		_w7465_,
		_w7565_,
		_w9065_,
		_w9069_,
		_w9211_
	);
	LUT4 #(
		.INIT('ha222)
	) name5164 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9212_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5165 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9213_
	);
	LUT2 #(
		.INIT('h1)
	) name5166 (
		_w8105_,
		_w9213_,
		_w9214_
	);
	LUT3 #(
		.INIT('h45)
	) name5167 (
		_w9084_,
		_w9212_,
		_w9214_,
		_w9215_
	);
	LUT3 #(
		.INIT('h08)
	) name5168 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9216_
	);
	LUT2 #(
		.INIT('h2)
	) name5169 (
		_w9067_,
		_w9216_,
		_w9217_
	);
	LUT2 #(
		.INIT('h4)
	) name5170 (
		_w9215_,
		_w9217_,
		_w9218_
	);
	LUT2 #(
		.INIT('h1)
	) name5171 (
		_w9211_,
		_w9218_,
		_w9219_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5172 (
		_w9208_,
		_w9209_,
		_w9210_,
		_w9219_,
		_w9220_
	);
	LUT4 #(
		.INIT('h0010)
	) name5173 (
		_w5327_,
		_w8157_,
		_w8162_,
		_w9065_,
		_w9221_
	);
	LUT4 #(
		.INIT('h335f)
	) name5174 (
		_w5025_,
		_w5041_,
		_w8137_,
		_w9064_,
		_w9222_
	);
	LUT4 #(
		.INIT('h00df)
	) name5175 (
		_w5041_,
		_w8132_,
		_w9064_,
		_w9067_,
		_w9223_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5176 (
		_w7140_,
		_w7240_,
		_w9065_,
		_w9069_,
		_w9224_
	);
	LUT4 #(
		.INIT('ha222)
	) name5177 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9225_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5178 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9226_
	);
	LUT2 #(
		.INIT('h1)
	) name5179 (
		_w8146_,
		_w9226_,
		_w9227_
	);
	LUT3 #(
		.INIT('h45)
	) name5180 (
		_w9084_,
		_w9225_,
		_w9227_,
		_w9228_
	);
	LUT3 #(
		.INIT('h08)
	) name5181 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9229_
	);
	LUT2 #(
		.INIT('h2)
	) name5182 (
		_w9067_,
		_w9229_,
		_w9230_
	);
	LUT2 #(
		.INIT('h4)
	) name5183 (
		_w9228_,
		_w9230_,
		_w9231_
	);
	LUT2 #(
		.INIT('h1)
	) name5184 (
		_w9224_,
		_w9231_,
		_w9232_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5185 (
		_w9221_,
		_w9222_,
		_w9223_,
		_w9232_,
		_w9233_
	);
	LUT2 #(
		.INIT('h8)
	) name5186 (
		_w4936_,
		_w4937_,
		_w9234_
	);
	LUT2 #(
		.INIT('h8)
	) name5187 (
		_w8191_,
		_w9234_,
		_w9235_
	);
	LUT4 #(
		.INIT('h0001)
	) name5188 (
		_w5785_,
		_w8608_,
		_w8610_,
		_w8606_,
		_w9236_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5189 (
		\bdma_BRdataBUF_reg[8]/P0001 ,
		_w5530_,
		_w9078_,
		_w9236_,
		_w9237_
	);
	LUT3 #(
		.INIT('hb8)
	) name5190 (
		\idma_DTMP_H_reg[0]/P0001 ,
		_w9235_,
		_w9237_,
		_w9238_
	);
	LUT4 #(
		.INIT('h0001)
	) name5191 (
		_w5938_,
		_w8655_,
		_w8656_,
		_w8654_,
		_w9239_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5192 (
		\bdma_BRdataBUF_reg[18]/P0001 ,
		_w5530_,
		_w9078_,
		_w9239_,
		_w9240_
	);
	LUT3 #(
		.INIT('hb8)
	) name5193 (
		\idma_DTMP_H_reg[10]/P0001 ,
		_w9235_,
		_w9240_,
		_w9241_
	);
	LUT4 #(
		.INIT('h0001)
	) name5194 (
		_w6264_,
		_w8678_,
		_w8679_,
		_w8677_,
		_w9242_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5195 (
		\bdma_BRdataBUF_reg[19]/P0001 ,
		_w5530_,
		_w9078_,
		_w9242_,
		_w9243_
	);
	LUT3 #(
		.INIT('hb8)
	) name5196 (
		\idma_DTMP_H_reg[11]/P0001 ,
		_w9235_,
		_w9243_,
		_w9244_
	);
	LUT4 #(
		.INIT('h0001)
	) name5197 (
		_w6660_,
		_w8702_,
		_w8703_,
		_w8701_,
		_w9245_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5198 (
		\bdma_BRdataBUF_reg[20]/P0001 ,
		_w5530_,
		_w9078_,
		_w9245_,
		_w9246_
	);
	LUT3 #(
		.INIT('hb8)
	) name5199 (
		\idma_DTMP_H_reg[12]/P0001 ,
		_w9235_,
		_w9246_,
		_w9247_
	);
	LUT4 #(
		.INIT('h0001)
	) name5200 (
		_w5626_,
		_w8725_,
		_w8726_,
		_w8724_,
		_w9248_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5201 (
		\bdma_BRdataBUF_reg[21]/P0001 ,
		_w5530_,
		_w9078_,
		_w9248_,
		_w9249_
	);
	LUT3 #(
		.INIT('hb8)
	) name5202 (
		\idma_DTMP_H_reg[13]/P0001 ,
		_w9235_,
		_w9249_,
		_w9250_
	);
	LUT4 #(
		.INIT('h0001)
	) name5203 (
		_w8237_,
		_w8765_,
		_w8766_,
		_w8764_,
		_w9251_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5204 (
		\bdma_BRdataBUF_reg[22]/P0001 ,
		_w5530_,
		_w9078_,
		_w9251_,
		_w9252_
	);
	LUT3 #(
		.INIT('hb8)
	) name5205 (
		\idma_DTMP_H_reg[14]/P0001 ,
		_w9235_,
		_w9252_,
		_w9253_
	);
	LUT4 #(
		.INIT('h0001)
	) name5206 (
		_w8318_,
		_w8805_,
		_w8806_,
		_w8804_,
		_w9254_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5207 (
		\bdma_BRdataBUF_reg[23]/P0001 ,
		_w5530_,
		_w9078_,
		_w9254_,
		_w9255_
	);
	LUT3 #(
		.INIT('hb8)
	) name5208 (
		\idma_DTMP_H_reg[15]/P0001 ,
		_w9235_,
		_w9255_,
		_w9256_
	);
	LUT4 #(
		.INIT('h0001)
	) name5209 (
		_w6775_,
		_w8826_,
		_w8827_,
		_w8825_,
		_w9257_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5210 (
		\bdma_BRdataBUF_reg[9]/P0001 ,
		_w5530_,
		_w9078_,
		_w9257_,
		_w9258_
	);
	LUT3 #(
		.INIT('hb8)
	) name5211 (
		\idma_DTMP_H_reg[1]/P0001 ,
		_w9235_,
		_w9258_,
		_w9259_
	);
	LUT4 #(
		.INIT('h0001)
	) name5212 (
		_w6379_,
		_w8848_,
		_w8849_,
		_w8847_,
		_w9260_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5213 (
		\bdma_BRdataBUF_reg[10]/P0001 ,
		_w5530_,
		_w9078_,
		_w9260_,
		_w9261_
	);
	LUT3 #(
		.INIT('hb8)
	) name5214 (
		\idma_DTMP_H_reg[2]/P0001 ,
		_w9235_,
		_w9261_,
		_w9262_
	);
	LUT4 #(
		.INIT('h0001)
	) name5215 (
		_w6055_,
		_w8870_,
		_w8871_,
		_w8869_,
		_w9263_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5216 (
		\bdma_BRdataBUF_reg[11]/P0001 ,
		_w5530_,
		_w9078_,
		_w9263_,
		_w9264_
	);
	LUT3 #(
		.INIT('hb8)
	) name5217 (
		\idma_DTMP_H_reg[3]/P0001 ,
		_w9235_,
		_w9264_,
		_w9265_
	);
	LUT4 #(
		.INIT('h0001)
	) name5218 (
		_w7258_,
		_w8892_,
		_w8893_,
		_w8891_,
		_w9266_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5219 (
		\bdma_BRdataBUF_reg[12]/P0001 ,
		_w5530_,
		_w9078_,
		_w9266_,
		_w9267_
	);
	LUT3 #(
		.INIT('hb8)
	) name5220 (
		\idma_DTMP_H_reg[4]/P0001 ,
		_w9235_,
		_w9267_,
		_w9268_
	);
	LUT4 #(
		.INIT('h0001)
	) name5221 (
		_w7593_,
		_w8914_,
		_w8915_,
		_w8913_,
		_w9269_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5222 (
		\bdma_BRdataBUF_reg[13]/P0001 ,
		_w5530_,
		_w9078_,
		_w9269_,
		_w9270_
	);
	LUT3 #(
		.INIT('hb8)
	) name5223 (
		\idma_DTMP_H_reg[5]/P0001 ,
		_w9235_,
		_w9270_,
		_w9271_
	);
	LUT4 #(
		.INIT('h1030)
	) name5224 (
		_w5530_,
		_w7928_,
		_w8949_,
		_w9078_,
		_w9272_
	);
	LUT3 #(
		.INIT('h40)
	) name5225 (
		\bdma_BRdataBUF_reg[14]/P0001 ,
		_w5530_,
		_w9078_,
		_w9273_
	);
	LUT4 #(
		.INIT('h888b)
	) name5226 (
		\idma_DTMP_H_reg[6]/P0001 ,
		_w9235_,
		_w9272_,
		_w9273_,
		_w9274_
	);
	LUT4 #(
		.INIT('h0001)
	) name5227 (
		_w7794_,
		_w8959_,
		_w8960_,
		_w8958_,
		_w9275_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5228 (
		\bdma_BRdataBUF_reg[15]/P0001 ,
		_w5530_,
		_w9078_,
		_w9275_,
		_w9276_
	);
	LUT3 #(
		.INIT('hb8)
	) name5229 (
		\idma_DTMP_H_reg[7]/P0001 ,
		_w9235_,
		_w9276_,
		_w9277_
	);
	LUT4 #(
		.INIT('h0001)
	) name5230 (
		_w7466_,
		_w8982_,
		_w8983_,
		_w8981_,
		_w9278_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5231 (
		\bdma_BRdataBUF_reg[16]/P0001 ,
		_w5530_,
		_w9078_,
		_w9278_,
		_w9279_
	);
	LUT3 #(
		.INIT('hb8)
	) name5232 (
		\idma_DTMP_H_reg[8]/P0001 ,
		_w9235_,
		_w9279_,
		_w9280_
	);
	LUT4 #(
		.INIT('h0001)
	) name5233 (
		_w7141_,
		_w9005_,
		_w9006_,
		_w9004_,
		_w9281_
	);
	LUT4 #(
		.INIT('h80bf)
	) name5234 (
		\bdma_BRdataBUF_reg[17]/P0001 ,
		_w5530_,
		_w9078_,
		_w9281_,
		_w9282_
	);
	LUT3 #(
		.INIT('hb8)
	) name5235 (
		\idma_DTMP_H_reg[9]/P0001 ,
		_w9235_,
		_w9282_,
		_w9283_
	);
	LUT4 #(
		.INIT('hc050)
	) name5236 (
		_w4966_,
		_w5041_,
		_w6608_,
		_w9064_,
		_w9284_
	);
	LUT3 #(
		.INIT('h04)
	) name5237 (
		_w9069_,
		_w9072_,
		_w9284_,
		_w9285_
	);
	LUT4 #(
		.INIT('hbf00)
	) name5238 (
		_w6576_,
		_w6580_,
		_w9068_,
		_w9285_,
		_w9286_
	);
	LUT3 #(
		.INIT('h20)
	) name5239 (
		_w6758_,
		_w9065_,
		_w9069_,
		_w9287_
	);
	LUT4 #(
		.INIT('h0008)
	) name5240 (
		_w4966_,
		_w5025_,
		_w6613_,
		_w9064_,
		_w9288_
	);
	LUT4 #(
		.INIT('ha222)
	) name5241 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9289_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5242 (
		\idma_DCTL_reg[12]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9290_
	);
	LUT4 #(
		.INIT('h0031)
	) name5243 (
		_w5530_,
		_w6620_,
		_w9083_,
		_w9290_,
		_w9291_
	);
	LUT3 #(
		.INIT('h04)
	) name5244 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9292_
	);
	LUT4 #(
		.INIT('h2022)
	) name5245 (
		_w9067_,
		_w9292_,
		_w9289_,
		_w9291_,
		_w9293_
	);
	LUT2 #(
		.INIT('h1)
	) name5246 (
		_w9288_,
		_w9293_,
		_w9294_
	);
	LUT2 #(
		.INIT('h4)
	) name5247 (
		_w9287_,
		_w9294_,
		_w9295_
	);
	LUT2 #(
		.INIT('hb)
	) name5248 (
		_w9286_,
		_w9295_,
		_w9296_
	);
	LUT3 #(
		.INIT('h10)
	) name5249 (
		PM_bdry_sel_pad,
		_w9286_,
		_w9295_,
		_w9297_
	);
	LUT4 #(
		.INIT('h0100)
	) name5250 (
		_w6909_,
		_w6910_,
		_w6911_,
		_w9068_,
		_w9298_
	);
	LUT4 #(
		.INIT('hc050)
	) name5251 (
		_w4966_,
		_w5041_,
		_w6918_,
		_w9064_,
		_w9299_
	);
	LUT3 #(
		.INIT('h04)
	) name5252 (
		_w9069_,
		_w9072_,
		_w9299_,
		_w9300_
	);
	LUT3 #(
		.INIT('h20)
	) name5253 (
		_w5760_,
		_w9065_,
		_w9069_,
		_w9301_
	);
	LUT4 #(
		.INIT('h0008)
	) name5254 (
		_w4966_,
		_w5025_,
		_w6923_,
		_w9064_,
		_w9302_
	);
	LUT4 #(
		.INIT('ha222)
	) name5255 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		_w5569_,
		_w5570_,
		_w9085_,
		_w9303_
	);
	LUT4 #(
		.INIT('h2a00)
	) name5256 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w4067_,
		_w4845_,
		_w4936_,
		_w9304_
	);
	LUT4 #(
		.INIT('h0031)
	) name5257 (
		_w5530_,
		_w6929_,
		_w9083_,
		_w9304_,
		_w9305_
	);
	LUT3 #(
		.INIT('h04)
	) name5258 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w5530_,
		_w9083_,
		_w9306_
	);
	LUT4 #(
		.INIT('h2022)
	) name5259 (
		_w9067_,
		_w9306_,
		_w9303_,
		_w9305_,
		_w9307_
	);
	LUT2 #(
		.INIT('h1)
	) name5260 (
		_w9302_,
		_w9307_,
		_w9308_
	);
	LUT2 #(
		.INIT('h4)
	) name5261 (
		_w9301_,
		_w9308_,
		_w9309_
	);
	LUT3 #(
		.INIT('hb0)
	) name5262 (
		_w9298_,
		_w9300_,
		_w9309_,
		_w9310_
	);
	LUT3 #(
		.INIT('h4f)
	) name5263 (
		_w9298_,
		_w9300_,
		_w9309_,
		_w9311_
	);
	LUT3 #(
		.INIT('h53)
	) name5264 (
		\bdma_BOVL_reg[9]/NET0131 ,
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		_w4519_,
		_w9312_
	);
	LUT3 #(
		.INIT('h74)
	) name5265 (
		\idma_DOVL_reg[9]/NET0131 ,
		_w4946_,
		_w9312_,
		_w9313_
	);
	LUT3 #(
		.INIT('h53)
	) name5266 (
		\bdma_BOVL_reg[11]/NET0131 ,
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w4519_,
		_w9314_
	);
	LUT3 #(
		.INIT('h74)
	) name5267 (
		\idma_DOVL_reg[11]/NET0131 ,
		_w4946_,
		_w9314_,
		_w9315_
	);
	LUT3 #(
		.INIT('h53)
	) name5268 (
		\bdma_BOVL_reg[10]/NET0131 ,
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		_w4519_,
		_w9316_
	);
	LUT3 #(
		.INIT('h74)
	) name5269 (
		\idma_DOVL_reg[10]/NET0131 ,
		_w4946_,
		_w9316_,
		_w9317_
	);
	LUT3 #(
		.INIT('h53)
	) name5270 (
		\bdma_BOVL_reg[8]/NET0131 ,
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		_w4519_,
		_w9318_
	);
	LUT3 #(
		.INIT('h74)
	) name5271 (
		\idma_DOVL_reg[8]/NET0131 ,
		_w4946_,
		_w9318_,
		_w9319_
	);
	LUT3 #(
		.INIT('h80)
	) name5272 (
		_w9315_,
		_w9317_,
		_w9319_,
		_w9320_
	);
	LUT4 #(
		.INIT('h1000)
	) name5273 (
		_w9297_,
		_w9310_,
		_w9313_,
		_w9320_,
		_w9321_
	);
	LUT4 #(
		.INIT('h4000)
	) name5274 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w5045_,
		_w5046_,
		_w9322_
	);
	LUT4 #(
		.INIT('h0010)
	) name5275 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w9323_
	);
	LUT3 #(
		.INIT('h23)
	) name5276 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w4967_,
		_w9323_,
		_w9324_
	);
	LUT2 #(
		.INIT('h4)
	) name5277 (
		_w9322_,
		_w9324_,
		_w9325_
	);
	LUT2 #(
		.INIT('h4)
	) name5278 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_RDcyc_reg/NET0131 ,
		_w9326_
	);
	LUT2 #(
		.INIT('h8)
	) name5279 (
		_w4937_,
		_w9326_,
		_w9327_
	);
	LUT4 #(
		.INIT('h135f)
	) name5280 (
		_w4519_,
		_w4520_,
		_w9082_,
		_w9327_,
		_w9328_
	);
	LUT4 #(
		.INIT('h00df)
	) name5281 (
		_w4067_,
		_w4068_,
		_w4845_,
		_w9328_,
		_w9329_
	);
	LUT4 #(
		.INIT('h2000)
	) name5282 (
		\memc_Pread_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w9330_
	);
	LUT2 #(
		.INIT('h1)
	) name5283 (
		_w9329_,
		_w9330_,
		_w9331_
	);
	LUT4 #(
		.INIT('hf700)
	) name5284 (
		_w8174_,
		_w9063_,
		_w9325_,
		_w9331_,
		_w9332_
	);
	LUT4 #(
		.INIT('h135f)
	) name5285 (
		_w5530_,
		_w8191_,
		_w9078_,
		_w9234_,
		_w9333_
	);
	LUT3 #(
		.INIT('h47)
	) name5286 (
		\memc_Pwrite_C_reg/NET0131 ,
		_w4971_,
		_w9085_,
		_w9334_
	);
	LUT2 #(
		.INIT('h8)
	) name5287 (
		_w9333_,
		_w9334_,
		_w9335_
	);
	LUT2 #(
		.INIT('h8)
	) name5288 (
		_w9332_,
		_w9335_,
		_w9336_
	);
	LUT2 #(
		.INIT('h2)
	) name5289 (
		_w9321_,
		_w9336_,
		_w9337_
	);
	LUT3 #(
		.INIT('h08)
	) name5290 (
		_w9315_,
		_w9317_,
		_w9319_,
		_w9338_
	);
	LUT4 #(
		.INIT('h1000)
	) name5291 (
		_w9297_,
		_w9310_,
		_w9313_,
		_w9338_,
		_w9339_
	);
	LUT2 #(
		.INIT('h4)
	) name5292 (
		_w9336_,
		_w9339_,
		_w9340_
	);
	LUT4 #(
		.INIT('h0100)
	) name5293 (
		_w9297_,
		_w9310_,
		_w9313_,
		_w9320_,
		_w9341_
	);
	LUT2 #(
		.INIT('h4)
	) name5294 (
		_w9336_,
		_w9341_,
		_w9342_
	);
	LUT4 #(
		.INIT('h0100)
	) name5295 (
		_w9297_,
		_w9310_,
		_w9313_,
		_w9338_,
		_w9343_
	);
	LUT2 #(
		.INIT('h4)
	) name5296 (
		_w9336_,
		_w9343_,
		_w9344_
	);
	LUT4 #(
		.INIT('h0010)
	) name5297 (
		_w9297_,
		_w9310_,
		_w9315_,
		_w9317_,
		_w9345_
	);
	LUT4 #(
		.INIT('h0800)
	) name5298 (
		_w9313_,
		_w9319_,
		_w9336_,
		_w9345_,
		_w9346_
	);
	LUT4 #(
		.INIT('h0200)
	) name5299 (
		_w9313_,
		_w9319_,
		_w9336_,
		_w9345_,
		_w9347_
	);
	LUT4 #(
		.INIT('h0400)
	) name5300 (
		_w9313_,
		_w9319_,
		_w9336_,
		_w9345_,
		_w9348_
	);
	LUT4 #(
		.INIT('h0100)
	) name5301 (
		_w9313_,
		_w9319_,
		_w9336_,
		_w9345_,
		_w9349_
	);
	LUT4 #(
		.INIT('h2a15)
	) name5302 (
		\sport0_cfg_FSi_reg/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w9350_
	);
	LUT4 #(
		.INIT('hd5ea)
	) name5303 (
		\sport0_cfg_FSi_reg/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w9351_
	);
	LUT4 #(
		.INIT('h2a15)
	) name5304 (
		\sport1_cfg_FSi_reg/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w9352_
	);
	LUT4 #(
		.INIT('hd5ea)
	) name5305 (
		\sport1_cfg_FSi_reg/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w9353_
	);
	LUT2 #(
		.INIT('h6)
	) name5306 (
		\sport0_cfg_SCLKi_h_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w9354_
	);
	LUT2 #(
		.INIT('h6)
	) name5307 (
		\sport1_cfg_SCLKi_h_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w9355_
	);
	LUT3 #(
		.INIT('h20)
	) name5308 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[2]/P0001 ,
		_w9356_
	);
	LUT4 #(
		.INIT('h5455)
	) name5309 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[0]/P0001 ,
		_w9357_
	);
	LUT3 #(
		.INIT('h20)
	) name5310 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[3]/P0001 ,
		_w9358_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5311 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[1]/P0001 ,
		_w9359_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5312 (
		_w9356_,
		_w9357_,
		_w9358_,
		_w9359_,
		_w9360_
	);
	LUT2 #(
		.INIT('h2)
	) name5313 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_txctl_TXSHT_reg[5]/P0001 ,
		_w9361_
	);
	LUT4 #(
		.INIT('h3020)
	) name5314 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[4]/P0001 ,
		_w9362_
	);
	LUT2 #(
		.INIT('h4)
	) name5315 (
		_w9361_,
		_w9362_,
		_w9363_
	);
	LUT2 #(
		.INIT('h2)
	) name5316 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_txctl_TXSHT_reg[7]/P0001 ,
		_w9364_
	);
	LUT4 #(
		.INIT('hc080)
	) name5317 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[6]/P0001 ,
		_w9365_
	);
	LUT3 #(
		.INIT('h45)
	) name5318 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w9364_,
		_w9365_,
		_w9366_
	);
	LUT3 #(
		.INIT('h10)
	) name5319 (
		_w9360_,
		_w9363_,
		_w9366_,
		_w9367_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5320 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[13]/P0001 ,
		_w9368_
	);
	LUT4 #(
		.INIT('hcedf)
	) name5321 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[11]/P0001 ,
		\sport0_txctl_TXSHT_reg[9]/P0001 ,
		_w9369_
	);
	LUT4 #(
		.INIT('h5455)
	) name5322 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[8]/P0001 ,
		_w9370_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name5323 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[10]/P0001 ,
		\sport0_txctl_TXSHT_reg[12]/P0001 ,
		_w9371_
	);
	LUT4 #(
		.INIT('h0777)
	) name5324 (
		_w9368_,
		_w9369_,
		_w9370_,
		_w9371_,
		_w9372_
	);
	LUT2 #(
		.INIT('h2)
	) name5325 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_txctl_TXSHT_reg[15]/P0001 ,
		_w9373_
	);
	LUT4 #(
		.INIT('hc080)
	) name5326 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_txctl_TXSHT_reg[14]/P0001 ,
		_w9374_
	);
	LUT3 #(
		.INIT('h8a)
	) name5327 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w9373_,
		_w9374_,
		_w9375_
	);
	LUT2 #(
		.INIT('h4)
	) name5328 (
		_w9372_,
		_w9375_,
		_w9376_
	);
	LUT4 #(
		.INIT('h888d)
	) name5329 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport0_txctl_TXSHT_reg[15]/P0001 ,
		_w9367_,
		_w9376_,
		_w9377_
	);
	LUT2 #(
		.INIT('h4)
	) name5330 (
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w9377_,
		_w9378_
	);
	LUT2 #(
		.INIT('h1)
	) name5331 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[2]/P0001 ,
		_w9379_
	);
	LUT4 #(
		.INIT('h0c04)
	) name5332 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_txctl_TXSHT_reg[3]/P0001 ,
		_w9380_
	);
	LUT3 #(
		.INIT('h45)
	) name5333 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w9379_,
		_w9380_,
		_w9381_
	);
	LUT2 #(
		.INIT('h2)
	) name5334 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[1]/P0001 ,
		_w9382_
	);
	LUT4 #(
		.INIT('h0302)
	) name5335 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_txctl_TXSHT_reg[0]/P0001 ,
		_w9383_
	);
	LUT2 #(
		.INIT('h4)
	) name5336 (
		_w9382_,
		_w9383_,
		_w9384_
	);
	LUT2 #(
		.INIT('h2)
	) name5337 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[7]/P0001 ,
		_w9385_
	);
	LUT4 #(
		.INIT('hc080)
	) name5338 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_txctl_TXSHT_reg[6]/P0001 ,
		_w9386_
	);
	LUT2 #(
		.INIT('h2)
	) name5339 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[5]/P0001 ,
		_w9387_
	);
	LUT4 #(
		.INIT('h3020)
	) name5340 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_txctl_TXSHT_reg[4]/P0001 ,
		_w9388_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5341 (
		_w9385_,
		_w9386_,
		_w9387_,
		_w9388_,
		_w9389_
	);
	LUT3 #(
		.INIT('h40)
	) name5342 (
		_w9384_,
		_w9381_,
		_w9389_,
		_w9390_
	);
	LUT2 #(
		.INIT('h2)
	) name5343 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[15]/P0001 ,
		_w9391_
	);
	LUT4 #(
		.INIT('hc080)
	) name5344 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_txctl_TXSHT_reg[14]/P0001 ,
		_w9392_
	);
	LUT3 #(
		.INIT('h8a)
	) name5345 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w9391_,
		_w9392_,
		_w9393_
	);
	LUT2 #(
		.INIT('h2)
	) name5346 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[13]/P0001 ,
		_w9394_
	);
	LUT4 #(
		.INIT('h3020)
	) name5347 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_txctl_TXSHT_reg[12]/P0001 ,
		_w9395_
	);
	LUT2 #(
		.INIT('h4)
	) name5348 (
		_w9394_,
		_w9395_,
		_w9396_
	);
	LUT2 #(
		.INIT('h2)
	) name5349 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[9]/P0001 ,
		_w9397_
	);
	LUT4 #(
		.INIT('h0302)
	) name5350 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_txctl_TXSHT_reg[8]/P0001 ,
		_w9398_
	);
	LUT2 #(
		.INIT('h2)
	) name5351 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[11]/P0001 ,
		_w9399_
	);
	LUT4 #(
		.INIT('h0c08)
	) name5352 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_txctl_TXSHT_reg[10]/P0001 ,
		_w9400_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5353 (
		_w9397_,
		_w9398_,
		_w9399_,
		_w9400_,
		_w9401_
	);
	LUT3 #(
		.INIT('h40)
	) name5354 (
		_w9396_,
		_w9393_,
		_w9401_,
		_w9402_
	);
	LUT4 #(
		.INIT('h888d)
	) name5355 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport1_txctl_TXSHT_reg[15]/P0001 ,
		_w9390_,
		_w9402_,
		_w9403_
	);
	LUT2 #(
		.INIT('h4)
	) name5356 (
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w9403_,
		_w9404_
	);
	LUT4 #(
		.INIT('h2a15)
	) name5357 (
		\sport0_cfg_FSi_reg/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w9405_
	);
	LUT4 #(
		.INIT('hd5ea)
	) name5358 (
		\sport0_cfg_FSi_reg/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w9406_
	);
	LUT4 #(
		.INIT('h2a15)
	) name5359 (
		\sport1_cfg_FSi_reg/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w9407_
	);
	LUT4 #(
		.INIT('hd5ea)
	) name5360 (
		\sport1_cfg_FSi_reg/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w9408_
	);
	LUT3 #(
		.INIT('hd8)
	) name5361 (
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWRn_reg/NET0131 ,
		\emc_WRn_h_reg/P0001 ,
		_w9409_
	);
	LUT3 #(
		.INIT('h10)
	) name5362 (
		T_BMODE_pad,
		T_MMAP_pad,
		\bdma_RST_pin_reg/P0001 ,
		_w9410_
	);
	LUT4 #(
		.INIT('hdbff)
	) name5363 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		\bdma_CMcnt_reg[1]/NET0131 ,
		_w4885_,
		_w4884_,
		_w9411_
	);
	LUT4 #(
		.INIT('h9fff)
	) name5364 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w9412_
	);
	LUT4 #(
		.INIT('h4000)
	) name5365 (
		_w4747_,
		_w4768_,
		_w4789_,
		_w4796_,
		_w9413_
	);
	LUT3 #(
		.INIT('h10)
	) name5366 (
		_w9411_,
		_w9412_,
		_w9413_,
		_w9414_
	);
	LUT4 #(
		.INIT('h0400)
	) name5367 (
		_w5532_,
		_w5531_,
		_w9412_,
		_w9413_,
		_w9415_
	);
	LUT2 #(
		.INIT('h1)
	) name5368 (
		\bdma_BWCOUNT_reg[3]/NET0131 ,
		\bdma_BWCOUNT_reg[4]/NET0131 ,
		_w9416_
	);
	LUT3 #(
		.INIT('h01)
	) name5369 (
		\bdma_BWCOUNT_reg[1]/NET0131 ,
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		\bdma_BWCOUNT_reg[6]/NET0131 ,
		_w9417_
	);
	LUT3 #(
		.INIT('h80)
	) name5370 (
		_w7610_,
		_w9416_,
		_w9417_,
		_w9418_
	);
	LUT3 #(
		.INIT('h01)
	) name5371 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		\bdma_BWCOUNT_reg[8]/NET0131 ,
		\bdma_BWCOUNT_reg[9]/NET0131 ,
		_w9419_
	);
	LUT4 #(
		.INIT('h0001)
	) name5372 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		\bdma_BWCOUNT_reg[11]/NET0131 ,
		\bdma_BWCOUNT_reg[12]/NET0131 ,
		\bdma_BWCOUNT_reg[13]/NET0131 ,
		_w9420_
	);
	LUT2 #(
		.INIT('h8)
	) name5373 (
		_w9419_,
		_w9420_,
		_w9421_
	);
	LUT2 #(
		.INIT('h8)
	) name5374 (
		_w9418_,
		_w9421_,
		_w9422_
	);
	LUT3 #(
		.INIT('h80)
	) name5375 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		_w9418_,
		_w9421_,
		_w9423_
	);
	LUT4 #(
		.INIT('h0155)
	) name5376 (
		_w4066_,
		_w9414_,
		_w9415_,
		_w9423_,
		_w9424_
	);
	LUT2 #(
		.INIT('he)
	) name5377 (
		_w9410_,
		_w9424_,
		_w9425_
	);
	LUT3 #(
		.INIT('h54)
	) name5378 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		_w9414_,
		_w9415_,
		_w9426_
	);
	LUT4 #(
		.INIT('h1110)
	) name5379 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		\bdma_BWCOUNT_reg[1]/NET0131 ,
		_w9414_,
		_w9415_,
		_w9427_
	);
	LUT3 #(
		.INIT('h40)
	) name5380 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		_w9416_,
		_w9427_,
		_w9428_
	);
	LUT4 #(
		.INIT('h4000)
	) name5381 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		_w7610_,
		_w9416_,
		_w9427_,
		_w9429_
	);
	LUT3 #(
		.INIT('h8a)
	) name5382 (
		\memc_Dwrite_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9430_
	);
	LUT4 #(
		.INIT('h4044)
	) name5383 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\memc_Dwrite_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9431_
	);
	LUT3 #(
		.INIT('h80)
	) name5384 (
		_w5657_,
		_w5658_,
		_w9431_,
		_w9432_
	);
	LUT4 #(
		.INIT('hba00)
	) name5385 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w9432_,
		_w9433_
	);
	LUT4 #(
		.INIT('h00ed)
	) name5386 (
		_w7610_,
		_w9432_,
		_w9428_,
		_w9433_,
		_w9434_
	);
	LUT2 #(
		.INIT('he)
	) name5387 (
		_w9410_,
		_w9434_,
		_w9435_
	);
	LUT2 #(
		.INIT('h8)
	) name5388 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w9436_
	);
	LUT3 #(
		.INIT('h08)
	) name5389 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w9437_
	);
	LUT2 #(
		.INIT('h8)
	) name5390 (
		\core_c_dec_MTCNTR_Eg_reg/P0001 ,
		\core_c_psq_CNTRval_reg/NET0131 ,
		_w9438_
	);
	LUT3 #(
		.INIT('hb0)
	) name5391 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9438_,
		_w9439_
	);
	LUT4 #(
		.INIT('h0b00)
	) name5392 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9437_,
		_w9438_,
		_w9440_
	);
	LUT4 #(
		.INIT('haccc)
	) name5393 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001 ,
		_w9436_,
		_w9440_,
		_w9441_
	);
	LUT2 #(
		.INIT('h1)
	) name5394 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w9442_
	);
	LUT4 #(
		.INIT('hb000)
	) name5395 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9438_,
		_w9442_,
		_w9443_
	);
	LUT3 #(
		.INIT('hac)
	) name5396 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001 ,
		_w9443_,
		_w9444_
	);
	LUT2 #(
		.INIT('h2)
	) name5397 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w9445_
	);
	LUT4 #(
		.INIT('hb000)
	) name5398 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9438_,
		_w9445_,
		_w9446_
	);
	LUT3 #(
		.INIT('hac)
	) name5399 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001 ,
		_w9446_,
		_w9447_
	);
	LUT2 #(
		.INIT('h4)
	) name5400 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w9448_
	);
	LUT4 #(
		.INIT('hb000)
	) name5401 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9438_,
		_w9448_,
		_w9449_
	);
	LUT3 #(
		.INIT('hac)
	) name5402 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001 ,
		_w9449_,
		_w9450_
	);
	LUT3 #(
		.INIT('h01)
	) name5403 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_c_dec_DIVS_E_reg/P0001 ,
		\core_c_dec_updAF_E_reg/P0001 ,
		_w9451_
	);
	LUT3 #(
		.INIT('h45)
	) name5404 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9452_
	);
	LUT4 #(
		.INIT('h0200)
	) name5405 (
		\core_c_dec_Usecond_E_reg/P0001 ,
		_w4160_,
		_w4158_,
		_w4167_,
		_w9453_
	);
	LUT4 #(
		.INIT('h0010)
	) name5406 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9451_,
		_w9452_,
		_w9453_,
		_w9454_
	);
	LUT3 #(
		.INIT('h0e)
	) name5407 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_c_dec_DIVS_E_reg/P0001 ,
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9455_
	);
	LUT4 #(
		.INIT('h7000)
	) name5408 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9456_
	);
	LUT3 #(
		.INIT('h80)
	) name5409 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9457_
	);
	LUT4 #(
		.INIT('h8000)
	) name5410 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9458_
	);
	LUT4 #(
		.INIT('h028a)
	) name5411 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001 ,
		_w9459_
	);
	LUT2 #(
		.INIT('h8)
	) name5412 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w9460_
	);
	LUT4 #(
		.INIT('h0145)
	) name5413 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001 ,
		_w9461_
	);
	LUT3 #(
		.INIT('h02)
	) name5414 (
		_w9460_,
		_w9461_,
		_w9459_,
		_w9462_
	);
	LUT3 #(
		.INIT('h08)
	) name5415 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w9463_
	);
	LUT3 #(
		.INIT('h10)
	) name5416 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w9464_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5417 (
		_w5713_,
		_w8349_,
		_w9463_,
		_w9464_,
		_w9465_
	);
	LUT3 #(
		.INIT('h40)
	) name5418 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w9466_
	);
	LUT3 #(
		.INIT('h02)
	) name5419 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w9467_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5420 (
		_w8375_,
		_w8371_,
		_w9466_,
		_w9467_,
		_w9468_
	);
	LUT4 #(
		.INIT('h028a)
	) name5421 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001 ,
		_w9469_
	);
	LUT2 #(
		.INIT('h1)
	) name5422 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w9470_
	);
	LUT4 #(
		.INIT('h0145)
	) name5423 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001 ,
		_w9471_
	);
	LUT3 #(
		.INIT('h02)
	) name5424 (
		_w9470_,
		_w9471_,
		_w9469_,
		_w9472_
	);
	LUT4 #(
		.INIT('h0040)
	) name5425 (
		_w9462_,
		_w9465_,
		_w9468_,
		_w9472_,
		_w9473_
	);
	LUT2 #(
		.INIT('h2)
	) name5426 (
		_w9458_,
		_w9473_,
		_w9474_
	);
	LUT3 #(
		.INIT('h01)
	) name5427 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w9475_
	);
	LUT4 #(
		.INIT('hfe32)
	) name5428 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_c_dec_DIVS_E_reg/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w9476_
	);
	LUT3 #(
		.INIT('h02)
	) name5429 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		_w9477_
	);
	LUT2 #(
		.INIT('h4)
	) name5430 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9478_
	);
	LUT3 #(
		.INIT('h8a)
	) name5431 (
		_w9476_,
		_w9477_,
		_w9478_,
		_w9479_
	);
	LUT3 #(
		.INIT('hd0)
	) name5432 (
		_w9458_,
		_w9473_,
		_w9479_,
		_w9480_
	);
	LUT4 #(
		.INIT('h028a)
	) name5433 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001 ,
		_w9481_
	);
	LUT4 #(
		.INIT('h0145)
	) name5434 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001 ,
		_w9482_
	);
	LUT3 #(
		.INIT('h02)
	) name5435 (
		_w9460_,
		_w9482_,
		_w9481_,
		_w9483_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5436 (
		_w6145_,
		_w6141_,
		_w9463_,
		_w9466_,
		_w9484_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5437 (
		_w6148_,
		_w6163_,
		_w9464_,
		_w9467_,
		_w9485_
	);
	LUT4 #(
		.INIT('h1000)
	) name5438 (
		_w9470_,
		_w9483_,
		_w9484_,
		_w9485_,
		_w9486_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5439 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9487_
	);
	LUT3 #(
		.INIT('h32)
	) name5440 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		_w9475_,
		_w9487_,
		_w9488_
	);
	LUT4 #(
		.INIT('ha820)
	) name5441 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001 ,
		_w9489_
	);
	LUT4 #(
		.INIT('h5410)
	) name5442 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001 ,
		_w9490_
	);
	LUT3 #(
		.INIT('h02)
	) name5443 (
		_w9470_,
		_w9490_,
		_w9489_,
		_w9491_
	);
	LUT2 #(
		.INIT('h2)
	) name5444 (
		_w9488_,
		_w9491_,
		_w9492_
	);
	LUT2 #(
		.INIT('h4)
	) name5445 (
		_w9486_,
		_w9492_,
		_w9493_
	);
	LUT2 #(
		.INIT('h2)
	) name5446 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9494_
	);
	LUT4 #(
		.INIT('h0001)
	) name5447 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w9495_
	);
	LUT2 #(
		.INIT('h2)
	) name5448 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w9495_,
		_w9496_
	);
	LUT2 #(
		.INIT('h2)
	) name5449 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001 ,
		_w9497_
	);
	LUT2 #(
		.INIT('h4)
	) name5450 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w9498_
	);
	LUT4 #(
		.INIT('h4440)
	) name5451 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001 ,
		_w9499_
	);
	LUT2 #(
		.INIT('h4)
	) name5452 (
		_w9497_,
		_w9499_,
		_w9500_
	);
	LUT4 #(
		.INIT('h028a)
	) name5453 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001 ,
		_w9501_
	);
	LUT4 #(
		.INIT('h0145)
	) name5454 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001 ,
		_w9502_
	);
	LUT3 #(
		.INIT('h01)
	) name5455 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w9502_,
		_w9501_,
		_w9503_
	);
	LUT4 #(
		.INIT('h4447)
	) name5456 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001 ,
		_w9496_,
		_w9500_,
		_w9503_,
		_w9504_
	);
	LUT2 #(
		.INIT('h1)
	) name5457 (
		_w9457_,
		_w9475_,
		_w9505_
	);
	LUT4 #(
		.INIT('h1145)
	) name5458 (
		_w9475_,
		_w9494_,
		_w9505_,
		_w9504_,
		_w9506_
	);
	LUT3 #(
		.INIT('h60)
	) name5459 (
		_w9480_,
		_w9493_,
		_w9506_,
		_w9507_
	);
	LUT4 #(
		.INIT('h028a)
	) name5460 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001 ,
		_w9508_
	);
	LUT4 #(
		.INIT('h0145)
	) name5461 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001 ,
		_w9509_
	);
	LUT3 #(
		.INIT('h02)
	) name5462 (
		_w9460_,
		_w9509_,
		_w9508_,
		_w9510_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5463 (
		_w6484_,
		_w6458_,
		_w9463_,
		_w9464_,
		_w9511_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5464 (
		_w6481_,
		_w6477_,
		_w9466_,
		_w9467_,
		_w9512_
	);
	LUT4 #(
		.INIT('h028a)
	) name5465 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001 ,
		_w9513_
	);
	LUT4 #(
		.INIT('h0145)
	) name5466 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001 ,
		_w9514_
	);
	LUT3 #(
		.INIT('h02)
	) name5467 (
		_w9470_,
		_w9514_,
		_w9513_,
		_w9515_
	);
	LUT4 #(
		.INIT('h0040)
	) name5468 (
		_w9510_,
		_w9511_,
		_w9512_,
		_w9515_,
		_w9516_
	);
	LUT2 #(
		.INIT('h2)
	) name5469 (
		_w9488_,
		_w9516_,
		_w9517_
	);
	LUT4 #(
		.INIT('h028a)
	) name5470 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001 ,
		_w9518_
	);
	LUT4 #(
		.INIT('h0145)
	) name5471 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001 ,
		_w9519_
	);
	LUT3 #(
		.INIT('h01)
	) name5472 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9519_,
		_w9518_,
		_w9520_
	);
	LUT2 #(
		.INIT('h2)
	) name5473 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w9521_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5474 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w6456_,
		_w9495_,
		_w9521_,
		_w9522_
	);
	LUT3 #(
		.INIT('h02)
	) name5475 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001 ,
		_w9495_,
		_w9523_
	);
	LUT4 #(
		.INIT('h2022)
	) name5476 (
		_w9505_,
		_w9523_,
		_w9520_,
		_w9522_,
		_w9524_
	);
	LUT3 #(
		.INIT('h3e)
	) name5477 (
		_w9475_,
		_w9494_,
		_w9524_,
		_w9525_
	);
	LUT3 #(
		.INIT('h06)
	) name5478 (
		_w9480_,
		_w9517_,
		_w9525_,
		_w9526_
	);
	LUT4 #(
		.INIT('h028a)
	) name5479 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001 ,
		_w9527_
	);
	LUT4 #(
		.INIT('h0145)
	) name5480 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001 ,
		_w9528_
	);
	LUT3 #(
		.INIT('h02)
	) name5481 (
		_w9460_,
		_w9528_,
		_w9527_,
		_w9529_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5482 (
		_w6860_,
		_w6848_,
		_w9463_,
		_w9464_,
		_w9530_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5483 (
		_w6867_,
		_w6864_,
		_w9466_,
		_w9467_,
		_w9531_
	);
	LUT4 #(
		.INIT('h028a)
	) name5484 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001 ,
		_w9532_
	);
	LUT4 #(
		.INIT('h0145)
	) name5485 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001 ,
		_w9533_
	);
	LUT3 #(
		.INIT('h02)
	) name5486 (
		_w9470_,
		_w9533_,
		_w9532_,
		_w9534_
	);
	LUT4 #(
		.INIT('h0040)
	) name5487 (
		_w9529_,
		_w9530_,
		_w9531_,
		_w9534_,
		_w9535_
	);
	LUT2 #(
		.INIT('h2)
	) name5488 (
		_w9488_,
		_w9535_,
		_w9536_
	);
	LUT4 #(
		.INIT('h028a)
	) name5489 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001 ,
		_w9537_
	);
	LUT4 #(
		.INIT('h0145)
	) name5490 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001 ,
		_w9538_
	);
	LUT3 #(
		.INIT('h01)
	) name5491 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9538_,
		_w9537_,
		_w9539_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5492 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w6852_,
		_w9495_,
		_w9521_,
		_w9540_
	);
	LUT3 #(
		.INIT('h02)
	) name5493 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001 ,
		_w9495_,
		_w9541_
	);
	LUT4 #(
		.INIT('h2022)
	) name5494 (
		_w9505_,
		_w9541_,
		_w9539_,
		_w9540_,
		_w9542_
	);
	LUT3 #(
		.INIT('h3e)
	) name5495 (
		_w9475_,
		_w9494_,
		_w9542_,
		_w9543_
	);
	LUT3 #(
		.INIT('h90)
	) name5496 (
		_w9480_,
		_w9536_,
		_w9543_,
		_w9544_
	);
	LUT4 #(
		.INIT('h028a)
	) name5497 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001 ,
		_w9545_
	);
	LUT4 #(
		.INIT('h0145)
	) name5498 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001 ,
		_w9546_
	);
	LUT3 #(
		.INIT('h02)
	) name5499 (
		_w9460_,
		_w9546_,
		_w9545_,
		_w9547_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5500 (
		_w5872_,
		_w5869_,
		_w9466_,
		_w9467_,
		_w9548_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5501 (
		_w5901_,
		_w5865_,
		_w9463_,
		_w9464_,
		_w9549_
	);
	LUT4 #(
		.INIT('h4555)
	) name5502 (
		_w9470_,
		_w9547_,
		_w9548_,
		_w9549_,
		_w9550_
	);
	LUT4 #(
		.INIT('h028a)
	) name5503 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001 ,
		_w9551_
	);
	LUT4 #(
		.INIT('h0145)
	) name5504 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001 ,
		_w9552_
	);
	LUT3 #(
		.INIT('h02)
	) name5505 (
		_w9470_,
		_w9552_,
		_w9551_,
		_w9553_
	);
	LUT3 #(
		.INIT('ha8)
	) name5506 (
		_w9488_,
		_w9550_,
		_w9553_,
		_w9554_
	);
	LUT2 #(
		.INIT('h9)
	) name5507 (
		_w9480_,
		_w9554_,
		_w9555_
	);
	LUT4 #(
		.INIT('h028a)
	) name5508 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001 ,
		_w9556_
	);
	LUT4 #(
		.INIT('h0145)
	) name5509 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001 ,
		_w9557_
	);
	LUT3 #(
		.INIT('h01)
	) name5510 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9557_,
		_w9556_,
		_w9558_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5511 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w5899_,
		_w9495_,
		_w9521_,
		_w9559_
	);
	LUT3 #(
		.INIT('h02)
	) name5512 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001 ,
		_w9495_,
		_w9560_
	);
	LUT4 #(
		.INIT('h2022)
	) name5513 (
		_w9505_,
		_w9560_,
		_w9558_,
		_w9559_,
		_w9561_
	);
	LUT3 #(
		.INIT('h3e)
	) name5514 (
		_w9475_,
		_w9494_,
		_w9561_,
		_w9562_
	);
	LUT3 #(
		.INIT('h15)
	) name5515 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w9563_
	);
	LUT4 #(
		.INIT('h0777)
	) name5516 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9564_
	);
	LUT4 #(
		.INIT('h0080)
	) name5517 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9565_
	);
	LUT4 #(
		.INIT('h008a)
	) name5518 (
		_w9476_,
		_w9563_,
		_w9564_,
		_w9565_,
		_w9566_
	);
	LUT3 #(
		.INIT('hd0)
	) name5519 (
		_w9458_,
		_w9473_,
		_w9566_,
		_w9567_
	);
	LUT4 #(
		.INIT('h00f9)
	) name5520 (
		_w9480_,
		_w9536_,
		_w9543_,
		_w9567_,
		_w9568_
	);
	LUT3 #(
		.INIT('h90)
	) name5521 (
		_w9480_,
		_w9554_,
		_w9562_,
		_w9569_
	);
	LUT4 #(
		.INIT('h0115)
	) name5522 (
		_w9544_,
		_w9555_,
		_w9562_,
		_w9568_,
		_w9570_
	);
	LUT3 #(
		.INIT('h09)
	) name5523 (
		_w9480_,
		_w9493_,
		_w9506_,
		_w9571_
	);
	LUT4 #(
		.INIT('h028a)
	) name5524 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001 ,
		_w9572_
	);
	LUT4 #(
		.INIT('h0145)
	) name5525 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001 ,
		_w9573_
	);
	LUT3 #(
		.INIT('h02)
	) name5526 (
		_w9460_,
		_w9573_,
		_w9572_,
		_w9574_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5527 (
		_w7671_,
		_w7668_,
		_w9466_,
		_w9467_,
		_w9575_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5528 (
		_w7686_,
		_w7664_,
		_w9463_,
		_w9464_,
		_w9576_
	);
	LUT4 #(
		.INIT('h028a)
	) name5529 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001 ,
		_w9577_
	);
	LUT4 #(
		.INIT('h0145)
	) name5530 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001 ,
		_w9578_
	);
	LUT3 #(
		.INIT('h02)
	) name5531 (
		_w9470_,
		_w9578_,
		_w9577_,
		_w9579_
	);
	LUT4 #(
		.INIT('h0040)
	) name5532 (
		_w9574_,
		_w9575_,
		_w9576_,
		_w9579_,
		_w9580_
	);
	LUT2 #(
		.INIT('h2)
	) name5533 (
		_w9488_,
		_w9580_,
		_w9581_
	);
	LUT2 #(
		.INIT('h2)
	) name5534 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001 ,
		_w9582_
	);
	LUT4 #(
		.INIT('h4440)
	) name5535 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001 ,
		_w9583_
	);
	LUT2 #(
		.INIT('h4)
	) name5536 (
		_w9582_,
		_w9583_,
		_w9584_
	);
	LUT4 #(
		.INIT('h028a)
	) name5537 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001 ,
		_w9585_
	);
	LUT4 #(
		.INIT('h0145)
	) name5538 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001 ,
		_w9586_
	);
	LUT3 #(
		.INIT('h01)
	) name5539 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w9586_,
		_w9585_,
		_w9587_
	);
	LUT4 #(
		.INIT('h4447)
	) name5540 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001 ,
		_w9496_,
		_w9584_,
		_w9587_,
		_w9588_
	);
	LUT4 #(
		.INIT('h1145)
	) name5541 (
		_w9475_,
		_w9494_,
		_w9505_,
		_w9588_,
		_w9589_
	);
	LUT3 #(
		.INIT('h60)
	) name5542 (
		_w9480_,
		_w9581_,
		_w9589_,
		_w9590_
	);
	LUT3 #(
		.INIT('h90)
	) name5543 (
		_w9480_,
		_w9517_,
		_w9525_,
		_w9591_
	);
	LUT3 #(
		.INIT('h45)
	) name5544 (
		_w9571_,
		_w9590_,
		_w9591_,
		_w9592_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5545 (
		_w9507_,
		_w9526_,
		_w9570_,
		_w9592_,
		_w9593_
	);
	LUT4 #(
		.INIT('h028a)
	) name5546 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001 ,
		_w9594_
	);
	LUT4 #(
		.INIT('h0145)
	) name5547 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001 ,
		_w9595_
	);
	LUT3 #(
		.INIT('h02)
	) name5548 (
		_w9460_,
		_w9595_,
		_w9594_,
		_w9596_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5549 (
		_w7346_,
		_w7342_,
		_w9463_,
		_w9466_,
		_w9597_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5550 (
		_w7349_,
		_w7365_,
		_w9464_,
		_w9467_,
		_w9598_
	);
	LUT4 #(
		.INIT('h028a)
	) name5551 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001 ,
		_w9599_
	);
	LUT4 #(
		.INIT('h0145)
	) name5552 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001 ,
		_w9600_
	);
	LUT3 #(
		.INIT('h02)
	) name5553 (
		_w9470_,
		_w9600_,
		_w9599_,
		_w9601_
	);
	LUT4 #(
		.INIT('h0040)
	) name5554 (
		_w9596_,
		_w9597_,
		_w9598_,
		_w9601_,
		_w9602_
	);
	LUT2 #(
		.INIT('h2)
	) name5555 (
		_w9488_,
		_w9602_,
		_w9603_
	);
	LUT4 #(
		.INIT('h028a)
	) name5556 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001 ,
		_w9604_
	);
	LUT4 #(
		.INIT('h0145)
	) name5557 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001 ,
		_w9605_
	);
	LUT3 #(
		.INIT('h01)
	) name5558 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9605_,
		_w9604_,
		_w9606_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5559 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w7363_,
		_w9495_,
		_w9521_,
		_w9607_
	);
	LUT3 #(
		.INIT('h02)
	) name5560 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001 ,
		_w9495_,
		_w9608_
	);
	LUT4 #(
		.INIT('h2022)
	) name5561 (
		_w9505_,
		_w9608_,
		_w9606_,
		_w9607_,
		_w9609_
	);
	LUT3 #(
		.INIT('h3e)
	) name5562 (
		_w9475_,
		_w9494_,
		_w9609_,
		_w9610_
	);
	LUT3 #(
		.INIT('h06)
	) name5563 (
		_w9480_,
		_w9603_,
		_w9610_,
		_w9611_
	);
	LUT2 #(
		.INIT('h1)
	) name5564 (
		_w9590_,
		_w9611_,
		_w9612_
	);
	LUT3 #(
		.INIT('h09)
	) name5565 (
		_w9480_,
		_w9581_,
		_w9589_,
		_w9613_
	);
	LUT3 #(
		.INIT('h90)
	) name5566 (
		_w9480_,
		_w9603_,
		_w9610_,
		_w9614_
	);
	LUT3 #(
		.INIT('h45)
	) name5567 (
		_w9613_,
		_w9507_,
		_w9614_,
		_w9615_
	);
	LUT4 #(
		.INIT('h028a)
	) name5568 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001 ,
		_w9616_
	);
	LUT4 #(
		.INIT('h0145)
	) name5569 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001 ,
		_w9617_
	);
	LUT3 #(
		.INIT('h02)
	) name5570 (
		_w9460_,
		_w9617_,
		_w9616_,
		_w9618_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5571 (
		_w5713_,
		_w7888_,
		_w9463_,
		_w9466_,
		_w9619_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5572 (
		_w7878_,
		_w7884_,
		_w9464_,
		_w9467_,
		_w9620_
	);
	LUT4 #(
		.INIT('h028a)
	) name5573 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001 ,
		_w9621_
	);
	LUT4 #(
		.INIT('h0145)
	) name5574 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001 ,
		_w9622_
	);
	LUT3 #(
		.INIT('h02)
	) name5575 (
		_w9470_,
		_w9622_,
		_w9621_,
		_w9623_
	);
	LUT4 #(
		.INIT('h0040)
	) name5576 (
		_w9618_,
		_w9619_,
		_w9620_,
		_w9623_,
		_w9624_
	);
	LUT2 #(
		.INIT('h2)
	) name5577 (
		_w9488_,
		_w9624_,
		_w9625_
	);
	LUT4 #(
		.INIT('h028a)
	) name5578 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001 ,
		_w9626_
	);
	LUT4 #(
		.INIT('h0145)
	) name5579 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001 ,
		_w9627_
	);
	LUT3 #(
		.INIT('h01)
	) name5580 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9627_,
		_w9626_,
		_w9628_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5581 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w7876_,
		_w9495_,
		_w9521_,
		_w9629_
	);
	LUT3 #(
		.INIT('h02)
	) name5582 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001 ,
		_w9495_,
		_w9630_
	);
	LUT4 #(
		.INIT('h2022)
	) name5583 (
		_w9505_,
		_w9630_,
		_w9628_,
		_w9629_,
		_w9631_
	);
	LUT3 #(
		.INIT('h3e)
	) name5584 (
		_w9475_,
		_w9494_,
		_w9631_,
		_w9632_
	);
	LUT3 #(
		.INIT('h06)
	) name5585 (
		_w9480_,
		_w9625_,
		_w9632_,
		_w9633_
	);
	LUT4 #(
		.INIT('h028a)
	) name5586 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001 ,
		_w9634_
	);
	LUT4 #(
		.INIT('h0145)
	) name5587 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001 ,
		_w9635_
	);
	LUT3 #(
		.INIT('h02)
	) name5588 (
		_w9460_,
		_w9635_,
		_w9634_,
		_w9636_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5589 (
		_w7934_,
		_w8026_,
		_w9463_,
		_w9464_,
		_w9637_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5590 (
		_w8023_,
		_w8019_,
		_w9466_,
		_w9467_,
		_w9638_
	);
	LUT4 #(
		.INIT('h028a)
	) name5591 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001 ,
		_w9639_
	);
	LUT4 #(
		.INIT('h0145)
	) name5592 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001 ,
		_w9640_
	);
	LUT3 #(
		.INIT('h02)
	) name5593 (
		_w9470_,
		_w9640_,
		_w9639_,
		_w9641_
	);
	LUT4 #(
		.INIT('h0040)
	) name5594 (
		_w9636_,
		_w9637_,
		_w9638_,
		_w9641_,
		_w9642_
	);
	LUT2 #(
		.INIT('h2)
	) name5595 (
		_w9488_,
		_w9642_,
		_w9643_
	);
	LUT4 #(
		.INIT('h028a)
	) name5596 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001 ,
		_w9644_
	);
	LUT4 #(
		.INIT('h0145)
	) name5597 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001 ,
		_w9645_
	);
	LUT3 #(
		.INIT('h01)
	) name5598 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9645_,
		_w9644_,
		_w9646_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5599 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w7936_,
		_w9495_,
		_w9521_,
		_w9647_
	);
	LUT3 #(
		.INIT('h02)
	) name5600 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001 ,
		_w9495_,
		_w9648_
	);
	LUT4 #(
		.INIT('h2022)
	) name5601 (
		_w9505_,
		_w9648_,
		_w9646_,
		_w9647_,
		_w9649_
	);
	LUT3 #(
		.INIT('h3e)
	) name5602 (
		_w9475_,
		_w9494_,
		_w9649_,
		_w9650_
	);
	LUT3 #(
		.INIT('h06)
	) name5603 (
		_w9480_,
		_w9643_,
		_w9650_,
		_w9651_
	);
	LUT2 #(
		.INIT('h1)
	) name5604 (
		_w9633_,
		_w9651_,
		_w9652_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5605 (
		_w9593_,
		_w9612_,
		_w9615_,
		_w9652_,
		_w9653_
	);
	LUT3 #(
		.INIT('h90)
	) name5606 (
		_w9480_,
		_w9625_,
		_w9632_,
		_w9654_
	);
	LUT3 #(
		.INIT('h90)
	) name5607 (
		_w9480_,
		_w9643_,
		_w9650_,
		_w9655_
	);
	LUT3 #(
		.INIT('h23)
	) name5608 (
		_w9633_,
		_w9654_,
		_w9655_,
		_w9656_
	);
	LUT4 #(
		.INIT('h028a)
	) name5609 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001 ,
		_w9657_
	);
	LUT4 #(
		.INIT('h0145)
	) name5610 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001 ,
		_w9658_
	);
	LUT3 #(
		.INIT('h02)
	) name5611 (
		_w9460_,
		_w9658_,
		_w9657_,
		_w9659_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5612 (
		_w5713_,
		_w7228_,
		_w9463_,
		_w9464_,
		_w9660_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5613 (
		_w7216_,
		_w7213_,
		_w9466_,
		_w9467_,
		_w9661_
	);
	LUT4 #(
		.INIT('h028a)
	) name5614 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001 ,
		_w9662_
	);
	LUT4 #(
		.INIT('h0145)
	) name5615 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001 ,
		_w9663_
	);
	LUT3 #(
		.INIT('h02)
	) name5616 (
		_w9470_,
		_w9663_,
		_w9662_,
		_w9664_
	);
	LUT4 #(
		.INIT('h0040)
	) name5617 (
		_w9659_,
		_w9660_,
		_w9661_,
		_w9664_,
		_w9665_
	);
	LUT2 #(
		.INIT('h2)
	) name5618 (
		_w9488_,
		_w9665_,
		_w9666_
	);
	LUT4 #(
		.INIT('h028a)
	) name5619 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001 ,
		_w9667_
	);
	LUT4 #(
		.INIT('h0145)
	) name5620 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001 ,
		_w9668_
	);
	LUT3 #(
		.INIT('h01)
	) name5621 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9668_,
		_w9667_,
		_w9669_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5622 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w7224_,
		_w9495_,
		_w9521_,
		_w9670_
	);
	LUT3 #(
		.INIT('h02)
	) name5623 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001 ,
		_w9495_,
		_w9671_
	);
	LUT4 #(
		.INIT('h4044)
	) name5624 (
		_w9671_,
		_w9505_,
		_w9669_,
		_w9670_,
		_w9672_
	);
	LUT3 #(
		.INIT('hc1)
	) name5625 (
		_w9475_,
		_w9494_,
		_w9672_,
		_w9673_
	);
	LUT3 #(
		.INIT('h60)
	) name5626 (
		_w9480_,
		_w9666_,
		_w9673_,
		_w9674_
	);
	LUT4 #(
		.INIT('h028a)
	) name5627 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001 ,
		_w9675_
	);
	LUT4 #(
		.INIT('h0145)
	) name5628 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001 ,
		_w9676_
	);
	LUT3 #(
		.INIT('h02)
	) name5629 (
		_w9460_,
		_w9676_,
		_w9675_,
		_w9677_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5630 (
		_w5713_,
		_w7538_,
		_w9463_,
		_w9464_,
		_w9678_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5631 (
		_w7549_,
		_w7545_,
		_w9466_,
		_w9467_,
		_w9679_
	);
	LUT4 #(
		.INIT('h028a)
	) name5632 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001 ,
		_w9680_
	);
	LUT4 #(
		.INIT('h0145)
	) name5633 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001 ,
		_w9681_
	);
	LUT3 #(
		.INIT('h02)
	) name5634 (
		_w9470_,
		_w9681_,
		_w9680_,
		_w9682_
	);
	LUT4 #(
		.INIT('h0040)
	) name5635 (
		_w9677_,
		_w9678_,
		_w9679_,
		_w9682_,
		_w9683_
	);
	LUT2 #(
		.INIT('h2)
	) name5636 (
		_w9488_,
		_w9683_,
		_w9684_
	);
	LUT4 #(
		.INIT('h028a)
	) name5637 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001 ,
		_w9685_
	);
	LUT4 #(
		.INIT('h0145)
	) name5638 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001 ,
		_w9686_
	);
	LUT3 #(
		.INIT('h01)
	) name5639 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9686_,
		_w9685_,
		_w9687_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5640 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w7534_,
		_w9495_,
		_w9521_,
		_w9688_
	);
	LUT3 #(
		.INIT('h02)
	) name5641 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001 ,
		_w9495_,
		_w9689_
	);
	LUT4 #(
		.INIT('h2022)
	) name5642 (
		_w9505_,
		_w9689_,
		_w9687_,
		_w9688_,
		_w9690_
	);
	LUT3 #(
		.INIT('h3e)
	) name5643 (
		_w9475_,
		_w9494_,
		_w9690_,
		_w9691_
	);
	LUT3 #(
		.INIT('h06)
	) name5644 (
		_w9480_,
		_w9684_,
		_w9691_,
		_w9692_
	);
	LUT2 #(
		.INIT('h1)
	) name5645 (
		_w9674_,
		_w9692_,
		_w9693_
	);
	LUT4 #(
		.INIT('h028a)
	) name5646 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001 ,
		_w9694_
	);
	LUT4 #(
		.INIT('h0145)
	) name5647 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001 ,
		_w9695_
	);
	LUT3 #(
		.INIT('h02)
	) name5648 (
		_w9460_,
		_w9695_,
		_w9694_,
		_w9696_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5649 (
		_w5713_,
		_w6335_,
		_w9463_,
		_w9466_,
		_w9697_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5650 (
		_w6331_,
		_w6349_,
		_w9464_,
		_w9467_,
		_w9698_
	);
	LUT4 #(
		.INIT('h028a)
	) name5651 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001 ,
		_w9699_
	);
	LUT4 #(
		.INIT('h0145)
	) name5652 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001 ,
		_w9700_
	);
	LUT3 #(
		.INIT('h02)
	) name5653 (
		_w9470_,
		_w9700_,
		_w9699_,
		_w9701_
	);
	LUT4 #(
		.INIT('h0040)
	) name5654 (
		_w9696_,
		_w9697_,
		_w9698_,
		_w9701_,
		_w9702_
	);
	LUT2 #(
		.INIT('h2)
	) name5655 (
		_w9488_,
		_w9702_,
		_w9703_
	);
	LUT4 #(
		.INIT('h028a)
	) name5656 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001 ,
		_w9704_
	);
	LUT4 #(
		.INIT('h0145)
	) name5657 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001 ,
		_w9705_
	);
	LUT3 #(
		.INIT('h01)
	) name5658 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9705_,
		_w9704_,
		_w9706_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5659 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w6353_,
		_w9495_,
		_w9521_,
		_w9707_
	);
	LUT3 #(
		.INIT('h02)
	) name5660 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001 ,
		_w9495_,
		_w9708_
	);
	LUT4 #(
		.INIT('h2022)
	) name5661 (
		_w9505_,
		_w9708_,
		_w9706_,
		_w9707_,
		_w9709_
	);
	LUT3 #(
		.INIT('hc1)
	) name5662 (
		_w9475_,
		_w9494_,
		_w9709_,
		_w9710_
	);
	LUT3 #(
		.INIT('h60)
	) name5663 (
		_w9480_,
		_w9703_,
		_w9710_,
		_w9711_
	);
	LUT3 #(
		.INIT('h90)
	) name5664 (
		_w9480_,
		_w9684_,
		_w9691_,
		_w9712_
	);
	LUT3 #(
		.INIT('h09)
	) name5665 (
		_w9480_,
		_w9666_,
		_w9673_,
		_w9713_
	);
	LUT3 #(
		.INIT('h0b)
	) name5666 (
		_w9711_,
		_w9712_,
		_w9713_,
		_w9714_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5667 (
		_w9653_,
		_w9656_,
		_w9693_,
		_w9714_,
		_w9715_
	);
	LUT4 #(
		.INIT('h028a)
	) name5668 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001 ,
		_w9716_
	);
	LUT4 #(
		.INIT('h0145)
	) name5669 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001 ,
		_w9717_
	);
	LUT3 #(
		.INIT('h02)
	) name5670 (
		_w9460_,
		_w9717_,
		_w9716_,
		_w9718_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5671 (
		_w5713_,
		_w6011_,
		_w9463_,
		_w9466_,
		_w9719_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5672 (
		_w6014_,
		_w6026_,
		_w9464_,
		_w9467_,
		_w9720_
	);
	LUT4 #(
		.INIT('h028a)
	) name5673 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001 ,
		_w9721_
	);
	LUT4 #(
		.INIT('h0145)
	) name5674 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001 ,
		_w9722_
	);
	LUT3 #(
		.INIT('h02)
	) name5675 (
		_w9470_,
		_w9722_,
		_w9721_,
		_w9723_
	);
	LUT4 #(
		.INIT('h0040)
	) name5676 (
		_w9718_,
		_w9719_,
		_w9720_,
		_w9723_,
		_w9724_
	);
	LUT2 #(
		.INIT('h2)
	) name5677 (
		_w9488_,
		_w9724_,
		_w9725_
	);
	LUT4 #(
		.INIT('h028a)
	) name5678 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001 ,
		_w9726_
	);
	LUT4 #(
		.INIT('h0145)
	) name5679 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001 ,
		_w9727_
	);
	LUT3 #(
		.INIT('h01)
	) name5680 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9727_,
		_w9726_,
		_w9728_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5681 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w6023_,
		_w9495_,
		_w9521_,
		_w9729_
	);
	LUT3 #(
		.INIT('h02)
	) name5682 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001 ,
		_w9495_,
		_w9730_
	);
	LUT4 #(
		.INIT('h2022)
	) name5683 (
		_w9505_,
		_w9730_,
		_w9728_,
		_w9729_,
		_w9731_
	);
	LUT3 #(
		.INIT('hc1)
	) name5684 (
		_w9475_,
		_w9494_,
		_w9731_,
		_w9732_
	);
	LUT3 #(
		.INIT('h60)
	) name5685 (
		_w9480_,
		_w9725_,
		_w9732_,
		_w9733_
	);
	LUT2 #(
		.INIT('h1)
	) name5686 (
		_w9711_,
		_w9733_,
		_w9734_
	);
	LUT3 #(
		.INIT('h09)
	) name5687 (
		_w9480_,
		_w9703_,
		_w9710_,
		_w9735_
	);
	LUT3 #(
		.INIT('h09)
	) name5688 (
		_w9480_,
		_w9725_,
		_w9732_,
		_w9736_
	);
	LUT3 #(
		.INIT('h23)
	) name5689 (
		_w9674_,
		_w9735_,
		_w9736_,
		_w9737_
	);
	LUT4 #(
		.INIT('h1055)
	) name5690 (
		_w9456_,
		_w9715_,
		_w9734_,
		_w9737_,
		_w9738_
	);
	LUT4 #(
		.INIT('h028a)
	) name5691 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001 ,
		_w9739_
	);
	LUT4 #(
		.INIT('h0145)
	) name5692 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001 ,
		_w9740_
	);
	LUT3 #(
		.INIT('h02)
	) name5693 (
		_w9460_,
		_w9740_,
		_w9739_,
		_w9741_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5694 (
		_w5713_,
		_w6731_,
		_w9463_,
		_w9466_,
		_w9742_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5695 (
		_w6734_,
		_w6746_,
		_w9464_,
		_w9467_,
		_w9743_
	);
	LUT4 #(
		.INIT('h028a)
	) name5696 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001 ,
		_w9744_
	);
	LUT4 #(
		.INIT('h0145)
	) name5697 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001 ,
		_w9745_
	);
	LUT3 #(
		.INIT('h02)
	) name5698 (
		_w9470_,
		_w9745_,
		_w9744_,
		_w9746_
	);
	LUT4 #(
		.INIT('h0040)
	) name5699 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9746_,
		_w9747_
	);
	LUT2 #(
		.INIT('h2)
	) name5700 (
		_w9488_,
		_w9747_,
		_w9748_
	);
	LUT4 #(
		.INIT('h028a)
	) name5701 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001 ,
		_w9749_
	);
	LUT4 #(
		.INIT('h0145)
	) name5702 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001 ,
		_w9750_
	);
	LUT3 #(
		.INIT('h01)
	) name5703 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9750_,
		_w9749_,
		_w9751_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5704 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w6742_,
		_w9495_,
		_w9521_,
		_w9752_
	);
	LUT3 #(
		.INIT('h02)
	) name5705 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001 ,
		_w9495_,
		_w9753_
	);
	LUT4 #(
		.INIT('h2022)
	) name5706 (
		_w9505_,
		_w9753_,
		_w9751_,
		_w9752_,
		_w9754_
	);
	LUT3 #(
		.INIT('h3e)
	) name5707 (
		_w9475_,
		_w9494_,
		_w9754_,
		_w9755_
	);
	LUT3 #(
		.INIT('h90)
	) name5708 (
		_w9480_,
		_w9748_,
		_w9755_,
		_w9756_
	);
	LUT3 #(
		.INIT('h40)
	) name5709 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9757_
	);
	LUT4 #(
		.INIT('h0090)
	) name5710 (
		_w9480_,
		_w9748_,
		_w9755_,
		_w9757_,
		_w9758_
	);
	LUT4 #(
		.INIT('h1000)
	) name5711 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w9759_
	);
	LUT3 #(
		.INIT('h06)
	) name5712 (
		_w9480_,
		_w9748_,
		_w9755_,
		_w9760_
	);
	LUT4 #(
		.INIT('h90f9)
	) name5713 (
		_w9480_,
		_w9748_,
		_w9755_,
		_w9759_,
		_w9761_
	);
	LUT2 #(
		.INIT('h4)
	) name5714 (
		_w9758_,
		_w9761_,
		_w9762_
	);
	LUT2 #(
		.INIT('h9)
	) name5715 (
		_w9738_,
		_w9762_,
		_w9763_
	);
	LUT4 #(
		.INIT('hf600)
	) name5716 (
		_w9480_,
		_w9703_,
		_w9710_,
		_w9759_,
		_w9764_
	);
	LUT4 #(
		.INIT('h9f96)
	) name5717 (
		_w9480_,
		_w9703_,
		_w9710_,
		_w9757_,
		_w9765_
	);
	LUT2 #(
		.INIT('h4)
	) name5718 (
		_w9764_,
		_w9765_,
		_w9766_
	);
	LUT4 #(
		.INIT('h4155)
	) name5719 (
		_w9456_,
		_w9480_,
		_w9725_,
		_w9732_,
		_w9767_
	);
	LUT4 #(
		.INIT('hd20f)
	) name5720 (
		_w9715_,
		_w9736_,
		_w9766_,
		_w9767_,
		_w9768_
	);
	LUT4 #(
		.INIT('h14be)
	) name5721 (
		_w9455_,
		_w9738_,
		_w9762_,
		_w9768_,
		_w9769_
	);
	LUT3 #(
		.INIT('he2)
	) name5722 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001 ,
		_w9454_,
		_w9769_,
		_w9770_
	);
	LUT4 #(
		.INIT('h028a)
	) name5723 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001 ,
		_w9771_
	);
	LUT4 #(
		.INIT('h0145)
	) name5724 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001 ,
		_w9772_
	);
	LUT3 #(
		.INIT('h02)
	) name5725 (
		_w9460_,
		_w9772_,
		_w9771_,
		_w9773_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5726 (
		_w5720_,
		_w5713_,
		_w9463_,
		_w9466_,
		_w9774_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5727 (
		_w5734_,
		_w5717_,
		_w9464_,
		_w9467_,
		_w9775_
	);
	LUT4 #(
		.INIT('h1000)
	) name5728 (
		_w9470_,
		_w9773_,
		_w9774_,
		_w9775_,
		_w9776_
	);
	LUT4 #(
		.INIT('ha820)
	) name5729 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001 ,
		_w9777_
	);
	LUT4 #(
		.INIT('h5410)
	) name5730 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001 ,
		_w9778_
	);
	LUT3 #(
		.INIT('h02)
	) name5731 (
		_w9470_,
		_w9778_,
		_w9777_,
		_w9779_
	);
	LUT2 #(
		.INIT('h2)
	) name5732 (
		_w9488_,
		_w9779_,
		_w9780_
	);
	LUT2 #(
		.INIT('h4)
	) name5733 (
		_w9776_,
		_w9780_,
		_w9781_
	);
	LUT2 #(
		.INIT('h2)
	) name5734 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001 ,
		_w9782_
	);
	LUT4 #(
		.INIT('h4440)
	) name5735 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001 ,
		_w9783_
	);
	LUT2 #(
		.INIT('h4)
	) name5736 (
		_w9782_,
		_w9783_,
		_w9784_
	);
	LUT4 #(
		.INIT('h028a)
	) name5737 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001 ,
		_w9785_
	);
	LUT4 #(
		.INIT('h0145)
	) name5738 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001 ,
		_w9786_
	);
	LUT3 #(
		.INIT('h01)
	) name5739 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w9786_,
		_w9785_,
		_w9787_
	);
	LUT4 #(
		.INIT('h4447)
	) name5740 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001 ,
		_w9496_,
		_w9784_,
		_w9787_,
		_w9788_
	);
	LUT4 #(
		.INIT('h1145)
	) name5741 (
		_w9475_,
		_w9494_,
		_w9505_,
		_w9788_,
		_w9789_
	);
	LUT3 #(
		.INIT('h60)
	) name5742 (
		_w9480_,
		_w9781_,
		_w9789_,
		_w9790_
	);
	LUT2 #(
		.INIT('h1)
	) name5743 (
		_w9760_,
		_w9790_,
		_w9791_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5744 (
		_w9715_,
		_w9734_,
		_w9737_,
		_w9791_,
		_w9792_
	);
	LUT3 #(
		.INIT('h09)
	) name5745 (
		_w9480_,
		_w9781_,
		_w9789_,
		_w9793_
	);
	LUT4 #(
		.INIT('h1c2f)
	) name5746 (
		_w9458_,
		_w9473_,
		_w9479_,
		_w9488_,
		_w9794_
	);
	LUT4 #(
		.INIT('h028a)
	) name5747 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001 ,
		_w9795_
	);
	LUT4 #(
		.INIT('h0145)
	) name5748 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001 ,
		_w9796_
	);
	LUT3 #(
		.INIT('h01)
	) name5749 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w9796_,
		_w9795_,
		_w9797_
	);
	LUT2 #(
		.INIT('h2)
	) name5750 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001 ,
		_w9798_
	);
	LUT4 #(
		.INIT('h4440)
	) name5751 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001 ,
		_w9799_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name5752 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w9495_,
		_w9798_,
		_w9799_,
		_w9800_
	);
	LUT3 #(
		.INIT('h02)
	) name5753 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001 ,
		_w9495_,
		_w9801_
	);
	LUT4 #(
		.INIT('h008a)
	) name5754 (
		_w9505_,
		_w9797_,
		_w9800_,
		_w9801_,
		_w9802_
	);
	LUT3 #(
		.INIT('hc1)
	) name5755 (
		_w9475_,
		_w9494_,
		_w9802_,
		_w9803_
	);
	LUT2 #(
		.INIT('h4)
	) name5756 (
		_w9794_,
		_w9803_,
		_w9804_
	);
	LUT3 #(
		.INIT('h31)
	) name5757 (
		_w9756_,
		_w9793_,
		_w9804_,
		_w9805_
	);
	LUT4 #(
		.INIT('h028a)
	) name5758 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001 ,
		_w9806_
	);
	LUT4 #(
		.INIT('h0145)
	) name5759 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001 ,
		_w9807_
	);
	LUT3 #(
		.INIT('h02)
	) name5760 (
		_w9460_,
		_w9807_,
		_w9806_,
		_w9808_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5761 (
		_w5713_,
		_w8267_,
		_w9463_,
		_w9464_,
		_w9809_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5762 (
		_w8296_,
		_w8292_,
		_w9466_,
		_w9467_,
		_w9810_
	);
	LUT4 #(
		.INIT('h028a)
	) name5763 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001 ,
		_w9811_
	);
	LUT4 #(
		.INIT('h0145)
	) name5764 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001 ,
		_w9812_
	);
	LUT3 #(
		.INIT('h02)
	) name5765 (
		_w9470_,
		_w9812_,
		_w9811_,
		_w9813_
	);
	LUT4 #(
		.INIT('h0040)
	) name5766 (
		_w9808_,
		_w9809_,
		_w9810_,
		_w9813_,
		_w9814_
	);
	LUT2 #(
		.INIT('h2)
	) name5767 (
		_w9488_,
		_w9814_,
		_w9815_
	);
	LUT4 #(
		.INIT('h028a)
	) name5768 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001 ,
		_w9816_
	);
	LUT4 #(
		.INIT('h0145)
	) name5769 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001 ,
		_w9817_
	);
	LUT3 #(
		.INIT('h01)
	) name5770 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9817_,
		_w9816_,
		_w9818_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5771 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w8271_,
		_w9495_,
		_w9521_,
		_w9819_
	);
	LUT3 #(
		.INIT('h02)
	) name5772 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001 ,
		_w9495_,
		_w9820_
	);
	LUT4 #(
		.INIT('h2022)
	) name5773 (
		_w9505_,
		_w9820_,
		_w9818_,
		_w9819_,
		_w9821_
	);
	LUT3 #(
		.INIT('h3e)
	) name5774 (
		_w9475_,
		_w9494_,
		_w9821_,
		_w9822_
	);
	LUT3 #(
		.INIT('h90)
	) name5775 (
		_w9480_,
		_w9815_,
		_w9822_,
		_w9823_
	);
	LUT4 #(
		.INIT('h8400)
	) name5776 (
		_w9480_,
		_w9757_,
		_w9815_,
		_w9822_,
		_w9824_
	);
	LUT3 #(
		.INIT('h06)
	) name5777 (
		_w9480_,
		_w9815_,
		_w9822_,
		_w9825_
	);
	LUT4 #(
		.INIT('h1221)
	) name5778 (
		_w9480_,
		_w9759_,
		_w9815_,
		_w9822_,
		_w9826_
	);
	LUT2 #(
		.INIT('h1)
	) name5779 (
		_w9824_,
		_w9826_,
		_w9827_
	);
	LUT4 #(
		.INIT('h45ba)
	) name5780 (
		_w9456_,
		_w9792_,
		_w9805_,
		_w9827_,
		_w9828_
	);
	LUT4 #(
		.INIT('h0021)
	) name5781 (
		_w9480_,
		_w9757_,
		_w9781_,
		_w9789_,
		_w9829_
	);
	LUT4 #(
		.INIT('h21b7)
	) name5782 (
		_w9480_,
		_w9759_,
		_w9781_,
		_w9789_,
		_w9830_
	);
	LUT2 #(
		.INIT('h4)
	) name5783 (
		_w9829_,
		_w9830_,
		_w9831_
	);
	LUT4 #(
		.INIT('h00b0)
	) name5784 (
		_w9715_,
		_w9734_,
		_w9737_,
		_w9756_,
		_w9832_
	);
	LUT4 #(
		.INIT('h5541)
	) name5785 (
		_w9456_,
		_w9480_,
		_w9748_,
		_w9755_,
		_w9833_
	);
	LUT3 #(
		.INIT('h65)
	) name5786 (
		_w9831_,
		_w9832_,
		_w9833_,
		_w9834_
	);
	LUT4 #(
		.INIT('h8a02)
	) name5787 (
		_w9454_,
		_w9455_,
		_w9828_,
		_w9834_,
		_w9835_
	);
	LUT2 #(
		.INIT('h1)
	) name5788 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001 ,
		_w9454_,
		_w9836_
	);
	LUT2 #(
		.INIT('h1)
	) name5789 (
		_w9835_,
		_w9836_,
		_w9837_
	);
	LUT4 #(
		.INIT('h0455)
	) name5790 (
		_w9456_,
		_w9458_,
		_w9473_,
		_w9566_,
		_w9838_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5791 (
		_w9480_,
		_w9554_,
		_w9562_,
		_w9759_,
		_w9839_
	);
	LUT4 #(
		.INIT('hf969)
	) name5792 (
		_w9480_,
		_w9554_,
		_w9562_,
		_w9757_,
		_w9840_
	);
	LUT3 #(
		.INIT('h65)
	) name5793 (
		_w9838_,
		_w9839_,
		_w9840_,
		_w9841_
	);
	LUT4 #(
		.INIT('h8288)
	) name5794 (
		_w9455_,
		_w9838_,
		_w9839_,
		_w9840_,
		_w9842_
	);
	LUT3 #(
		.INIT('h54)
	) name5795 (
		_w9456_,
		_w9568_,
		_w9569_,
		_w9843_
	);
	LUT4 #(
		.INIT('h9000)
	) name5796 (
		_w9480_,
		_w9536_,
		_w9543_,
		_w9757_,
		_w9844_
	);
	LUT4 #(
		.INIT('h0069)
	) name5797 (
		_w9480_,
		_w9536_,
		_w9543_,
		_w9759_,
		_w9845_
	);
	LUT2 #(
		.INIT('h1)
	) name5798 (
		_w9844_,
		_w9845_,
		_w9846_
	);
	LUT2 #(
		.INIT('h9)
	) name5799 (
		_w9843_,
		_w9846_,
		_w9847_
	);
	LUT4 #(
		.INIT('h2332)
	) name5800 (
		_w9455_,
		_w9842_,
		_w9843_,
		_w9846_,
		_w9848_
	);
	LUT3 #(
		.INIT('h2e)
	) name5801 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001 ,
		_w9454_,
		_w9848_,
		_w9849_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5802 (
		_w9480_,
		_w9517_,
		_w9525_,
		_w9759_,
		_w9850_
	);
	LUT4 #(
		.INIT('hf969)
	) name5803 (
		_w9480_,
		_w9517_,
		_w9525_,
		_w9757_,
		_w9851_
	);
	LUT2 #(
		.INIT('h4)
	) name5804 (
		_w9850_,
		_w9851_,
		_w9852_
	);
	LUT3 #(
		.INIT('h1e)
	) name5805 (
		_w9456_,
		_w9570_,
		_w9852_,
		_w9853_
	);
	LUT4 #(
		.INIT('h5401)
	) name5806 (
		_w9455_,
		_w9456_,
		_w9570_,
		_w9852_,
		_w9854_
	);
	LUT3 #(
		.INIT('h82)
	) name5807 (
		_w9455_,
		_w9843_,
		_w9846_,
		_w9855_
	);
	LUT4 #(
		.INIT('heee2)
	) name5808 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001 ,
		_w9454_,
		_w9854_,
		_w9855_,
		_w9856_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5809 (
		_w9480_,
		_w9603_,
		_w9610_,
		_w9759_,
		_w9857_
	);
	LUT4 #(
		.INIT('hf969)
	) name5810 (
		_w9480_,
		_w9603_,
		_w9610_,
		_w9757_,
		_w9858_
	);
	LUT2 #(
		.INIT('h4)
	) name5811 (
		_w9857_,
		_w9858_,
		_w9859_
	);
	LUT3 #(
		.INIT('h1e)
	) name5812 (
		_w9456_,
		_w9593_,
		_w9859_,
		_w9860_
	);
	LUT4 #(
		.INIT('h5401)
	) name5813 (
		_w9455_,
		_w9456_,
		_w9593_,
		_w9859_,
		_w9861_
	);
	LUT4 #(
		.INIT('h5501)
	) name5814 (
		_w9456_,
		_w9526_,
		_w9570_,
		_w9591_,
		_w9862_
	);
	LUT4 #(
		.INIT('hf600)
	) name5815 (
		_w9480_,
		_w9493_,
		_w9506_,
		_w9759_,
		_w9863_
	);
	LUT4 #(
		.INIT('h9f96)
	) name5816 (
		_w9480_,
		_w9493_,
		_w9506_,
		_w9757_,
		_w9864_
	);
	LUT2 #(
		.INIT('h4)
	) name5817 (
		_w9863_,
		_w9864_,
		_w9865_
	);
	LUT2 #(
		.INIT('h9)
	) name5818 (
		_w9862_,
		_w9865_,
		_w9866_
	);
	LUT3 #(
		.INIT('h28)
	) name5819 (
		_w9455_,
		_w9862_,
		_w9865_,
		_w9867_
	);
	LUT4 #(
		.INIT('heee2)
	) name5820 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001 ,
		_w9454_,
		_w9861_,
		_w9867_,
		_w9868_
	);
	LUT4 #(
		.INIT('h1055)
	) name5821 (
		_w9456_,
		_w9593_,
		_w9612_,
		_w9615_,
		_w9869_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5822 (
		_w9480_,
		_w9643_,
		_w9650_,
		_w9759_,
		_w9870_
	);
	LUT4 #(
		.INIT('hf969)
	) name5823 (
		_w9480_,
		_w9643_,
		_w9650_,
		_w9757_,
		_w9871_
	);
	LUT2 #(
		.INIT('h4)
	) name5824 (
		_w9870_,
		_w9871_,
		_w9872_
	);
	LUT2 #(
		.INIT('h9)
	) name5825 (
		_w9869_,
		_w9872_,
		_w9873_
	);
	LUT4 #(
		.INIT('hf600)
	) name5826 (
		_w9480_,
		_w9581_,
		_w9589_,
		_w9759_,
		_w9874_
	);
	LUT4 #(
		.INIT('h9f96)
	) name5827 (
		_w9480_,
		_w9581_,
		_w9589_,
		_w9757_,
		_w9875_
	);
	LUT2 #(
		.INIT('h4)
	) name5828 (
		_w9874_,
		_w9875_,
		_w9876_
	);
	LUT4 #(
		.INIT('h5541)
	) name5829 (
		_w9456_,
		_w9480_,
		_w9603_,
		_w9610_,
		_w9877_
	);
	LUT4 #(
		.INIT('hb40f)
	) name5830 (
		_w9614_,
		_w9593_,
		_w9876_,
		_w9877_,
		_w9878_
	);
	LUT4 #(
		.INIT('heb41)
	) name5831 (
		_w9455_,
		_w9869_,
		_w9872_,
		_w9878_,
		_w9879_
	);
	LUT3 #(
		.INIT('h2e)
	) name5832 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001 ,
		_w9454_,
		_w9879_,
		_w9880_
	);
	LUT4 #(
		.INIT('hf600)
	) name5833 (
		_w9480_,
		_w9666_,
		_w9673_,
		_w9759_,
		_w9881_
	);
	LUT4 #(
		.INIT('h9f96)
	) name5834 (
		_w9480_,
		_w9666_,
		_w9673_,
		_w9757_,
		_w9882_
	);
	LUT2 #(
		.INIT('h4)
	) name5835 (
		_w9881_,
		_w9882_,
		_w9883_
	);
	LUT4 #(
		.INIT('h5541)
	) name5836 (
		_w9456_,
		_w9480_,
		_w9684_,
		_w9691_,
		_w9884_
	);
	LUT4 #(
		.INIT('hfb00)
	) name5837 (
		_w9653_,
		_w9656_,
		_w9712_,
		_w9884_,
		_w9885_
	);
	LUT2 #(
		.INIT('h9)
	) name5838 (
		_w9883_,
		_w9885_,
		_w9886_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5839 (
		_w9480_,
		_w9684_,
		_w9691_,
		_w9759_,
		_w9887_
	);
	LUT4 #(
		.INIT('hf969)
	) name5840 (
		_w9480_,
		_w9684_,
		_w9691_,
		_w9757_,
		_w9888_
	);
	LUT2 #(
		.INIT('h4)
	) name5841 (
		_w9887_,
		_w9888_,
		_w9889_
	);
	LUT4 #(
		.INIT('h45ba)
	) name5842 (
		_w9456_,
		_w9653_,
		_w9656_,
		_w9889_,
		_w9890_
	);
	LUT4 #(
		.INIT('heb41)
	) name5843 (
		_w9455_,
		_w9883_,
		_w9885_,
		_w9890_,
		_w9891_
	);
	LUT3 #(
		.INIT('h2e)
	) name5844 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001 ,
		_w9454_,
		_w9891_,
		_w9892_
	);
	LUT3 #(
		.INIT('h8a)
	) name5845 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9893_
	);
	LUT4 #(
		.INIT('h4044)
	) name5846 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9894_
	);
	LUT3 #(
		.INIT('h10)
	) name5847 (
		_w9451_,
		_w9453_,
		_w9894_,
		_w9895_
	);
	LUT3 #(
		.INIT('hca)
	) name5848 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001 ,
		_w9769_,
		_w9895_,
		_w9896_
	);
	LUT4 #(
		.INIT('hb100)
	) name5849 (
		_w9455_,
		_w9828_,
		_w9834_,
		_w9895_,
		_w9897_
	);
	LUT4 #(
		.INIT('h5455)
	) name5850 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001 ,
		_w9451_,
		_w9453_,
		_w9894_,
		_w9898_
	);
	LUT2 #(
		.INIT('h1)
	) name5851 (
		_w9897_,
		_w9898_,
		_w9899_
	);
	LUT3 #(
		.INIT('h3a)
	) name5852 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001 ,
		_w9848_,
		_w9895_,
		_w9900_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5853 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001 ,
		_w9854_,
		_w9855_,
		_w9895_,
		_w9901_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5854 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001 ,
		_w9861_,
		_w9867_,
		_w9895_,
		_w9902_
	);
	LUT3 #(
		.INIT('h3a)
	) name5855 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001 ,
		_w9879_,
		_w9895_,
		_w9903_
	);
	LUT3 #(
		.INIT('h3a)
	) name5856 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001 ,
		_w9891_,
		_w9895_,
		_w9904_
	);
	LUT4 #(
		.INIT('h2022)
	) name5857 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w7927_,
		_w8040_,
		_w8042_,
		_w9905_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5858 (
		\core_c_dec_RTI_Ed_reg/P0001 ,
		_w4160_,
		_w4158_,
		_w4167_,
		_w9906_
	);
	LUT2 #(
		.INIT('h8)
	) name5859 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w9907_
	);
	LUT2 #(
		.INIT('h8)
	) name5860 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		_w9908_
	);
	LUT3 #(
		.INIT('h80)
	) name5861 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9909_
	);
	LUT3 #(
		.INIT('h0e)
	) name5862 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w9906_,
		_w9909_,
		_w9910_
	);
	LUT4 #(
		.INIT('h00ec)
	) name5863 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w9906_,
		_w9907_,
		_w9909_,
		_w9911_
	);
	LUT3 #(
		.INIT('h04)
	) name5864 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9912_
	);
	LUT4 #(
		.INIT('h0400)
	) name5865 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001 ,
		_w9913_
	);
	LUT3 #(
		.INIT('h02)
	) name5866 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9914_
	);
	LUT4 #(
		.INIT('h0200)
	) name5867 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001 ,
		_w9915_
	);
	LUT3 #(
		.INIT('h40)
	) name5868 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9916_
	);
	LUT4 #(
		.INIT('h4000)
	) name5869 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001 ,
		_w9917_
	);
	LUT3 #(
		.INIT('h01)
	) name5870 (
		_w9915_,
		_w9917_,
		_w9913_,
		_w9918_
	);
	LUT3 #(
		.INIT('h20)
	) name5871 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9919_
	);
	LUT4 #(
		.INIT('h2000)
	) name5872 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001 ,
		_w9920_
	);
	LUT2 #(
		.INIT('h1)
	) name5873 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		_w9921_
	);
	LUT3 #(
		.INIT('h01)
	) name5874 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9922_
	);
	LUT4 #(
		.INIT('h0100)
	) name5875 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001 ,
		_w9923_
	);
	LUT4 #(
		.INIT('h0800)
	) name5876 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001 ,
		_w9924_
	);
	LUT3 #(
		.INIT('h10)
	) name5877 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9925_
	);
	LUT4 #(
		.INIT('h1000)
	) name5878 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001 ,
		_w9926_
	);
	LUT4 #(
		.INIT('h0001)
	) name5879 (
		_w9920_,
		_w9923_,
		_w9924_,
		_w9926_,
		_w9927_
	);
	LUT2 #(
		.INIT('h8)
	) name5880 (
		_w9918_,
		_w9927_,
		_w9928_
	);
	LUT2 #(
		.INIT('h2)
	) name5881 (
		_w9911_,
		_w9928_,
		_w9929_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name5882 (
		\core_eu_ec_cun_MVi_pre_C_reg/P0001 ,
		_w4971_,
		_w9905_,
		_w9929_,
		_w9930_
	);
	LUT4 #(
		.INIT('h0004)
	) name5883 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w9931_
	);
	LUT2 #(
		.INIT('h4)
	) name5884 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w9931_,
		_w9932_
	);
	LUT4 #(
		.INIT('h00bf)
	) name5885 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w9932_,
		_w9933_
	);
	LUT4 #(
		.INIT('h1000)
	) name5886 (
		\core_eu_em_mac_em_reg_Sq_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w9934_
	);
	LUT3 #(
		.INIT('h01)
	) name5887 (
		_w4516_,
		_w9934_,
		_w9933_,
		_w9935_
	);
	LUT4 #(
		.INIT('h0145)
	) name5888 (
		\emc_EXTC_Eg_syn_reg/P0001 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		_w9936_
	);
	LUT4 #(
		.INIT('h0080)
	) name5889 (
		_w4738_,
		_w4729_,
		_w4745_,
		_w9936_,
		_w9937_
	);
	LUT2 #(
		.INIT('h1)
	) name5890 (
		\memc_Dread_E_reg/NET0131 ,
		\memc_IOcmd_E_reg/NET0131 ,
		_w9938_
	);
	LUT2 #(
		.INIT('h2)
	) name5891 (
		_w4719_,
		_w9938_,
		_w9939_
	);
	LUT2 #(
		.INIT('h8)
	) name5892 (
		_w9937_,
		_w9939_,
		_w9940_
	);
	LUT4 #(
		.INIT('hcacc)
	) name5893 (
		\T_ED[8]_pad ,
		\emc_DMDreg_reg[8]/P0001 ,
		_w8594_,
		_w9940_,
		_w9941_
	);
	LUT4 #(
		.INIT('hcacc)
	) name5894 (
		\T_ED[9]_pad ,
		\emc_DMDreg_reg[9]/P0001 ,
		_w8594_,
		_w9940_,
		_w9942_
	);
	LUT2 #(
		.INIT('h8)
	) name5895 (
		\memc_Pread_E_reg/NET0131 ,
		_w4721_,
		_w9943_
	);
	LUT4 #(
		.INIT('haccc)
	) name5896 (
		\T_ED[8]_pad ,
		\emc_PMDreg_reg[8]/P0001 ,
		_w9937_,
		_w9943_,
		_w9944_
	);
	LUT4 #(
		.INIT('haccc)
	) name5897 (
		\T_ED[9]_pad ,
		\emc_PMDreg_reg[9]/P0001 ,
		_w9937_,
		_w9943_,
		_w9945_
	);
	LUT4 #(
		.INIT('h0040)
	) name5898 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_updMR_E_reg/P0001 ,
		_w9452_,
		_w9453_,
		_w9946_
	);
	LUT2 #(
		.INIT('h4)
	) name5899 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9947_
	);
	LUT4 #(
		.INIT('hebd7)
	) name5900 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w9948_
	);
	LUT4 #(
		.INIT('hd7eb)
	) name5901 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w9949_
	);
	LUT3 #(
		.INIT('he4)
	) name5902 (
		_w9947_,
		_w9948_,
		_w9949_,
		_w9950_
	);
	LUT4 #(
		.INIT('h0180)
	) name5903 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w9951_
	);
	LUT4 #(
		.INIT('h0240)
	) name5904 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w9952_
	);
	LUT3 #(
		.INIT('h1b)
	) name5905 (
		_w9947_,
		_w9951_,
		_w9952_,
		_w9953_
	);
	LUT2 #(
		.INIT('h8)
	) name5906 (
		_w9950_,
		_w9953_,
		_w9954_
	);
	LUT4 #(
		.INIT('hebd7)
	) name5907 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w9955_
	);
	LUT4 #(
		.INIT('hd7eb)
	) name5908 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w9956_
	);
	LUT3 #(
		.INIT('he4)
	) name5909 (
		_w9947_,
		_w9955_,
		_w9956_,
		_w9957_
	);
	LUT4 #(
		.INIT('h0180)
	) name5910 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w9958_
	);
	LUT4 #(
		.INIT('h0240)
	) name5911 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w9959_
	);
	LUT3 #(
		.INIT('h1b)
	) name5912 (
		_w9947_,
		_w9958_,
		_w9959_,
		_w9960_
	);
	LUT2 #(
		.INIT('h8)
	) name5913 (
		_w9957_,
		_w9960_,
		_w9961_
	);
	LUT4 #(
		.INIT('h8000)
	) name5914 (
		_w9950_,
		_w9953_,
		_w9957_,
		_w9960_,
		_w9962_
	);
	LUT4 #(
		.INIT('hebd7)
	) name5915 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w9963_
	);
	LUT4 #(
		.INIT('hd7eb)
	) name5916 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w9964_
	);
	LUT3 #(
		.INIT('he4)
	) name5917 (
		_w9947_,
		_w9963_,
		_w9964_,
		_w9965_
	);
	LUT4 #(
		.INIT('h0180)
	) name5918 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w9966_
	);
	LUT4 #(
		.INIT('h0240)
	) name5919 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w9967_
	);
	LUT3 #(
		.INIT('h1b)
	) name5920 (
		_w9947_,
		_w9966_,
		_w9967_,
		_w9968_
	);
	LUT2 #(
		.INIT('h8)
	) name5921 (
		_w9965_,
		_w9968_,
		_w9969_
	);
	LUT3 #(
		.INIT('hb7)
	) name5922 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w9970_
	);
	LUT3 #(
		.INIT('h7b)
	) name5923 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w9971_
	);
	LUT3 #(
		.INIT('h10)
	) name5924 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w9972_
	);
	LUT4 #(
		.INIT('h5ba7)
	) name5925 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w9947_,
		_w9973_
	);
	LUT3 #(
		.INIT('h80)
	) name5926 (
		_w9962_,
		_w9969_,
		_w9973_,
		_w9974_
	);
	LUT4 #(
		.INIT('hebd7)
	) name5927 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w9975_
	);
	LUT4 #(
		.INIT('hd7eb)
	) name5928 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w9976_
	);
	LUT3 #(
		.INIT('he4)
	) name5929 (
		_w9947_,
		_w9975_,
		_w9976_,
		_w9977_
	);
	LUT4 #(
		.INIT('h0180)
	) name5930 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w9978_
	);
	LUT4 #(
		.INIT('h0240)
	) name5931 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w9979_
	);
	LUT3 #(
		.INIT('h1b)
	) name5932 (
		_w9947_,
		_w9978_,
		_w9979_,
		_w9980_
	);
	LUT2 #(
		.INIT('h8)
	) name5933 (
		_w9977_,
		_w9980_,
		_w9981_
	);
	LUT4 #(
		.INIT('hedb7)
	) name5934 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w9982_
	);
	LUT4 #(
		.INIT('hde7b)
	) name5935 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w9983_
	);
	LUT3 #(
		.INIT('he4)
	) name5936 (
		_w9947_,
		_w9982_,
		_w9983_,
		_w9984_
	);
	LUT4 #(
		.INIT('h0810)
	) name5937 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w9985_
	);
	LUT4 #(
		.INIT('h0420)
	) name5938 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w9986_
	);
	LUT3 #(
		.INIT('h1b)
	) name5939 (
		_w9947_,
		_w9985_,
		_w9986_,
		_w9987_
	);
	LUT2 #(
		.INIT('h8)
	) name5940 (
		_w9984_,
		_w9987_,
		_w9988_
	);
	LUT4 #(
		.INIT('h8000)
	) name5941 (
		_w9977_,
		_w9980_,
		_w9984_,
		_w9987_,
		_w9989_
	);
	LUT4 #(
		.INIT('hebd7)
	) name5942 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w9990_
	);
	LUT4 #(
		.INIT('hd7eb)
	) name5943 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w9991_
	);
	LUT3 #(
		.INIT('he4)
	) name5944 (
		_w9947_,
		_w9990_,
		_w9991_,
		_w9992_
	);
	LUT4 #(
		.INIT('h0180)
	) name5945 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w9993_
	);
	LUT4 #(
		.INIT('h0240)
	) name5946 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w9994_
	);
	LUT3 #(
		.INIT('h1b)
	) name5947 (
		_w9947_,
		_w9993_,
		_w9994_,
		_w9995_
	);
	LUT2 #(
		.INIT('h8)
	) name5948 (
		_w9992_,
		_w9995_,
		_w9996_
	);
	LUT2 #(
		.INIT('h8)
	) name5949 (
		_w9989_,
		_w9996_,
		_w9997_
	);
	LUT4 #(
		.INIT('ha820)
	) name5950 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 ,
		_w9998_
	);
	LUT4 #(
		.INIT('ha820)
	) name5951 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 ,
		_w9999_
	);
	LUT4 #(
		.INIT('h3120)
	) name5952 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9999_,
		_w9998_,
		_w10000_
	);
	LUT4 #(
		.INIT('hebd7)
	) name5953 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10001_
	);
	LUT4 #(
		.INIT('hd7eb)
	) name5954 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10002_
	);
	LUT3 #(
		.INIT('he4)
	) name5955 (
		_w9947_,
		_w10001_,
		_w10002_,
		_w10003_
	);
	LUT4 #(
		.INIT('h0180)
	) name5956 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10004_
	);
	LUT4 #(
		.INIT('h0240)
	) name5957 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10005_
	);
	LUT3 #(
		.INIT('h1b)
	) name5958 (
		_w9947_,
		_w10004_,
		_w10005_,
		_w10006_
	);
	LUT2 #(
		.INIT('h8)
	) name5959 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10007_
	);
	LUT3 #(
		.INIT('h80)
	) name5960 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10008_
	);
	LUT3 #(
		.INIT('h9f)
	) name5961 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w9947_,
		_w10007_,
		_w10009_
	);
	LUT3 #(
		.INIT('h80)
	) name5962 (
		_w10003_,
		_w10006_,
		_w10009_,
		_w10010_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5963 (
		_w10000_,
		_w10003_,
		_w10006_,
		_w10009_,
		_w10011_
	);
	LUT4 #(
		.INIT('h9555)
	) name5964 (
		_w10000_,
		_w10003_,
		_w10006_,
		_w10009_,
		_w10012_
	);
	LUT4 #(
		.INIT('h4800)
	) name5965 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10013_
	);
	LUT4 #(
		.INIT('ha820)
	) name5966 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 ,
		_w10014_
	);
	LUT4 #(
		.INIT('h3210)
	) name5967 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9999_,
		_w10014_,
		_w10015_
	);
	LUT4 #(
		.INIT('hf770)
	) name5968 (
		_w10003_,
		_w10006_,
		_w10013_,
		_w10015_,
		_w10016_
	);
	LUT4 #(
		.INIT('h7770)
	) name5969 (
		_w9989_,
		_w9996_,
		_w10012_,
		_w10016_,
		_w10017_
	);
	LUT4 #(
		.INIT('h0777)
	) name5970 (
		_w9977_,
		_w9980_,
		_w9984_,
		_w9987_,
		_w10018_
	);
	LUT2 #(
		.INIT('h4)
	) name5971 (
		_w9996_,
		_w10018_,
		_w10019_
	);
	LUT3 #(
		.INIT('h7e)
	) name5972 (
		_w9981_,
		_w9988_,
		_w9996_,
		_w10020_
	);
	LUT4 #(
		.INIT('hfd75)
	) name5973 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w6484_,
		_w6860_,
		_w10021_
	);
	LUT2 #(
		.INIT('h1)
	) name5974 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10021_,
		_w10022_
	);
	LUT3 #(
		.INIT('h12)
	) name5975 (
		_w10010_,
		_w10011_,
		_w10022_,
		_w10023_
	);
	LUT3 #(
		.INIT('he1)
	) name5976 (
		_w10000_,
		_w10010_,
		_w10022_,
		_w10024_
	);
	LUT3 #(
		.INIT('h69)
	) name5977 (
		_w10017_,
		_w10020_,
		_w10024_,
		_w10025_
	);
	LUT4 #(
		.INIT('h8778)
	) name5978 (
		_w10003_,
		_w10006_,
		_w10013_,
		_w10015_,
		_w10026_
	);
	LUT4 #(
		.INIT('h4800)
	) name5979 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10027_
	);
	LUT3 #(
		.INIT('h1b)
	) name5980 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w10004_,
		_w10005_,
		_w10028_
	);
	LUT4 #(
		.INIT('ha820)
	) name5981 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 ,
		_w10029_
	);
	LUT4 #(
		.INIT('h3210)
	) name5982 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10014_,
		_w10029_,
		_w10030_
	);
	LUT4 #(
		.INIT('hdf4c)
	) name5983 (
		_w10003_,
		_w10027_,
		_w10028_,
		_w10030_,
		_w10031_
	);
	LUT4 #(
		.INIT('h7707)
	) name5984 (
		_w9989_,
		_w9996_,
		_w10026_,
		_w10031_,
		_w10032_
	);
	LUT2 #(
		.INIT('h6)
	) name5985 (
		_w10012_,
		_w10016_,
		_w10033_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name5986 (
		_w9996_,
		_w10012_,
		_w10016_,
		_w10018_,
		_w10034_
	);
	LUT4 #(
		.INIT('h48ed)
	) name5987 (
		_w10020_,
		_w10032_,
		_w10033_,
		_w10034_,
		_w10035_
	);
	LUT2 #(
		.INIT('h2)
	) name5988 (
		_w10025_,
		_w10035_,
		_w10036_
	);
	LUT3 #(
		.INIT('h51)
	) name5989 (
		_w9974_,
		_w10025_,
		_w10035_,
		_w10037_
	);
	LUT4 #(
		.INIT('hfd75)
	) name5990 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w6145_,
		_w6484_,
		_w10038_
	);
	LUT2 #(
		.INIT('h1)
	) name5991 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10038_,
		_w10039_
	);
	LUT3 #(
		.INIT('h1a)
	) name5992 (
		_w10010_,
		_w10022_,
		_w10039_,
		_w10040_
	);
	LUT3 #(
		.INIT('h40)
	) name5993 (
		_w10010_,
		_w10022_,
		_w10038_,
		_w10041_
	);
	LUT4 #(
		.INIT('h0376)
	) name5994 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10010_,
		_w10022_,
		_w10038_,
		_w10042_
	);
	LUT4 #(
		.INIT('h32c8)
	) name5995 (
		_w9997_,
		_w10020_,
		_w10023_,
		_w10042_,
		_w10043_
	);
	LUT4 #(
		.INIT('hc936)
	) name5996 (
		_w9997_,
		_w10020_,
		_w10023_,
		_w10042_,
		_w10044_
	);
	LUT4 #(
		.INIT('haf23)
	) name5997 (
		_w9996_,
		_w10011_,
		_w10018_,
		_w10022_,
		_w10045_
	);
	LUT4 #(
		.INIT('h28eb)
	) name5998 (
		_w10017_,
		_w10020_,
		_w10024_,
		_w10045_,
		_w10046_
	);
	LUT2 #(
		.INIT('h9)
	) name5999 (
		_w10044_,
		_w10046_,
		_w10047_
	);
	LUT3 #(
		.INIT('h96)
	) name6000 (
		_w9974_,
		_w10044_,
		_w10046_,
		_w10048_
	);
	LUT3 #(
		.INIT('h4b)
	) name6001 (
		_w9974_,
		_w10036_,
		_w10047_,
		_w10049_
	);
	LUT3 #(
		.INIT('h69)
	) name6002 (
		_w10020_,
		_w10032_,
		_w10033_,
		_w10050_
	);
	LUT4 #(
		.INIT('h936c)
	) name6003 (
		_w10003_,
		_w10027_,
		_w10028_,
		_w10030_,
		_w10051_
	);
	LUT4 #(
		.INIT('h4800)
	) name6004 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10052_
	);
	LUT2 #(
		.INIT('h2)
	) name6005 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w10002_,
		_w10053_
	);
	LUT2 #(
		.INIT('h1)
	) name6006 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w10001_,
		_w10054_
	);
	LUT3 #(
		.INIT('h1b)
	) name6007 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w10004_,
		_w10005_,
		_w10055_
	);
	LUT3 #(
		.INIT('h10)
	) name6008 (
		_w10054_,
		_w10053_,
		_w10055_,
		_w10056_
	);
	LUT4 #(
		.INIT('h0100)
	) name6009 (
		_w10052_,
		_w10054_,
		_w10053_,
		_w10055_,
		_w10057_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6010 (
		_w10052_,
		_w10054_,
		_w10053_,
		_w10055_,
		_w10058_
	);
	LUT4 #(
		.INIT('ha820)
	) name6011 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 ,
		_w10059_
	);
	LUT4 #(
		.INIT('h3210)
	) name6012 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10029_,
		_w10059_,
		_w10060_
	);
	LUT3 #(
		.INIT('h54)
	) name6013 (
		_w10057_,
		_w10058_,
		_w10060_,
		_w10061_
	);
	LUT4 #(
		.INIT('h20a2)
	) name6014 (
		_w10051_,
		_w10052_,
		_w10056_,
		_w10060_,
		_w10062_
	);
	LUT2 #(
		.INIT('h9)
	) name6015 (
		_w10026_,
		_w10031_,
		_w10063_
	);
	LUT4 #(
		.INIT('h32c8)
	) name6016 (
		_w9997_,
		_w10020_,
		_w10062_,
		_w10063_,
		_w10064_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6017 (
		_w9996_,
		_w10018_,
		_w10026_,
		_w10031_,
		_w10065_
	);
	LUT3 #(
		.INIT('h90)
	) name6018 (
		_w10020_,
		_w10063_,
		_w10065_,
		_w10066_
	);
	LUT3 #(
		.INIT('ha8)
	) name6019 (
		_w10050_,
		_w10064_,
		_w10066_,
		_w10067_
	);
	LUT4 #(
		.INIT('h1115)
	) name6020 (
		_w9974_,
		_w10050_,
		_w10064_,
		_w10066_,
		_w10068_
	);
	LUT2 #(
		.INIT('h9)
	) name6021 (
		_w10025_,
		_w10035_,
		_w10069_
	);
	LUT3 #(
		.INIT('h69)
	) name6022 (
		_w9974_,
		_w10025_,
		_w10035_,
		_w10070_
	);
	LUT3 #(
		.INIT('h49)
	) name6023 (
		_w9974_,
		_w10025_,
		_w10035_,
		_w10071_
	);
	LUT3 #(
		.INIT('h0e)
	) name6024 (
		_w10068_,
		_w10070_,
		_w10071_,
		_w10072_
	);
	LUT2 #(
		.INIT('h9)
	) name6025 (
		_w10049_,
		_w10072_,
		_w10073_
	);
	LUT4 #(
		.INIT('hc936)
	) name6026 (
		_w9997_,
		_w10020_,
		_w10062_,
		_w10063_,
		_w10074_
	);
	LUT3 #(
		.INIT('h1b)
	) name6027 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9993_,
		_w9994_,
		_w10075_
	);
	LUT2 #(
		.INIT('h8)
	) name6028 (
		_w9992_,
		_w10075_,
		_w10076_
	);
	LUT3 #(
		.INIT('h32)
	) name6029 (
		_w9989_,
		_w10018_,
		_w10076_,
		_w10077_
	);
	LUT4 #(
		.INIT('h7888)
	) name6030 (
		_w9977_,
		_w9980_,
		_w9984_,
		_w9987_,
		_w10078_
	);
	LUT2 #(
		.INIT('h9)
	) name6031 (
		_w9996_,
		_w10078_,
		_w10079_
	);
	LUT4 #(
		.INIT('h8680)
	) name6032 (
		_w9981_,
		_w9988_,
		_w9996_,
		_w10076_,
		_w10080_
	);
	LUT4 #(
		.INIT('h5655)
	) name6033 (
		_w10052_,
		_w10054_,
		_w10053_,
		_w10055_,
		_w10081_
	);
	LUT2 #(
		.INIT('h9)
	) name6034 (
		_w10060_,
		_w10081_,
		_w10082_
	);
	LUT4 #(
		.INIT('ha820)
	) name6035 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 ,
		_w10083_
	);
	LUT4 #(
		.INIT('h3210)
	) name6036 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10059_,
		_w10083_,
		_w10084_
	);
	LUT2 #(
		.INIT('h2)
	) name6037 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w10002_,
		_w10085_
	);
	LUT2 #(
		.INIT('h1)
	) name6038 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w10001_,
		_w10086_
	);
	LUT3 #(
		.INIT('h1b)
	) name6039 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w10004_,
		_w10005_,
		_w10087_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6040 (
		_w10084_,
		_w10086_,
		_w10085_,
		_w10087_,
		_w10088_
	);
	LUT4 #(
		.INIT('h0100)
	) name6041 (
		_w10084_,
		_w10086_,
		_w10085_,
		_w10087_,
		_w10089_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name6042 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10090_
	);
	LUT3 #(
		.INIT('h54)
	) name6043 (
		_w10088_,
		_w10089_,
		_w10090_,
		_w10091_
	);
	LUT3 #(
		.INIT('h15)
	) name6044 (
		_w10080_,
		_w10082_,
		_w10091_,
		_w10092_
	);
	LUT4 #(
		.INIT('h4504)
	) name6045 (
		_w10051_,
		_w10052_,
		_w10056_,
		_w10060_,
		_w10093_
	);
	LUT4 #(
		.INIT('h6665)
	) name6046 (
		_w10051_,
		_w10057_,
		_w10058_,
		_w10060_,
		_w10094_
	);
	LUT2 #(
		.INIT('h9)
	) name6047 (
		_w10020_,
		_w10094_,
		_w10095_
	);
	LUT2 #(
		.INIT('h1)
	) name6048 (
		_w10019_,
		_w10093_,
		_w10096_
	);
	LUT4 #(
		.INIT('h4014)
	) name6049 (
		_w10019_,
		_w10020_,
		_w10051_,
		_w10061_,
		_w10097_
	);
	LUT4 #(
		.INIT('ha202)
	) name6050 (
		_w10074_,
		_w10092_,
		_w10095_,
		_w10096_,
		_w10098_
	);
	LUT3 #(
		.INIT('h56)
	) name6051 (
		_w10050_,
		_w10064_,
		_w10066_,
		_w10099_
	);
	LUT4 #(
		.INIT('h9994)
	) name6052 (
		_w9974_,
		_w10050_,
		_w10064_,
		_w10066_,
		_w10100_
	);
	LUT4 #(
		.INIT('h005b)
	) name6053 (
		_w9974_,
		_w10098_,
		_w10099_,
		_w10100_,
		_w10101_
	);
	LUT3 #(
		.INIT('h4b)
	) name6054 (
		_w9974_,
		_w10067_,
		_w10069_,
		_w10102_
	);
	LUT2 #(
		.INIT('h2)
	) name6055 (
		_w10101_,
		_w10102_,
		_w10103_
	);
	LUT2 #(
		.INIT('h4)
	) name6056 (
		_w10101_,
		_w10102_,
		_w10104_
	);
	LUT2 #(
		.INIT('h6)
	) name6057 (
		_w10092_,
		_w10095_,
		_w10105_
	);
	LUT2 #(
		.INIT('h2)
	) name6058 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9991_,
		_w10106_
	);
	LUT2 #(
		.INIT('h1)
	) name6059 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9990_,
		_w10107_
	);
	LUT3 #(
		.INIT('h1b)
	) name6060 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9993_,
		_w9994_,
		_w10108_
	);
	LUT3 #(
		.INIT('h10)
	) name6061 (
		_w10107_,
		_w10106_,
		_w10108_,
		_w10109_
	);
	LUT3 #(
		.INIT('h32)
	) name6062 (
		_w9989_,
		_w10018_,
		_w10109_,
		_w10110_
	);
	LUT2 #(
		.INIT('h9)
	) name6063 (
		_w10076_,
		_w10078_,
		_w10111_
	);
	LUT4 #(
		.INIT('h8680)
	) name6064 (
		_w9981_,
		_w9988_,
		_w10076_,
		_w10109_,
		_w10112_
	);
	LUT4 #(
		.INIT('h4800)
	) name6065 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10113_
	);
	LUT2 #(
		.INIT('h2)
	) name6066 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w10002_,
		_w10114_
	);
	LUT2 #(
		.INIT('h1)
	) name6067 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w10001_,
		_w10115_
	);
	LUT3 #(
		.INIT('h1b)
	) name6068 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w10004_,
		_w10005_,
		_w10116_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6069 (
		_w10113_,
		_w10115_,
		_w10114_,
		_w10116_,
		_w10117_
	);
	LUT4 #(
		.INIT('h0100)
	) name6070 (
		_w10113_,
		_w10115_,
		_w10114_,
		_w10116_,
		_w10118_
	);
	LUT4 #(
		.INIT('ha820)
	) name6071 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 ,
		_w10119_
	);
	LUT4 #(
		.INIT('h3210)
	) name6072 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10083_,
		_w10119_,
		_w10120_
	);
	LUT3 #(
		.INIT('h45)
	) name6073 (
		_w10117_,
		_w10118_,
		_w10120_,
		_w10121_
	);
	LUT4 #(
		.INIT('h5655)
	) name6074 (
		_w10084_,
		_w10086_,
		_w10085_,
		_w10087_,
		_w10122_
	);
	LUT2 #(
		.INIT('h9)
	) name6075 (
		_w10090_,
		_w10122_,
		_w10123_
	);
	LUT3 #(
		.INIT('h51)
	) name6076 (
		_w10112_,
		_w10121_,
		_w10123_,
		_w10124_
	);
	LUT4 #(
		.INIT('hc6c3)
	) name6077 (
		_w9989_,
		_w9996_,
		_w10018_,
		_w10076_,
		_w10125_
	);
	LUT3 #(
		.INIT('h96)
	) name6078 (
		_w10082_,
		_w10091_,
		_w10125_,
		_w10126_
	);
	LUT4 #(
		.INIT('h2990)
	) name6079 (
		_w10077_,
		_w10079_,
		_w10082_,
		_w10091_,
		_w10127_
	);
	LUT3 #(
		.INIT('h0b)
	) name6080 (
		_w10124_,
		_w10126_,
		_w10127_,
		_w10128_
	);
	LUT4 #(
		.INIT('h0454)
	) name6081 (
		_w10074_,
		_w10092_,
		_w10095_,
		_w10096_,
		_w10129_
	);
	LUT4 #(
		.INIT('h55a9)
	) name6082 (
		_w10074_,
		_w10092_,
		_w10095_,
		_w10097_,
		_w10130_
	);
	LUT4 #(
		.INIT('haa04)
	) name6083 (
		_w9974_,
		_w10105_,
		_w10128_,
		_w10130_,
		_w10131_
	);
	LUT4 #(
		.INIT('h04fb)
	) name6084 (
		_w9974_,
		_w10105_,
		_w10128_,
		_w10130_,
		_w10132_
	);
	LUT3 #(
		.INIT('h4b)
	) name6085 (
		_w9974_,
		_w10098_,
		_w10099_,
		_w10133_
	);
	LUT2 #(
		.INIT('h1)
	) name6086 (
		_w10132_,
		_w10133_,
		_w10134_
	);
	LUT2 #(
		.INIT('h9)
	) name6087 (
		_w10124_,
		_w10126_,
		_w10135_
	);
	LUT4 #(
		.INIT('h5655)
	) name6088 (
		_w10113_,
		_w10115_,
		_w10114_,
		_w10116_,
		_w10136_
	);
	LUT2 #(
		.INIT('h6)
	) name6089 (
		_w10120_,
		_w10136_,
		_w10137_
	);
	LUT4 #(
		.INIT('ha820)
	) name6090 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 ,
		_w10138_
	);
	LUT4 #(
		.INIT('h3210)
	) name6091 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10119_,
		_w10138_,
		_w10139_
	);
	LUT2 #(
		.INIT('h2)
	) name6092 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w10002_,
		_w10140_
	);
	LUT2 #(
		.INIT('h1)
	) name6093 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w10001_,
		_w10141_
	);
	LUT3 #(
		.INIT('h1b)
	) name6094 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w10004_,
		_w10005_,
		_w10142_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6095 (
		_w10139_,
		_w10141_,
		_w10140_,
		_w10142_,
		_w10143_
	);
	LUT4 #(
		.INIT('h0100)
	) name6096 (
		_w10139_,
		_w10141_,
		_w10140_,
		_w10142_,
		_w10144_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name6097 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10145_
	);
	LUT3 #(
		.INIT('h54)
	) name6098 (
		_w10143_,
		_w10144_,
		_w10145_,
		_w10146_
	);
	LUT2 #(
		.INIT('h2)
	) name6099 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9991_,
		_w10147_
	);
	LUT2 #(
		.INIT('h1)
	) name6100 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9990_,
		_w10148_
	);
	LUT3 #(
		.INIT('h1b)
	) name6101 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9993_,
		_w9994_,
		_w10149_
	);
	LUT3 #(
		.INIT('h10)
	) name6102 (
		_w10148_,
		_w10147_,
		_w10149_,
		_w10150_
	);
	LUT3 #(
		.INIT('h1b)
	) name6103 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9985_,
		_w9986_,
		_w10151_
	);
	LUT2 #(
		.INIT('h8)
	) name6104 (
		_w9984_,
		_w10151_,
		_w10152_
	);
	LUT3 #(
		.INIT('he8)
	) name6105 (
		_w9981_,
		_w10150_,
		_w10152_,
		_w10153_
	);
	LUT2 #(
		.INIT('h9)
	) name6106 (
		_w10078_,
		_w10109_,
		_w10154_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name6107 (
		_w10137_,
		_w10146_,
		_w10153_,
		_w10154_,
		_w10155_
	);
	LUT4 #(
		.INIT('hd2c3)
	) name6108 (
		_w9989_,
		_w10018_,
		_w10076_,
		_w10109_,
		_w10156_
	);
	LUT3 #(
		.INIT('h69)
	) name6109 (
		_w10121_,
		_w10123_,
		_w10156_,
		_w10157_
	);
	LUT4 #(
		.INIT('h9029)
	) name6110 (
		_w10110_,
		_w10111_,
		_w10121_,
		_w10123_,
		_w10158_
	);
	LUT3 #(
		.INIT('h0b)
	) name6111 (
		_w10155_,
		_w10157_,
		_w10158_,
		_w10159_
	);
	LUT2 #(
		.INIT('h2)
	) name6112 (
		_w10135_,
		_w10159_,
		_w10160_
	);
	LUT3 #(
		.INIT('h51)
	) name6113 (
		_w9974_,
		_w10135_,
		_w10159_,
		_w10161_
	);
	LUT2 #(
		.INIT('h9)
	) name6114 (
		_w10105_,
		_w10128_,
		_w10162_
	);
	LUT3 #(
		.INIT('h69)
	) name6115 (
		_w9974_,
		_w10105_,
		_w10128_,
		_w10163_
	);
	LUT3 #(
		.INIT('h49)
	) name6116 (
		_w9974_,
		_w10105_,
		_w10128_,
		_w10164_
	);
	LUT3 #(
		.INIT('h0e)
	) name6117 (
		_w10161_,
		_w10163_,
		_w10164_,
		_w10165_
	);
	LUT3 #(
		.INIT('h09)
	) name6118 (
		_w9974_,
		_w10098_,
		_w10129_,
		_w10166_
	);
	LUT3 #(
		.INIT('hc8)
	) name6119 (
		_w10131_,
		_w10133_,
		_w10166_,
		_w10167_
	);
	LUT3 #(
		.INIT('h51)
	) name6120 (
		_w10134_,
		_w10165_,
		_w10167_,
		_w10168_
	);
	LUT2 #(
		.INIT('h2)
	) name6121 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9956_,
		_w10169_
	);
	LUT2 #(
		.INIT('h1)
	) name6122 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9955_,
		_w10170_
	);
	LUT3 #(
		.INIT('h1b)
	) name6123 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9958_,
		_w9959_,
		_w10171_
	);
	LUT3 #(
		.INIT('h10)
	) name6124 (
		_w10170_,
		_w10169_,
		_w10171_,
		_w10172_
	);
	LUT2 #(
		.INIT('h2)
	) name6125 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9949_,
		_w10173_
	);
	LUT2 #(
		.INIT('h1)
	) name6126 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9948_,
		_w10174_
	);
	LUT3 #(
		.INIT('h1b)
	) name6127 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9951_,
		_w9952_,
		_w10175_
	);
	LUT3 #(
		.INIT('h10)
	) name6128 (
		_w10174_,
		_w10173_,
		_w10175_,
		_w10176_
	);
	LUT2 #(
		.INIT('h2)
	) name6129 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9956_,
		_w10177_
	);
	LUT2 #(
		.INIT('h1)
	) name6130 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9955_,
		_w10178_
	);
	LUT3 #(
		.INIT('h1b)
	) name6131 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9958_,
		_w9959_,
		_w10179_
	);
	LUT3 #(
		.INIT('h10)
	) name6132 (
		_w10178_,
		_w10177_,
		_w10179_,
		_w10180_
	);
	LUT3 #(
		.INIT('he4)
	) name6133 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9963_,
		_w9964_,
		_w10181_
	);
	LUT2 #(
		.INIT('h2)
	) name6134 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9949_,
		_w10182_
	);
	LUT2 #(
		.INIT('h1)
	) name6135 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9948_,
		_w10183_
	);
	LUT3 #(
		.INIT('h1b)
	) name6136 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9951_,
		_w9952_,
		_w10184_
	);
	LUT4 #(
		.INIT('h5455)
	) name6137 (
		_w10181_,
		_w10183_,
		_w10182_,
		_w10184_,
		_w10185_
	);
	LUT4 #(
		.INIT('h0200)
	) name6138 (
		_w10181_,
		_w10183_,
		_w10182_,
		_w10184_,
		_w10186_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6139 (
		_w10181_,
		_w10183_,
		_w10182_,
		_w10184_,
		_w10187_
	);
	LUT4 #(
		.INIT('h54a8)
	) name6140 (
		_w10180_,
		_w10172_,
		_w10176_,
		_w10187_,
		_w10188_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name6141 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w7668_,
		_w8023_,
		_w10189_
	);
	LUT4 #(
		.INIT('h8040)
	) name6142 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10190_
	);
	LUT4 #(
		.INIT('h1020)
	) name6143 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10191_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6144 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10192_
	);
	LUT3 #(
		.INIT('h10)
	) name6145 (
		_w10191_,
		_w10190_,
		_w10192_,
		_w10193_
	);
	LUT4 #(
		.INIT('h04cd)
	) name6146 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9958_,
		_w10189_,
		_w10193_,
		_w10194_
	);
	LUT4 #(
		.INIT('h8040)
	) name6147 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10195_
	);
	LUT4 #(
		.INIT('h1020)
	) name6148 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10196_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6149 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10197_
	);
	LUT3 #(
		.INIT('h10)
	) name6150 (
		_w10196_,
		_w10195_,
		_w10197_,
		_w10198_
	);
	LUT4 #(
		.INIT('hfd75)
	) name6151 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w7888_,
		_w8023_,
		_w10199_
	);
	LUT4 #(
		.INIT('hc936)
	) name6152 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9963_,
		_w10199_,
		_w10198_,
		_w10200_
	);
	LUT2 #(
		.INIT('h4)
	) name6153 (
		_w10194_,
		_w10200_,
		_w10201_
	);
	LUT2 #(
		.INIT('h1)
	) name6154 (
		_w10188_,
		_w10201_,
		_w10202_
	);
	LUT3 #(
		.INIT('h54)
	) name6155 (
		_w10185_,
		_w10186_,
		_w10180_,
		_w10203_
	);
	LUT2 #(
		.INIT('h2)
	) name6156 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9964_,
		_w10204_
	);
	LUT2 #(
		.INIT('h1)
	) name6157 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9963_,
		_w10205_
	);
	LUT3 #(
		.INIT('h1b)
	) name6158 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9966_,
		_w9967_,
		_w10206_
	);
	LUT3 #(
		.INIT('h10)
	) name6159 (
		_w10205_,
		_w10204_,
		_w10206_,
		_w10207_
	);
	LUT2 #(
		.INIT('h2)
	) name6160 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9949_,
		_w10208_
	);
	LUT2 #(
		.INIT('h1)
	) name6161 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9948_,
		_w10209_
	);
	LUT3 #(
		.INIT('h1b)
	) name6162 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9951_,
		_w9952_,
		_w10210_
	);
	LUT3 #(
		.INIT('h10)
	) name6163 (
		_w10209_,
		_w10208_,
		_w10210_,
		_w10211_
	);
	LUT2 #(
		.INIT('h2)
	) name6164 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9956_,
		_w10212_
	);
	LUT2 #(
		.INIT('h1)
	) name6165 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9955_,
		_w10213_
	);
	LUT3 #(
		.INIT('h1b)
	) name6166 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9958_,
		_w9959_,
		_w10214_
	);
	LUT3 #(
		.INIT('h10)
	) name6167 (
		_w10213_,
		_w10212_,
		_w10214_,
		_w10215_
	);
	LUT3 #(
		.INIT('h69)
	) name6168 (
		_w10211_,
		_w10215_,
		_w10207_,
		_w10216_
	);
	LUT4 #(
		.INIT('hfd75)
	) name6169 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w7549_,
		_w7888_,
		_w10217_
	);
	LUT4 #(
		.INIT('h8040)
	) name6170 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10218_
	);
	LUT4 #(
		.INIT('h1020)
	) name6171 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10219_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6172 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10220_
	);
	LUT4 #(
		.INIT('h0100)
	) name6173 (
		_w9966_,
		_w10219_,
		_w10218_,
		_w10220_,
		_w10221_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6174 (
		_w9966_,
		_w10219_,
		_w10218_,
		_w10220_,
		_w10222_
	);
	LUT4 #(
		.INIT('h5655)
	) name6175 (
		_w9966_,
		_w10219_,
		_w10218_,
		_w10220_,
		_w10223_
	);
	LUT3 #(
		.INIT('he1)
	) name6176 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10217_,
		_w10223_,
		_w10224_
	);
	LUT4 #(
		.INIT('hfec8)
	) name6177 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9963_,
		_w10199_,
		_w10198_,
		_w10225_
	);
	LUT2 #(
		.INIT('h4)
	) name6178 (
		_w10224_,
		_w10225_,
		_w10226_
	);
	LUT2 #(
		.INIT('h2)
	) name6179 (
		_w10224_,
		_w10225_,
		_w10227_
	);
	LUT2 #(
		.INIT('h9)
	) name6180 (
		_w10224_,
		_w10225_,
		_w10228_
	);
	LUT3 #(
		.INIT('h96)
	) name6181 (
		_w10203_,
		_w10216_,
		_w10228_,
		_w10229_
	);
	LUT2 #(
		.INIT('h6)
	) name6182 (
		_w10202_,
		_w10229_,
		_w10230_
	);
	LUT3 #(
		.INIT('he4)
	) name6183 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9955_,
		_w9956_,
		_w10231_
	);
	LUT2 #(
		.INIT('h2)
	) name6184 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9949_,
		_w10232_
	);
	LUT2 #(
		.INIT('h1)
	) name6185 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9948_,
		_w10233_
	);
	LUT3 #(
		.INIT('h1b)
	) name6186 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9951_,
		_w9952_,
		_w10234_
	);
	LUT4 #(
		.INIT('h5455)
	) name6187 (
		_w10231_,
		_w10233_,
		_w10232_,
		_w10234_,
		_w10235_
	);
	LUT2 #(
		.INIT('h6)
	) name6188 (
		_w10172_,
		_w10176_,
		_w10236_
	);
	LUT3 #(
		.INIT('h09)
	) name6189 (
		_w10172_,
		_w10176_,
		_w10235_,
		_w10237_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name6190 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w7342_,
		_w7668_,
		_w10238_
	);
	LUT4 #(
		.INIT('h8040)
	) name6191 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10239_
	);
	LUT4 #(
		.INIT('h1020)
	) name6192 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10240_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6193 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10241_
	);
	LUT3 #(
		.INIT('h10)
	) name6194 (
		_w10240_,
		_w10239_,
		_w10241_,
		_w10242_
	);
	LUT4 #(
		.INIT('hfec8)
	) name6195 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9955_,
		_w10238_,
		_w10242_,
		_w10243_
	);
	LUT4 #(
		.INIT('h36c9)
	) name6196 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9958_,
		_w10189_,
		_w10193_,
		_w10244_
	);
	LUT2 #(
		.INIT('h8)
	) name6197 (
		_w10243_,
		_w10244_,
		_w10245_
	);
	LUT4 #(
		.INIT('h0201)
	) name6198 (
		_w10180_,
		_w10172_,
		_w10176_,
		_w10187_,
		_w10246_
	);
	LUT4 #(
		.INIT('ha956)
	) name6199 (
		_w10180_,
		_w10172_,
		_w10176_,
		_w10187_,
		_w10247_
	);
	LUT2 #(
		.INIT('h2)
	) name6200 (
		_w10194_,
		_w10200_,
		_w10248_
	);
	LUT2 #(
		.INIT('h9)
	) name6201 (
		_w10194_,
		_w10200_,
		_w10249_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name6202 (
		_w10237_,
		_w10245_,
		_w10247_,
		_w10249_,
		_w10250_
	);
	LUT4 #(
		.INIT('h0012)
	) name6203 (
		_w10201_,
		_w10246_,
		_w10247_,
		_w10248_,
		_w10251_
	);
	LUT2 #(
		.INIT('h1)
	) name6204 (
		_w10250_,
		_w10251_,
		_w10252_
	);
	LUT4 #(
		.INIT('h0009)
	) name6205 (
		_w10202_,
		_w10229_,
		_w10250_,
		_w10251_,
		_w10253_
	);
	LUT4 #(
		.INIT('h6660)
	) name6206 (
		_w10202_,
		_w10229_,
		_w10250_,
		_w10251_,
		_w10254_
	);
	LUT4 #(
		.INIT('h9996)
	) name6207 (
		_w10202_,
		_w10229_,
		_w10250_,
		_w10251_,
		_w10255_
	);
	LUT4 #(
		.INIT('he11e)
	) name6208 (
		_w10237_,
		_w10245_,
		_w10247_,
		_w10249_,
		_w10256_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name6209 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w6141_,
		_w7342_,
		_w10257_
	);
	LUT4 #(
		.INIT('h1020)
	) name6210 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10258_
	);
	LUT4 #(
		.INIT('h8040)
	) name6211 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10259_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6212 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10260_
	);
	LUT3 #(
		.INIT('h10)
	) name6213 (
		_w10259_,
		_w10258_,
		_w10260_,
		_w10261_
	);
	LUT4 #(
		.INIT('h04cd)
	) name6214 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9951_,
		_w10257_,
		_w10261_,
		_w10262_
	);
	LUT4 #(
		.INIT('h36c9)
	) name6215 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9955_,
		_w10238_,
		_w10242_,
		_w10263_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6216 (
		_w10231_,
		_w10233_,
		_w10232_,
		_w10234_,
		_w10264_
	);
	LUT3 #(
		.INIT('he0)
	) name6217 (
		_w10262_,
		_w10263_,
		_w10264_,
		_w10265_
	);
	LUT2 #(
		.INIT('h1)
	) name6218 (
		_w10243_,
		_w10244_,
		_w10266_
	);
	LUT2 #(
		.INIT('h6)
	) name6219 (
		_w10243_,
		_w10244_,
		_w10267_
	);
	LUT3 #(
		.INIT('h96)
	) name6220 (
		_w10172_,
		_w10176_,
		_w10235_,
		_w10268_
	);
	LUT3 #(
		.INIT('h14)
	) name6221 (
		_w10265_,
		_w10267_,
		_w10268_,
		_w10269_
	);
	LUT4 #(
		.INIT('h0601)
	) name6222 (
		_w10235_,
		_w10236_,
		_w10266_,
		_w10267_,
		_w10270_
	);
	LUT3 #(
		.INIT('h01)
	) name6223 (
		_w10256_,
		_w10269_,
		_w10270_,
		_w10271_
	);
	LUT3 #(
		.INIT('ha8)
	) name6224 (
		_w10256_,
		_w10269_,
		_w10270_,
		_w10272_
	);
	LUT4 #(
		.INIT('hfd75)
	) name6225 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w6141_,
		_w6481_,
		_w10273_
	);
	LUT4 #(
		.INIT('h8040)
	) name6226 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10274_
	);
	LUT4 #(
		.INIT('h1020)
	) name6227 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10275_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6228 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10276_
	);
	LUT3 #(
		.INIT('h10)
	) name6229 (
		_w10275_,
		_w10274_,
		_w10276_,
		_w10277_
	);
	LUT4 #(
		.INIT('h0137)
	) name6230 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9948_,
		_w10273_,
		_w10277_,
		_w10278_
	);
	LUT4 #(
		.INIT('h36c9)
	) name6231 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9951_,
		_w10257_,
		_w10261_,
		_w10279_
	);
	LUT2 #(
		.INIT('h2)
	) name6232 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9949_,
		_w10280_
	);
	LUT2 #(
		.INIT('h1)
	) name6233 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9948_,
		_w10281_
	);
	LUT3 #(
		.INIT('h1b)
	) name6234 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9951_,
		_w9952_,
		_w10282_
	);
	LUT3 #(
		.INIT('h10)
	) name6235 (
		_w10281_,
		_w10280_,
		_w10282_,
		_w10283_
	);
	LUT3 #(
		.INIT('h0b)
	) name6236 (
		_w10278_,
		_w10279_,
		_w10283_,
		_w10284_
	);
	LUT3 #(
		.INIT('h96)
	) name6237 (
		_w10262_,
		_w10263_,
		_w10264_,
		_w10285_
	);
	LUT3 #(
		.INIT('h61)
	) name6238 (
		_w10262_,
		_w10263_,
		_w10264_,
		_w10286_
	);
	LUT3 #(
		.INIT('h0b)
	) name6239 (
		_w10284_,
		_w10285_,
		_w10286_,
		_w10287_
	);
	LUT3 #(
		.INIT('h69)
	) name6240 (
		_w10265_,
		_w10267_,
		_w10268_,
		_w10288_
	);
	LUT2 #(
		.INIT('h2)
	) name6241 (
		_w10287_,
		_w10288_,
		_w10289_
	);
	LUT2 #(
		.INIT('h9)
	) name6242 (
		_w10287_,
		_w10288_,
		_w10290_
	);
	LUT2 #(
		.INIT('h9)
	) name6243 (
		_w10284_,
		_w10285_,
		_w10291_
	);
	LUT4 #(
		.INIT('hfd75)
	) name6244 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w6481_,
		_w6864_,
		_w10292_
	);
	LUT4 #(
		.INIT('h8040)
	) name6245 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10293_
	);
	LUT4 #(
		.INIT('h1020)
	) name6246 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10294_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6247 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10295_
	);
	LUT3 #(
		.INIT('h10)
	) name6248 (
		_w10294_,
		_w10293_,
		_w10295_,
		_w10296_
	);
	LUT4 #(
		.INIT('hfb32)
	) name6249 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9972_,
		_w10292_,
		_w10296_,
		_w10297_
	);
	LUT4 #(
		.INIT('hc936)
	) name6250 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9948_,
		_w10273_,
		_w10277_,
		_w10298_
	);
	LUT3 #(
		.INIT('he4)
	) name6251 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9948_,
		_w9949_,
		_w10299_
	);
	LUT3 #(
		.INIT('h07)
	) name6252 (
		_w10297_,
		_w10298_,
		_w10299_,
		_w10300_
	);
	LUT3 #(
		.INIT('h96)
	) name6253 (
		_w10278_,
		_w10279_,
		_w10283_,
		_w10301_
	);
	LUT3 #(
		.INIT('h49)
	) name6254 (
		_w10278_,
		_w10279_,
		_w10283_,
		_w10302_
	);
	LUT3 #(
		.INIT('h0b)
	) name6255 (
		_w10300_,
		_w10301_,
		_w10302_,
		_w10303_
	);
	LUT2 #(
		.INIT('h4)
	) name6256 (
		_w10291_,
		_w10303_,
		_w10304_
	);
	LUT2 #(
		.INIT('h9)
	) name6257 (
		_w10291_,
		_w10303_,
		_w10305_
	);
	LUT4 #(
		.INIT('hc936)
	) name6258 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9972_,
		_w10292_,
		_w10296_,
		_w10306_
	);
	LUT4 #(
		.INIT('h1020)
	) name6259 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10307_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name6260 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w5869_,
		_w6864_,
		_w10308_
	);
	LUT4 #(
		.INIT('h2f1f)
	) name6261 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10309_
	);
	LUT4 #(
		.INIT('h3332)
	) name6262 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10307_,
		_w10308_,
		_w10309_,
		_w10310_
	);
	LUT2 #(
		.INIT('h2)
	) name6263 (
		_w10306_,
		_w10310_,
		_w10311_
	);
	LUT3 #(
		.INIT('h69)
	) name6264 (
		_w10297_,
		_w10298_,
		_w10299_,
		_w10312_
	);
	LUT2 #(
		.INIT('h8)
	) name6265 (
		_w10311_,
		_w10312_,
		_w10313_
	);
	LUT3 #(
		.INIT('h10)
	) name6266 (
		_w10297_,
		_w10298_,
		_w10299_,
		_w10314_
	);
	LUT3 #(
		.INIT('h09)
	) name6267 (
		_w10300_,
		_w10301_,
		_w10314_,
		_w10315_
	);
	LUT2 #(
		.INIT('h8)
	) name6268 (
		_w10301_,
		_w10314_,
		_w10316_
	);
	LUT3 #(
		.INIT('h0d)
	) name6269 (
		_w10313_,
		_w10315_,
		_w10316_,
		_w10317_
	);
	LUT4 #(
		.INIT('h20a2)
	) name6270 (
		_w10290_,
		_w10291_,
		_w10303_,
		_w10317_,
		_w10318_
	);
	LUT4 #(
		.INIT('h4445)
	) name6271 (
		_w10271_,
		_w10272_,
		_w10289_,
		_w10318_,
		_w10319_
	);
	LUT3 #(
		.INIT('h54)
	) name6272 (
		_w10253_,
		_w10254_,
		_w10319_,
		_w10320_
	);
	LUT3 #(
		.INIT('h0d)
	) name6273 (
		_w10203_,
		_w10216_,
		_w10226_,
		_w10321_
	);
	LUT3 #(
		.INIT('he8)
	) name6274 (
		_w10211_,
		_w10215_,
		_w10207_,
		_w10322_
	);
	LUT2 #(
		.INIT('h2)
	) name6275 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9964_,
		_w10323_
	);
	LUT2 #(
		.INIT('h1)
	) name6276 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9963_,
		_w10324_
	);
	LUT3 #(
		.INIT('h1b)
	) name6277 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9966_,
		_w9967_,
		_w10325_
	);
	LUT3 #(
		.INIT('h10)
	) name6278 (
		_w10324_,
		_w10323_,
		_w10325_,
		_w10326_
	);
	LUT2 #(
		.INIT('h2)
	) name6279 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9949_,
		_w10327_
	);
	LUT2 #(
		.INIT('h1)
	) name6280 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9948_,
		_w10328_
	);
	LUT3 #(
		.INIT('h1b)
	) name6281 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9951_,
		_w9952_,
		_w10329_
	);
	LUT3 #(
		.INIT('h10)
	) name6282 (
		_w10328_,
		_w10327_,
		_w10329_,
		_w10330_
	);
	LUT2 #(
		.INIT('h2)
	) name6283 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9956_,
		_w10331_
	);
	LUT2 #(
		.INIT('h1)
	) name6284 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9955_,
		_w10332_
	);
	LUT3 #(
		.INIT('h1b)
	) name6285 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9958_,
		_w9959_,
		_w10333_
	);
	LUT3 #(
		.INIT('h10)
	) name6286 (
		_w10332_,
		_w10331_,
		_w10333_,
		_w10334_
	);
	LUT3 #(
		.INIT('h69)
	) name6287 (
		_w10330_,
		_w10334_,
		_w10326_,
		_w10335_
	);
	LUT4 #(
		.INIT('hfd75)
	) name6288 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w7213_,
		_w7549_,
		_w10336_
	);
	LUT4 #(
		.INIT('h8040)
	) name6289 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10337_
	);
	LUT4 #(
		.INIT('h1020)
	) name6290 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10338_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6291 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10339_
	);
	LUT3 #(
		.INIT('h10)
	) name6292 (
		_w10338_,
		_w10337_,
		_w10339_,
		_w10340_
	);
	LUT4 #(
		.INIT('h36c9)
	) name6293 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9975_,
		_w10336_,
		_w10340_,
		_w10341_
	);
	LUT4 #(
		.INIT('h3301)
	) name6294 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10221_,
		_w10217_,
		_w10222_,
		_w10342_
	);
	LUT2 #(
		.INIT('h1)
	) name6295 (
		_w10341_,
		_w10342_,
		_w10343_
	);
	LUT2 #(
		.INIT('h8)
	) name6296 (
		_w10341_,
		_w10342_,
		_w10344_
	);
	LUT2 #(
		.INIT('h6)
	) name6297 (
		_w10341_,
		_w10342_,
		_w10345_
	);
	LUT3 #(
		.INIT('h69)
	) name6298 (
		_w10322_,
		_w10335_,
		_w10345_,
		_w10346_
	);
	LUT2 #(
		.INIT('h9)
	) name6299 (
		_w10321_,
		_w10346_,
		_w10347_
	);
	LUT4 #(
		.INIT('h0029)
	) name6300 (
		_w10203_,
		_w10216_,
		_w10226_,
		_w10227_,
		_w10348_
	);
	LUT3 #(
		.INIT('h0e)
	) name6301 (
		_w10202_,
		_w10229_,
		_w10348_,
		_w10349_
	);
	LUT3 #(
		.INIT('he4)
	) name6302 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9975_,
		_w9976_,
		_w10350_
	);
	LUT3 #(
		.INIT('h96)
	) name6303 (
		_w10347_,
		_w10349_,
		_w10350_,
		_w10351_
	);
	LUT4 #(
		.INIT('h4d00)
	) name6304 (
		_w10230_,
		_w10252_,
		_w10319_,
		_w10351_,
		_w10352_
	);
	LUT3 #(
		.INIT('h0d)
	) name6305 (
		_w10347_,
		_w10349_,
		_w10350_,
		_w10353_
	);
	LUT2 #(
		.INIT('h2)
	) name6306 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9976_,
		_w10354_
	);
	LUT2 #(
		.INIT('h1)
	) name6307 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9975_,
		_w10355_
	);
	LUT3 #(
		.INIT('h1b)
	) name6308 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9978_,
		_w9979_,
		_w10356_
	);
	LUT3 #(
		.INIT('h10)
	) name6309 (
		_w10355_,
		_w10354_,
		_w10356_,
		_w10357_
	);
	LUT3 #(
		.INIT('h0d)
	) name6310 (
		_w10322_,
		_w10335_,
		_w10343_,
		_w10358_
	);
	LUT3 #(
		.INIT('he8)
	) name6311 (
		_w10330_,
		_w10334_,
		_w10326_,
		_w10359_
	);
	LUT2 #(
		.INIT('h2)
	) name6312 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9964_,
		_w10360_
	);
	LUT2 #(
		.INIT('h1)
	) name6313 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9963_,
		_w10361_
	);
	LUT3 #(
		.INIT('h1b)
	) name6314 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9966_,
		_w9967_,
		_w10362_
	);
	LUT3 #(
		.INIT('h10)
	) name6315 (
		_w10361_,
		_w10360_,
		_w10362_,
		_w10363_
	);
	LUT2 #(
		.INIT('h2)
	) name6316 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9956_,
		_w10364_
	);
	LUT2 #(
		.INIT('h1)
	) name6317 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9955_,
		_w10365_
	);
	LUT3 #(
		.INIT('h1b)
	) name6318 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9958_,
		_w9959_,
		_w10366_
	);
	LUT3 #(
		.INIT('h10)
	) name6319 (
		_w10365_,
		_w10364_,
		_w10366_,
		_w10367_
	);
	LUT2 #(
		.INIT('h2)
	) name6320 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9949_,
		_w10368_
	);
	LUT2 #(
		.INIT('h1)
	) name6321 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9948_,
		_w10369_
	);
	LUT3 #(
		.INIT('h1b)
	) name6322 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9951_,
		_w9952_,
		_w10370_
	);
	LUT3 #(
		.INIT('h10)
	) name6323 (
		_w10369_,
		_w10368_,
		_w10370_,
		_w10371_
	);
	LUT3 #(
		.INIT('h69)
	) name6324 (
		_w10367_,
		_w10371_,
		_w10363_,
		_w10372_
	);
	LUT4 #(
		.INIT('h0137)
	) name6325 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9975_,
		_w10336_,
		_w10340_,
		_w10373_
	);
	LUT4 #(
		.INIT('hfd75)
	) name6326 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w6011_,
		_w7213_,
		_w10374_
	);
	LUT4 #(
		.INIT('h8040)
	) name6327 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10375_
	);
	LUT4 #(
		.INIT('h1020)
	) name6328 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10376_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6329 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10377_
	);
	LUT3 #(
		.INIT('h10)
	) name6330 (
		_w10376_,
		_w10375_,
		_w10377_,
		_w10378_
	);
	LUT4 #(
		.INIT('hc936)
	) name6331 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9978_,
		_w10374_,
		_w10378_,
		_w10379_
	);
	LUT2 #(
		.INIT('h1)
	) name6332 (
		_w10373_,
		_w10379_,
		_w10380_
	);
	LUT2 #(
		.INIT('h8)
	) name6333 (
		_w10373_,
		_w10379_,
		_w10381_
	);
	LUT2 #(
		.INIT('h6)
	) name6334 (
		_w10373_,
		_w10379_,
		_w10382_
	);
	LUT3 #(
		.INIT('h69)
	) name6335 (
		_w10359_,
		_w10372_,
		_w10382_,
		_w10383_
	);
	LUT2 #(
		.INIT('h9)
	) name6336 (
		_w10358_,
		_w10383_,
		_w10384_
	);
	LUT4 #(
		.INIT('h0029)
	) name6337 (
		_w10322_,
		_w10335_,
		_w10343_,
		_w10344_,
		_w10385_
	);
	LUT3 #(
		.INIT('h0b)
	) name6338 (
		_w10321_,
		_w10346_,
		_w10385_,
		_w10386_
	);
	LUT3 #(
		.INIT('h96)
	) name6339 (
		_w10384_,
		_w10386_,
		_w10357_,
		_w10387_
	);
	LUT3 #(
		.INIT('h29)
	) name6340 (
		_w10384_,
		_w10386_,
		_w10357_,
		_w10388_
	);
	LUT3 #(
		.INIT('h0b)
	) name6341 (
		_w10353_,
		_w10387_,
		_w10388_,
		_w10389_
	);
	LUT3 #(
		.INIT('h0d)
	) name6342 (
		_w10384_,
		_w10386_,
		_w10357_,
		_w10390_
	);
	LUT3 #(
		.INIT('he4)
	) name6343 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9982_,
		_w9983_,
		_w10391_
	);
	LUT2 #(
		.INIT('h2)
	) name6344 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9976_,
		_w10392_
	);
	LUT2 #(
		.INIT('h1)
	) name6345 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9975_,
		_w10393_
	);
	LUT3 #(
		.INIT('h1b)
	) name6346 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9978_,
		_w9979_,
		_w10394_
	);
	LUT4 #(
		.INIT('h5455)
	) name6347 (
		_w10391_,
		_w10393_,
		_w10392_,
		_w10394_,
		_w10395_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6348 (
		_w10391_,
		_w10393_,
		_w10392_,
		_w10394_,
		_w10396_
	);
	LUT3 #(
		.INIT('h0d)
	) name6349 (
		_w10359_,
		_w10372_,
		_w10380_,
		_w10397_
	);
	LUT3 #(
		.INIT('he8)
	) name6350 (
		_w10367_,
		_w10371_,
		_w10363_,
		_w10398_
	);
	LUT2 #(
		.INIT('h2)
	) name6351 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9964_,
		_w10399_
	);
	LUT2 #(
		.INIT('h1)
	) name6352 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9963_,
		_w10400_
	);
	LUT3 #(
		.INIT('h1b)
	) name6353 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9966_,
		_w9967_,
		_w10401_
	);
	LUT3 #(
		.INIT('h10)
	) name6354 (
		_w10400_,
		_w10399_,
		_w10401_,
		_w10402_
	);
	LUT2 #(
		.INIT('h2)
	) name6355 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9956_,
		_w10403_
	);
	LUT2 #(
		.INIT('h1)
	) name6356 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9955_,
		_w10404_
	);
	LUT3 #(
		.INIT('h1b)
	) name6357 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9958_,
		_w9959_,
		_w10405_
	);
	LUT3 #(
		.INIT('h10)
	) name6358 (
		_w10404_,
		_w10403_,
		_w10405_,
		_w10406_
	);
	LUT2 #(
		.INIT('h2)
	) name6359 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9949_,
		_w10407_
	);
	LUT2 #(
		.INIT('h1)
	) name6360 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9948_,
		_w10408_
	);
	LUT3 #(
		.INIT('h1b)
	) name6361 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9951_,
		_w9952_,
		_w10409_
	);
	LUT3 #(
		.INIT('h10)
	) name6362 (
		_w10408_,
		_w10407_,
		_w10409_,
		_w10410_
	);
	LUT3 #(
		.INIT('h69)
	) name6363 (
		_w10406_,
		_w10410_,
		_w10402_,
		_w10411_
	);
	LUT4 #(
		.INIT('h04cd)
	) name6364 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9978_,
		_w10374_,
		_w10378_,
		_w10412_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name6365 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w6011_,
		_w6335_,
		_w10413_
	);
	LUT4 #(
		.INIT('h8040)
	) name6366 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10414_
	);
	LUT4 #(
		.INIT('h1020)
	) name6367 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10415_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6368 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10416_
	);
	LUT3 #(
		.INIT('h10)
	) name6369 (
		_w10415_,
		_w10414_,
		_w10416_,
		_w10417_
	);
	LUT4 #(
		.INIT('h36c9)
	) name6370 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9982_,
		_w10413_,
		_w10417_,
		_w10418_
	);
	LUT2 #(
		.INIT('h1)
	) name6371 (
		_w10412_,
		_w10418_,
		_w10419_
	);
	LUT2 #(
		.INIT('h8)
	) name6372 (
		_w10412_,
		_w10418_,
		_w10420_
	);
	LUT2 #(
		.INIT('h6)
	) name6373 (
		_w10412_,
		_w10418_,
		_w10421_
	);
	LUT3 #(
		.INIT('h69)
	) name6374 (
		_w10398_,
		_w10411_,
		_w10421_,
		_w10422_
	);
	LUT2 #(
		.INIT('h9)
	) name6375 (
		_w10397_,
		_w10422_,
		_w10423_
	);
	LUT4 #(
		.INIT('h0029)
	) name6376 (
		_w10359_,
		_w10372_,
		_w10380_,
		_w10381_,
		_w10424_
	);
	LUT3 #(
		.INIT('h0b)
	) name6377 (
		_w10358_,
		_w10383_,
		_w10424_,
		_w10425_
	);
	LUT3 #(
		.INIT('h69)
	) name6378 (
		_w10396_,
		_w10423_,
		_w10425_,
		_w10426_
	);
	LUT2 #(
		.INIT('h9)
	) name6379 (
		_w10390_,
		_w10426_,
		_w10427_
	);
	LUT3 #(
		.INIT('h40)
	) name6380 (
		_w10347_,
		_w10349_,
		_w10350_,
		_w10428_
	);
	LUT3 #(
		.INIT('h09)
	) name6381 (
		_w10353_,
		_w10387_,
		_w10428_,
		_w10429_
	);
	LUT3 #(
		.INIT('h0b)
	) name6382 (
		_w10389_,
		_w10427_,
		_w10429_,
		_w10430_
	);
	LUT2 #(
		.INIT('h8)
	) name6383 (
		_w10387_,
		_w10428_,
		_w10431_
	);
	LUT3 #(
		.INIT('h4d)
	) name6384 (
		_w10389_,
		_w10427_,
		_w10431_,
		_w10432_
	);
	LUT3 #(
		.INIT('h70)
	) name6385 (
		_w10352_,
		_w10430_,
		_w10432_,
		_w10433_
	);
	LUT4 #(
		.INIT('h0137)
	) name6386 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9982_,
		_w10413_,
		_w10417_,
		_w10434_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name6387 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w6335_,
		_w6731_,
		_w10435_
	);
	LUT4 #(
		.INIT('h8040)
	) name6388 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10436_
	);
	LUT4 #(
		.INIT('h1020)
	) name6389 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10437_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6390 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10438_
	);
	LUT3 #(
		.INIT('h10)
	) name6391 (
		_w10437_,
		_w10436_,
		_w10438_,
		_w10439_
	);
	LUT4 #(
		.INIT('hc936)
	) name6392 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9985_,
		_w10435_,
		_w10439_,
		_w10440_
	);
	LUT2 #(
		.INIT('h1)
	) name6393 (
		_w10434_,
		_w10440_,
		_w10441_
	);
	LUT3 #(
		.INIT('he8)
	) name6394 (
		_w10406_,
		_w10410_,
		_w10402_,
		_w10442_
	);
	LUT2 #(
		.INIT('h2)
	) name6395 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9956_,
		_w10443_
	);
	LUT2 #(
		.INIT('h1)
	) name6396 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9955_,
		_w10444_
	);
	LUT3 #(
		.INIT('h1b)
	) name6397 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9958_,
		_w9959_,
		_w10445_
	);
	LUT3 #(
		.INIT('h10)
	) name6398 (
		_w10444_,
		_w10443_,
		_w10445_,
		_w10446_
	);
	LUT2 #(
		.INIT('h2)
	) name6399 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9949_,
		_w10447_
	);
	LUT2 #(
		.INIT('h1)
	) name6400 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9948_,
		_w10448_
	);
	LUT3 #(
		.INIT('h1b)
	) name6401 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9951_,
		_w9952_,
		_w10449_
	);
	LUT3 #(
		.INIT('h10)
	) name6402 (
		_w10448_,
		_w10447_,
		_w10449_,
		_w10450_
	);
	LUT2 #(
		.INIT('h2)
	) name6403 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9964_,
		_w10451_
	);
	LUT2 #(
		.INIT('h1)
	) name6404 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9963_,
		_w10452_
	);
	LUT3 #(
		.INIT('h1b)
	) name6405 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9966_,
		_w9967_,
		_w10453_
	);
	LUT3 #(
		.INIT('h10)
	) name6406 (
		_w10452_,
		_w10451_,
		_w10453_,
		_w10454_
	);
	LUT3 #(
		.INIT('h69)
	) name6407 (
		_w10446_,
		_w10450_,
		_w10454_,
		_w10455_
	);
	LUT3 #(
		.INIT('h51)
	) name6408 (
		_w10441_,
		_w10442_,
		_w10455_,
		_w10456_
	);
	LUT3 #(
		.INIT('he8)
	) name6409 (
		_w10446_,
		_w10450_,
		_w10454_,
		_w10457_
	);
	LUT2 #(
		.INIT('h2)
	) name6410 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9949_,
		_w10458_
	);
	LUT2 #(
		.INIT('h1)
	) name6411 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9948_,
		_w10459_
	);
	LUT3 #(
		.INIT('h1b)
	) name6412 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9951_,
		_w9952_,
		_w10460_
	);
	LUT3 #(
		.INIT('h10)
	) name6413 (
		_w10459_,
		_w10458_,
		_w10460_,
		_w10461_
	);
	LUT2 #(
		.INIT('h2)
	) name6414 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9956_,
		_w10462_
	);
	LUT2 #(
		.INIT('h1)
	) name6415 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9955_,
		_w10463_
	);
	LUT3 #(
		.INIT('h1b)
	) name6416 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9958_,
		_w9959_,
		_w10464_
	);
	LUT3 #(
		.INIT('h10)
	) name6417 (
		_w10463_,
		_w10462_,
		_w10464_,
		_w10465_
	);
	LUT2 #(
		.INIT('h2)
	) name6418 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9964_,
		_w10466_
	);
	LUT2 #(
		.INIT('h1)
	) name6419 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9963_,
		_w10467_
	);
	LUT3 #(
		.INIT('h1b)
	) name6420 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9966_,
		_w9967_,
		_w10468_
	);
	LUT3 #(
		.INIT('h10)
	) name6421 (
		_w10467_,
		_w10466_,
		_w10468_,
		_w10469_
	);
	LUT3 #(
		.INIT('h69)
	) name6422 (
		_w10461_,
		_w10465_,
		_w10469_,
		_w10470_
	);
	LUT4 #(
		.INIT('h04cd)
	) name6423 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9985_,
		_w10435_,
		_w10439_,
		_w10471_
	);
	LUT4 #(
		.INIT('hfd75)
	) name6424 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w5720_,
		_w6731_,
		_w10472_
	);
	LUT4 #(
		.INIT('h8040)
	) name6425 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10473_
	);
	LUT4 #(
		.INIT('h1020)
	) name6426 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10474_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6427 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10475_
	);
	LUT3 #(
		.INIT('h10)
	) name6428 (
		_w10474_,
		_w10473_,
		_w10475_,
		_w10476_
	);
	LUT4 #(
		.INIT('h36c9)
	) name6429 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9990_,
		_w10472_,
		_w10476_,
		_w10477_
	);
	LUT2 #(
		.INIT('h1)
	) name6430 (
		_w10471_,
		_w10477_,
		_w10478_
	);
	LUT2 #(
		.INIT('h8)
	) name6431 (
		_w10471_,
		_w10477_,
		_w10479_
	);
	LUT2 #(
		.INIT('h6)
	) name6432 (
		_w10471_,
		_w10477_,
		_w10480_
	);
	LUT3 #(
		.INIT('h69)
	) name6433 (
		_w10457_,
		_w10470_,
		_w10480_,
		_w10481_
	);
	LUT2 #(
		.INIT('h9)
	) name6434 (
		_w10456_,
		_w10481_,
		_w10482_
	);
	LUT3 #(
		.INIT('h0d)
	) name6435 (
		_w10398_,
		_w10411_,
		_w10419_,
		_w10483_
	);
	LUT2 #(
		.INIT('h8)
	) name6436 (
		_w10434_,
		_w10440_,
		_w10484_
	);
	LUT2 #(
		.INIT('h6)
	) name6437 (
		_w10434_,
		_w10440_,
		_w10485_
	);
	LUT3 #(
		.INIT('h69)
	) name6438 (
		_w10442_,
		_w10455_,
		_w10485_,
		_w10486_
	);
	LUT4 #(
		.INIT('h3c20)
	) name6439 (
		_w10441_,
		_w10442_,
		_w10455_,
		_w10484_,
		_w10487_
	);
	LUT3 #(
		.INIT('h07)
	) name6440 (
		_w10483_,
		_w10486_,
		_w10487_,
		_w10488_
	);
	LUT2 #(
		.INIT('h2)
	) name6441 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9983_,
		_w10489_
	);
	LUT2 #(
		.INIT('h1)
	) name6442 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9982_,
		_w10490_
	);
	LUT3 #(
		.INIT('h1b)
	) name6443 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9985_,
		_w9986_,
		_w10491_
	);
	LUT3 #(
		.INIT('h10)
	) name6444 (
		_w10490_,
		_w10489_,
		_w10491_,
		_w10492_
	);
	LUT2 #(
		.INIT('h2)
	) name6445 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9976_,
		_w10493_
	);
	LUT2 #(
		.INIT('h1)
	) name6446 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9975_,
		_w10494_
	);
	LUT3 #(
		.INIT('h1b)
	) name6447 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9978_,
		_w9979_,
		_w10495_
	);
	LUT3 #(
		.INIT('h10)
	) name6448 (
		_w10494_,
		_w10493_,
		_w10495_,
		_w10496_
	);
	LUT2 #(
		.INIT('h1)
	) name6449 (
		_w10492_,
		_w10496_,
		_w10497_
	);
	LUT3 #(
		.INIT('h28)
	) name6450 (
		_w10395_,
		_w10492_,
		_w10496_,
		_w10498_
	);
	LUT3 #(
		.INIT('he4)
	) name6451 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9990_,
		_w9991_,
		_w10499_
	);
	LUT2 #(
		.INIT('h2)
	) name6452 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9983_,
		_w10500_
	);
	LUT2 #(
		.INIT('h1)
	) name6453 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9982_,
		_w10501_
	);
	LUT3 #(
		.INIT('h1b)
	) name6454 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9985_,
		_w9986_,
		_w10502_
	);
	LUT4 #(
		.INIT('h0200)
	) name6455 (
		_w10499_,
		_w10501_,
		_w10500_,
		_w10502_,
		_w10503_
	);
	LUT4 #(
		.INIT('h5455)
	) name6456 (
		_w10499_,
		_w10501_,
		_w10500_,
		_w10502_,
		_w10504_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6457 (
		_w10499_,
		_w10501_,
		_w10500_,
		_w10502_,
		_w10505_
	);
	LUT2 #(
		.INIT('h2)
	) name6458 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9976_,
		_w10506_
	);
	LUT2 #(
		.INIT('h1)
	) name6459 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9975_,
		_w10507_
	);
	LUT3 #(
		.INIT('h1b)
	) name6460 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9978_,
		_w9979_,
		_w10508_
	);
	LUT3 #(
		.INIT('h10)
	) name6461 (
		_w10507_,
		_w10506_,
		_w10508_,
		_w10509_
	);
	LUT2 #(
		.INIT('h9)
	) name6462 (
		_w10505_,
		_w10509_,
		_w10510_
	);
	LUT4 #(
		.INIT('h1001)
	) name6463 (
		_w10492_,
		_w10496_,
		_w10505_,
		_w10509_,
		_w10511_
	);
	LUT4 #(
		.INIT('he11e)
	) name6464 (
		_w10492_,
		_w10496_,
		_w10505_,
		_w10509_,
		_w10512_
	);
	LUT2 #(
		.INIT('h1)
	) name6465 (
		_w10498_,
		_w10512_,
		_w10513_
	);
	LUT3 #(
		.INIT('h07)
	) name6466 (
		_w10482_,
		_w10488_,
		_w10513_,
		_w10514_
	);
	LUT3 #(
		.INIT('h0d)
	) name6467 (
		_w10457_,
		_w10470_,
		_w10478_,
		_w10515_
	);
	LUT3 #(
		.INIT('he8)
	) name6468 (
		_w10461_,
		_w10465_,
		_w10469_,
		_w10516_
	);
	LUT2 #(
		.INIT('h2)
	) name6469 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9956_,
		_w10517_
	);
	LUT2 #(
		.INIT('h1)
	) name6470 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9955_,
		_w10518_
	);
	LUT3 #(
		.INIT('h1b)
	) name6471 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9958_,
		_w9959_,
		_w10519_
	);
	LUT3 #(
		.INIT('h10)
	) name6472 (
		_w10518_,
		_w10517_,
		_w10519_,
		_w10520_
	);
	LUT2 #(
		.INIT('h2)
	) name6473 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9949_,
		_w10521_
	);
	LUT2 #(
		.INIT('h1)
	) name6474 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9948_,
		_w10522_
	);
	LUT3 #(
		.INIT('h1b)
	) name6475 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9951_,
		_w9952_,
		_w10523_
	);
	LUT3 #(
		.INIT('h10)
	) name6476 (
		_w10522_,
		_w10521_,
		_w10523_,
		_w10524_
	);
	LUT2 #(
		.INIT('h2)
	) name6477 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9964_,
		_w10525_
	);
	LUT2 #(
		.INIT('h1)
	) name6478 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9963_,
		_w10526_
	);
	LUT3 #(
		.INIT('h1b)
	) name6479 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9966_,
		_w9967_,
		_w10527_
	);
	LUT3 #(
		.INIT('h10)
	) name6480 (
		_w10526_,
		_w10525_,
		_w10527_,
		_w10528_
	);
	LUT3 #(
		.INIT('h69)
	) name6481 (
		_w10520_,
		_w10524_,
		_w10528_,
		_w10529_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name6482 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w5720_,
		_w8296_,
		_w10530_
	);
	LUT4 #(
		.INIT('h8040)
	) name6483 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10531_
	);
	LUT4 #(
		.INIT('h1020)
	) name6484 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10532_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6485 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10533_
	);
	LUT3 #(
		.INIT('h10)
	) name6486 (
		_w10532_,
		_w10531_,
		_w10533_,
		_w10534_
	);
	LUT4 #(
		.INIT('hc936)
	) name6487 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9993_,
		_w10530_,
		_w10534_,
		_w10535_
	);
	LUT4 #(
		.INIT('h0137)
	) name6488 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9990_,
		_w10472_,
		_w10476_,
		_w10536_
	);
	LUT2 #(
		.INIT('h1)
	) name6489 (
		_w10535_,
		_w10536_,
		_w10537_
	);
	LUT2 #(
		.INIT('h8)
	) name6490 (
		_w10535_,
		_w10536_,
		_w10538_
	);
	LUT2 #(
		.INIT('h6)
	) name6491 (
		_w10535_,
		_w10536_,
		_w10539_
	);
	LUT3 #(
		.INIT('h69)
	) name6492 (
		_w10516_,
		_w10529_,
		_w10539_,
		_w10540_
	);
	LUT2 #(
		.INIT('h9)
	) name6493 (
		_w10515_,
		_w10540_,
		_w10541_
	);
	LUT4 #(
		.INIT('h0029)
	) name6494 (
		_w10457_,
		_w10470_,
		_w10478_,
		_w10479_,
		_w10542_
	);
	LUT3 #(
		.INIT('h0b)
	) name6495 (
		_w10456_,
		_w10481_,
		_w10542_,
		_w10543_
	);
	LUT3 #(
		.INIT('h32)
	) name6496 (
		_w10503_,
		_w10504_,
		_w10509_,
		_w10544_
	);
	LUT2 #(
		.INIT('h2)
	) name6497 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9976_,
		_w10545_
	);
	LUT2 #(
		.INIT('h1)
	) name6498 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9975_,
		_w10546_
	);
	LUT3 #(
		.INIT('h1b)
	) name6499 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9978_,
		_w9979_,
		_w10547_
	);
	LUT3 #(
		.INIT('h10)
	) name6500 (
		_w10546_,
		_w10545_,
		_w10547_,
		_w10548_
	);
	LUT2 #(
		.INIT('h2)
	) name6501 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9991_,
		_w10549_
	);
	LUT2 #(
		.INIT('h1)
	) name6502 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9990_,
		_w10550_
	);
	LUT3 #(
		.INIT('h1b)
	) name6503 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w9993_,
		_w9994_,
		_w10551_
	);
	LUT3 #(
		.INIT('h10)
	) name6504 (
		_w10550_,
		_w10549_,
		_w10551_,
		_w10552_
	);
	LUT2 #(
		.INIT('h2)
	) name6505 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9983_,
		_w10553_
	);
	LUT2 #(
		.INIT('h1)
	) name6506 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9982_,
		_w10554_
	);
	LUT3 #(
		.INIT('h1b)
	) name6507 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9985_,
		_w9986_,
		_w10555_
	);
	LUT3 #(
		.INIT('h10)
	) name6508 (
		_w10554_,
		_w10553_,
		_w10555_,
		_w10556_
	);
	LUT3 #(
		.INIT('h69)
	) name6509 (
		_w10548_,
		_w10552_,
		_w10556_,
		_w10557_
	);
	LUT2 #(
		.INIT('h4)
	) name6510 (
		_w10544_,
		_w10557_,
		_w10558_
	);
	LUT2 #(
		.INIT('h9)
	) name6511 (
		_w10544_,
		_w10557_,
		_w10559_
	);
	LUT3 #(
		.INIT('h14)
	) name6512 (
		_w10511_,
		_w10544_,
		_w10557_,
		_w10560_
	);
	LUT3 #(
		.INIT('h69)
	) name6513 (
		_w10511_,
		_w10544_,
		_w10557_,
		_w10561_
	);
	LUT3 #(
		.INIT('h69)
	) name6514 (
		_w10541_,
		_w10543_,
		_w10561_,
		_w10562_
	);
	LUT2 #(
		.INIT('h9)
	) name6515 (
		_w10514_,
		_w10562_,
		_w10563_
	);
	LUT3 #(
		.INIT('h96)
	) name6516 (
		_w10395_,
		_w10492_,
		_w10496_,
		_w10564_
	);
	LUT2 #(
		.INIT('h6)
	) name6517 (
		_w10483_,
		_w10486_,
		_w10565_
	);
	LUT4 #(
		.INIT('h0029)
	) name6518 (
		_w10398_,
		_w10411_,
		_w10419_,
		_w10420_,
		_w10566_
	);
	LUT3 #(
		.INIT('h0b)
	) name6519 (
		_w10397_,
		_w10422_,
		_w10566_,
		_w10567_
	);
	LUT3 #(
		.INIT('ha8)
	) name6520 (
		_w10564_,
		_w10565_,
		_w10567_,
		_w10568_
	);
	LUT2 #(
		.INIT('h8)
	) name6521 (
		_w10498_,
		_w10510_,
		_w10569_
	);
	LUT3 #(
		.INIT('h1e)
	) name6522 (
		_w10497_,
		_w10498_,
		_w10510_,
		_w10570_
	);
	LUT3 #(
		.INIT('h96)
	) name6523 (
		_w10482_,
		_w10488_,
		_w10570_,
		_w10571_
	);
	LUT4 #(
		.INIT('h0608)
	) name6524 (
		_w10482_,
		_w10488_,
		_w10569_,
		_w10570_,
		_w10572_
	);
	LUT3 #(
		.INIT('h0b)
	) name6525 (
		_w10568_,
		_w10571_,
		_w10572_,
		_w10573_
	);
	LUT2 #(
		.INIT('h2)
	) name6526 (
		_w10563_,
		_w10573_,
		_w10574_
	);
	LUT3 #(
		.INIT('h0d)
	) name6527 (
		_w10541_,
		_w10543_,
		_w10560_,
		_w10575_
	);
	LUT2 #(
		.INIT('h4)
	) name6528 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 ,
		_w10576_
	);
	LUT4 #(
		.INIT('h1b00)
	) name6529 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w10001_,
		_w10002_,
		_w10576_,
		_w10577_
	);
	LUT4 #(
		.INIT('he41b)
	) name6530 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w10001_,
		_w10002_,
		_w10576_,
		_w10578_
	);
	LUT3 #(
		.INIT('he8)
	) name6531 (
		_w10548_,
		_w10552_,
		_w10556_,
		_w10579_
	);
	LUT2 #(
		.INIT('h2)
	) name6532 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9983_,
		_w10580_
	);
	LUT2 #(
		.INIT('h1)
	) name6533 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9982_,
		_w10581_
	);
	LUT3 #(
		.INIT('h1b)
	) name6534 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9985_,
		_w9986_,
		_w10582_
	);
	LUT3 #(
		.INIT('h10)
	) name6535 (
		_w10581_,
		_w10580_,
		_w10582_,
		_w10583_
	);
	LUT2 #(
		.INIT('h2)
	) name6536 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9976_,
		_w10584_
	);
	LUT2 #(
		.INIT('h1)
	) name6537 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9975_,
		_w10585_
	);
	LUT3 #(
		.INIT('h1b)
	) name6538 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9978_,
		_w9979_,
		_w10586_
	);
	LUT3 #(
		.INIT('h10)
	) name6539 (
		_w10585_,
		_w10584_,
		_w10586_,
		_w10587_
	);
	LUT2 #(
		.INIT('h2)
	) name6540 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9991_,
		_w10588_
	);
	LUT2 #(
		.INIT('h1)
	) name6541 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9990_,
		_w10589_
	);
	LUT3 #(
		.INIT('h1b)
	) name6542 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w9993_,
		_w9994_,
		_w10590_
	);
	LUT3 #(
		.INIT('h10)
	) name6543 (
		_w10589_,
		_w10588_,
		_w10590_,
		_w10591_
	);
	LUT3 #(
		.INIT('h69)
	) name6544 (
		_w10583_,
		_w10587_,
		_w10591_,
		_w10592_
	);
	LUT3 #(
		.INIT('h69)
	) name6545 (
		_w10578_,
		_w10579_,
		_w10592_,
		_w10593_
	);
	LUT2 #(
		.INIT('h1)
	) name6546 (
		_w10558_,
		_w10593_,
		_w10594_
	);
	LUT2 #(
		.INIT('h6)
	) name6547 (
		_w10558_,
		_w10593_,
		_w10595_
	);
	LUT3 #(
		.INIT('h0d)
	) name6548 (
		_w10516_,
		_w10529_,
		_w10537_,
		_w10596_
	);
	LUT3 #(
		.INIT('he8)
	) name6549 (
		_w10520_,
		_w10524_,
		_w10528_,
		_w10597_
	);
	LUT2 #(
		.INIT('h2)
	) name6550 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9956_,
		_w10598_
	);
	LUT2 #(
		.INIT('h1)
	) name6551 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9955_,
		_w10599_
	);
	LUT3 #(
		.INIT('h1b)
	) name6552 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9958_,
		_w9959_,
		_w10600_
	);
	LUT3 #(
		.INIT('h10)
	) name6553 (
		_w10599_,
		_w10598_,
		_w10600_,
		_w10601_
	);
	LUT2 #(
		.INIT('h2)
	) name6554 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9949_,
		_w10602_
	);
	LUT2 #(
		.INIT('h1)
	) name6555 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9948_,
		_w10603_
	);
	LUT3 #(
		.INIT('h1b)
	) name6556 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9951_,
		_w9952_,
		_w10604_
	);
	LUT3 #(
		.INIT('h10)
	) name6557 (
		_w10603_,
		_w10602_,
		_w10604_,
		_w10605_
	);
	LUT2 #(
		.INIT('h2)
	) name6558 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9964_,
		_w10606_
	);
	LUT2 #(
		.INIT('h1)
	) name6559 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9963_,
		_w10607_
	);
	LUT3 #(
		.INIT('h1b)
	) name6560 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9966_,
		_w9967_,
		_w10608_
	);
	LUT3 #(
		.INIT('h10)
	) name6561 (
		_w10607_,
		_w10606_,
		_w10608_,
		_w10609_
	);
	LUT3 #(
		.INIT('h69)
	) name6562 (
		_w10601_,
		_w10605_,
		_w10609_,
		_w10610_
	);
	LUT4 #(
		.INIT('hfb32)
	) name6563 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w9993_,
		_w10530_,
		_w10534_,
		_w10611_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name6564 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w8296_,
		_w8375_,
		_w10612_
	);
	LUT4 #(
		.INIT('h8040)
	) name6565 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10613_
	);
	LUT4 #(
		.INIT('h1020)
	) name6566 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10614_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6567 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w10615_
	);
	LUT3 #(
		.INIT('h10)
	) name6568 (
		_w10614_,
		_w10613_,
		_w10615_,
		_w10616_
	);
	LUT4 #(
		.INIT('hc936)
	) name6569 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10001_,
		_w10612_,
		_w10616_,
		_w10617_
	);
	LUT2 #(
		.INIT('h8)
	) name6570 (
		_w10611_,
		_w10617_,
		_w10618_
	);
	LUT2 #(
		.INIT('h1)
	) name6571 (
		_w10611_,
		_w10617_,
		_w10619_
	);
	LUT2 #(
		.INIT('h6)
	) name6572 (
		_w10611_,
		_w10617_,
		_w10620_
	);
	LUT3 #(
		.INIT('h69)
	) name6573 (
		_w10597_,
		_w10610_,
		_w10620_,
		_w10621_
	);
	LUT2 #(
		.INIT('h9)
	) name6574 (
		_w10596_,
		_w10621_,
		_w10622_
	);
	LUT4 #(
		.INIT('h0029)
	) name6575 (
		_w10516_,
		_w10529_,
		_w10537_,
		_w10538_,
		_w10623_
	);
	LUT3 #(
		.INIT('h0b)
	) name6576 (
		_w10515_,
		_w10540_,
		_w10623_,
		_w10624_
	);
	LUT3 #(
		.INIT('h69)
	) name6577 (
		_w10595_,
		_w10622_,
		_w10624_,
		_w10625_
	);
	LUT2 #(
		.INIT('h9)
	) name6578 (
		_w10575_,
		_w10625_,
		_w10626_
	);
	LUT4 #(
		.INIT('h4186)
	) name6579 (
		_w10511_,
		_w10541_,
		_w10543_,
		_w10559_,
		_w10627_
	);
	LUT3 #(
		.INIT('h0b)
	) name6580 (
		_w10514_,
		_w10562_,
		_w10627_,
		_w10628_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name6581 (
		_w10563_,
		_w10573_,
		_w10626_,
		_w10628_,
		_w10629_
	);
	LUT3 #(
		.INIT('ha2)
	) name6582 (
		_w10396_,
		_w10423_,
		_w10425_,
		_w10630_
	);
	LUT3 #(
		.INIT('h69)
	) name6583 (
		_w10564_,
		_w10565_,
		_w10567_,
		_w10631_
	);
	LUT3 #(
		.INIT('h29)
	) name6584 (
		_w10564_,
		_w10565_,
		_w10567_,
		_w10632_
	);
	LUT3 #(
		.INIT('h0e)
	) name6585 (
		_w10630_,
		_w10631_,
		_w10632_,
		_w10633_
	);
	LUT2 #(
		.INIT('h9)
	) name6586 (
		_w10568_,
		_w10571_,
		_w10634_
	);
	LUT3 #(
		.INIT('h86)
	) name6587 (
		_w10396_,
		_w10423_,
		_w10425_,
		_w10635_
	);
	LUT3 #(
		.INIT('h0b)
	) name6588 (
		_w10390_,
		_w10426_,
		_w10635_,
		_w10636_
	);
	LUT2 #(
		.INIT('h6)
	) name6589 (
		_w10630_,
		_w10631_,
		_w10637_
	);
	LUT2 #(
		.INIT('h4)
	) name6590 (
		_w10636_,
		_w10637_,
		_w10638_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6591 (
		_w10633_,
		_w10634_,
		_w10636_,
		_w10637_,
		_w10639_
	);
	LUT2 #(
		.INIT('h8)
	) name6592 (
		_w10629_,
		_w10639_,
		_w10640_
	);
	LUT2 #(
		.INIT('h2)
	) name6593 (
		_w10636_,
		_w10637_,
		_w10641_
	);
	LUT4 #(
		.INIT('hdd4d)
	) name6594 (
		_w10633_,
		_w10634_,
		_w10636_,
		_w10637_,
		_w10642_
	);
	LUT2 #(
		.INIT('h4)
	) name6595 (
		_w10563_,
		_w10573_,
		_w10643_
	);
	LUT4 #(
		.INIT('hb0fb)
	) name6596 (
		_w10563_,
		_w10573_,
		_w10626_,
		_w10628_,
		_w10644_
	);
	LUT3 #(
		.INIT('hd0)
	) name6597 (
		_w10629_,
		_w10642_,
		_w10644_,
		_w10645_
	);
	LUT3 #(
		.INIT('hb0)
	) name6598 (
		_w10433_,
		_w10640_,
		_w10645_,
		_w10646_
	);
	LUT4 #(
		.INIT('h0777)
	) name6599 (
		_w9950_,
		_w9953_,
		_w9957_,
		_w9960_,
		_w10647_
	);
	LUT2 #(
		.INIT('h2)
	) name6600 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9964_,
		_w10648_
	);
	LUT2 #(
		.INIT('h1)
	) name6601 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9963_,
		_w10649_
	);
	LUT3 #(
		.INIT('h1b)
	) name6602 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9966_,
		_w9967_,
		_w10650_
	);
	LUT3 #(
		.INIT('h10)
	) name6603 (
		_w10649_,
		_w10648_,
		_w10650_,
		_w10651_
	);
	LUT4 #(
		.INIT('h7888)
	) name6604 (
		_w9950_,
		_w9953_,
		_w9957_,
		_w9960_,
		_w10652_
	);
	LUT3 #(
		.INIT('h1b)
	) name6605 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9966_,
		_w9967_,
		_w10653_
	);
	LUT2 #(
		.INIT('h8)
	) name6606 (
		_w9965_,
		_w10653_,
		_w10654_
	);
	LUT4 #(
		.INIT('h8860)
	) name6607 (
		_w9954_,
		_w9961_,
		_w10651_,
		_w10654_,
		_w10655_
	);
	LUT4 #(
		.INIT('h0161)
	) name6608 (
		_w9954_,
		_w9961_,
		_w9969_,
		_w10654_,
		_w10656_
	);
	LUT4 #(
		.INIT('h8680)
	) name6609 (
		_w9954_,
		_w9961_,
		_w9969_,
		_w10654_,
		_w10657_
	);
	LUT4 #(
		.INIT('hc6c3)
	) name6610 (
		_w9962_,
		_w9969_,
		_w10647_,
		_w10654_,
		_w10658_
	);
	LUT3 #(
		.INIT('h4b)
	) name6611 (
		_w9973_,
		_w10655_,
		_w10658_,
		_w10659_
	);
	LUT3 #(
		.INIT('h1b)
	) name6612 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9958_,
		_w9959_,
		_w10660_
	);
	LUT2 #(
		.INIT('h8)
	) name6613 (
		_w9957_,
		_w10660_,
		_w10661_
	);
	LUT2 #(
		.INIT('h2)
	) name6614 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9964_,
		_w10662_
	);
	LUT2 #(
		.INIT('h1)
	) name6615 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9963_,
		_w10663_
	);
	LUT3 #(
		.INIT('h1b)
	) name6616 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9966_,
		_w9967_,
		_w10664_
	);
	LUT3 #(
		.INIT('h10)
	) name6617 (
		_w10663_,
		_w10662_,
		_w10664_,
		_w10665_
	);
	LUT3 #(
		.INIT('he8)
	) name6618 (
		_w9954_,
		_w10661_,
		_w10665_,
		_w10666_
	);
	LUT2 #(
		.INIT('h9)
	) name6619 (
		_w10651_,
		_w10652_,
		_w10667_
	);
	LUT3 #(
		.INIT('h51)
	) name6620 (
		_w9973_,
		_w10666_,
		_w10667_,
		_w10668_
	);
	LUT4 #(
		.INIT('h0611)
	) name6621 (
		_w9954_,
		_w9961_,
		_w10651_,
		_w10654_,
		_w10669_
	);
	LUT4 #(
		.INIT('hdc23)
	) name6622 (
		_w9962_,
		_w10647_,
		_w10651_,
		_w10654_,
		_w10670_
	);
	LUT3 #(
		.INIT('h56)
	) name6623 (
		_w9973_,
		_w10655_,
		_w10669_,
		_w10671_
	);
	LUT3 #(
		.INIT('h09)
	) name6624 (
		_w9973_,
		_w10655_,
		_w10669_,
		_w10672_
	);
	LUT3 #(
		.INIT('h0b)
	) name6625 (
		_w10668_,
		_w10671_,
		_w10672_,
		_w10673_
	);
	LUT4 #(
		.INIT('h220a)
	) name6626 (
		_w10659_,
		_w10668_,
		_w10669_,
		_w10671_,
		_w10674_
	);
	LUT2 #(
		.INIT('h1)
	) name6627 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9975_,
		_w10675_
	);
	LUT2 #(
		.INIT('h2)
	) name6628 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9976_,
		_w10676_
	);
	LUT3 #(
		.INIT('h1b)
	) name6629 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9978_,
		_w9979_,
		_w10677_
	);
	LUT3 #(
		.INIT('h10)
	) name6630 (
		_w10676_,
		_w10675_,
		_w10677_,
		_w10678_
	);
	LUT2 #(
		.INIT('h2)
	) name6631 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9983_,
		_w10679_
	);
	LUT2 #(
		.INIT('h1)
	) name6632 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9982_,
		_w10680_
	);
	LUT3 #(
		.INIT('h1b)
	) name6633 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9985_,
		_w9986_,
		_w10681_
	);
	LUT3 #(
		.INIT('h10)
	) name6634 (
		_w10680_,
		_w10679_,
		_w10681_,
		_w10682_
	);
	LUT2 #(
		.INIT('h2)
	) name6635 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9991_,
		_w10683_
	);
	LUT2 #(
		.INIT('h1)
	) name6636 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9990_,
		_w10684_
	);
	LUT3 #(
		.INIT('h1b)
	) name6637 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9993_,
		_w9994_,
		_w10685_
	);
	LUT3 #(
		.INIT('h10)
	) name6638 (
		_w10684_,
		_w10683_,
		_w10685_,
		_w10686_
	);
	LUT3 #(
		.INIT('he8)
	) name6639 (
		_w10678_,
		_w10682_,
		_w10686_,
		_w10687_
	);
	LUT2 #(
		.INIT('h2)
	) name6640 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9976_,
		_w10688_
	);
	LUT2 #(
		.INIT('h1)
	) name6641 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9975_,
		_w10689_
	);
	LUT3 #(
		.INIT('h1b)
	) name6642 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9978_,
		_w9979_,
		_w10690_
	);
	LUT3 #(
		.INIT('h10)
	) name6643 (
		_w10689_,
		_w10688_,
		_w10690_,
		_w10691_
	);
	LUT2 #(
		.INIT('h2)
	) name6644 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9983_,
		_w10692_
	);
	LUT2 #(
		.INIT('h1)
	) name6645 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9982_,
		_w10693_
	);
	LUT3 #(
		.INIT('h1b)
	) name6646 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9985_,
		_w9986_,
		_w10694_
	);
	LUT3 #(
		.INIT('h10)
	) name6647 (
		_w10693_,
		_w10692_,
		_w10694_,
		_w10695_
	);
	LUT2 #(
		.INIT('h2)
	) name6648 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9991_,
		_w10696_
	);
	LUT2 #(
		.INIT('h1)
	) name6649 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9990_,
		_w10697_
	);
	LUT3 #(
		.INIT('h1b)
	) name6650 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9993_,
		_w9994_,
		_w10698_
	);
	LUT3 #(
		.INIT('h10)
	) name6651 (
		_w10697_,
		_w10696_,
		_w10698_,
		_w10699_
	);
	LUT3 #(
		.INIT('h69)
	) name6652 (
		_w10691_,
		_w10695_,
		_w10699_,
		_w10700_
	);
	LUT4 #(
		.INIT('h4800)
	) name6653 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10701_
	);
	LUT2 #(
		.INIT('h2)
	) name6654 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w10002_,
		_w10702_
	);
	LUT2 #(
		.INIT('h1)
	) name6655 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w10001_,
		_w10703_
	);
	LUT3 #(
		.INIT('h1b)
	) name6656 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w10004_,
		_w10005_,
		_w10704_
	);
	LUT4 #(
		.INIT('h0100)
	) name6657 (
		_w10701_,
		_w10703_,
		_w10702_,
		_w10704_,
		_w10705_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6658 (
		_w10701_,
		_w10703_,
		_w10702_,
		_w10704_,
		_w10706_
	);
	LUT4 #(
		.INIT('h5655)
	) name6659 (
		_w10701_,
		_w10703_,
		_w10702_,
		_w10704_,
		_w10707_
	);
	LUT4 #(
		.INIT('ha820)
	) name6660 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 ,
		_w10708_
	);
	LUT4 #(
		.INIT('ha820)
	) name6661 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 ,
		_w10709_
	);
	LUT4 #(
		.INIT('h3120)
	) name6662 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10709_,
		_w10708_,
		_w10710_
	);
	LUT2 #(
		.INIT('h9)
	) name6663 (
		_w10707_,
		_w10710_,
		_w10711_
	);
	LUT4 #(
		.INIT('h4800)
	) name6664 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10712_
	);
	LUT2 #(
		.INIT('h2)
	) name6665 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w10002_,
		_w10713_
	);
	LUT2 #(
		.INIT('h1)
	) name6666 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w10001_,
		_w10714_
	);
	LUT3 #(
		.INIT('h1b)
	) name6667 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w10004_,
		_w10005_,
		_w10715_
	);
	LUT4 #(
		.INIT('h0100)
	) name6668 (
		_w10712_,
		_w10714_,
		_w10713_,
		_w10715_,
		_w10716_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6669 (
		_w10712_,
		_w10714_,
		_w10713_,
		_w10715_,
		_w10717_
	);
	LUT4 #(
		.INIT('ha820)
	) name6670 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 ,
		_w10718_
	);
	LUT4 #(
		.INIT('h3210)
	) name6671 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10709_,
		_w10718_,
		_w10719_
	);
	LUT3 #(
		.INIT('h54)
	) name6672 (
		_w10716_,
		_w10717_,
		_w10719_,
		_w10720_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name6673 (
		_w10687_,
		_w10700_,
		_w10711_,
		_w10720_,
		_w10721_
	);
	LUT3 #(
		.INIT('h23)
	) name6674 (
		_w10705_,
		_w10706_,
		_w10710_,
		_w10722_
	);
	LUT4 #(
		.INIT('ha820)
	) name6675 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 ,
		_w10723_
	);
	LUT4 #(
		.INIT('h3120)
	) name6676 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10708_,
		_w10723_,
		_w10724_
	);
	LUT2 #(
		.INIT('h2)
	) name6677 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w10002_,
		_w10725_
	);
	LUT2 #(
		.INIT('h1)
	) name6678 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w10001_,
		_w10726_
	);
	LUT3 #(
		.INIT('h1b)
	) name6679 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w10004_,
		_w10005_,
		_w10727_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6680 (
		_w10724_,
		_w10726_,
		_w10725_,
		_w10727_,
		_w10728_
	);
	LUT4 #(
		.INIT('h0100)
	) name6681 (
		_w10724_,
		_w10726_,
		_w10725_,
		_w10727_,
		_w10729_
	);
	LUT4 #(
		.INIT('h5655)
	) name6682 (
		_w10724_,
		_w10726_,
		_w10725_,
		_w10727_,
		_w10730_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name6683 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10731_
	);
	LUT2 #(
		.INIT('h6)
	) name6684 (
		_w10730_,
		_w10731_,
		_w10732_
	);
	LUT3 #(
		.INIT('he8)
	) name6685 (
		_w10691_,
		_w10695_,
		_w10699_,
		_w10733_
	);
	LUT2 #(
		.INIT('h2)
	) name6686 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9983_,
		_w10734_
	);
	LUT2 #(
		.INIT('h1)
	) name6687 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9982_,
		_w10735_
	);
	LUT3 #(
		.INIT('h1b)
	) name6688 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9985_,
		_w9986_,
		_w10736_
	);
	LUT3 #(
		.INIT('h10)
	) name6689 (
		_w10735_,
		_w10734_,
		_w10736_,
		_w10737_
	);
	LUT2 #(
		.INIT('h2)
	) name6690 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9976_,
		_w10738_
	);
	LUT2 #(
		.INIT('h1)
	) name6691 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9975_,
		_w10739_
	);
	LUT3 #(
		.INIT('h1b)
	) name6692 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9978_,
		_w9979_,
		_w10740_
	);
	LUT3 #(
		.INIT('h10)
	) name6693 (
		_w10739_,
		_w10738_,
		_w10740_,
		_w10741_
	);
	LUT2 #(
		.INIT('h2)
	) name6694 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9991_,
		_w10742_
	);
	LUT2 #(
		.INIT('h1)
	) name6695 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9990_,
		_w10743_
	);
	LUT3 #(
		.INIT('h1b)
	) name6696 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9993_,
		_w9994_,
		_w10744_
	);
	LUT3 #(
		.INIT('h10)
	) name6697 (
		_w10743_,
		_w10742_,
		_w10744_,
		_w10745_
	);
	LUT3 #(
		.INIT('h69)
	) name6698 (
		_w10737_,
		_w10741_,
		_w10745_,
		_w10746_
	);
	LUT4 #(
		.INIT('h6996)
	) name6699 (
		_w10722_,
		_w10732_,
		_w10733_,
		_w10746_,
		_w10747_
	);
	LUT2 #(
		.INIT('h6)
	) name6700 (
		_w10721_,
		_w10747_,
		_w10748_
	);
	LUT4 #(
		.INIT('h5655)
	) name6701 (
		_w10712_,
		_w10714_,
		_w10713_,
		_w10715_,
		_w10749_
	);
	LUT2 #(
		.INIT('h9)
	) name6702 (
		_w10719_,
		_w10749_,
		_w10750_
	);
	LUT4 #(
		.INIT('ha820)
	) name6703 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 ,
		_w10751_
	);
	LUT4 #(
		.INIT('h3210)
	) name6704 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10718_,
		_w10751_,
		_w10752_
	);
	LUT2 #(
		.INIT('h2)
	) name6705 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w10002_,
		_w10753_
	);
	LUT2 #(
		.INIT('h1)
	) name6706 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w10001_,
		_w10754_
	);
	LUT3 #(
		.INIT('h1b)
	) name6707 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w10004_,
		_w10005_,
		_w10755_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6708 (
		_w10752_,
		_w10754_,
		_w10753_,
		_w10755_,
		_w10756_
	);
	LUT4 #(
		.INIT('h0100)
	) name6709 (
		_w10752_,
		_w10754_,
		_w10753_,
		_w10755_,
		_w10757_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name6710 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10758_
	);
	LUT3 #(
		.INIT('h54)
	) name6711 (
		_w10756_,
		_w10757_,
		_w10758_,
		_w10759_
	);
	LUT2 #(
		.INIT('h2)
	) name6712 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9983_,
		_w10760_
	);
	LUT2 #(
		.INIT('h1)
	) name6713 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9982_,
		_w10761_
	);
	LUT3 #(
		.INIT('h1b)
	) name6714 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9985_,
		_w9986_,
		_w10762_
	);
	LUT3 #(
		.INIT('h10)
	) name6715 (
		_w10761_,
		_w10760_,
		_w10762_,
		_w10763_
	);
	LUT2 #(
		.INIT('h2)
	) name6716 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9976_,
		_w10764_
	);
	LUT2 #(
		.INIT('h1)
	) name6717 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9975_,
		_w10765_
	);
	LUT3 #(
		.INIT('h1b)
	) name6718 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9978_,
		_w9979_,
		_w10766_
	);
	LUT3 #(
		.INIT('h10)
	) name6719 (
		_w10765_,
		_w10764_,
		_w10766_,
		_w10767_
	);
	LUT2 #(
		.INIT('h2)
	) name6720 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9991_,
		_w10768_
	);
	LUT2 #(
		.INIT('h1)
	) name6721 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9990_,
		_w10769_
	);
	LUT3 #(
		.INIT('h1b)
	) name6722 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9993_,
		_w9994_,
		_w10770_
	);
	LUT3 #(
		.INIT('h10)
	) name6723 (
		_w10769_,
		_w10768_,
		_w10770_,
		_w10771_
	);
	LUT3 #(
		.INIT('he8)
	) name6724 (
		_w10763_,
		_w10767_,
		_w10771_,
		_w10772_
	);
	LUT3 #(
		.INIT('h69)
	) name6725 (
		_w10678_,
		_w10682_,
		_w10686_,
		_w10773_
	);
	LUT4 #(
		.INIT('h7707)
	) name6726 (
		_w10750_,
		_w10759_,
		_w10772_,
		_w10773_,
		_w10774_
	);
	LUT4 #(
		.INIT('h6996)
	) name6727 (
		_w10687_,
		_w10700_,
		_w10711_,
		_w10720_,
		_w10775_
	);
	LUT4 #(
		.INIT('h9029)
	) name6728 (
		_w10687_,
		_w10700_,
		_w10711_,
		_w10720_,
		_w10776_
	);
	LUT3 #(
		.INIT('h0b)
	) name6729 (
		_w10774_,
		_w10775_,
		_w10776_,
		_w10777_
	);
	LUT3 #(
		.INIT('h51)
	) name6730 (
		_w10674_,
		_w10748_,
		_w10777_,
		_w10778_
	);
	LUT4 #(
		.INIT('h7707)
	) name6731 (
		_w10722_,
		_w10732_,
		_w10733_,
		_w10746_,
		_w10779_
	);
	LUT3 #(
		.INIT('he8)
	) name6732 (
		_w10737_,
		_w10741_,
		_w10745_,
		_w10780_
	);
	LUT3 #(
		.INIT('h1b)
	) name6733 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9978_,
		_w9979_,
		_w10781_
	);
	LUT2 #(
		.INIT('h8)
	) name6734 (
		_w9977_,
		_w10781_,
		_w10782_
	);
	LUT2 #(
		.INIT('h2)
	) name6735 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9983_,
		_w10783_
	);
	LUT2 #(
		.INIT('h1)
	) name6736 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9982_,
		_w10784_
	);
	LUT3 #(
		.INIT('h1b)
	) name6737 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9985_,
		_w9986_,
		_w10785_
	);
	LUT3 #(
		.INIT('h10)
	) name6738 (
		_w10784_,
		_w10783_,
		_w10785_,
		_w10786_
	);
	LUT2 #(
		.INIT('h2)
	) name6739 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9991_,
		_w10787_
	);
	LUT2 #(
		.INIT('h1)
	) name6740 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9990_,
		_w10788_
	);
	LUT3 #(
		.INIT('h1b)
	) name6741 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9993_,
		_w9994_,
		_w10789_
	);
	LUT3 #(
		.INIT('h10)
	) name6742 (
		_w10788_,
		_w10787_,
		_w10789_,
		_w10790_
	);
	LUT3 #(
		.INIT('h69)
	) name6743 (
		_w10782_,
		_w10786_,
		_w10790_,
		_w10791_
	);
	LUT4 #(
		.INIT('h4800)
	) name6744 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10792_
	);
	LUT2 #(
		.INIT('h2)
	) name6745 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w10002_,
		_w10793_
	);
	LUT2 #(
		.INIT('h1)
	) name6746 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w10001_,
		_w10794_
	);
	LUT3 #(
		.INIT('h1b)
	) name6747 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w10004_,
		_w10005_,
		_w10795_
	);
	LUT4 #(
		.INIT('h0100)
	) name6748 (
		_w10792_,
		_w10794_,
		_w10793_,
		_w10795_,
		_w10796_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6749 (
		_w10792_,
		_w10794_,
		_w10793_,
		_w10795_,
		_w10797_
	);
	LUT4 #(
		.INIT('h5655)
	) name6750 (
		_w10792_,
		_w10794_,
		_w10793_,
		_w10795_,
		_w10798_
	);
	LUT4 #(
		.INIT('ha820)
	) name6751 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 ,
		_w10799_
	);
	LUT4 #(
		.INIT('h3120)
	) name6752 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10723_,
		_w10799_,
		_w10800_
	);
	LUT2 #(
		.INIT('h6)
	) name6753 (
		_w10798_,
		_w10800_,
		_w10801_
	);
	LUT3 #(
		.INIT('h54)
	) name6754 (
		_w10728_,
		_w10729_,
		_w10731_,
		_w10802_
	);
	LUT4 #(
		.INIT('h6996)
	) name6755 (
		_w10780_,
		_w10791_,
		_w10801_,
		_w10802_,
		_w10803_
	);
	LUT2 #(
		.INIT('h9)
	) name6756 (
		_w10779_,
		_w10803_,
		_w10804_
	);
	LUT4 #(
		.INIT('h6086)
	) name6757 (
		_w10722_,
		_w10732_,
		_w10733_,
		_w10746_,
		_w10805_
	);
	LUT3 #(
		.INIT('h0e)
	) name6758 (
		_w10721_,
		_w10747_,
		_w10805_,
		_w10806_
	);
	LUT4 #(
		.INIT('hb1b0)
	) name6759 (
		_w9973_,
		_w10655_,
		_w10656_,
		_w10657_,
		_w10807_
	);
	LUT3 #(
		.INIT('h7e)
	) name6760 (
		_w9954_,
		_w9961_,
		_w9969_,
		_w10808_
	);
	LUT3 #(
		.INIT('h4b)
	) name6761 (
		_w9973_,
		_w10657_,
		_w10808_,
		_w10809_
	);
	LUT2 #(
		.INIT('h2)
	) name6762 (
		_w10807_,
		_w10809_,
		_w10810_
	);
	LUT2 #(
		.INIT('h4)
	) name6763 (
		_w10807_,
		_w10809_,
		_w10811_
	);
	LUT2 #(
		.INIT('h9)
	) name6764 (
		_w10807_,
		_w10809_,
		_w10812_
	);
	LUT3 #(
		.INIT('h69)
	) name6765 (
		_w10804_,
		_w10806_,
		_w10812_,
		_w10813_
	);
	LUT2 #(
		.INIT('h9)
	) name6766 (
		_w10778_,
		_w10813_,
		_w10814_
	);
	LUT4 #(
		.INIT('h5100)
	) name6767 (
		_w9973_,
		_w10666_,
		_w10667_,
		_w10670_,
		_w10815_
	);
	LUT3 #(
		.INIT('h0b)
	) name6768 (
		_w10668_,
		_w10671_,
		_w10815_,
		_w10816_
	);
	LUT2 #(
		.INIT('h2)
	) name6769 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9956_,
		_w10817_
	);
	LUT2 #(
		.INIT('h1)
	) name6770 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9955_,
		_w10818_
	);
	LUT3 #(
		.INIT('h1b)
	) name6771 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9958_,
		_w9959_,
		_w10819_
	);
	LUT3 #(
		.INIT('h10)
	) name6772 (
		_w10818_,
		_w10817_,
		_w10819_,
		_w10820_
	);
	LUT2 #(
		.INIT('h2)
	) name6773 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9964_,
		_w10821_
	);
	LUT2 #(
		.INIT('h1)
	) name6774 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9963_,
		_w10822_
	);
	LUT3 #(
		.INIT('h1b)
	) name6775 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9966_,
		_w9967_,
		_w10823_
	);
	LUT3 #(
		.INIT('h10)
	) name6776 (
		_w10822_,
		_w10821_,
		_w10823_,
		_w10824_
	);
	LUT3 #(
		.INIT('he8)
	) name6777 (
		_w9954_,
		_w10820_,
		_w10824_,
		_w10825_
	);
	LUT4 #(
		.INIT('h7888)
	) name6778 (
		_w9950_,
		_w9953_,
		_w9957_,
		_w10660_,
		_w10826_
	);
	LUT2 #(
		.INIT('h9)
	) name6779 (
		_w10665_,
		_w10826_,
		_w10827_
	);
	LUT2 #(
		.INIT('h2)
	) name6780 (
		_w10825_,
		_w10827_,
		_w10828_
	);
	LUT3 #(
		.INIT('h51)
	) name6781 (
		_w9973_,
		_w10825_,
		_w10827_,
		_w10829_
	);
	LUT2 #(
		.INIT('h9)
	) name6782 (
		_w10666_,
		_w10667_,
		_w10830_
	);
	LUT3 #(
		.INIT('h96)
	) name6783 (
		_w9973_,
		_w10666_,
		_w10667_,
		_w10831_
	);
	LUT3 #(
		.INIT('h49)
	) name6784 (
		_w9973_,
		_w10666_,
		_w10667_,
		_w10832_
	);
	LUT3 #(
		.INIT('h0b)
	) name6785 (
		_w10829_,
		_w10831_,
		_w10832_,
		_w10833_
	);
	LUT2 #(
		.INIT('h9)
	) name6786 (
		_w10774_,
		_w10775_,
		_w10834_
	);
	LUT4 #(
		.INIT('h4800)
	) name6787 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10835_
	);
	LUT2 #(
		.INIT('h2)
	) name6788 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w10002_,
		_w10836_
	);
	LUT2 #(
		.INIT('h1)
	) name6789 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w10001_,
		_w10837_
	);
	LUT3 #(
		.INIT('h1b)
	) name6790 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w10004_,
		_w10005_,
		_w10838_
	);
	LUT4 #(
		.INIT('h0100)
	) name6791 (
		_w10835_,
		_w10837_,
		_w10836_,
		_w10838_,
		_w10839_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6792 (
		_w10835_,
		_w10837_,
		_w10836_,
		_w10838_,
		_w10840_
	);
	LUT4 #(
		.INIT('ha820)
	) name6793 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 ,
		_w10841_
	);
	LUT4 #(
		.INIT('h3210)
	) name6794 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10751_,
		_w10841_,
		_w10842_
	);
	LUT3 #(
		.INIT('h54)
	) name6795 (
		_w10839_,
		_w10840_,
		_w10842_,
		_w10843_
	);
	LUT4 #(
		.INIT('h5655)
	) name6796 (
		_w10752_,
		_w10754_,
		_w10753_,
		_w10755_,
		_w10844_
	);
	LUT2 #(
		.INIT('h9)
	) name6797 (
		_w10758_,
		_w10844_,
		_w10845_
	);
	LUT2 #(
		.INIT('h2)
	) name6798 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9976_,
		_w10846_
	);
	LUT2 #(
		.INIT('h1)
	) name6799 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9975_,
		_w10847_
	);
	LUT3 #(
		.INIT('h1b)
	) name6800 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9978_,
		_w9979_,
		_w10848_
	);
	LUT3 #(
		.INIT('h10)
	) name6801 (
		_w10847_,
		_w10846_,
		_w10848_,
		_w10849_
	);
	LUT2 #(
		.INIT('h2)
	) name6802 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9983_,
		_w10850_
	);
	LUT2 #(
		.INIT('h1)
	) name6803 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9982_,
		_w10851_
	);
	LUT3 #(
		.INIT('h1b)
	) name6804 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9985_,
		_w9986_,
		_w10852_
	);
	LUT3 #(
		.INIT('h10)
	) name6805 (
		_w10851_,
		_w10850_,
		_w10852_,
		_w10853_
	);
	LUT2 #(
		.INIT('h2)
	) name6806 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9991_,
		_w10854_
	);
	LUT2 #(
		.INIT('h1)
	) name6807 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9990_,
		_w10855_
	);
	LUT3 #(
		.INIT('h1b)
	) name6808 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9993_,
		_w9994_,
		_w10856_
	);
	LUT3 #(
		.INIT('h10)
	) name6809 (
		_w10855_,
		_w10854_,
		_w10856_,
		_w10857_
	);
	LUT3 #(
		.INIT('he8)
	) name6810 (
		_w10849_,
		_w10853_,
		_w10857_,
		_w10858_
	);
	LUT3 #(
		.INIT('h69)
	) name6811 (
		_w10763_,
		_w10767_,
		_w10771_,
		_w10859_
	);
	LUT4 #(
		.INIT('hee0e)
	) name6812 (
		_w10843_,
		_w10845_,
		_w10858_,
		_w10859_,
		_w10860_
	);
	LUT4 #(
		.INIT('h6996)
	) name6813 (
		_w10750_,
		_w10759_,
		_w10772_,
		_w10773_,
		_w10861_
	);
	LUT4 #(
		.INIT('h6086)
	) name6814 (
		_w10750_,
		_w10759_,
		_w10772_,
		_w10773_,
		_w10862_
	);
	LUT3 #(
		.INIT('h0e)
	) name6815 (
		_w10860_,
		_w10861_,
		_w10862_,
		_w10863_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name6816 (
		_w10816_,
		_w10833_,
		_w10834_,
		_w10863_,
		_w10864_
	);
	LUT4 #(
		.INIT('h559a)
	) name6817 (
		_w10659_,
		_w10668_,
		_w10671_,
		_w10672_,
		_w10865_
	);
	LUT3 #(
		.INIT('h69)
	) name6818 (
		_w10748_,
		_w10777_,
		_w10865_,
		_w10866_
	);
	LUT4 #(
		.INIT('h0640)
	) name6819 (
		_w10659_,
		_w10673_,
		_w10748_,
		_w10777_,
		_w10867_
	);
	LUT3 #(
		.INIT('h07)
	) name6820 (
		_w10864_,
		_w10866_,
		_w10867_,
		_w10868_
	);
	LUT2 #(
		.INIT('h6)
	) name6821 (
		_w10864_,
		_w10866_,
		_w10869_
	);
	LUT2 #(
		.INIT('h6)
	) name6822 (
		_w10860_,
		_w10861_,
		_w10870_
	);
	LUT2 #(
		.INIT('h2)
	) name6823 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9976_,
		_w10871_
	);
	LUT2 #(
		.INIT('h1)
	) name6824 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9975_,
		_w10872_
	);
	LUT3 #(
		.INIT('h1b)
	) name6825 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9978_,
		_w9979_,
		_w10873_
	);
	LUT3 #(
		.INIT('h10)
	) name6826 (
		_w10872_,
		_w10871_,
		_w10873_,
		_w10874_
	);
	LUT2 #(
		.INIT('h2)
	) name6827 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9983_,
		_w10875_
	);
	LUT2 #(
		.INIT('h1)
	) name6828 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9982_,
		_w10876_
	);
	LUT3 #(
		.INIT('h1b)
	) name6829 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9985_,
		_w9986_,
		_w10877_
	);
	LUT3 #(
		.INIT('h10)
	) name6830 (
		_w10876_,
		_w10875_,
		_w10877_,
		_w10878_
	);
	LUT2 #(
		.INIT('h2)
	) name6831 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9991_,
		_w10879_
	);
	LUT2 #(
		.INIT('h1)
	) name6832 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9990_,
		_w10880_
	);
	LUT3 #(
		.INIT('h1b)
	) name6833 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9993_,
		_w9994_,
		_w10881_
	);
	LUT3 #(
		.INIT('h10)
	) name6834 (
		_w10880_,
		_w10879_,
		_w10881_,
		_w10882_
	);
	LUT3 #(
		.INIT('he8)
	) name6835 (
		_w10874_,
		_w10878_,
		_w10882_,
		_w10883_
	);
	LUT3 #(
		.INIT('h69)
	) name6836 (
		_w10849_,
		_w10853_,
		_w10857_,
		_w10884_
	);
	LUT4 #(
		.INIT('h5655)
	) name6837 (
		_w10835_,
		_w10837_,
		_w10836_,
		_w10838_,
		_w10885_
	);
	LUT2 #(
		.INIT('h9)
	) name6838 (
		_w10842_,
		_w10885_,
		_w10886_
	);
	LUT4 #(
		.INIT('ha820)
	) name6839 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 ,
		_w10887_
	);
	LUT4 #(
		.INIT('h3210)
	) name6840 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10841_,
		_w10887_,
		_w10888_
	);
	LUT2 #(
		.INIT('h2)
	) name6841 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w10002_,
		_w10889_
	);
	LUT2 #(
		.INIT('h1)
	) name6842 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w10001_,
		_w10890_
	);
	LUT3 #(
		.INIT('h1b)
	) name6843 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w10004_,
		_w10005_,
		_w10891_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6844 (
		_w10888_,
		_w10890_,
		_w10889_,
		_w10891_,
		_w10892_
	);
	LUT4 #(
		.INIT('h0100)
	) name6845 (
		_w10888_,
		_w10890_,
		_w10889_,
		_w10891_,
		_w10893_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name6846 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10894_
	);
	LUT3 #(
		.INIT('h54)
	) name6847 (
		_w10892_,
		_w10893_,
		_w10894_,
		_w10895_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name6848 (
		_w10883_,
		_w10884_,
		_w10886_,
		_w10895_,
		_w10896_
	);
	LUT4 #(
		.INIT('h6996)
	) name6849 (
		_w10843_,
		_w10845_,
		_w10858_,
		_w10859_,
		_w10897_
	);
	LUT4 #(
		.INIT('h0980)
	) name6850 (
		_w10843_,
		_w10845_,
		_w10858_,
		_w10859_,
		_w10898_
	);
	LUT3 #(
		.INIT('h0d)
	) name6851 (
		_w10896_,
		_w10897_,
		_w10898_,
		_w10899_
	);
	LUT2 #(
		.INIT('h2)
	) name6852 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9964_,
		_w10900_
	);
	LUT2 #(
		.INIT('h1)
	) name6853 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9963_,
		_w10901_
	);
	LUT3 #(
		.INIT('h1b)
	) name6854 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9966_,
		_w9967_,
		_w10902_
	);
	LUT3 #(
		.INIT('h10)
	) name6855 (
		_w10901_,
		_w10900_,
		_w10902_,
		_w10903_
	);
	LUT2 #(
		.INIT('h2)
	) name6856 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9956_,
		_w10904_
	);
	LUT2 #(
		.INIT('h1)
	) name6857 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9955_,
		_w10905_
	);
	LUT3 #(
		.INIT('h1b)
	) name6858 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9958_,
		_w9959_,
		_w10906_
	);
	LUT3 #(
		.INIT('h10)
	) name6859 (
		_w10905_,
		_w10904_,
		_w10906_,
		_w10907_
	);
	LUT3 #(
		.INIT('h1b)
	) name6860 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9951_,
		_w9952_,
		_w10908_
	);
	LUT2 #(
		.INIT('h8)
	) name6861 (
		_w9950_,
		_w10908_,
		_w10909_
	);
	LUT3 #(
		.INIT('he8)
	) name6862 (
		_w10903_,
		_w10907_,
		_w10909_,
		_w10910_
	);
	LUT3 #(
		.INIT('h69)
	) name6863 (
		_w9954_,
		_w10820_,
		_w10824_,
		_w10911_
	);
	LUT3 #(
		.INIT('h51)
	) name6864 (
		_w9973_,
		_w10910_,
		_w10911_,
		_w10912_
	);
	LUT2 #(
		.INIT('h9)
	) name6865 (
		_w10825_,
		_w10827_,
		_w10913_
	);
	LUT3 #(
		.INIT('h96)
	) name6866 (
		_w9973_,
		_w10825_,
		_w10827_,
		_w10914_
	);
	LUT3 #(
		.INIT('h49)
	) name6867 (
		_w9973_,
		_w10825_,
		_w10827_,
		_w10915_
	);
	LUT3 #(
		.INIT('h0b)
	) name6868 (
		_w10912_,
		_w10914_,
		_w10915_,
		_w10916_
	);
	LUT3 #(
		.INIT('h4b)
	) name6869 (
		_w9973_,
		_w10828_,
		_w10830_,
		_w10917_
	);
	LUT4 #(
		.INIT('h7077)
	) name6870 (
		_w10870_,
		_w10899_,
		_w10916_,
		_w10917_,
		_w10918_
	);
	LUT4 #(
		.INIT('h6996)
	) name6871 (
		_w10816_,
		_w10833_,
		_w10834_,
		_w10863_,
		_w10919_
	);
	LUT4 #(
		.INIT('h9029)
	) name6872 (
		_w10816_,
		_w10833_,
		_w10834_,
		_w10863_,
		_w10920_
	);
	LUT3 #(
		.INIT('h0b)
	) name6873 (
		_w10918_,
		_w10919_,
		_w10920_,
		_w10921_
	);
	LUT2 #(
		.INIT('h1)
	) name6874 (
		_w10869_,
		_w10921_,
		_w10922_
	);
	LUT4 #(
		.INIT('h7770)
	) name6875 (
		_w10814_,
		_w10868_,
		_w10869_,
		_w10921_,
		_w10923_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name6876 (
		_w10780_,
		_w10791_,
		_w10801_,
		_w10802_,
		_w10924_
	);
	LUT3 #(
		.INIT('he8)
	) name6877 (
		_w10782_,
		_w10786_,
		_w10790_,
		_w10925_
	);
	LUT2 #(
		.INIT('h2)
	) name6878 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9991_,
		_w10926_
	);
	LUT2 #(
		.INIT('h1)
	) name6879 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9990_,
		_w10927_
	);
	LUT3 #(
		.INIT('h1b)
	) name6880 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9993_,
		_w9994_,
		_w10928_
	);
	LUT3 #(
		.INIT('h10)
	) name6881 (
		_w10927_,
		_w10926_,
		_w10928_,
		_w10929_
	);
	LUT2 #(
		.INIT('h1)
	) name6882 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9982_,
		_w10930_
	);
	LUT2 #(
		.INIT('h2)
	) name6883 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9983_,
		_w10931_
	);
	LUT3 #(
		.INIT('h1b)
	) name6884 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9985_,
		_w9986_,
		_w10932_
	);
	LUT3 #(
		.INIT('h10)
	) name6885 (
		_w10931_,
		_w10930_,
		_w10932_,
		_w10933_
	);
	LUT3 #(
		.INIT('h69)
	) name6886 (
		_w9981_,
		_w10929_,
		_w10933_,
		_w10934_
	);
	LUT4 #(
		.INIT('h4800)
	) name6887 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w10935_
	);
	LUT2 #(
		.INIT('h2)
	) name6888 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w10002_,
		_w10936_
	);
	LUT2 #(
		.INIT('h1)
	) name6889 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w10001_,
		_w10937_
	);
	LUT3 #(
		.INIT('h1b)
	) name6890 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w10004_,
		_w10005_,
		_w10938_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6891 (
		_w10935_,
		_w10937_,
		_w10936_,
		_w10938_,
		_w10939_
	);
	LUT4 #(
		.INIT('h0100)
	) name6892 (
		_w10935_,
		_w10937_,
		_w10936_,
		_w10938_,
		_w10940_
	);
	LUT4 #(
		.INIT('h5655)
	) name6893 (
		_w10935_,
		_w10937_,
		_w10936_,
		_w10938_,
		_w10941_
	);
	LUT4 #(
		.INIT('h3210)
	) name6894 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10138_,
		_w10799_,
		_w10942_
	);
	LUT2 #(
		.INIT('h9)
	) name6895 (
		_w10941_,
		_w10942_,
		_w10943_
	);
	LUT3 #(
		.INIT('h54)
	) name6896 (
		_w10796_,
		_w10797_,
		_w10800_,
		_w10944_
	);
	LUT4 #(
		.INIT('h6996)
	) name6897 (
		_w10925_,
		_w10934_,
		_w10943_,
		_w10944_,
		_w10945_
	);
	LUT2 #(
		.INIT('h9)
	) name6898 (
		_w10924_,
		_w10945_,
		_w10946_
	);
	LUT4 #(
		.INIT('h9209)
	) name6899 (
		_w10780_,
		_w10791_,
		_w10801_,
		_w10802_,
		_w10947_
	);
	LUT3 #(
		.INIT('h0b)
	) name6900 (
		_w10779_,
		_w10803_,
		_w10947_,
		_w10948_
	);
	LUT2 #(
		.INIT('h2)
	) name6901 (
		_w10946_,
		_w10948_,
		_w10949_
	);
	LUT3 #(
		.INIT('h51)
	) name6902 (
		_w9974_,
		_w10946_,
		_w10948_,
		_w10950_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name6903 (
		_w10925_,
		_w10934_,
		_w10943_,
		_w10944_,
		_w10951_
	);
	LUT3 #(
		.INIT('he8)
	) name6904 (
		_w9981_,
		_w10929_,
		_w10933_,
		_w10952_
	);
	LUT3 #(
		.INIT('h69)
	) name6905 (
		_w9981_,
		_w10150_,
		_w10152_,
		_w10953_
	);
	LUT4 #(
		.INIT('h5655)
	) name6906 (
		_w10139_,
		_w10141_,
		_w10140_,
		_w10142_,
		_w10954_
	);
	LUT2 #(
		.INIT('h9)
	) name6907 (
		_w10145_,
		_w10954_,
		_w10955_
	);
	LUT3 #(
		.INIT('h45)
	) name6908 (
		_w10939_,
		_w10940_,
		_w10942_,
		_w10956_
	);
	LUT4 #(
		.INIT('h6996)
	) name6909 (
		_w10952_,
		_w10953_,
		_w10955_,
		_w10956_,
		_w10957_
	);
	LUT2 #(
		.INIT('h9)
	) name6910 (
		_w10951_,
		_w10957_,
		_w10958_
	);
	LUT4 #(
		.INIT('h9029)
	) name6911 (
		_w10925_,
		_w10934_,
		_w10943_,
		_w10944_,
		_w10959_
	);
	LUT3 #(
		.INIT('h0b)
	) name6912 (
		_w10924_,
		_w10945_,
		_w10959_,
		_w10960_
	);
	LUT2 #(
		.INIT('h2)
	) name6913 (
		_w10958_,
		_w10960_,
		_w10961_
	);
	LUT2 #(
		.INIT('h9)
	) name6914 (
		_w10958_,
		_w10960_,
		_w10962_
	);
	LUT3 #(
		.INIT('h69)
	) name6915 (
		_w9974_,
		_w10958_,
		_w10960_,
		_w10963_
	);
	LUT3 #(
		.INIT('h4b)
	) name6916 (
		_w9974_,
		_w10949_,
		_w10962_,
		_w10964_
	);
	LUT3 #(
		.INIT('h0d)
	) name6917 (
		_w10804_,
		_w10806_,
		_w10811_,
		_w10965_
	);
	LUT3 #(
		.INIT('h69)
	) name6918 (
		_w9974_,
		_w10946_,
		_w10948_,
		_w10966_
	);
	LUT2 #(
		.INIT('h6)
	) name6919 (
		_w10965_,
		_w10966_,
		_w10967_
	);
	LUT4 #(
		.INIT('h0209)
	) name6920 (
		_w10804_,
		_w10806_,
		_w10810_,
		_w10811_,
		_w10968_
	);
	LUT3 #(
		.INIT('h0b)
	) name6921 (
		_w10778_,
		_w10813_,
		_w10968_,
		_w10969_
	);
	LUT2 #(
		.INIT('h2)
	) name6922 (
		_w10967_,
		_w10969_,
		_w10970_
	);
	LUT3 #(
		.INIT('h49)
	) name6923 (
		_w9974_,
		_w10946_,
		_w10948_,
		_w10971_
	);
	LUT3 #(
		.INIT('h0e)
	) name6924 (
		_w10965_,
		_w10966_,
		_w10971_,
		_w10972_
	);
	LUT4 #(
		.INIT('h0eae)
	) name6925 (
		_w10964_,
		_w10967_,
		_w10969_,
		_w10972_,
		_w10973_
	);
	LUT2 #(
		.INIT('h2)
	) name6926 (
		_w10923_,
		_w10973_,
		_w10974_
	);
	LUT2 #(
		.INIT('h2)
	) name6927 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9956_,
		_w10975_
	);
	LUT2 #(
		.INIT('h1)
	) name6928 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9955_,
		_w10976_
	);
	LUT3 #(
		.INIT('h1b)
	) name6929 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9958_,
		_w9959_,
		_w10977_
	);
	LUT3 #(
		.INIT('h10)
	) name6930 (
		_w10976_,
		_w10975_,
		_w10977_,
		_w10978_
	);
	LUT2 #(
		.INIT('h2)
	) name6931 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9949_,
		_w10979_
	);
	LUT2 #(
		.INIT('h1)
	) name6932 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w9948_,
		_w10980_
	);
	LUT3 #(
		.INIT('h1b)
	) name6933 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9951_,
		_w9952_,
		_w10981_
	);
	LUT3 #(
		.INIT('h10)
	) name6934 (
		_w10980_,
		_w10979_,
		_w10981_,
		_w10982_
	);
	LUT2 #(
		.INIT('h2)
	) name6935 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9964_,
		_w10983_
	);
	LUT2 #(
		.INIT('h1)
	) name6936 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9963_,
		_w10984_
	);
	LUT3 #(
		.INIT('h1b)
	) name6937 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9966_,
		_w9967_,
		_w10985_
	);
	LUT3 #(
		.INIT('h10)
	) name6938 (
		_w10984_,
		_w10983_,
		_w10985_,
		_w10986_
	);
	LUT3 #(
		.INIT('he8)
	) name6939 (
		_w10978_,
		_w10982_,
		_w10986_,
		_w10987_
	);
	LUT3 #(
		.INIT('h69)
	) name6940 (
		_w10903_,
		_w10907_,
		_w10909_,
		_w10988_
	);
	LUT2 #(
		.INIT('h2)
	) name6941 (
		_w10987_,
		_w10988_,
		_w10989_
	);
	LUT3 #(
		.INIT('h51)
	) name6942 (
		_w9973_,
		_w10987_,
		_w10988_,
		_w10990_
	);
	LUT2 #(
		.INIT('h9)
	) name6943 (
		_w10910_,
		_w10911_,
		_w10991_
	);
	LUT3 #(
		.INIT('h96)
	) name6944 (
		_w9973_,
		_w10910_,
		_w10911_,
		_w10992_
	);
	LUT3 #(
		.INIT('h4b)
	) name6945 (
		_w9973_,
		_w10989_,
		_w10991_,
		_w10993_
	);
	LUT2 #(
		.INIT('h2)
	) name6946 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9956_,
		_w10994_
	);
	LUT2 #(
		.INIT('h1)
	) name6947 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9955_,
		_w10995_
	);
	LUT3 #(
		.INIT('h1b)
	) name6948 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9958_,
		_w9959_,
		_w10996_
	);
	LUT3 #(
		.INIT('h10)
	) name6949 (
		_w10995_,
		_w10994_,
		_w10996_,
		_w10997_
	);
	LUT2 #(
		.INIT('h2)
	) name6950 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9949_,
		_w10998_
	);
	LUT2 #(
		.INIT('h1)
	) name6951 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w9948_,
		_w10999_
	);
	LUT3 #(
		.INIT('h1b)
	) name6952 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9951_,
		_w9952_,
		_w11000_
	);
	LUT3 #(
		.INIT('h10)
	) name6953 (
		_w10999_,
		_w10998_,
		_w11000_,
		_w11001_
	);
	LUT2 #(
		.INIT('h2)
	) name6954 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9964_,
		_w11002_
	);
	LUT2 #(
		.INIT('h1)
	) name6955 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9963_,
		_w11003_
	);
	LUT3 #(
		.INIT('h1b)
	) name6956 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9966_,
		_w9967_,
		_w11004_
	);
	LUT3 #(
		.INIT('h10)
	) name6957 (
		_w11003_,
		_w11002_,
		_w11004_,
		_w11005_
	);
	LUT3 #(
		.INIT('he8)
	) name6958 (
		_w10997_,
		_w11001_,
		_w11005_,
		_w11006_
	);
	LUT3 #(
		.INIT('h69)
	) name6959 (
		_w10978_,
		_w10982_,
		_w10986_,
		_w11007_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6960 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w11008_
	);
	LUT4 #(
		.INIT('he400)
	) name6961 (
		_w9947_,
		_w9970_,
		_w9971_,
		_w11008_,
		_w11009_
	);
	LUT3 #(
		.INIT('ha2)
	) name6962 (
		_w9973_,
		_w10008_,
		_w11009_,
		_w11010_
	);
	LUT3 #(
		.INIT('h0d)
	) name6963 (
		_w11006_,
		_w11007_,
		_w11010_,
		_w11011_
	);
	LUT3 #(
		.INIT('h96)
	) name6964 (
		_w9973_,
		_w10987_,
		_w10988_,
		_w11012_
	);
	LUT3 #(
		.INIT('h20)
	) name6965 (
		_w9973_,
		_w10987_,
		_w10988_,
		_w11013_
	);
	LUT3 #(
		.INIT('h07)
	) name6966 (
		_w11011_,
		_w11012_,
		_w11013_,
		_w11014_
	);
	LUT2 #(
		.INIT('h2)
	) name6967 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9976_,
		_w11015_
	);
	LUT2 #(
		.INIT('h1)
	) name6968 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9975_,
		_w11016_
	);
	LUT3 #(
		.INIT('h1b)
	) name6969 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9978_,
		_w9979_,
		_w11017_
	);
	LUT3 #(
		.INIT('h10)
	) name6970 (
		_w11016_,
		_w11015_,
		_w11017_,
		_w11018_
	);
	LUT2 #(
		.INIT('h2)
	) name6971 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9991_,
		_w11019_
	);
	LUT2 #(
		.INIT('h1)
	) name6972 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9990_,
		_w11020_
	);
	LUT3 #(
		.INIT('h1b)
	) name6973 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9993_,
		_w9994_,
		_w11021_
	);
	LUT3 #(
		.INIT('h10)
	) name6974 (
		_w11020_,
		_w11019_,
		_w11021_,
		_w11022_
	);
	LUT2 #(
		.INIT('h2)
	) name6975 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9983_,
		_w11023_
	);
	LUT2 #(
		.INIT('h1)
	) name6976 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9982_,
		_w11024_
	);
	LUT3 #(
		.INIT('h1b)
	) name6977 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9985_,
		_w9986_,
		_w11025_
	);
	LUT3 #(
		.INIT('h10)
	) name6978 (
		_w11024_,
		_w11023_,
		_w11025_,
		_w11026_
	);
	LUT3 #(
		.INIT('he8)
	) name6979 (
		_w11018_,
		_w11022_,
		_w11026_,
		_w11027_
	);
	LUT3 #(
		.INIT('h69)
	) name6980 (
		_w10874_,
		_w10878_,
		_w10882_,
		_w11028_
	);
	LUT4 #(
		.INIT('h5655)
	) name6981 (
		_w10888_,
		_w10890_,
		_w10889_,
		_w10891_,
		_w11029_
	);
	LUT2 #(
		.INIT('h9)
	) name6982 (
		_w10894_,
		_w11029_,
		_w11030_
	);
	LUT4 #(
		.INIT('ha820)
	) name6983 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 ,
		_w11031_
	);
	LUT4 #(
		.INIT('h3210)
	) name6984 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10887_,
		_w11031_,
		_w11032_
	);
	LUT2 #(
		.INIT('h2)
	) name6985 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w10002_,
		_w11033_
	);
	LUT2 #(
		.INIT('h1)
	) name6986 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w10001_,
		_w11034_
	);
	LUT3 #(
		.INIT('h1b)
	) name6987 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w10004_,
		_w10005_,
		_w11035_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6988 (
		_w11032_,
		_w11034_,
		_w11033_,
		_w11035_,
		_w11036_
	);
	LUT4 #(
		.INIT('h0100)
	) name6989 (
		_w11032_,
		_w11034_,
		_w11033_,
		_w11035_,
		_w11037_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name6990 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w11038_
	);
	LUT3 #(
		.INIT('h54)
	) name6991 (
		_w11036_,
		_w11037_,
		_w11038_,
		_w11039_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name6992 (
		_w11027_,
		_w11028_,
		_w11030_,
		_w11039_,
		_w11040_
	);
	LUT4 #(
		.INIT('h9669)
	) name6993 (
		_w10883_,
		_w10884_,
		_w10886_,
		_w10895_,
		_w11041_
	);
	LUT2 #(
		.INIT('h9)
	) name6994 (
		_w11040_,
		_w11041_,
		_w11042_
	);
	LUT2 #(
		.INIT('h2)
	) name6995 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9983_,
		_w11043_
	);
	LUT2 #(
		.INIT('h1)
	) name6996 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9982_,
		_w11044_
	);
	LUT3 #(
		.INIT('h1b)
	) name6997 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9985_,
		_w9986_,
		_w11045_
	);
	LUT3 #(
		.INIT('h10)
	) name6998 (
		_w11044_,
		_w11043_,
		_w11045_,
		_w11046_
	);
	LUT2 #(
		.INIT('h2)
	) name6999 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9976_,
		_w11047_
	);
	LUT2 #(
		.INIT('h1)
	) name7000 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9975_,
		_w11048_
	);
	LUT3 #(
		.INIT('h1b)
	) name7001 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9978_,
		_w9979_,
		_w11049_
	);
	LUT3 #(
		.INIT('h10)
	) name7002 (
		_w11048_,
		_w11047_,
		_w11049_,
		_w11050_
	);
	LUT2 #(
		.INIT('h2)
	) name7003 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9991_,
		_w11051_
	);
	LUT2 #(
		.INIT('h1)
	) name7004 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9990_,
		_w11052_
	);
	LUT3 #(
		.INIT('h1b)
	) name7005 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9993_,
		_w9994_,
		_w11053_
	);
	LUT3 #(
		.INIT('h10)
	) name7006 (
		_w11052_,
		_w11051_,
		_w11053_,
		_w11054_
	);
	LUT3 #(
		.INIT('he8)
	) name7007 (
		_w11046_,
		_w11050_,
		_w11054_,
		_w11055_
	);
	LUT3 #(
		.INIT('h69)
	) name7008 (
		_w11018_,
		_w11022_,
		_w11026_,
		_w11056_
	);
	LUT4 #(
		.INIT('h5655)
	) name7009 (
		_w11032_,
		_w11034_,
		_w11033_,
		_w11035_,
		_w11057_
	);
	LUT2 #(
		.INIT('h9)
	) name7010 (
		_w11038_,
		_w11057_,
		_w11058_
	);
	LUT4 #(
		.INIT('ha820)
	) name7011 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 ,
		_w11059_
	);
	LUT4 #(
		.INIT('h3210)
	) name7012 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w11031_,
		_w11059_,
		_w11060_
	);
	LUT2 #(
		.INIT('h2)
	) name7013 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w10002_,
		_w11061_
	);
	LUT2 #(
		.INIT('h1)
	) name7014 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w10001_,
		_w11062_
	);
	LUT3 #(
		.INIT('h1b)
	) name7015 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w10004_,
		_w10005_,
		_w11063_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7016 (
		_w11060_,
		_w11062_,
		_w11061_,
		_w11063_,
		_w11064_
	);
	LUT4 #(
		.INIT('h0100)
	) name7017 (
		_w11060_,
		_w11062_,
		_w11061_,
		_w11063_,
		_w11065_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name7018 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w11066_
	);
	LUT3 #(
		.INIT('h54)
	) name7019 (
		_w11064_,
		_w11065_,
		_w11066_,
		_w11067_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name7020 (
		_w11055_,
		_w11056_,
		_w11058_,
		_w11067_,
		_w11068_
	);
	LUT4 #(
		.INIT('h6996)
	) name7021 (
		_w11027_,
		_w11028_,
		_w11030_,
		_w11039_,
		_w11069_
	);
	LUT4 #(
		.INIT('h9209)
	) name7022 (
		_w11027_,
		_w11028_,
		_w11030_,
		_w11039_,
		_w11070_
	);
	LUT3 #(
		.INIT('h0b)
	) name7023 (
		_w11068_,
		_w11069_,
		_w11070_,
		_w11071_
	);
	LUT4 #(
		.INIT('h7707)
	) name7024 (
		_w10993_,
		_w11014_,
		_w11042_,
		_w11071_,
		_w11072_
	);
	LUT2 #(
		.INIT('h9)
	) name7025 (
		_w10896_,
		_w10897_,
		_w11073_
	);
	LUT4 #(
		.INIT('h2990)
	) name7026 (
		_w10883_,
		_w10884_,
		_w10886_,
		_w10895_,
		_w11074_
	);
	LUT3 #(
		.INIT('h0b)
	) name7027 (
		_w11040_,
		_w11041_,
		_w11074_,
		_w11075_
	);
	LUT3 #(
		.INIT('h27)
	) name7028 (
		_w10912_,
		_w10913_,
		_w10914_,
		_w11076_
	);
	LUT3 #(
		.INIT('h49)
	) name7029 (
		_w9973_,
		_w10910_,
		_w10911_,
		_w11077_
	);
	LUT3 #(
		.INIT('h0b)
	) name7030 (
		_w10990_,
		_w10992_,
		_w11077_,
		_w11078_
	);
	LUT4 #(
		.INIT('h9669)
	) name7031 (
		_w11073_,
		_w11075_,
		_w11076_,
		_w11078_,
		_w11079_
	);
	LUT2 #(
		.INIT('h6)
	) name7032 (
		_w11072_,
		_w11079_,
		_w11080_
	);
	LUT2 #(
		.INIT('h9)
	) name7033 (
		_w11068_,
		_w11069_,
		_w11081_
	);
	LUT2 #(
		.INIT('h8)
	) name7034 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 ,
		_w11082_
	);
	LUT2 #(
		.INIT('h1)
	) name7035 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w11083_
	);
	LUT3 #(
		.INIT('h13)
	) name7036 (
		_w11059_,
		_w11082_,
		_w11083_,
		_w11084_
	);
	LUT2 #(
		.INIT('h1)
	) name7037 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w10001_,
		_w11085_
	);
	LUT2 #(
		.INIT('h2)
	) name7038 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w10002_,
		_w11086_
	);
	LUT3 #(
		.INIT('h1b)
	) name7039 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w10004_,
		_w10005_,
		_w11087_
	);
	LUT4 #(
		.INIT('h5455)
	) name7040 (
		_w11084_,
		_w11086_,
		_w11085_,
		_w11087_,
		_w11088_
	);
	LUT4 #(
		.INIT('h5655)
	) name7041 (
		_w11060_,
		_w11062_,
		_w11061_,
		_w11063_,
		_w11089_
	);
	LUT2 #(
		.INIT('h9)
	) name7042 (
		_w11066_,
		_w11089_,
		_w11090_
	);
	LUT3 #(
		.INIT('h12)
	) name7043 (
		_w11066_,
		_w11088_,
		_w11089_,
		_w11091_
	);
	LUT2 #(
		.INIT('h2)
	) name7044 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9983_,
		_w11092_
	);
	LUT2 #(
		.INIT('h1)
	) name7045 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w9982_,
		_w11093_
	);
	LUT3 #(
		.INIT('h1b)
	) name7046 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w9985_,
		_w9986_,
		_w11094_
	);
	LUT3 #(
		.INIT('h10)
	) name7047 (
		_w11093_,
		_w11092_,
		_w11094_,
		_w11095_
	);
	LUT2 #(
		.INIT('h2)
	) name7048 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9976_,
		_w11096_
	);
	LUT2 #(
		.INIT('h1)
	) name7049 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w9975_,
		_w11097_
	);
	LUT3 #(
		.INIT('h1b)
	) name7050 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w9978_,
		_w9979_,
		_w11098_
	);
	LUT3 #(
		.INIT('h10)
	) name7051 (
		_w11097_,
		_w11096_,
		_w11098_,
		_w11099_
	);
	LUT2 #(
		.INIT('h2)
	) name7052 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9991_,
		_w11100_
	);
	LUT2 #(
		.INIT('h1)
	) name7053 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w9990_,
		_w11101_
	);
	LUT3 #(
		.INIT('h1b)
	) name7054 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w9993_,
		_w9994_,
		_w11102_
	);
	LUT3 #(
		.INIT('h10)
	) name7055 (
		_w11101_,
		_w11100_,
		_w11102_,
		_w11103_
	);
	LUT3 #(
		.INIT('he8)
	) name7056 (
		_w11095_,
		_w11099_,
		_w11103_,
		_w11104_
	);
	LUT3 #(
		.INIT('h69)
	) name7057 (
		_w11046_,
		_w11050_,
		_w11054_,
		_w11105_
	);
	LUT3 #(
		.INIT('h51)
	) name7058 (
		_w11091_,
		_w11104_,
		_w11105_,
		_w11106_
	);
	LUT4 #(
		.INIT('h9669)
	) name7059 (
		_w11055_,
		_w11056_,
		_w11058_,
		_w11067_,
		_w11107_
	);
	LUT4 #(
		.INIT('h0460)
	) name7060 (
		_w11055_,
		_w11056_,
		_w11058_,
		_w11067_,
		_w11108_
	);
	LUT3 #(
		.INIT('h0d)
	) name7061 (
		_w11106_,
		_w11107_,
		_w11108_,
		_w11109_
	);
	LUT2 #(
		.INIT('h6)
	) name7062 (
		_w11011_,
		_w11012_,
		_w11110_
	);
	LUT2 #(
		.INIT('h2)
	) name7063 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9956_,
		_w11111_
	);
	LUT2 #(
		.INIT('h1)
	) name7064 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w9955_,
		_w11112_
	);
	LUT3 #(
		.INIT('h1b)
	) name7065 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w9958_,
		_w9959_,
		_w11113_
	);
	LUT3 #(
		.INIT('h10)
	) name7066 (
		_w11112_,
		_w11111_,
		_w11113_,
		_w11114_
	);
	LUT2 #(
		.INIT('h2)
	) name7067 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9949_,
		_w11115_
	);
	LUT2 #(
		.INIT('h1)
	) name7068 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w9948_,
		_w11116_
	);
	LUT3 #(
		.INIT('h1b)
	) name7069 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w9951_,
		_w9952_,
		_w11117_
	);
	LUT3 #(
		.INIT('h10)
	) name7070 (
		_w11116_,
		_w11115_,
		_w11117_,
		_w11118_
	);
	LUT2 #(
		.INIT('h2)
	) name7071 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9964_,
		_w11119_
	);
	LUT2 #(
		.INIT('h1)
	) name7072 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w9963_,
		_w11120_
	);
	LUT3 #(
		.INIT('h1b)
	) name7073 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w9966_,
		_w9967_,
		_w11121_
	);
	LUT3 #(
		.INIT('h10)
	) name7074 (
		_w11120_,
		_w11119_,
		_w11121_,
		_w11122_
	);
	LUT3 #(
		.INIT('he8)
	) name7075 (
		_w11114_,
		_w11118_,
		_w11122_,
		_w11123_
	);
	LUT3 #(
		.INIT('h69)
	) name7076 (
		_w10997_,
		_w11001_,
		_w11005_,
		_w11124_
	);
	LUT2 #(
		.INIT('h9)
	) name7077 (
		_w10008_,
		_w11009_,
		_w11125_
	);
	LUT4 #(
		.INIT('h8040)
	) name7078 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w11126_
	);
	LUT4 #(
		.INIT('h1020)
	) name7079 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w11127_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name7080 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w11128_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7081 (
		_w10004_,
		_w11127_,
		_w11126_,
		_w11128_,
		_w11129_
	);
	LUT4 #(
		.INIT('h0100)
	) name7082 (
		_w10004_,
		_w11127_,
		_w11126_,
		_w11128_,
		_w11130_
	);
	LUT2 #(
		.INIT('h2)
	) name7083 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w11131_
	);
	LUT3 #(
		.INIT('h08)
	) name7084 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w11132_
	);
	LUT2 #(
		.INIT('h4)
	) name7085 (
		_w8375_,
		_w11132_,
		_w11133_
	);
	LUT3 #(
		.INIT('h45)
	) name7086 (
		_w11129_,
		_w11130_,
		_w11133_,
		_w11134_
	);
	LUT2 #(
		.INIT('h4)
	) name7087 (
		_w11125_,
		_w11134_,
		_w11135_
	);
	LUT3 #(
		.INIT('h0d)
	) name7088 (
		_w11123_,
		_w11124_,
		_w11135_,
		_w11136_
	);
	LUT3 #(
		.INIT('h04)
	) name7089 (
		_w9973_,
		_w10008_,
		_w11009_,
		_w11137_
	);
	LUT3 #(
		.INIT('h59)
	) name7090 (
		_w9973_,
		_w10008_,
		_w11009_,
		_w11138_
	);
	LUT3 #(
		.INIT('h69)
	) name7091 (
		_w11006_,
		_w11007_,
		_w11138_,
		_w11139_
	);
	LUT4 #(
		.INIT('h6640)
	) name7092 (
		_w11006_,
		_w11007_,
		_w11010_,
		_w11137_,
		_w11140_
	);
	LUT3 #(
		.INIT('h07)
	) name7093 (
		_w11136_,
		_w11139_,
		_w11140_,
		_w11141_
	);
	LUT4 #(
		.INIT('h7077)
	) name7094 (
		_w11081_,
		_w11109_,
		_w11110_,
		_w11141_,
		_w11142_
	);
	LUT4 #(
		.INIT('h6996)
	) name7095 (
		_w10993_,
		_w11014_,
		_w11042_,
		_w11071_,
		_w11143_
	);
	LUT4 #(
		.INIT('h6086)
	) name7096 (
		_w10993_,
		_w11014_,
		_w11042_,
		_w11071_,
		_w11144_
	);
	LUT3 #(
		.INIT('h0e)
	) name7097 (
		_w11142_,
		_w11143_,
		_w11144_,
		_w11145_
	);
	LUT2 #(
		.INIT('h6)
	) name7098 (
		_w11142_,
		_w11143_,
		_w11146_
	);
	LUT2 #(
		.INIT('h6)
	) name7099 (
		_w11136_,
		_w11139_,
		_w11147_
	);
	LUT4 #(
		.INIT('hfec8)
	) name7100 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10001_,
		_w10612_,
		_w10616_,
		_w11148_
	);
	LUT4 #(
		.INIT('h5655)
	) name7101 (
		_w10004_,
		_w11127_,
		_w11126_,
		_w11128_,
		_w11149_
	);
	LUT2 #(
		.INIT('h6)
	) name7102 (
		_w11133_,
		_w11149_,
		_w11150_
	);
	LUT2 #(
		.INIT('h2)
	) name7103 (
		_w11148_,
		_w11150_,
		_w11151_
	);
	LUT3 #(
		.INIT('he8)
	) name7104 (
		_w10601_,
		_w10605_,
		_w10609_,
		_w11152_
	);
	LUT3 #(
		.INIT('h69)
	) name7105 (
		_w11114_,
		_w11118_,
		_w11122_,
		_w11153_
	);
	LUT3 #(
		.INIT('h51)
	) name7106 (
		_w11151_,
		_w11152_,
		_w11153_,
		_w11154_
	);
	LUT2 #(
		.INIT('h2)
	) name7107 (
		_w11125_,
		_w11134_,
		_w11155_
	);
	LUT2 #(
		.INIT('h9)
	) name7108 (
		_w11125_,
		_w11134_,
		_w11156_
	);
	LUT3 #(
		.INIT('h69)
	) name7109 (
		_w11123_,
		_w11124_,
		_w11156_,
		_w11157_
	);
	LUT4 #(
		.INIT('h6640)
	) name7110 (
		_w11123_,
		_w11124_,
		_w11135_,
		_w11155_,
		_w11158_
	);
	LUT3 #(
		.INIT('h07)
	) name7111 (
		_w11154_,
		_w11157_,
		_w11158_,
		_w11159_
	);
	LUT2 #(
		.INIT('h9)
	) name7112 (
		_w11106_,
		_w11107_,
		_w11160_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name7113 (
		_w11084_,
		_w11086_,
		_w11085_,
		_w11087_,
		_w11161_
	);
	LUT2 #(
		.INIT('h1)
	) name7114 (
		_w10577_,
		_w11161_,
		_w11162_
	);
	LUT3 #(
		.INIT('he8)
	) name7115 (
		_w10583_,
		_w10587_,
		_w10591_,
		_w11163_
	);
	LUT3 #(
		.INIT('h69)
	) name7116 (
		_w11095_,
		_w11099_,
		_w11103_,
		_w11164_
	);
	LUT3 #(
		.INIT('h51)
	) name7117 (
		_w11162_,
		_w11163_,
		_w11164_,
		_w11165_
	);
	LUT3 #(
		.INIT('h69)
	) name7118 (
		_w11066_,
		_w11088_,
		_w11089_,
		_w11166_
	);
	LUT3 #(
		.INIT('h69)
	) name7119 (
		_w11104_,
		_w11105_,
		_w11166_,
		_w11167_
	);
	LUT4 #(
		.INIT('h0980)
	) name7120 (
		_w11088_,
		_w11090_,
		_w11104_,
		_w11105_,
		_w11168_
	);
	LUT3 #(
		.INIT('h07)
	) name7121 (
		_w11165_,
		_w11167_,
		_w11168_,
		_w11169_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name7122 (
		_w11147_,
		_w11159_,
		_w11160_,
		_w11169_,
		_w11170_
	);
	LUT4 #(
		.INIT('h9669)
	) name7123 (
		_w11081_,
		_w11109_,
		_w11110_,
		_w11141_,
		_w11171_
	);
	LUT4 #(
		.INIT('h0190)
	) name7124 (
		_w11081_,
		_w11109_,
		_w11110_,
		_w11141_,
		_w11172_
	);
	LUT3 #(
		.INIT('h07)
	) name7125 (
		_w11170_,
		_w11171_,
		_w11172_,
		_w11173_
	);
	LUT2 #(
		.INIT('h8)
	) name7126 (
		_w11146_,
		_w11173_,
		_w11174_
	);
	LUT4 #(
		.INIT('h0eee)
	) name7127 (
		_w11080_,
		_w11145_,
		_w11146_,
		_w11173_,
		_w11175_
	);
	LUT4 #(
		.INIT('hee0e)
	) name7128 (
		_w11073_,
		_w11075_,
		_w11076_,
		_w11078_,
		_w11176_
	);
	LUT4 #(
		.INIT('h9669)
	) name7129 (
		_w10870_,
		_w10899_,
		_w10916_,
		_w10917_,
		_w11177_
	);
	LUT2 #(
		.INIT('h6)
	) name7130 (
		_w11176_,
		_w11177_,
		_w11178_
	);
	LUT4 #(
		.INIT('h0980)
	) name7131 (
		_w11073_,
		_w11075_,
		_w11076_,
		_w11078_,
		_w11179_
	);
	LUT3 #(
		.INIT('h07)
	) name7132 (
		_w11072_,
		_w11079_,
		_w11179_,
		_w11180_
	);
	LUT2 #(
		.INIT('h4)
	) name7133 (
		_w11178_,
		_w11180_,
		_w11181_
	);
	LUT4 #(
		.INIT('h0190)
	) name7134 (
		_w10870_,
		_w10899_,
		_w10916_,
		_w10917_,
		_w11182_
	);
	LUT3 #(
		.INIT('h07)
	) name7135 (
		_w11176_,
		_w11177_,
		_w11182_,
		_w11183_
	);
	LUT2 #(
		.INIT('h9)
	) name7136 (
		_w10918_,
		_w10919_,
		_w11184_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7137 (
		_w11178_,
		_w11180_,
		_w11183_,
		_w11184_,
		_w11185_
	);
	LUT2 #(
		.INIT('h8)
	) name7138 (
		_w11175_,
		_w11185_,
		_w11186_
	);
	LUT4 #(
		.INIT('h2000)
	) name7139 (
		_w10923_,
		_w10973_,
		_w11175_,
		_w11185_,
		_w11187_
	);
	LUT2 #(
		.INIT('h6)
	) name7140 (
		_w11170_,
		_w11171_,
		_w11188_
	);
	LUT2 #(
		.INIT('h6)
	) name7141 (
		_w11154_,
		_w11157_,
		_w11189_
	);
	LUT3 #(
		.INIT('h0d)
	) name7142 (
		_w10597_,
		_w10610_,
		_w10618_,
		_w11190_
	);
	LUT2 #(
		.INIT('h4)
	) name7143 (
		_w11148_,
		_w11150_,
		_w11191_
	);
	LUT2 #(
		.INIT('h9)
	) name7144 (
		_w11148_,
		_w11150_,
		_w11192_
	);
	LUT3 #(
		.INIT('h96)
	) name7145 (
		_w11152_,
		_w11153_,
		_w11192_,
		_w11193_
	);
	LUT4 #(
		.INIT('h0049)
	) name7146 (
		_w11151_,
		_w11152_,
		_w11153_,
		_w11191_,
		_w11194_
	);
	LUT3 #(
		.INIT('h0e)
	) name7147 (
		_w11190_,
		_w11193_,
		_w11194_,
		_w11195_
	);
	LUT2 #(
		.INIT('h6)
	) name7148 (
		_w11165_,
		_w11167_,
		_w11196_
	);
	LUT3 #(
		.INIT('ha2)
	) name7149 (
		_w10578_,
		_w10579_,
		_w10592_,
		_w11197_
	);
	LUT2 #(
		.INIT('h8)
	) name7150 (
		_w10577_,
		_w11161_,
		_w11198_
	);
	LUT2 #(
		.INIT('h6)
	) name7151 (
		_w10577_,
		_w11161_,
		_w11199_
	);
	LUT3 #(
		.INIT('h96)
	) name7152 (
		_w11163_,
		_w11164_,
		_w11199_,
		_w11200_
	);
	LUT4 #(
		.INIT('h0049)
	) name7153 (
		_w11162_,
		_w11163_,
		_w11164_,
		_w11198_,
		_w11201_
	);
	LUT3 #(
		.INIT('h0e)
	) name7154 (
		_w11197_,
		_w11200_,
		_w11201_,
		_w11202_
	);
	LUT4 #(
		.INIT('heee0)
	) name7155 (
		_w11189_,
		_w11195_,
		_w11196_,
		_w11202_,
		_w11203_
	);
	LUT4 #(
		.INIT('h6996)
	) name7156 (
		_w11147_,
		_w11159_,
		_w11160_,
		_w11169_,
		_w11204_
	);
	LUT4 #(
		.INIT('h0260)
	) name7157 (
		_w11147_,
		_w11159_,
		_w11160_,
		_w11169_,
		_w11205_
	);
	LUT3 #(
		.INIT('h07)
	) name7158 (
		_w11203_,
		_w11204_,
		_w11205_,
		_w11206_
	);
	LUT2 #(
		.INIT('h6)
	) name7159 (
		_w11203_,
		_w11204_,
		_w11207_
	);
	LUT2 #(
		.INIT('h6)
	) name7160 (
		_w11190_,
		_w11193_,
		_w11208_
	);
	LUT4 #(
		.INIT('h0029)
	) name7161 (
		_w10597_,
		_w10610_,
		_w10618_,
		_w10619_,
		_w11209_
	);
	LUT3 #(
		.INIT('h0b)
	) name7162 (
		_w10596_,
		_w10621_,
		_w11209_,
		_w11210_
	);
	LUT3 #(
		.INIT('h10)
	) name7163 (
		_w10578_,
		_w10579_,
		_w10592_,
		_w11211_
	);
	LUT3 #(
		.INIT('h06)
	) name7164 (
		_w11197_,
		_w11200_,
		_w11211_,
		_w11212_
	);
	LUT3 #(
		.INIT('h0d)
	) name7165 (
		_w11208_,
		_w11210_,
		_w11212_,
		_w11213_
	);
	LUT4 #(
		.INIT('h9669)
	) name7166 (
		_w11189_,
		_w11195_,
		_w11196_,
		_w11202_,
		_w11214_
	);
	LUT4 #(
		.INIT('h0661)
	) name7167 (
		_w11189_,
		_w11195_,
		_w11196_,
		_w11202_,
		_w11215_
	);
	LUT3 #(
		.INIT('h0e)
	) name7168 (
		_w11213_,
		_w11214_,
		_w11215_,
		_w11216_
	);
	LUT2 #(
		.INIT('h1)
	) name7169 (
		_w11207_,
		_w11216_,
		_w11217_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name7170 (
		_w11188_,
		_w11206_,
		_w11207_,
		_w11216_,
		_w11218_
	);
	LUT2 #(
		.INIT('h6)
	) name7171 (
		_w11213_,
		_w11214_,
		_w11219_
	);
	LUT3 #(
		.INIT('h51)
	) name7172 (
		_w10594_,
		_w10622_,
		_w10624_,
		_w11220_
	);
	LUT2 #(
		.INIT('h4)
	) name7173 (
		_w11200_,
		_w11211_,
		_w11221_
	);
	LUT3 #(
		.INIT('hc9)
	) name7174 (
		_w11197_,
		_w11200_,
		_w11211_,
		_w11222_
	);
	LUT3 #(
		.INIT('h69)
	) name7175 (
		_w11208_,
		_w11210_,
		_w11222_,
		_w11223_
	);
	LUT4 #(
		.INIT('h0029)
	) name7176 (
		_w11208_,
		_w11210_,
		_w11212_,
		_w11221_,
		_w11224_
	);
	LUT3 #(
		.INIT('h0b)
	) name7177 (
		_w11220_,
		_w11223_,
		_w11224_,
		_w11225_
	);
	LUT2 #(
		.INIT('h9)
	) name7178 (
		_w11220_,
		_w11223_,
		_w11226_
	);
	LUT4 #(
		.INIT('h6016)
	) name7179 (
		_w10558_,
		_w10593_,
		_w10622_,
		_w10624_,
		_w11227_
	);
	LUT3 #(
		.INIT('h0b)
	) name7180 (
		_w10575_,
		_w10625_,
		_w11227_,
		_w11228_
	);
	LUT2 #(
		.INIT('h2)
	) name7181 (
		_w11226_,
		_w11228_,
		_w11229_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name7182 (
		_w11219_,
		_w11225_,
		_w11226_,
		_w11228_,
		_w11230_
	);
	LUT2 #(
		.INIT('h8)
	) name7183 (
		_w11218_,
		_w11230_,
		_w11231_
	);
	LUT2 #(
		.INIT('h8)
	) name7184 (
		_w11187_,
		_w11231_,
		_w11232_
	);
	LUT2 #(
		.INIT('h1)
	) name7185 (
		_w11146_,
		_w11173_,
		_w11233_
	);
	LUT4 #(
		.INIT('h888e)
	) name7186 (
		_w11080_,
		_w11145_,
		_w11146_,
		_w11173_,
		_w11234_
	);
	LUT2 #(
		.INIT('h2)
	) name7187 (
		_w11178_,
		_w11180_,
		_w11235_
	);
	LUT4 #(
		.INIT('hfdd0)
	) name7188 (
		_w11178_,
		_w11180_,
		_w11183_,
		_w11184_,
		_w11236_
	);
	LUT3 #(
		.INIT('h70)
	) name7189 (
		_w11185_,
		_w11234_,
		_w11236_,
		_w11237_
	);
	LUT2 #(
		.INIT('h2)
	) name7190 (
		_w10974_,
		_w11237_,
		_w11238_
	);
	LUT2 #(
		.INIT('h4)
	) name7191 (
		_w11226_,
		_w11228_,
		_w11239_
	);
	LUT4 #(
		.INIT('h4d44)
	) name7192 (
		_w11219_,
		_w11225_,
		_w11226_,
		_w11228_,
		_w11240_
	);
	LUT2 #(
		.INIT('h8)
	) name7193 (
		_w11207_,
		_w11216_,
		_w11241_
	);
	LUT4 #(
		.INIT('h4ddd)
	) name7194 (
		_w11188_,
		_w11206_,
		_w11207_,
		_w11216_,
		_w11242_
	);
	LUT3 #(
		.INIT('h70)
	) name7195 (
		_w11218_,
		_w11240_,
		_w11242_,
		_w11243_
	);
	LUT2 #(
		.INIT('h8)
	) name7196 (
		_w10869_,
		_w10921_,
		_w11244_
	);
	LUT4 #(
		.INIT('h8eee)
	) name7197 (
		_w10814_,
		_w10868_,
		_w10869_,
		_w10921_,
		_w11245_
	);
	LUT2 #(
		.INIT('h4)
	) name7198 (
		_w10967_,
		_w10969_,
		_w11246_
	);
	LUT4 #(
		.INIT('h5510)
	) name7199 (
		_w10964_,
		_w10967_,
		_w10969_,
		_w10972_,
		_w11247_
	);
	LUT3 #(
		.INIT('h0e)
	) name7200 (
		_w10973_,
		_w11245_,
		_w11247_,
		_w11248_
	);
	LUT3 #(
		.INIT('hd0)
	) name7201 (
		_w11187_,
		_w11243_,
		_w11248_,
		_w11249_
	);
	LUT4 #(
		.INIT('h0b00)
	) name7202 (
		_w10646_,
		_w11232_,
		_w11238_,
		_w11249_,
		_w11250_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name7203 (
		_w10952_,
		_w10953_,
		_w10955_,
		_w10956_,
		_w11251_
	);
	LUT4 #(
		.INIT('h9669)
	) name7204 (
		_w10137_,
		_w10146_,
		_w10153_,
		_w10154_,
		_w11252_
	);
	LUT2 #(
		.INIT('h6)
	) name7205 (
		_w11251_,
		_w11252_,
		_w11253_
	);
	LUT4 #(
		.INIT('h9209)
	) name7206 (
		_w10952_,
		_w10953_,
		_w10955_,
		_w10956_,
		_w11254_
	);
	LUT3 #(
		.INIT('h0b)
	) name7207 (
		_w10951_,
		_w10957_,
		_w11254_,
		_w11255_
	);
	LUT2 #(
		.INIT('h2)
	) name7208 (
		_w11253_,
		_w11255_,
		_w11256_
	);
	LUT3 #(
		.INIT('h51)
	) name7209 (
		_w9974_,
		_w11253_,
		_w11255_,
		_w11257_
	);
	LUT2 #(
		.INIT('h9)
	) name7210 (
		_w10155_,
		_w10157_,
		_w11258_
	);
	LUT4 #(
		.INIT('h9049)
	) name7211 (
		_w10137_,
		_w10146_,
		_w10153_,
		_w10154_,
		_w11259_
	);
	LUT3 #(
		.INIT('h0e)
	) name7212 (
		_w11251_,
		_w11252_,
		_w11259_,
		_w11260_
	);
	LUT2 #(
		.INIT('h2)
	) name7213 (
		_w11258_,
		_w11260_,
		_w11261_
	);
	LUT2 #(
		.INIT('h9)
	) name7214 (
		_w11258_,
		_w11260_,
		_w11262_
	);
	LUT3 #(
		.INIT('h69)
	) name7215 (
		_w9974_,
		_w11258_,
		_w11260_,
		_w11263_
	);
	LUT3 #(
		.INIT('h4b)
	) name7216 (
		_w9974_,
		_w11256_,
		_w11262_,
		_w11264_
	);
	LUT3 #(
		.INIT('h51)
	) name7217 (
		_w9974_,
		_w10958_,
		_w10960_,
		_w11265_
	);
	LUT2 #(
		.INIT('h9)
	) name7218 (
		_w11253_,
		_w11255_,
		_w11266_
	);
	LUT3 #(
		.INIT('h69)
	) name7219 (
		_w9974_,
		_w11253_,
		_w11255_,
		_w11267_
	);
	LUT3 #(
		.INIT('h4b)
	) name7220 (
		_w9974_,
		_w10961_,
		_w11266_,
		_w11268_
	);
	LUT3 #(
		.INIT('h49)
	) name7221 (
		_w9974_,
		_w11253_,
		_w11255_,
		_w11269_
	);
	LUT3 #(
		.INIT('h0e)
	) name7222 (
		_w11265_,
		_w11267_,
		_w11269_,
		_w11270_
	);
	LUT3 #(
		.INIT('h49)
	) name7223 (
		_w9974_,
		_w10958_,
		_w10960_,
		_w11271_
	);
	LUT3 #(
		.INIT('h0e)
	) name7224 (
		_w10950_,
		_w10963_,
		_w11271_,
		_w11272_
	);
	LUT4 #(
		.INIT('h0aee)
	) name7225 (
		_w11264_,
		_w11268_,
		_w11270_,
		_w11272_,
		_w11273_
	);
	LUT3 #(
		.INIT('h4b)
	) name7226 (
		_w9974_,
		_w10160_,
		_w10162_,
		_w11274_
	);
	LUT3 #(
		.INIT('h49)
	) name7227 (
		_w9974_,
		_w11258_,
		_w11260_,
		_w11275_
	);
	LUT3 #(
		.INIT('h0e)
	) name7228 (
		_w11257_,
		_w11263_,
		_w11275_,
		_w11276_
	);
	LUT3 #(
		.INIT('h51)
	) name7229 (
		_w9974_,
		_w11258_,
		_w11260_,
		_w11277_
	);
	LUT2 #(
		.INIT('h9)
	) name7230 (
		_w10135_,
		_w10159_,
		_w11278_
	);
	LUT3 #(
		.INIT('h69)
	) name7231 (
		_w9974_,
		_w10135_,
		_w10159_,
		_w11279_
	);
	LUT3 #(
		.INIT('h4b)
	) name7232 (
		_w9974_,
		_w11261_,
		_w11278_,
		_w11280_
	);
	LUT2 #(
		.INIT('h4)
	) name7233 (
		_w11276_,
		_w11280_,
		_w11281_
	);
	LUT3 #(
		.INIT('h49)
	) name7234 (
		_w9974_,
		_w10135_,
		_w10159_,
		_w11282_
	);
	LUT3 #(
		.INIT('h0e)
	) name7235 (
		_w11277_,
		_w11279_,
		_w11282_,
		_w11283_
	);
	LUT4 #(
		.INIT('h32ba)
	) name7236 (
		_w11274_,
		_w11276_,
		_w11280_,
		_w11283_,
		_w11284_
	);
	LUT2 #(
		.INIT('h1)
	) name7237 (
		_w11273_,
		_w11284_,
		_w11285_
	);
	LUT4 #(
		.INIT('haeaf)
	) name7238 (
		_w11264_,
		_w11268_,
		_w11270_,
		_w11272_,
		_w11286_
	);
	LUT2 #(
		.INIT('h2)
	) name7239 (
		_w11276_,
		_w11280_,
		_w11287_
	);
	LUT4 #(
		.INIT('ha2fb)
	) name7240 (
		_w11274_,
		_w11276_,
		_w11280_,
		_w11283_,
		_w11288_
	);
	LUT3 #(
		.INIT('he0)
	) name7241 (
		_w11284_,
		_w11286_,
		_w11288_,
		_w11289_
	);
	LUT4 #(
		.INIT('h4500)
	) name7242 (
		_w10165_,
		_w11250_,
		_w11285_,
		_w11289_,
		_w11290_
	);
	LUT3 #(
		.INIT('h01)
	) name7243 (
		_w10131_,
		_w10133_,
		_w10166_,
		_w11291_
	);
	LUT3 #(
		.INIT('h07)
	) name7244 (
		_w10134_,
		_w10165_,
		_w11291_,
		_w11292_
	);
	LUT4 #(
		.INIT('hfe00)
	) name7245 (
		_w10132_,
		_w10168_,
		_w11290_,
		_w11292_,
		_w11293_
	);
	LUT4 #(
		.INIT('h6665)
	) name7246 (
		_w10073_,
		_w10103_,
		_w10104_,
		_w11293_,
		_w11294_
	);
	LUT2 #(
		.INIT('h9)
	) name7247 (
		_w10101_,
		_w10102_,
		_w11295_
	);
	LUT2 #(
		.INIT('h6)
	) name7248 (
		_w11293_,
		_w11295_,
		_w11296_
	);
	LUT3 #(
		.INIT('h14)
	) name7249 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11293_,
		_w11295_,
		_w11297_
	);
	LUT3 #(
		.INIT('h0d)
	) name7250 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11294_,
		_w11297_,
		_w11298_
	);
	LUT4 #(
		.INIT('h4c08)
	) name7251 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w11294_,
		_w11296_,
		_w11299_
	);
	LUT4 #(
		.INIT('h1011)
	) name7252 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w11300_
	);
	LUT2 #(
		.INIT('h8)
	) name7253 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		_w11300_,
		_w11301_
	);
	LUT3 #(
		.INIT('h13)
	) name7254 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001 ,
		_w11300_,
		_w11302_
	);
	LUT2 #(
		.INIT('h4)
	) name7255 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR2_E_reg/P0001 ,
		_w11303_
	);
	LUT2 #(
		.INIT('h4)
	) name7256 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w11304_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name7257 (
		\core_c_dec_satMR_E_reg/P0001 ,
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4145_,
		_w4154_,
		_w11305_
	);
	LUT2 #(
		.INIT('h4)
	) name7258 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w11305_,
		_w11306_
	);
	LUT3 #(
		.INIT('hab)
	) name7259 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w11305_,
		_w11307_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name7260 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_c_dec_updMR_E_reg/P0001 ,
		_w11305_,
		_w11308_
	);
	LUT3 #(
		.INIT('h45)
	) name7261 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11303_,
		_w11308_,
		_w11309_
	);
	LUT4 #(
		.INIT('h5040)
	) name7262 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w9452_,
		_w11305_,
		_w11310_
	);
	LUT2 #(
		.INIT('h1)
	) name7263 (
		_w11301_,
		_w11310_,
		_w11311_
	);
	LUT2 #(
		.INIT('h2)
	) name7264 (
		_w11309_,
		_w11311_,
		_w11312_
	);
	LUT4 #(
		.INIT('h4544)
	) name7265 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6378_,
		_w6498_,
		_w6500_,
		_w11313_
	);
	LUT2 #(
		.INIT('h2)
	) name7266 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8863_,
		_w11314_
	);
	LUT2 #(
		.INIT('h1)
	) name7267 (
		_w11313_,
		_w11314_,
		_w11315_
	);
	LUT4 #(
		.INIT('hccc8)
	) name7268 (
		_w11310_,
		_w11312_,
		_w11313_,
		_w11314_,
		_w11316_
	);
	LUT2 #(
		.INIT('h2)
	) name7269 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8821_,
		_w11317_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7270 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8798_,
		_w8801_,
		_w11317_,
		_w11318_
	);
	LUT2 #(
		.INIT('h2)
	) name7271 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w11305_,
		_w11319_
	);
	LUT3 #(
		.INIT('h80)
	) name7272 (
		_w11300_,
		_w11318_,
		_w11319_,
		_w11320_
	);
	LUT4 #(
		.INIT('h2322)
	) name7273 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001 ,
		_w11303_,
		_w11308_,
		_w11321_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7274 (
		_w11302_,
		_w11316_,
		_w11320_,
		_w11321_,
		_w11322_
	);
	LUT2 #(
		.INIT('h8)
	) name7275 (
		_w11300_,
		_w11305_,
		_w11323_
	);
	LUT3 #(
		.INIT('h80)
	) name7276 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 ,
		_w11300_,
		_w11305_,
		_w11324_
	);
	LUT2 #(
		.INIT('h1)
	) name7277 (
		_w9946_,
		_w11324_,
		_w11325_
	);
	LUT2 #(
		.INIT('h4)
	) name7278 (
		_w11322_,
		_w11325_,
		_w11326_
	);
	LUT2 #(
		.INIT('h1)
	) name7279 (
		_w11299_,
		_w11326_,
		_w11327_
	);
	LUT2 #(
		.INIT('h1)
	) name7280 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		\core_c_dec_updSR_E_reg/P0001 ,
		_w11328_
	);
	LUT4 #(
		.INIT('h0004)
	) name7281 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9452_,
		_w9453_,
		_w11328_,
		_w11329_
	);
	LUT2 #(
		.INIT('h2)
	) name7282 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8740_,
		_w11330_
	);
	LUT3 #(
		.INIT('h0e)
	) name7283 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w11330_,
		_w11331_
	);
	LUT4 #(
		.INIT('h028a)
	) name7284 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w11332_
	);
	LUT3 #(
		.INIT('h70)
	) name7285 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_SHTop_E_reg/P0001 ,
		_w11333_
	);
	LUT2 #(
		.INIT('h4)
	) name7286 (
		_w8367_,
		_w9470_,
		_w11334_
	);
	LUT4 #(
		.INIT('h0040)
	) name7287 (
		_w9462_,
		_w9465_,
		_w9468_,
		_w11334_,
		_w11335_
	);
	LUT2 #(
		.INIT('h2)
	) name7288 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w11336_
	);
	LUT2 #(
		.INIT('h4)
	) name7289 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w11337_
	);
	LUT3 #(
		.INIT('h40)
	) name7290 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w11338_
	);
	LUT2 #(
		.INIT('h8)
	) name7291 (
		_w11337_,
		_w11338_,
		_w11339_
	);
	LUT3 #(
		.INIT('h0b)
	) name7292 (
		_w11335_,
		_w11336_,
		_w11339_,
		_w11340_
	);
	LUT4 #(
		.INIT('haa20)
	) name7293 (
		_w11333_,
		_w11335_,
		_w11336_,
		_w11339_,
		_w11341_
	);
	LUT4 #(
		.INIT('h8000)
	) name7294 (
		_w5889_,
		_w6133_,
		_w6469_,
		_w6884_,
		_w11342_
	);
	LUT4 #(
		.INIT('h8000)
	) name7295 (
		_w7331_,
		_w7692_,
		_w8008_,
		_w11342_,
		_w11343_
	);
	LUT4 #(
		.INIT('h78f0)
	) name7296 (
		_w7331_,
		_w7692_,
		_w8008_,
		_w11342_,
		_w11344_
	);
	LUT4 #(
		.INIT('h5410)
	) name7297 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001 ,
		_w11345_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7298 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w11346_
	);
	LUT2 #(
		.INIT('h4)
	) name7299 (
		_w11345_,
		_w11346_,
		_w11347_
	);
	LUT3 #(
		.INIT('h0d)
	) name7300 (
		_w11337_,
		_w11344_,
		_w11347_,
		_w11348_
	);
	LUT4 #(
		.INIT('h9030)
	) name7301 (
		_w7331_,
		_w7692_,
		_w11337_,
		_w11342_,
		_w11349_
	);
	LUT4 #(
		.INIT('h5410)
	) name7302 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001 ,
		_w11350_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7303 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w11351_
	);
	LUT2 #(
		.INIT('h4)
	) name7304 (
		_w11350_,
		_w11351_,
		_w11352_
	);
	LUT2 #(
		.INIT('h1)
	) name7305 (
		_w11349_,
		_w11352_,
		_w11353_
	);
	LUT4 #(
		.INIT('h5410)
	) name7306 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001 ,
		_w11354_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7307 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_IRE_reg[7]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w11355_
	);
	LUT2 #(
		.INIT('h4)
	) name7308 (
		_w11354_,
		_w11355_,
		_w11356_
	);
	LUT4 #(
		.INIT('h007b)
	) name7309 (
		_w5744_,
		_w11337_,
		_w11343_,
		_w11356_,
		_w11357_
	);
	LUT4 #(
		.INIT('h8000)
	) name7310 (
		_w11333_,
		_w11348_,
		_w11357_,
		_w11353_,
		_w11358_
	);
	LUT3 #(
		.INIT('h90)
	) name7311 (
		_w5889_,
		_w6884_,
		_w11337_,
		_w11359_
	);
	LUT4 #(
		.INIT('h5410)
	) name7312 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001 ,
		_w11360_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7313 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_IRE_reg[1]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w11361_
	);
	LUT2 #(
		.INIT('h4)
	) name7314 (
		_w11360_,
		_w11361_,
		_w11362_
	);
	LUT2 #(
		.INIT('h1)
	) name7315 (
		_w11359_,
		_w11362_,
		_w11363_
	);
	LUT3 #(
		.INIT('h02)
	) name7316 (
		_w11333_,
		_w11359_,
		_w11362_,
		_w11364_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name7317 (
		_w5889_,
		_w6133_,
		_w6469_,
		_w6884_,
		_w11365_
	);
	LUT4 #(
		.INIT('h5410)
	) name7318 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001 ,
		_w11366_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7319 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w11367_
	);
	LUT2 #(
		.INIT('h4)
	) name7320 (
		_w11366_,
		_w11367_,
		_w11368_
	);
	LUT3 #(
		.INIT('h0d)
	) name7321 (
		_w11337_,
		_w11365_,
		_w11368_,
		_w11369_
	);
	LUT4 #(
		.INIT('h00a2)
	) name7322 (
		_w11333_,
		_w11337_,
		_w11365_,
		_w11368_,
		_w11370_
	);
	LUT2 #(
		.INIT('h1)
	) name7323 (
		_w11364_,
		_w11370_,
		_w11371_
	);
	LUT4 #(
		.INIT('h5410)
	) name7324 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001 ,
		_w11372_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7325 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w11373_
	);
	LUT2 #(
		.INIT('h4)
	) name7326 (
		_w11372_,
		_w11373_,
		_w11374_
	);
	LUT4 #(
		.INIT('h007b)
	) name7327 (
		_w7331_,
		_w11337_,
		_w11342_,
		_w11374_,
		_w11375_
	);
	LUT4 #(
		.INIT('h9300)
	) name7328 (
		_w5889_,
		_w6469_,
		_w6884_,
		_w11337_,
		_w11376_
	);
	LUT4 #(
		.INIT('h5410)
	) name7329 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001 ,
		_w11377_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7330 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w11378_
	);
	LUT2 #(
		.INIT('h4)
	) name7331 (
		_w11377_,
		_w11378_,
		_w11379_
	);
	LUT2 #(
		.INIT('h1)
	) name7332 (
		_w11376_,
		_w11379_,
		_w11380_
	);
	LUT3 #(
		.INIT('h02)
	) name7333 (
		_w11333_,
		_w11376_,
		_w11379_,
		_w11381_
	);
	LUT4 #(
		.INIT('h1000)
	) name7334 (
		_w11364_,
		_w11370_,
		_w11375_,
		_w11381_,
		_w11382_
	);
	LUT3 #(
		.INIT('h40)
	) name7335 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11382_,
		_w11383_
	);
	LUT3 #(
		.INIT('hb0)
	) name7336 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w11384_
	);
	LUT3 #(
		.INIT('ha3)
	) name7337 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w5889_,
		_w11384_,
		_w11385_
	);
	LUT4 #(
		.INIT('ha030)
	) name7338 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w5889_,
		_w11333_,
		_w11384_,
		_w11386_
	);
	LUT4 #(
		.INIT('h2a00)
	) name7339 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_SHTop_E_reg/P0001 ,
		_w11387_
	);
	LUT3 #(
		.INIT('he0)
	) name7340 (
		_w11349_,
		_w11352_,
		_w11387_,
		_w11388_
	);
	LUT3 #(
		.INIT('h10)
	) name7341 (
		_w11348_,
		_w11357_,
		_w11388_,
		_w11389_
	);
	LUT3 #(
		.INIT('h07)
	) name7342 (
		_w11333_,
		_w11375_,
		_w11381_,
		_w11390_
	);
	LUT2 #(
		.INIT('h2)
	) name7343 (
		_w11364_,
		_w11369_,
		_w11391_
	);
	LUT2 #(
		.INIT('h8)
	) name7344 (
		_w11390_,
		_w11391_,
		_w11392_
	);
	LUT2 #(
		.INIT('h8)
	) name7345 (
		_w11389_,
		_w11392_,
		_w11393_
	);
	LUT3 #(
		.INIT('h20)
	) name7346 (
		_w11389_,
		_w11386_,
		_w11392_,
		_w11394_
	);
	LUT4 #(
		.INIT('h2000)
	) name7347 (
		_w11364_,
		_w11369_,
		_w11375_,
		_w11381_,
		_w11395_
	);
	LUT3 #(
		.INIT('h80)
	) name7348 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11395_,
		_w11396_
	);
	LUT4 #(
		.INIT('h8000)
	) name7349 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11385_,
		_w11358_,
		_w11395_,
		_w11397_
	);
	LUT4 #(
		.INIT('h0103)
	) name7350 (
		_w11333_,
		_w11383_,
		_w11394_,
		_w11397_,
		_w11398_
	);
	LUT2 #(
		.INIT('h2)
	) name7351 (
		_w11341_,
		_w11398_,
		_w11399_
	);
	LUT3 #(
		.INIT('h08)
	) name7352 (
		_w11333_,
		_w11375_,
		_w11380_,
		_w11400_
	);
	LUT2 #(
		.INIT('h8)
	) name7353 (
		_w11371_,
		_w11400_,
		_w11401_
	);
	LUT4 #(
		.INIT('haa20)
	) name7354 (
		_w11386_,
		_w11335_,
		_w11336_,
		_w11339_,
		_w11402_
	);
	LUT4 #(
		.INIT('h8000)
	) name7355 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11401_,
		_w11358_,
		_w11402_,
		_w11403_
	);
	LUT2 #(
		.INIT('h8)
	) name7356 (
		_w11363_,
		_w11370_,
		_w11404_
	);
	LUT4 #(
		.INIT('h0800)
	) name7357 (
		_w11363_,
		_w11370_,
		_w11375_,
		_w11381_,
		_w11405_
	);
	LUT2 #(
		.INIT('h4)
	) name7358 (
		_w11385_,
		_w11341_,
		_w11406_
	);
	LUT4 #(
		.INIT('h4000)
	) name7359 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11406_,
		_w11405_,
		_w11407_
	);
	LUT2 #(
		.INIT('h1)
	) name7360 (
		_w11403_,
		_w11407_,
		_w11408_
	);
	LUT4 #(
		.INIT('h4000)
	) name7361 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11395_,
		_w11409_
	);
	LUT4 #(
		.INIT('h2000)
	) name7362 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11395_,
		_w11410_
	);
	LUT4 #(
		.INIT('h9fff)
	) name7363 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11395_,
		_w11411_
	);
	LUT4 #(
		.INIT('h0301)
	) name7364 (
		_w11341_,
		_w11403_,
		_w11407_,
		_w11411_,
		_w11412_
	);
	LUT2 #(
		.INIT('h4)
	) name7365 (
		_w11363_,
		_w11370_,
		_w11413_
	);
	LUT4 #(
		.INIT('h0400)
	) name7366 (
		_w11363_,
		_w11370_,
		_w11375_,
		_w11381_,
		_w11414_
	);
	LUT4 #(
		.INIT('h1000)
	) name7367 (
		_w11348_,
		_w11357_,
		_w11388_,
		_w11414_,
		_w11415_
	);
	LUT2 #(
		.INIT('h8)
	) name7368 (
		_w11406_,
		_w11415_,
		_w11416_
	);
	LUT2 #(
		.INIT('h2)
	) name7369 (
		_w11412_,
		_w11416_,
		_w11417_
	);
	LUT4 #(
		.INIT('h4000)
	) name7370 (
		_w11363_,
		_w11370_,
		_w11375_,
		_w11381_,
		_w11418_
	);
	LUT3 #(
		.INIT('h80)
	) name7371 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11418_,
		_w11419_
	);
	LUT4 #(
		.INIT('h8000)
	) name7372 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11418_,
		_w11420_
	);
	LUT4 #(
		.INIT('h4000)
	) name7373 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11414_,
		_w11421_
	);
	LUT3 #(
		.INIT('ha8)
	) name7374 (
		_w11341_,
		_w11420_,
		_w11421_,
		_w11422_
	);
	LUT4 #(
		.INIT('h0200)
	) name7375 (
		_w11364_,
		_w11369_,
		_w11375_,
		_w11381_,
		_w11423_
	);
	LUT4 #(
		.INIT('h1000)
	) name7376 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11423_,
		_w11424_
	);
	LUT4 #(
		.INIT('h2000)
	) name7377 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11382_,
		_w11425_
	);
	LUT3 #(
		.INIT('ha8)
	) name7378 (
		_w11341_,
		_w11424_,
		_w11425_,
		_w11426_
	);
	LUT4 #(
		.INIT('h8000)
	) name7379 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11406_,
		_w11418_,
		_w11427_
	);
	LUT4 #(
		.INIT('h0100)
	) name7380 (
		_w11364_,
		_w11370_,
		_w11375_,
		_w11381_,
		_w11428_
	);
	LUT4 #(
		.INIT('h1000)
	) name7381 (
		_w11348_,
		_w11357_,
		_w11388_,
		_w11428_,
		_w11429_
	);
	LUT2 #(
		.INIT('h8)
	) name7382 (
		_w11402_,
		_w11429_,
		_w11430_
	);
	LUT2 #(
		.INIT('h1)
	) name7383 (
		_w11427_,
		_w11430_,
		_w11431_
	);
	LUT3 #(
		.INIT('h10)
	) name7384 (
		_w11426_,
		_w11422_,
		_w11431_,
		_w11432_
	);
	LUT3 #(
		.INIT('h40)
	) name7385 (
		_w11399_,
		_w11417_,
		_w11432_,
		_w11433_
	);
	LUT2 #(
		.INIT('h8)
	) name7386 (
		_w11400_,
		_w11413_,
		_w11434_
	);
	LUT4 #(
		.INIT('h1000)
	) name7387 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11434_,
		_w11435_
	);
	LUT3 #(
		.INIT('h80)
	) name7388 (
		_w11389_,
		_w11392_,
		_w11402_,
		_w11436_
	);
	LUT3 #(
		.INIT('h07)
	) name7389 (
		_w11341_,
		_w11435_,
		_w11436_,
		_w11437_
	);
	LUT4 #(
		.INIT('h8000)
	) name7390 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11401_,
		_w11358_,
		_w11406_,
		_w11438_
	);
	LUT4 #(
		.INIT('h8000)
	) name7391 (
		_w11363_,
		_w11370_,
		_w11375_,
		_w11381_,
		_w11439_
	);
	LUT4 #(
		.INIT('h8000)
	) name7392 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11402_,
		_w11439_,
		_w11440_
	);
	LUT2 #(
		.INIT('h1)
	) name7393 (
		_w11438_,
		_w11440_,
		_w11441_
	);
	LUT2 #(
		.INIT('h8)
	) name7394 (
		_w11437_,
		_w11441_,
		_w11442_
	);
	LUT3 #(
		.INIT('h54)
	) name7395 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11349_,
		_w11352_,
		_w11443_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7396 (
		_w11333_,
		_w11348_,
		_w11357_,
		_w11443_,
		_w11444_
	);
	LUT2 #(
		.INIT('h8)
	) name7397 (
		_w11390_,
		_w11413_,
		_w11445_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7398 (
		_w11444_,
		_w11389_,
		_w11434_,
		_w11445_,
		_w11446_
	);
	LUT2 #(
		.INIT('h4)
	) name7399 (
		_w7697_,
		_w9470_,
		_w11447_
	);
	LUT4 #(
		.INIT('h0040)
	) name7400 (
		_w9574_,
		_w9575_,
		_w9576_,
		_w11447_,
		_w11448_
	);
	LUT2 #(
		.INIT('h2)
	) name7401 (
		_w11333_,
		_w11448_,
		_w11449_
	);
	LUT3 #(
		.INIT('h02)
	) name7402 (
		_w11333_,
		_w11385_,
		_w11448_,
		_w11450_
	);
	LUT2 #(
		.INIT('h4)
	) name7403 (
		_w7336_,
		_w9470_,
		_w11451_
	);
	LUT4 #(
		.INIT('h0040)
	) name7404 (
		_w9596_,
		_w9597_,
		_w9598_,
		_w11451_,
		_w11452_
	);
	LUT2 #(
		.INIT('h2)
	) name7405 (
		_w11386_,
		_w11452_,
		_w11453_
	);
	LUT4 #(
		.INIT('hfd75)
	) name7406 (
		_w11333_,
		_w11385_,
		_w11448_,
		_w11452_,
		_w11454_
	);
	LUT4 #(
		.INIT('h1000)
	) name7407 (
		_w11348_,
		_w11357_,
		_w11388_,
		_w11382_,
		_w11455_
	);
	LUT2 #(
		.INIT('h4)
	) name7408 (
		_w7205_,
		_w9470_,
		_w11456_
	);
	LUT4 #(
		.INIT('h0040)
	) name7409 (
		_w9659_,
		_w9660_,
		_w9661_,
		_w11456_,
		_w11457_
	);
	LUT2 #(
		.INIT('h2)
	) name7410 (
		_w11333_,
		_w11457_,
		_w11458_
	);
	LUT3 #(
		.INIT('h02)
	) name7411 (
		_w11333_,
		_w11385_,
		_w11457_,
		_w11459_
	);
	LUT4 #(
		.INIT('hf400)
	) name7412 (
		_w11444_,
		_w11428_,
		_w11455_,
		_w11459_,
		_w11460_
	);
	LUT3 #(
		.INIT('h0e)
	) name7413 (
		_w11446_,
		_w11454_,
		_w11460_,
		_w11461_
	);
	LUT4 #(
		.INIT('h1000)
	) name7414 (
		_w11348_,
		_w11357_,
		_w11388_,
		_w11395_,
		_w11462_
	);
	LUT2 #(
		.INIT('h4)
	) name7415 (
		_w7868_,
		_w9470_,
		_w11463_
	);
	LUT4 #(
		.INIT('h0040)
	) name7416 (
		_w9618_,
		_w9619_,
		_w9620_,
		_w11463_,
		_w11464_
	);
	LUT2 #(
		.INIT('h2)
	) name7417 (
		_w11333_,
		_w11464_,
		_w11465_
	);
	LUT3 #(
		.INIT('h02)
	) name7418 (
		_w11333_,
		_w11385_,
		_w11464_,
		_w11466_
	);
	LUT2 #(
		.INIT('h4)
	) name7419 (
		_w8013_,
		_w9470_,
		_w11467_
	);
	LUT4 #(
		.INIT('h0040)
	) name7420 (
		_w9636_,
		_w9637_,
		_w9638_,
		_w11467_,
		_w11468_
	);
	LUT2 #(
		.INIT('h2)
	) name7421 (
		_w11333_,
		_w11468_,
		_w11469_
	);
	LUT3 #(
		.INIT('h08)
	) name7422 (
		_w11333_,
		_w11385_,
		_w11468_,
		_w11470_
	);
	LUT4 #(
		.INIT('hfd75)
	) name7423 (
		_w11333_,
		_w11385_,
		_w11464_,
		_w11468_,
		_w11471_
	);
	LUT4 #(
		.INIT('h00f4)
	) name7424 (
		_w11444_,
		_w11423_,
		_w11462_,
		_w11471_,
		_w11472_
	);
	LUT2 #(
		.INIT('h8)
	) name7425 (
		_w11371_,
		_w11390_,
		_w11473_
	);
	LUT2 #(
		.INIT('h8)
	) name7426 (
		_w11473_,
		_w11389_,
		_w11474_
	);
	LUT3 #(
		.INIT('h80)
	) name7427 (
		_w11473_,
		_w11389_,
		_w11341_,
		_w11475_
	);
	LUT2 #(
		.INIT('h8)
	) name7428 (
		_w11390_,
		_w11404_,
		_w11476_
	);
	LUT3 #(
		.INIT('h13)
	) name7429 (
		_w11390_,
		_w11395_,
		_w11404_,
		_w11477_
	);
	LUT4 #(
		.INIT('h0040)
	) name7430 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11406_,
		_w11477_,
		_w11478_
	);
	LUT2 #(
		.INIT('h1)
	) name7431 (
		_w11475_,
		_w11478_,
		_w11479_
	);
	LUT3 #(
		.INIT('h01)
	) name7432 (
		_w11472_,
		_w11475_,
		_w11478_,
		_w11480_
	);
	LUT4 #(
		.INIT('h1000)
	) name7433 (
		_w11348_,
		_w11357_,
		_w11388_,
		_w11418_,
		_w11481_
	);
	LUT2 #(
		.INIT('h4)
	) name7434 (
		_w6877_,
		_w9470_,
		_w11482_
	);
	LUT4 #(
		.INIT('h0040)
	) name7435 (
		_w9529_,
		_w9530_,
		_w9531_,
		_w11482_,
		_w11483_
	);
	LUT2 #(
		.INIT('h2)
	) name7436 (
		_w11333_,
		_w11483_,
		_w11484_
	);
	LUT3 #(
		.INIT('h02)
	) name7437 (
		_w11333_,
		_w11385_,
		_w11483_,
		_w11485_
	);
	LUT2 #(
		.INIT('h4)
	) name7438 (
		_w5884_,
		_w9470_,
		_w11486_
	);
	LUT2 #(
		.INIT('h1)
	) name7439 (
		_w9550_,
		_w11486_,
		_w11487_
	);
	LUT3 #(
		.INIT('hc8)
	) name7440 (
		_w9550_,
		_w11386_,
		_w11486_,
		_w11488_
	);
	LUT2 #(
		.INIT('h1)
	) name7441 (
		_w11485_,
		_w11488_,
		_w11489_
	);
	LUT4 #(
		.INIT('h00f4)
	) name7442 (
		_w11444_,
		_w11414_,
		_w11481_,
		_w11489_,
		_w11490_
	);
	LUT2 #(
		.INIT('h8)
	) name7443 (
		_w11400_,
		_w11391_,
		_w11491_
	);
	LUT4 #(
		.INIT('h23af)
	) name7444 (
		_w11444_,
		_w11389_,
		_w11392_,
		_w11491_,
		_w11492_
	);
	LUT2 #(
		.INIT('h4)
	) name7445 (
		_w6327_,
		_w9470_,
		_w11493_
	);
	LUT4 #(
		.INIT('h0040)
	) name7446 (
		_w9696_,
		_w9697_,
		_w9698_,
		_w11493_,
		_w11494_
	);
	LUT2 #(
		.INIT('h2)
	) name7447 (
		_w11333_,
		_w11494_,
		_w11495_
	);
	LUT3 #(
		.INIT('h02)
	) name7448 (
		_w11333_,
		_w11385_,
		_w11494_,
		_w11496_
	);
	LUT2 #(
		.INIT('h4)
	) name7449 (
		_w6003_,
		_w9470_,
		_w11497_
	);
	LUT4 #(
		.INIT('h0040)
	) name7450 (
		_w9718_,
		_w9719_,
		_w9720_,
		_w11497_,
		_w11498_
	);
	LUT2 #(
		.INIT('h2)
	) name7451 (
		_w11333_,
		_w11498_,
		_w11499_
	);
	LUT3 #(
		.INIT('h08)
	) name7452 (
		_w11333_,
		_w11385_,
		_w11498_,
		_w11500_
	);
	LUT4 #(
		.INIT('hfd75)
	) name7453 (
		_w11333_,
		_w11385_,
		_w11494_,
		_w11498_,
		_w11501_
	);
	LUT3 #(
		.INIT('h54)
	) name7454 (
		_w11490_,
		_w11492_,
		_w11501_,
		_w11502_
	);
	LUT2 #(
		.INIT('h8)
	) name7455 (
		_w11400_,
		_w11404_,
		_w11503_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name7456 (
		_w11444_,
		_w11389_,
		_w11503_,
		_w11476_,
		_w11504_
	);
	LUT2 #(
		.INIT('h4)
	) name7457 (
		_w6128_,
		_w9470_,
		_w11505_
	);
	LUT4 #(
		.INIT('h0040)
	) name7458 (
		_w9483_,
		_w9484_,
		_w9485_,
		_w11505_,
		_w11506_
	);
	LUT2 #(
		.INIT('h2)
	) name7459 (
		_w11333_,
		_w11506_,
		_w11507_
	);
	LUT3 #(
		.INIT('h02)
	) name7460 (
		_w11333_,
		_w11385_,
		_w11506_,
		_w11508_
	);
	LUT2 #(
		.INIT('h4)
	) name7461 (
		_w6464_,
		_w9470_,
		_w11509_
	);
	LUT4 #(
		.INIT('h0040)
	) name7462 (
		_w9510_,
		_w9511_,
		_w9512_,
		_w11509_,
		_w11510_
	);
	LUT2 #(
		.INIT('h2)
	) name7463 (
		_w11386_,
		_w11510_,
		_w11511_
	);
	LUT4 #(
		.INIT('hfd75)
	) name7464 (
		_w11333_,
		_w11385_,
		_w11506_,
		_w11510_,
		_w11512_
	);
	LUT2 #(
		.INIT('h4)
	) name7465 (
		_w7530_,
		_w9470_,
		_w11513_
	);
	LUT4 #(
		.INIT('h0040)
	) name7466 (
		_w9677_,
		_w9678_,
		_w9679_,
		_w11513_,
		_w11514_
	);
	LUT2 #(
		.INIT('h2)
	) name7467 (
		_w11386_,
		_w11514_,
		_w11515_
	);
	LUT4 #(
		.INIT('hf400)
	) name7468 (
		_w11444_,
		_w11428_,
		_w11455_,
		_w11515_,
		_w11516_
	);
	LUT3 #(
		.INIT('h0e)
	) name7469 (
		_w11504_,
		_w11512_,
		_w11516_,
		_w11517_
	);
	LUT4 #(
		.INIT('h8000)
	) name7470 (
		_w11502_,
		_w11517_,
		_w11461_,
		_w11480_,
		_w11518_
	);
	LUT4 #(
		.INIT('h4000)
	) name7471 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11423_,
		_w11519_
	);
	LUT4 #(
		.INIT('h1000)
	) name7472 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11428_,
		_w11520_
	);
	LUT2 #(
		.INIT('h1)
	) name7473 (
		_w11519_,
		_w11520_,
		_w11521_
	);
	LUT4 #(
		.INIT('h4000)
	) name7474 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11418_,
		_w11522_
	);
	LUT2 #(
		.INIT('h8)
	) name7475 (
		_w11386_,
		_w11415_,
		_w11523_
	);
	LUT2 #(
		.INIT('h8)
	) name7476 (
		_w11389_,
		_w11476_,
		_w11524_
	);
	LUT3 #(
		.INIT('h01)
	) name7477 (
		_w11522_,
		_w11523_,
		_w11524_,
		_w11525_
	);
	LUT3 #(
		.INIT('h2a)
	) name7478 (
		_w11341_,
		_w11521_,
		_w11525_,
		_w11526_
	);
	LUT2 #(
		.INIT('h4)
	) name7479 (
		_w8288_,
		_w9470_,
		_w11527_
	);
	LUT4 #(
		.INIT('h0040)
	) name7480 (
		_w9808_,
		_w9809_,
		_w9810_,
		_w11527_,
		_w11528_
	);
	LUT4 #(
		.INIT('h1000)
	) name7481 (
		_w11348_,
		_w11357_,
		_w11388_,
		_w11405_,
		_w11529_
	);
	LUT4 #(
		.INIT('h00bf)
	) name7482 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11439_,
		_w11529_,
		_w11530_
	);
	LUT3 #(
		.INIT('h02)
	) name7483 (
		_w11386_,
		_w11530_,
		_w11528_,
		_w11531_
	);
	LUT2 #(
		.INIT('h2)
	) name7484 (
		_w11333_,
		_w11335_,
		_w11532_
	);
	LUT3 #(
		.INIT('h04)
	) name7485 (
		_w11386_,
		_w11532_,
		_w11530_,
		_w11533_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name7486 (
		_w11473_,
		_w11444_,
		_w11401_,
		_w11389_,
		_w11534_
	);
	LUT2 #(
		.INIT('h4)
	) name7487 (
		_w5751_,
		_w9470_,
		_w11535_
	);
	LUT4 #(
		.INIT('h0040)
	) name7488 (
		_w9773_,
		_w9774_,
		_w9775_,
		_w11535_,
		_w11536_
	);
	LUT2 #(
		.INIT('h2)
	) name7489 (
		_w11333_,
		_w11536_,
		_w11537_
	);
	LUT3 #(
		.INIT('h02)
	) name7490 (
		_w11333_,
		_w11536_,
		_w11385_,
		_w11538_
	);
	LUT2 #(
		.INIT('h4)
	) name7491 (
		_w6723_,
		_w9470_,
		_w11539_
	);
	LUT4 #(
		.INIT('h0040)
	) name7492 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w11539_,
		_w11540_
	);
	LUT2 #(
		.INIT('h2)
	) name7493 (
		_w11386_,
		_w11540_,
		_w11541_
	);
	LUT4 #(
		.INIT('hfd5d)
	) name7494 (
		_w11333_,
		_w11536_,
		_w11385_,
		_w11540_,
		_w11542_
	);
	LUT4 #(
		.INIT('ha820)
	) name7495 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001 ,
		_w11543_
	);
	LUT3 #(
		.INIT('h0e)
	) name7496 (
		_w11534_,
		_w11542_,
		_w11543_,
		_w11544_
	);
	LUT3 #(
		.INIT('h10)
	) name7497 (
		_w11533_,
		_w11531_,
		_w11544_,
		_w11545_
	);
	LUT4 #(
		.INIT('h2000)
	) name7498 (
		_w11442_,
		_w11526_,
		_w11545_,
		_w11518_,
		_w11546_
	);
	LUT4 #(
		.INIT('h1000)
	) name7499 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11414_,
		_w11547_
	);
	LUT4 #(
		.INIT('h2000)
	) name7500 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11434_,
		_w11548_
	);
	LUT3 #(
		.INIT('ha8)
	) name7501 (
		_w11341_,
		_w11547_,
		_w11548_,
		_w11549_
	);
	LUT4 #(
		.INIT('h4000)
	) name7502 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11402_,
		_w11405_,
		_w11550_
	);
	LUT4 #(
		.INIT('h4000)
	) name7503 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11341_,
		_w11358_,
		_w11445_,
		_w11551_
	);
	LUT3 #(
		.INIT('h40)
	) name7504 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11401_,
		_w11358_,
		_w11552_
	);
	LUT4 #(
		.INIT('h4000)
	) name7505 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11401_,
		_w11358_,
		_w11402_,
		_w11553_
	);
	LUT3 #(
		.INIT('h01)
	) name7506 (
		_w11550_,
		_w11551_,
		_w11553_,
		_w11554_
	);
	LUT4 #(
		.INIT('h1000)
	) name7507 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11418_,
		_w11555_
	);
	LUT3 #(
		.INIT('h80)
	) name7508 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11491_,
		_w11556_
	);
	LUT4 #(
		.INIT('h2000)
	) name7509 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11491_,
		_w11557_
	);
	LUT4 #(
		.INIT('h4000)
	) name7510 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11503_,
		_w11558_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7511 (
		_w11341_,
		_w11555_,
		_w11557_,
		_w11558_,
		_w11559_
	);
	LUT3 #(
		.INIT('h04)
	) name7512 (
		_w11549_,
		_w11554_,
		_w11559_,
		_w11560_
	);
	LUT4 #(
		.INIT('haa08)
	) name7513 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11337_,
		_w11344_,
		_w11347_,
		_w11561_
	);
	LUT2 #(
		.INIT('h8)
	) name7514 (
		_w11357_,
		_w11341_,
		_w11562_
	);
	LUT3 #(
		.INIT('h80)
	) name7515 (
		_w11357_,
		_w11341_,
		_w11561_,
		_w11563_
	);
	LUT2 #(
		.INIT('h4)
	) name7516 (
		_w11375_,
		_w11341_,
		_w11564_
	);
	LUT3 #(
		.INIT('h80)
	) name7517 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11564_,
		_w11565_
	);
	LUT3 #(
		.INIT('h1d)
	) name7518 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11348_,
		_w11353_,
		_w11566_
	);
	LUT2 #(
		.INIT('h8)
	) name7519 (
		_w11562_,
		_w11566_,
		_w11567_
	);
	LUT2 #(
		.INIT('h1)
	) name7520 (
		_w11565_,
		_w11567_,
		_w11568_
	);
	LUT3 #(
		.INIT('h01)
	) name7521 (
		_w11563_,
		_w11565_,
		_w11567_,
		_w11569_
	);
	LUT4 #(
		.INIT('h4000)
	) name7522 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11473_,
		_w11341_,
		_w11358_,
		_w11570_
	);
	LUT4 #(
		.INIT('h0001)
	) name7523 (
		_w11563_,
		_w11565_,
		_w11567_,
		_w11570_,
		_w11571_
	);
	LUT4 #(
		.INIT('h8000)
	) name7524 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11491_,
		_w11572_
	);
	LUT2 #(
		.INIT('h4)
	) name7525 (
		_w11340_,
		_w11572_,
		_w11573_
	);
	LUT2 #(
		.INIT('h2)
	) name7526 (
		_w11571_,
		_w11573_,
		_w11574_
	);
	LUT4 #(
		.INIT('h8000)
	) name7527 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11406_,
		_w11503_,
		_w11575_
	);
	LUT4 #(
		.INIT('h8000)
	) name7528 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11402_,
		_w11434_,
		_w11576_
	);
	LUT2 #(
		.INIT('h1)
	) name7529 (
		_w11575_,
		_w11576_,
		_w11577_
	);
	LUT4 #(
		.INIT('h1000)
	) name7530 (
		_w11348_,
		_w11357_,
		_w11388_,
		_w11423_,
		_w11578_
	);
	LUT4 #(
		.INIT('h8880)
	) name7531 (
		_w11389_,
		_w11406_,
		_w11423_,
		_w11445_,
		_w11579_
	);
	LUT3 #(
		.INIT('h01)
	) name7532 (
		_w11575_,
		_w11576_,
		_w11579_,
		_w11580_
	);
	LUT4 #(
		.INIT('h4000)
	) name7533 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11341_,
		_w11358_,
		_w11392_,
		_w11581_
	);
	LUT2 #(
		.INIT('h8)
	) name7534 (
		_w11406_,
		_w11429_,
		_w11582_
	);
	LUT2 #(
		.INIT('h1)
	) name7535 (
		_w11581_,
		_w11582_,
		_w11583_
	);
	LUT4 #(
		.INIT('h2000)
	) name7536 (
		_w11571_,
		_w11573_,
		_w11580_,
		_w11583_,
		_w11584_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name7537 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11401_,
		_w11358_,
		_w11439_,
		_w11585_
	);
	LUT2 #(
		.INIT('h2)
	) name7538 (
		_w11406_,
		_w11585_,
		_w11586_
	);
	LUT4 #(
		.INIT('h4000)
	) name7539 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11434_,
		_w11587_
	);
	LUT4 #(
		.INIT('h1000)
	) name7540 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11503_,
		_w11588_
	);
	LUT3 #(
		.INIT('h40)
	) name7541 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11491_,
		_w11589_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7542 (
		_w11341_,
		_w11588_,
		_w11587_,
		_w11589_,
		_w11590_
	);
	LUT4 #(
		.INIT('h8880)
	) name7543 (
		_w11389_,
		_w11402_,
		_w11423_,
		_w11445_,
		_w11591_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name7544 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11503_,
		_w11476_,
		_w11592_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name7545 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11382_,
		_w11428_,
		_w11593_
	);
	LUT3 #(
		.INIT('hd5)
	) name7546 (
		_w11386_,
		_w11592_,
		_w11593_,
		_w11594_
	);
	LUT4 #(
		.INIT('h0888)
	) name7547 (
		_w11386_,
		_w11341_,
		_w11592_,
		_w11593_,
		_w11595_
	);
	LUT4 #(
		.INIT('h0001)
	) name7548 (
		_w11591_,
		_w11586_,
		_w11590_,
		_w11595_,
		_w11596_
	);
	LUT3 #(
		.INIT('h80)
	) name7549 (
		_w11560_,
		_w11584_,
		_w11596_,
		_w11597_
	);
	LUT4 #(
		.INIT('h4000)
	) name7550 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11433_,
		_w11546_,
		_w11597_,
		_w11598_
	);
	LUT4 #(
		.INIT('h222e)
	) name7551 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001 ,
		_w11329_,
		_w11332_,
		_w11598_,
		_w11599_
	);
	LUT3 #(
		.INIT('h8a)
	) name7552 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4094_,
		_w4097_,
		_w11600_
	);
	LUT3 #(
		.INIT('h40)
	) name7553 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		\core_c_dec_IRE_reg[1]/NET0131 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w11601_
	);
	LUT4 #(
		.INIT('h040f)
	) name7554 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w11600_,
		_w11601_,
		_w11602_
	);
	LUT4 #(
		.INIT('haaca)
	) name7555 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w9912_,
		_w11602_,
		_w11603_
	);
	LUT4 #(
		.INIT('h8000)
	) name7556 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w5053_,
		_w5052_,
		_w5054_,
		_w11604_
	);
	LUT2 #(
		.INIT('h8)
	) name7557 (
		_w9431_,
		_w11604_,
		_w11605_
	);
	LUT4 #(
		.INIT('h0040)
	) name7558 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w11606_
	);
	LUT4 #(
		.INIT('h4000)
	) name7559 (
		\memc_MMR_web_reg/NET0131 ,
		_w9431_,
		_w11604_,
		_w11606_,
		_w11607_
	);
	LUT4 #(
		.INIT('h0080)
	) name7560 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w11608_
	);
	LUT4 #(
		.INIT('h4000)
	) name7561 (
		\memc_MMR_web_reg/NET0131 ,
		_w9431_,
		_w11604_,
		_w11608_,
		_w11609_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name7562 (
		_w8757_,
		_w8760_,
		_w11607_,
		_w11609_,
		_w11610_
	);
	LUT4 #(
		.INIT('hf1f0)
	) name7563 (
		_w8757_,
		_w8760_,
		_w11607_,
		_w11609_,
		_w11611_
	);
	LUT2 #(
		.INIT('h8)
	) name7564 (
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w11610_,
		_w11612_
	);
	LUT4 #(
		.INIT('h1000)
	) name7565 (
		_w8757_,
		_w8760_,
		_w11605_,
		_w11608_,
		_w11613_
	);
	LUT2 #(
		.INIT('h2)
	) name7566 (
		_w11607_,
		_w11613_,
		_w11614_
	);
	LUT3 #(
		.INIT('h08)
	) name7567 (
		_w6758_,
		_w11607_,
		_w11613_,
		_w11615_
	);
	LUT2 #(
		.INIT('he)
	) name7568 (
		_w11612_,
		_w11615_,
		_w11616_
	);
	LUT4 #(
		.INIT('hccac)
	) name7569 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001 ,
		_w9914_,
		_w11602_,
		_w11617_
	);
	LUT4 #(
		.INIT('hccac)
	) name7570 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001 ,
		_w9914_,
		_w11602_,
		_w11618_
	);
	LUT4 #(
		.INIT('haaca)
	) name7571 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001 ,
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w9914_,
		_w11602_,
		_w11619_
	);
	LUT4 #(
		.INIT('haa3a)
	) name7572 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001 ,
		_w4155_,
		_w9914_,
		_w11602_,
		_w11620_
	);
	LUT4 #(
		.INIT('haaca)
	) name7573 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w9914_,
		_w11602_,
		_w11621_
	);
	LUT4 #(
		.INIT('haaca)
	) name7574 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w9914_,
		_w11602_,
		_w11622_
	);
	LUT4 #(
		.INIT('haaca)
	) name7575 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w9914_,
		_w11602_,
		_w11623_
	);
	LUT3 #(
		.INIT('h20)
	) name7576 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w9453_,
		_w9894_,
		_w11624_
	);
	LUT2 #(
		.INIT('h8)
	) name7577 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		_w9894_,
		_w11625_
	);
	LUT4 #(
		.INIT('h4544)
	) name7578 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w7927_,
		_w8040_,
		_w8042_,
		_w11626_
	);
	LUT2 #(
		.INIT('h2)
	) name7579 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8952_,
		_w11627_
	);
	LUT2 #(
		.INIT('h1)
	) name7580 (
		_w11626_,
		_w11627_,
		_w11628_
	);
	LUT3 #(
		.INIT('h13)
	) name7581 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001 ,
		_w9894_,
		_w11629_
	);
	LUT2 #(
		.INIT('h4)
	) name7582 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR0_E_reg/P0001 ,
		_w11630_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name7583 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_c_dec_updMR_E_reg/P0001 ,
		_w11305_,
		_w11631_
	);
	LUT2 #(
		.INIT('h8)
	) name7584 (
		_w9894_,
		_w11305_,
		_w11632_
	);
	LUT4 #(
		.INIT('h0002)
	) name7585 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w11629_,
		_w11633_
	);
	LUT4 #(
		.INIT('h5700)
	) name7586 (
		_w11625_,
		_w11626_,
		_w11627_,
		_w11633_,
		_w11634_
	);
	LUT3 #(
		.INIT('h40)
	) name7587 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 ,
		_w9894_,
		_w11305_,
		_w11635_
	);
	LUT4 #(
		.INIT('h313b)
	) name7588 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001 ,
		_w11631_,
		_w11635_,
		_w11636_
	);
	LUT4 #(
		.INIT('h6656)
	) name7589 (
		_w10290_,
		_w10304_,
		_w10305_,
		_w10317_,
		_w11637_
	);
	LUT2 #(
		.INIT('h1)
	) name7590 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11637_,
		_w11638_
	);
	LUT3 #(
		.INIT('h56)
	) name7591 (
		_w10256_,
		_w10269_,
		_w10270_,
		_w11639_
	);
	LUT4 #(
		.INIT('ha802)
	) name7592 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10289_,
		_w10318_,
		_w11639_,
		_w11640_
	);
	LUT3 #(
		.INIT('h02)
	) name7593 (
		_w11624_,
		_w11638_,
		_w11640_,
		_w11641_
	);
	LUT4 #(
		.INIT('hff45)
	) name7594 (
		_w11624_,
		_w11634_,
		_w11636_,
		_w11641_,
		_w11642_
	);
	LUT4 #(
		.INIT('haaca)
	) name7595 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w9914_,
		_w11602_,
		_w11643_
	);
	LUT4 #(
		.INIT('hccac)
	) name7596 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001 ,
		_w9914_,
		_w11602_,
		_w11644_
	);
	LUT4 #(
		.INIT('hccac)
	) name7597 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001 ,
		_w9914_,
		_w11602_,
		_w11645_
	);
	LUT4 #(
		.INIT('hccac)
	) name7598 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001 ,
		_w9914_,
		_w11602_,
		_w11646_
	);
	LUT4 #(
		.INIT('hccac)
	) name7599 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001 ,
		_w9914_,
		_w11602_,
		_w11647_
	);
	LUT4 #(
		.INIT('hccac)
	) name7600 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001 ,
		_w9914_,
		_w11602_,
		_w11648_
	);
	LUT4 #(
		.INIT('haaca)
	) name7601 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001 ,
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w9914_,
		_w11602_,
		_w11649_
	);
	LUT4 #(
		.INIT('hccac)
	) name7602 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001 ,
		_w9914_,
		_w11602_,
		_w11650_
	);
	LUT4 #(
		.INIT('hccac)
	) name7603 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001 ,
		_w9914_,
		_w11602_,
		_w11651_
	);
	LUT4 #(
		.INIT('hccac)
	) name7604 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001 ,
		_w9914_,
		_w11602_,
		_w11652_
	);
	LUT3 #(
		.INIT('ha8)
	) name7605 (
		_w9946_,
		_w11638_,
		_w11640_,
		_w11653_
	);
	LUT4 #(
		.INIT('h0040)
	) name7606 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR0_E_reg/P0001 ,
		_w9452_,
		_w11305_,
		_w11654_
	);
	LUT3 #(
		.INIT('h10)
	) name7607 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11654_,
		_w11655_
	);
	LUT4 #(
		.INIT('h5040)
	) name7608 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR0_E_reg/P0001 ,
		_w9452_,
		_w11305_,
		_w11656_
	);
	LUT2 #(
		.INIT('h2)
	) name7609 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001 ,
		_w11656_,
		_w11657_
	);
	LUT3 #(
		.INIT('h40)
	) name7610 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 ,
		_w11300_,
		_w11305_,
		_w11658_
	);
	LUT3 #(
		.INIT('h10)
	) name7611 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11658_,
		_w11659_
	);
	LUT3 #(
		.INIT('h01)
	) name7612 (
		_w9946_,
		_w11657_,
		_w11659_,
		_w11660_
	);
	LUT4 #(
		.INIT('hef00)
	) name7613 (
		_w11626_,
		_w11627_,
		_w11655_,
		_w11660_,
		_w11661_
	);
	LUT2 #(
		.INIT('h1)
	) name7614 (
		_w11653_,
		_w11661_,
		_w11662_
	);
	LUT4 #(
		.INIT('hccac)
	) name7615 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001 ,
		_w9914_,
		_w11602_,
		_w11663_
	);
	LUT4 #(
		.INIT('hccac)
	) name7616 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001 ,
		_w9914_,
		_w11602_,
		_w11664_
	);
	LUT4 #(
		.INIT('hccac)
	) name7617 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001 ,
		_w9914_,
		_w11602_,
		_w11665_
	);
	LUT4 #(
		.INIT('hccac)
	) name7618 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001 ,
		_w9914_,
		_w11602_,
		_w11666_
	);
	LUT4 #(
		.INIT('hccac)
	) name7619 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001 ,
		_w9914_,
		_w11602_,
		_w11667_
	);
	LUT4 #(
		.INIT('hccac)
	) name7620 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001 ,
		_w9914_,
		_w11602_,
		_w11668_
	);
	LUT4 #(
		.INIT('hccac)
	) name7621 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001 ,
		_w9914_,
		_w11602_,
		_w11669_
	);
	LUT4 #(
		.INIT('haaca)
	) name7622 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w9914_,
		_w11602_,
		_w11670_
	);
	LUT4 #(
		.INIT('hccac)
	) name7623 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001 ,
		_w9922_,
		_w11602_,
		_w11671_
	);
	LUT4 #(
		.INIT('hccac)
	) name7624 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001 ,
		_w9922_,
		_w11602_,
		_w11672_
	);
	LUT4 #(
		.INIT('h0001)
	) name7625 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		\sport0_txctl_TX_reg[2]/P0001 ,
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w11673_
	);
	LUT4 #(
		.INIT('h0100)
	) name7626 (
		\sport0_txctl_TX_reg[4]/P0001 ,
		\sport0_txctl_TX_reg[5]/P0001 ,
		\sport0_txctl_TX_reg[6]/P0001 ,
		_w11673_,
		_w11674_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7627 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[7]/P0001 ,
		\sport0_txctl_TX_reg[8]/P0001 ,
		_w11674_,
		_w11675_
	);
	LUT2 #(
		.INIT('h6)
	) name7628 (
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w11675_,
		_w11676_
	);
	LUT4 #(
		.INIT('h785a)
	) name7629 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[4]/P0001 ,
		\sport0_txctl_TX_reg[5]/P0001 ,
		_w11673_,
		_w11677_
	);
	LUT3 #(
		.INIT('h87)
	) name7630 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w11678_
	);
	LUT4 #(
		.INIT('h0440)
	) name7631 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w11679_
	);
	LUT4 #(
		.INIT('hc837)
	) name7632 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		\sport0_txctl_TX_reg[2]/P0001 ,
		_w11680_
	);
	LUT4 #(
		.INIT('hccc8)
	) name7633 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		\sport0_txctl_TX_reg[2]/P0001 ,
		_w11681_
	);
	LUT4 #(
		.INIT('h0408)
	) name7634 (
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w11679_,
		_w11680_,
		_w11681_,
		_w11682_
	);
	LUT3 #(
		.INIT('h39)
	) name7635 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[4]/P0001 ,
		_w11673_,
		_w11683_
	);
	LUT2 #(
		.INIT('h2)
	) name7636 (
		_w11682_,
		_w11683_,
		_w11684_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name7637 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11677_,
		_w11682_,
		_w11683_,
		_w11685_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7638 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[4]/P0001 ,
		\sport0_txctl_TX_reg[5]/P0001 ,
		_w11673_,
		_w11686_
	);
	LUT2 #(
		.INIT('h6)
	) name7639 (
		\sport0_txctl_TX_reg[6]/P0001 ,
		_w11686_,
		_w11687_
	);
	LUT3 #(
		.INIT('hc6)
	) name7640 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[7]/P0001 ,
		_w11674_,
		_w11688_
	);
	LUT4 #(
		.INIT('h785a)
	) name7641 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[7]/P0001 ,
		\sport0_txctl_TX_reg[8]/P0001 ,
		_w11674_,
		_w11689_
	);
	LUT4 #(
		.INIT('h4000)
	) name7642 (
		_w11685_,
		_w11687_,
		_w11688_,
		_w11689_,
		_w11690_
	);
	LUT4 #(
		.INIT('h0100)
	) name7643 (
		\sport0_txctl_TX_reg[7]/P0001 ,
		\sport0_txctl_TX_reg[8]/P0001 ,
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w11674_,
		_w11691_
	);
	LUT3 #(
		.INIT('ha6)
	) name7644 (
		\sport0_txctl_TX_reg[10]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w11691_,
		_w11692_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name7645 (
		\sport0_txctl_TX_reg[10]/P0001 ,
		\sport0_txctl_TX_reg[11]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w11691_,
		_w11693_
	);
	LUT4 #(
		.INIT('h8000)
	) name7646 (
		_w11676_,
		_w11690_,
		_w11692_,
		_w11693_,
		_w11694_
	);
	LUT3 #(
		.INIT('he0)
	) name7647 (
		\sport0_txctl_TX_reg[10]/P0001 ,
		\sport0_txctl_TX_reg[11]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w11695_
	);
	LUT4 #(
		.INIT('h55a6)
	) name7648 (
		\sport0_txctl_TX_reg[12]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w11691_,
		_w11695_,
		_w11696_
	);
	LUT2 #(
		.INIT('h6)
	) name7649 (
		_w11694_,
		_w11696_,
		_w11697_
	);
	LUT3 #(
		.INIT('h28)
	) name7650 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11694_,
		_w11696_,
		_w11698_
	);
	LUT2 #(
		.INIT('h2)
	) name7651 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11677_,
		_w11699_
	);
	LUT3 #(
		.INIT('h01)
	) name7652 (
		\sport0_txctl_TX_reg[10]/P0001 ,
		\sport0_txctl_TX_reg[11]/P0001 ,
		\sport0_txctl_TX_reg[12]/P0001 ,
		_w11700_
	);
	LUT2 #(
		.INIT('h8)
	) name7653 (
		\sport0_txctl_TX_reg[13]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w11701_
	);
	LUT4 #(
		.INIT('h80aa)
	) name7654 (
		\sport0_txctl_TX_reg[14]/P0001 ,
		_w11691_,
		_w11700_,
		_w11701_,
		_w11702_
	);
	LUT3 #(
		.INIT('h32)
	) name7655 (
		\sport0_txctl_TX_reg[13]/P0001 ,
		\sport0_txctl_TX_reg[14]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w11703_
	);
	LUT2 #(
		.INIT('h1)
	) name7656 (
		_w11702_,
		_w11703_,
		_w11704_
	);
	LUT4 #(
		.INIT('hf700)
	) name7657 (
		_w11694_,
		_w11696_,
		_w11699_,
		_w11704_,
		_w11705_
	);
	LUT2 #(
		.INIT('h4)
	) name7658 (
		_w11698_,
		_w11705_,
		_w11706_
	);
	LUT4 #(
		.INIT('h0080)
	) name7659 (
		_w11676_,
		_w11690_,
		_w11692_,
		_w11699_,
		_w11707_
	);
	LUT4 #(
		.INIT('h2a80)
	) name7660 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11676_,
		_w11690_,
		_w11692_,
		_w11708_
	);
	LUT4 #(
		.INIT('h00eb)
	) name7661 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11693_,
		_w11707_,
		_w11708_,
		_w11709_
	);
	LUT3 #(
		.INIT('h40)
	) name7662 (
		_w11698_,
		_w11705_,
		_w11709_,
		_w11710_
	);
	LUT3 #(
		.INIT('h28)
	) name7663 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11693_,
		_w11707_,
		_w11711_
	);
	LUT4 #(
		.INIT('h9100)
	) name7664 (
		_w11694_,
		_w11696_,
		_w11699_,
		_w11704_,
		_w11712_
	);
	LUT2 #(
		.INIT('h4)
	) name7665 (
		_w11711_,
		_w11712_,
		_w11713_
	);
	LUT2 #(
		.INIT('h8)
	) name7666 (
		_w11710_,
		_w11713_,
		_w11714_
	);
	LUT4 #(
		.INIT('h1540)
	) name7667 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11676_,
		_w11690_,
		_w11692_,
		_w11715_
	);
	LUT4 #(
		.INIT('h2888)
	) name7668 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11676_,
		_w11677_,
		_w11690_,
		_w11716_
	);
	LUT2 #(
		.INIT('h1)
	) name7669 (
		_w11715_,
		_w11716_,
		_w11717_
	);
	LUT3 #(
		.INIT('h40)
	) name7670 (
		_w11698_,
		_w11705_,
		_w11717_,
		_w11718_
	);
	LUT3 #(
		.INIT('h3b)
	) name7671 (
		_w11710_,
		_w11713_,
		_w11718_,
		_w11719_
	);
	LUT4 #(
		.INIT('h297c)
	) name7672 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11677_,
		_w11684_,
		_w11687_,
		_w11720_
	);
	LUT3 #(
		.INIT('h40)
	) name7673 (
		_w11698_,
		_w11705_,
		_w11720_,
		_w11721_
	);
	LUT4 #(
		.INIT('h0f4b)
	) name7674 (
		_w11685_,
		_w11687_,
		_w11688_,
		_w11699_,
		_w11722_
	);
	LUT3 #(
		.INIT('h82)
	) name7675 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11685_,
		_w11687_,
		_w11723_
	);
	LUT3 #(
		.INIT('h0e)
	) name7676 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11722_,
		_w11723_,
		_w11724_
	);
	LUT3 #(
		.INIT('h40)
	) name7677 (
		_w11698_,
		_w11705_,
		_w11724_,
		_w11725_
	);
	LUT4 #(
		.INIT('h4000)
	) name7678 (
		_w11698_,
		_w11705_,
		_w11720_,
		_w11724_,
		_w11726_
	);
	LUT4 #(
		.INIT('hbf40)
	) name7679 (
		_w11685_,
		_w11687_,
		_w11688_,
		_w11689_,
		_w11727_
	);
	LUT3 #(
		.INIT('h8d)
	) name7680 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11722_,
		_w11727_,
		_w11728_
	);
	LUT3 #(
		.INIT('h40)
	) name7681 (
		_w11698_,
		_w11705_,
		_w11728_,
		_w11729_
	);
	LUT2 #(
		.INIT('h4)
	) name7682 (
		_w11726_,
		_w11729_,
		_w11730_
	);
	LUT4 #(
		.INIT('h1144)
	) name7683 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11676_,
		_w11677_,
		_w11690_,
		_w11731_
	);
	LUT2 #(
		.INIT('h8)
	) name7684 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11727_,
		_w11732_
	);
	LUT2 #(
		.INIT('h1)
	) name7685 (
		_w11731_,
		_w11732_,
		_w11733_
	);
	LUT3 #(
		.INIT('h40)
	) name7686 (
		_w11698_,
		_w11705_,
		_w11733_,
		_w11734_
	);
	LUT4 #(
		.INIT('h4000)
	) name7687 (
		_w11698_,
		_w11705_,
		_w11717_,
		_w11733_,
		_w11735_
	);
	LUT3 #(
		.INIT('h80)
	) name7688 (
		_w11710_,
		_w11713_,
		_w11735_,
		_w11736_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7689 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11719_,
		_w11730_,
		_w11736_,
		_w11737_
	);
	LUT4 #(
		.INIT('h4044)
	) name7690 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTTX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w11738_
	);
	LUT2 #(
		.INIT('h1)
	) name7691 (
		\auctl_T0Sack_reg/NET0131 ,
		_w11738_,
		_w11739_
	);
	LUT2 #(
		.INIT('he)
	) name7692 (
		\auctl_T0Sack_reg/NET0131 ,
		_w11738_,
		_w11740_
	);
	LUT4 #(
		.INIT('h0045)
	) name7693 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w11739_,
		_w11741_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name7694 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[4]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w11742_
	);
	LUT2 #(
		.INIT('h4)
	) name7695 (
		_w11741_,
		_w11742_,
		_w11743_
	);
	LUT2 #(
		.INIT('h1)
	) name7696 (
		_w11737_,
		_w11743_,
		_w11744_
	);
	LUT4 #(
		.INIT('haaca)
	) name7697 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001 ,
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w9922_,
		_w11602_,
		_w11745_
	);
	LUT4 #(
		.INIT('haa3a)
	) name7698 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001 ,
		_w4155_,
		_w9922_,
		_w11602_,
		_w11746_
	);
	LUT4 #(
		.INIT('haaca)
	) name7699 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w9922_,
		_w11602_,
		_w11747_
	);
	LUT4 #(
		.INIT('haaca)
	) name7700 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w9922_,
		_w11602_,
		_w11748_
	);
	LUT4 #(
		.INIT('haaca)
	) name7701 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w9922_,
		_w11602_,
		_w11749_
	);
	LUT4 #(
		.INIT('haaca)
	) name7702 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w9922_,
		_w11602_,
		_w11750_
	);
	LUT4 #(
		.INIT('hccac)
	) name7703 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001 ,
		_w9922_,
		_w11602_,
		_w11751_
	);
	LUT4 #(
		.INIT('hccac)
	) name7704 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001 ,
		_w9922_,
		_w11602_,
		_w11752_
	);
	LUT4 #(
		.INIT('hccac)
	) name7705 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001 ,
		_w9922_,
		_w11602_,
		_w11753_
	);
	LUT4 #(
		.INIT('hccac)
	) name7706 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001 ,
		_w9922_,
		_w11602_,
		_w11754_
	);
	LUT4 #(
		.INIT('hccac)
	) name7707 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001 ,
		_w9922_,
		_w11602_,
		_w11755_
	);
	LUT4 #(
		.INIT('haaca)
	) name7708 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001 ,
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w9922_,
		_w11602_,
		_w11756_
	);
	LUT4 #(
		.INIT('hccac)
	) name7709 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001 ,
		_w9922_,
		_w11602_,
		_w11757_
	);
	LUT4 #(
		.INIT('hccac)
	) name7710 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001 ,
		_w9922_,
		_w11602_,
		_w11758_
	);
	LUT4 #(
		.INIT('hccac)
	) name7711 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001 ,
		_w9922_,
		_w11602_,
		_w11759_
	);
	LUT4 #(
		.INIT('hccac)
	) name7712 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001 ,
		_w9922_,
		_w11602_,
		_w11760_
	);
	LUT4 #(
		.INIT('hccac)
	) name7713 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001 ,
		_w9922_,
		_w11602_,
		_w11761_
	);
	LUT4 #(
		.INIT('hccac)
	) name7714 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001 ,
		_w9922_,
		_w11602_,
		_w11762_
	);
	LUT4 #(
		.INIT('hccac)
	) name7715 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001 ,
		_w9922_,
		_w11602_,
		_w11763_
	);
	LUT4 #(
		.INIT('hccac)
	) name7716 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001 ,
		_w9922_,
		_w11602_,
		_w11764_
	);
	LUT4 #(
		.INIT('hccac)
	) name7717 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001 ,
		_w9922_,
		_w11602_,
		_w11765_
	);
	LUT4 #(
		.INIT('hccac)
	) name7718 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001 ,
		_w9922_,
		_w11602_,
		_w11766_
	);
	LUT4 #(
		.INIT('haaca)
	) name7719 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w9922_,
		_w11602_,
		_w11767_
	);
	LUT4 #(
		.INIT('hccac)
	) name7720 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001 ,
		_w9909_,
		_w11602_,
		_w11768_
	);
	LUT4 #(
		.INIT('hccac)
	) name7721 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001 ,
		_w9909_,
		_w11602_,
		_w11769_
	);
	LUT4 #(
		.INIT('haaca)
	) name7722 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001 ,
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w9909_,
		_w11602_,
		_w11770_
	);
	LUT4 #(
		.INIT('haa3a)
	) name7723 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001 ,
		_w4155_,
		_w9909_,
		_w11602_,
		_w11771_
	);
	LUT4 #(
		.INIT('haaca)
	) name7724 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w9909_,
		_w11602_,
		_w11772_
	);
	LUT4 #(
		.INIT('haaca)
	) name7725 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w9909_,
		_w11602_,
		_w11773_
	);
	LUT4 #(
		.INIT('haaca)
	) name7726 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w9909_,
		_w11602_,
		_w11774_
	);
	LUT4 #(
		.INIT('haaca)
	) name7727 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w9909_,
		_w11602_,
		_w11775_
	);
	LUT4 #(
		.INIT('hccac)
	) name7728 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001 ,
		_w9909_,
		_w11602_,
		_w11776_
	);
	LUT4 #(
		.INIT('hccac)
	) name7729 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001 ,
		_w9909_,
		_w11602_,
		_w11777_
	);
	LUT4 #(
		.INIT('hccac)
	) name7730 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001 ,
		_w9909_,
		_w11602_,
		_w11778_
	);
	LUT4 #(
		.INIT('hccac)
	) name7731 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001 ,
		_w9909_,
		_w11602_,
		_w11779_
	);
	LUT4 #(
		.INIT('hccac)
	) name7732 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001 ,
		_w9909_,
		_w11602_,
		_w11780_
	);
	LUT4 #(
		.INIT('haaca)
	) name7733 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001 ,
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w9909_,
		_w11602_,
		_w11781_
	);
	LUT4 #(
		.INIT('hccac)
	) name7734 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001 ,
		_w9909_,
		_w11602_,
		_w11782_
	);
	LUT4 #(
		.INIT('hccac)
	) name7735 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001 ,
		_w9909_,
		_w11602_,
		_w11783_
	);
	LUT4 #(
		.INIT('hccac)
	) name7736 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001 ,
		_w9909_,
		_w11602_,
		_w11784_
	);
	LUT4 #(
		.INIT('hccac)
	) name7737 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001 ,
		_w9909_,
		_w11602_,
		_w11785_
	);
	LUT4 #(
		.INIT('hccac)
	) name7738 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001 ,
		_w9909_,
		_w11602_,
		_w11786_
	);
	LUT4 #(
		.INIT('h4000)
	) name7739 (
		\memc_MMR_web_reg/NET0131 ,
		_w5657_,
		_w9431_,
		_w11604_,
		_w11787_
	);
	LUT4 #(
		.INIT('h00ef)
	) name7740 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w11787_,
		_w11788_
	);
	LUT2 #(
		.INIT('h8)
	) name7741 (
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w11788_,
		_w11789_
	);
	LUT4 #(
		.INIT('h0100)
	) name7742 (
		_w7140_,
		_w7240_,
		_w11613_,
		_w11787_,
		_w11790_
	);
	LUT2 #(
		.INIT('he)
	) name7743 (
		_w11789_,
		_w11790_,
		_w11791_
	);
	LUT4 #(
		.INIT('hccac)
	) name7744 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001 ,
		_w9909_,
		_w11602_,
		_w11792_
	);
	LUT4 #(
		.INIT('hccac)
	) name7745 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001 ,
		_w9909_,
		_w11602_,
		_w11793_
	);
	LUT4 #(
		.INIT('hccac)
	) name7746 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001 ,
		_w9909_,
		_w11602_,
		_w11794_
	);
	LUT4 #(
		.INIT('hccac)
	) name7747 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001 ,
		_w9909_,
		_w11602_,
		_w11795_
	);
	LUT2 #(
		.INIT('h8)
	) name7748 (
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w11788_,
		_w11796_
	);
	LUT4 #(
		.INIT('h0100)
	) name7749 (
		_w7465_,
		_w7565_,
		_w11613_,
		_w11787_,
		_w11797_
	);
	LUT2 #(
		.INIT('he)
	) name7750 (
		_w11796_,
		_w11797_,
		_w11798_
	);
	LUT4 #(
		.INIT('hccac)
	) name7751 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001 ,
		_w9909_,
		_w11602_,
		_w11799_
	);
	LUT4 #(
		.INIT('haaca)
	) name7752 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w9909_,
		_w11602_,
		_w11800_
	);
	LUT2 #(
		.INIT('h2)
	) name7753 (
		_w9908_,
		_w11602_,
		_w11801_
	);
	LUT3 #(
		.INIT('h54)
	) name7754 (
		_w4971_,
		_w9906_,
		_w9907_,
		_w11802_
	);
	LUT2 #(
		.INIT('h8)
	) name7755 (
		_w9921_,
		_w11602_,
		_w11803_
	);
	LUT4 #(
		.INIT('h1333)
	) name7756 (
		_w9910_,
		_w11801_,
		_w11802_,
		_w11803_,
		_w11804_
	);
	LUT2 #(
		.INIT('h9)
	) name7757 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w11804_,
		_w11805_
	);
	LUT2 #(
		.INIT('h1)
	) name7758 (
		_w9916_,
		_w11602_,
		_w11806_
	);
	LUT3 #(
		.INIT('hf8)
	) name7759 (
		_w9910_,
		_w11802_,
		_w11806_,
		_w11807_
	);
	LUT4 #(
		.INIT('h556a)
	) name7760 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		_w9910_,
		_w11802_,
		_w11806_,
		_w11808_
	);
	LUT2 #(
		.INIT('h8)
	) name7761 (
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w11788_,
		_w11809_
	);
	LUT3 #(
		.INIT('h20)
	) name7762 (
		_w8761_,
		_w11613_,
		_w11787_,
		_w11810_
	);
	LUT2 #(
		.INIT('he)
	) name7763 (
		_w11809_,
		_w11810_,
		_w11811_
	);
	LUT4 #(
		.INIT('h4144)
	) name7764 (
		_w9455_,
		_w9831_,
		_w9832_,
		_w9833_,
		_w11812_
	);
	LUT3 #(
		.INIT('h28)
	) name7765 (
		_w9455_,
		_w9738_,
		_w9762_,
		_w11813_
	);
	LUT4 #(
		.INIT('heee2)
	) name7766 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001 ,
		_w9895_,
		_w11812_,
		_w11813_,
		_w11814_
	);
	LUT2 #(
		.INIT('h8)
	) name7767 (
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w11788_,
		_w11815_
	);
	LUT3 #(
		.INIT('h20)
	) name7768 (
		_w5760_,
		_w11613_,
		_w11787_,
		_w11816_
	);
	LUT2 #(
		.INIT('he)
	) name7769 (
		_w11815_,
		_w11816_,
		_w11817_
	);
	LUT2 #(
		.INIT('h8)
	) name7770 (
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w11788_,
		_w11818_
	);
	LUT3 #(
		.INIT('h20)
	) name7771 (
		_w8802_,
		_w11613_,
		_w11787_,
		_w11819_
	);
	LUT2 #(
		.INIT('he)
	) name7772 (
		_w11818_,
		_w11819_,
		_w11820_
	);
	LUT2 #(
		.INIT('h8)
	) name7773 (
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w11788_,
		_w11821_
	);
	LUT3 #(
		.INIT('h20)
	) name7774 (
		_w6758_,
		_w11613_,
		_w11787_,
		_w11822_
	);
	LUT2 #(
		.INIT('he)
	) name7775 (
		_w11821_,
		_w11822_,
		_w11823_
	);
	LUT2 #(
		.INIT('h8)
	) name7776 (
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w11788_,
		_w11824_
	);
	LUT4 #(
		.INIT('h0100)
	) name7777 (
		_w6263_,
		_w6362_,
		_w11613_,
		_w11787_,
		_w11825_
	);
	LUT2 #(
		.INIT('he)
	) name7778 (
		_w11824_,
		_w11825_,
		_w11826_
	);
	LUT2 #(
		.INIT('h8)
	) name7779 (
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w11788_,
		_w11827_
	);
	LUT4 #(
		.INIT('h0100)
	) name7780 (
		_w5937_,
		_w6038_,
		_w11613_,
		_w11787_,
		_w11828_
	);
	LUT2 #(
		.INIT('he)
	) name7781 (
		_w11827_,
		_w11828_,
		_w11829_
	);
	LUT3 #(
		.INIT('h04)
	) name7782 (
		_w9453_,
		_w9894_,
		_w11328_,
		_w11830_
	);
	LUT4 #(
		.INIT('h4000)
	) name7783 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11392_,
		_w11831_
	);
	LUT3 #(
		.INIT('ha8)
	) name7784 (
		_w11341_,
		_w11520_,
		_w11831_,
		_w11832_
	);
	LUT2 #(
		.INIT('h2)
	) name7785 (
		_w11568_,
		_w11832_,
		_w11833_
	);
	LUT3 #(
		.INIT('h02)
	) name7786 (
		_w11568_,
		_w11570_,
		_w11832_,
		_w11834_
	);
	LUT3 #(
		.INIT('h0d)
	) name7787 (
		_w11341_,
		_w11398_,
		_w11595_,
		_w11835_
	);
	LUT2 #(
		.INIT('h8)
	) name7788 (
		_w11834_,
		_w11835_,
		_w11836_
	);
	LUT3 #(
		.INIT('h40)
	) name7789 (
		_w11582_,
		_w11834_,
		_w11835_,
		_w11837_
	);
	LUT2 #(
		.INIT('h2)
	) name7790 (
		_w11386_,
		_w11448_,
		_w11838_
	);
	LUT4 #(
		.INIT('h4000)
	) name7791 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11439_,
		_w11839_
	);
	LUT4 #(
		.INIT('h8caf)
	) name7792 (
		_w11534_,
		_w11464_,
		_w11838_,
		_w11839_,
		_w11840_
	);
	LUT2 #(
		.INIT('h2)
	) name7793 (
		_w11333_,
		_w11510_,
		_w11841_
	);
	LUT3 #(
		.INIT('h02)
	) name7794 (
		_w11333_,
		_w11385_,
		_w11510_,
		_w11842_
	);
	LUT2 #(
		.INIT('h2)
	) name7795 (
		_w11386_,
		_w11483_,
		_w11843_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name7796 (
		_w11333_,
		_w11385_,
		_w11483_,
		_w11510_,
		_w11844_
	);
	LUT4 #(
		.INIT('h00f4)
	) name7797 (
		_w11444_,
		_w11428_,
		_w11455_,
		_w11844_,
		_w11845_
	);
	LUT3 #(
		.INIT('h0d)
	) name7798 (
		_w11522_,
		_w11457_,
		_w11845_,
		_w11846_
	);
	LUT2 #(
		.INIT('h8)
	) name7799 (
		_w11840_,
		_w11846_,
		_w11847_
	);
	LUT3 #(
		.INIT('h08)
	) name7800 (
		_w11333_,
		_w11385_,
		_w11464_,
		_w11848_
	);
	LUT2 #(
		.INIT('h8)
	) name7801 (
		_w11529_,
		_w11848_,
		_w11849_
	);
	LUT3 #(
		.INIT('h02)
	) name7802 (
		_w11333_,
		_w11385_,
		_w11468_,
		_w11850_
	);
	LUT3 #(
		.INIT('h80)
	) name7803 (
		_w11401_,
		_w11389_,
		_w11850_,
		_w11851_
	);
	LUT3 #(
		.INIT('h08)
	) name7804 (
		_w11333_,
		_w11385_,
		_w11506_,
		_w11852_
	);
	LUT3 #(
		.INIT('h80)
	) name7805 (
		_w11389_,
		_w11491_,
		_w11852_,
		_w11853_
	);
	LUT2 #(
		.INIT('h2)
	) name7806 (
		_w11333_,
		_w11528_,
		_w11854_
	);
	LUT3 #(
		.INIT('h02)
	) name7807 (
		_w11333_,
		_w11385_,
		_w11528_,
		_w11855_
	);
	LUT3 #(
		.INIT('h80)
	) name7808 (
		_w11389_,
		_w11445_,
		_w11855_,
		_w11856_
	);
	LUT4 #(
		.INIT('h0001)
	) name7809 (
		_w11849_,
		_w11851_,
		_w11853_,
		_w11856_,
		_w11857_
	);
	LUT4 #(
		.INIT('ha820)
	) name7810 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001 ,
		_w11858_
	);
	LUT3 #(
		.INIT('h07)
	) name7811 (
		_w11402_,
		_w11429_,
		_w11858_,
		_w11859_
	);
	LUT2 #(
		.INIT('h2)
	) name7812 (
		_w11333_,
		_w11540_,
		_w11860_
	);
	LUT3 #(
		.INIT('h02)
	) name7813 (
		_w11333_,
		_w11385_,
		_w11540_,
		_w11861_
	);
	LUT3 #(
		.INIT('h80)
	) name7814 (
		_w11389_,
		_w11476_,
		_w11861_,
		_w11862_
	);
	LUT3 #(
		.INIT('hc8)
	) name7815 (
		_w9550_,
		_w11333_,
		_w11486_,
		_w11863_
	);
	LUT4 #(
		.INIT('h0c08)
	) name7816 (
		_w9550_,
		_w11333_,
		_w11385_,
		_w11486_,
		_w11864_
	);
	LUT2 #(
		.INIT('h8)
	) name7817 (
		_w11462_,
		_w11864_,
		_w11865_
	);
	LUT3 #(
		.INIT('h10)
	) name7818 (
		_w11862_,
		_w11865_,
		_w11859_,
		_w11866_
	);
	LUT4 #(
		.INIT('h0001)
	) name7819 (
		_w11403_,
		_w11407_,
		_w11575_,
		_w11576_,
		_w11867_
	);
	LUT3 #(
		.INIT('h80)
	) name7820 (
		_w11857_,
		_w11866_,
		_w11867_,
		_w11868_
	);
	LUT3 #(
		.INIT('ha8)
	) name7821 (
		_w11341_,
		_w11424_,
		_w11421_,
		_w11869_
	);
	LUT3 #(
		.INIT('ha8)
	) name7822 (
		_w11341_,
		_w11419_,
		_w11425_,
		_w11870_
	);
	LUT2 #(
		.INIT('h1)
	) name7823 (
		_w11869_,
		_w11870_,
		_w11871_
	);
	LUT2 #(
		.INIT('h2)
	) name7824 (
		_w11333_,
		_w11452_,
		_w11872_
	);
	LUT3 #(
		.INIT('h02)
	) name7825 (
		_w11333_,
		_w11385_,
		_w11452_,
		_w11873_
	);
	LUT2 #(
		.INIT('h2)
	) name7826 (
		_w11333_,
		_w11514_,
		_w11874_
	);
	LUT3 #(
		.INIT('h02)
	) name7827 (
		_w11333_,
		_w11385_,
		_w11514_,
		_w11875_
	);
	LUT4 #(
		.INIT('h8acf)
	) name7828 (
		_w11530_,
		_w11492_,
		_w11873_,
		_w11875_,
		_w11876_
	);
	LUT4 #(
		.INIT('h0777)
	) name7829 (
		_w11555_,
		_w11499_,
		_w11435_,
		_w11854_,
		_w11877_
	);
	LUT4 #(
		.INIT('h1000)
	) name7830 (
		_w11869_,
		_w11870_,
		_w11876_,
		_w11877_,
		_w11878_
	);
	LUT3 #(
		.INIT('h80)
	) name7831 (
		_w11847_,
		_w11868_,
		_w11878_,
		_w11879_
	);
	LUT3 #(
		.INIT('h80)
	) name7832 (
		_w11389_,
		_w11385_,
		_w11445_,
		_w11880_
	);
	LUT3 #(
		.INIT('h54)
	) name7833 (
		_w11536_,
		_w11587_,
		_w11880_,
		_w11881_
	);
	LUT2 #(
		.INIT('h4)
	) name7834 (
		_w11540_,
		_w11588_,
		_w11882_
	);
	LUT3 #(
		.INIT('ha8)
	) name7835 (
		_w11333_,
		_w11881_,
		_w11882_,
		_w11883_
	);
	LUT3 #(
		.INIT('h08)
	) name7836 (
		_w11386_,
		_w11415_,
		_w11457_,
		_w11884_
	);
	LUT4 #(
		.INIT('h8000)
	) name7837 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11406_,
		_w11491_,
		_w11885_
	);
	LUT3 #(
		.INIT('h40)
	) name7838 (
		_w11444_,
		_w11423_,
		_w11864_,
		_w11886_
	);
	LUT3 #(
		.INIT('h01)
	) name7839 (
		_w11885_,
		_w11886_,
		_w11884_,
		_w11887_
	);
	LUT2 #(
		.INIT('h4)
	) name7840 (
		_w11385_,
		_w11415_,
		_w11888_
	);
	LUT3 #(
		.INIT('h40)
	) name7841 (
		_w11385_,
		_w11415_,
		_w11499_,
		_w11889_
	);
	LUT4 #(
		.INIT('h8000)
	) name7842 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11395_,
		_w11496_,
		_w11890_
	);
	LUT3 #(
		.INIT('h20)
	) name7843 (
		_w11473_,
		_w11444_,
		_w11850_,
		_w11891_
	);
	LUT3 #(
		.INIT('h40)
	) name7844 (
		_w11444_,
		_w11392_,
		_w11852_,
		_w11892_
	);
	LUT4 #(
		.INIT('h0001)
	) name7845 (
		_w11889_,
		_w11890_,
		_w11891_,
		_w11892_,
		_w11893_
	);
	LUT3 #(
		.INIT('h80)
	) name7846 (
		_w11389_,
		_w11386_,
		_w11476_,
		_w11894_
	);
	LUT3 #(
		.INIT('hc8)
	) name7847 (
		_w11558_,
		_w11495_,
		_w11894_,
		_w11895_
	);
	LUT2 #(
		.INIT('h8)
	) name7848 (
		_w11386_,
		_w11578_,
		_w11896_
	);
	LUT3 #(
		.INIT('hc8)
	) name7849 (
		_w11409_,
		_w11532_,
		_w11896_,
		_w11897_
	);
	LUT4 #(
		.INIT('h1000)
	) name7850 (
		_w11895_,
		_w11897_,
		_w11887_,
		_w11893_,
		_w11898_
	);
	LUT2 #(
		.INIT('h4)
	) name7851 (
		_w11883_,
		_w11898_,
		_w11899_
	);
	LUT2 #(
		.INIT('h4)
	) name7852 (
		_w11549_,
		_w11441_,
		_w11900_
	);
	LUT4 #(
		.INIT('h4000)
	) name7853 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11341_,
		_w11358_,
		_w11491_,
		_w11901_
	);
	LUT3 #(
		.INIT('h04)
	) name7854 (
		_w11549_,
		_w11441_,
		_w11901_,
		_w11902_
	);
	LUT3 #(
		.INIT('h01)
	) name7855 (
		_w11550_,
		_w11551_,
		_w11436_,
		_w11903_
	);
	LUT3 #(
		.INIT('h31)
	) name7856 (
		_w11406_,
		_w11553_,
		_w11585_,
		_w11904_
	);
	LUT3 #(
		.INIT('h80)
	) name7857 (
		_w11479_,
		_w11903_,
		_w11904_,
		_w11905_
	);
	LUT2 #(
		.INIT('h8)
	) name7858 (
		_w11406_,
		_w11578_,
		_w11906_
	);
	LUT2 #(
		.INIT('h8)
	) name7859 (
		_w11341_,
		_w11519_,
		_w11907_
	);
	LUT2 #(
		.INIT('h4)
	) name7860 (
		_w11385_,
		_w11581_,
		_w11908_
	);
	LUT3 #(
		.INIT('h23)
	) name7861 (
		_w11340_,
		_w11563_,
		_w11572_,
		_w11909_
	);
	LUT3 #(
		.INIT('h10)
	) name7862 (
		_w11907_,
		_w11908_,
		_w11909_,
		_w11910_
	);
	LUT4 #(
		.INIT('h0100)
	) name7863 (
		_w11906_,
		_w11907_,
		_w11908_,
		_w11909_,
		_w11911_
	);
	LUT3 #(
		.INIT('h80)
	) name7864 (
		_w11902_,
		_w11905_,
		_w11911_,
		_w11912_
	);
	LUT4 #(
		.INIT('h8000)
	) name7865 (
		_w11837_,
		_w11879_,
		_w11899_,
		_w11912_,
		_w11913_
	);
	LUT4 #(
		.INIT('h7020)
	) name7866 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11628_,
		_w11830_,
		_w11913_,
		_w11914_
	);
	LUT4 #(
		.INIT('h5545)
	) name7867 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w11915_
	);
	LUT2 #(
		.INIT('h1)
	) name7868 (
		_w11914_,
		_w11915_,
		_w11916_
	);
	LUT3 #(
		.INIT('h0d)
	) name7869 (
		_w4090_,
		_w4091_,
		_w4967_,
		_w11917_
	);
	LUT4 #(
		.INIT('h0008)
	) name7870 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w11918_
	);
	LUT4 #(
		.INIT('hffe7)
	) name7871 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w11919_
	);
	LUT3 #(
		.INIT('hb0)
	) name7872 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w9931_,
		_w11919_,
		_w11920_
	);
	LUT2 #(
		.INIT('h8)
	) name7873 (
		_w11917_,
		_w11920_,
		_w11921_
	);
	LUT2 #(
		.INIT('h1)
	) name7874 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w11922_
	);
	LUT4 #(
		.INIT('h0001)
	) name7875 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\core_c_dec_IR_reg[14]/NET0131 ,
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w11923_
	);
	LUT2 #(
		.INIT('h1)
	) name7876 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w11923_,
		_w11924_
	);
	LUT3 #(
		.INIT('h70)
	) name7877 (
		_w11917_,
		_w11920_,
		_w11924_,
		_w11925_
	);
	LUT4 #(
		.INIT('hbf00)
	) name7878 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w11925_,
		_w11926_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name7879 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w11927_
	);
	LUT4 #(
		.INIT('h0004)
	) name7880 (
		_w4094_,
		_w4097_,
		_w4101_,
		_w11927_,
		_w11928_
	);
	LUT4 #(
		.INIT('hf888)
	) name7881 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w4106_,
		_w11926_,
		_w11928_,
		_w11929_
	);
	LUT4 #(
		.INIT('heee2)
	) name7882 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001 ,
		_w9454_,
		_w11812_,
		_w11813_,
		_w11930_
	);
	LUT4 #(
		.INIT('h8000)
	) name7883 (
		\sice_ICYC_reg[0]/NET0131 ,
		\sice_ICYC_reg[1]/NET0131 ,
		\sice_ICYC_reg[2]/NET0131 ,
		\sice_ICYC_reg[3]/NET0131 ,
		_w11931_
	);
	LUT4 #(
		.INIT('h8000)
	) name7884 (
		\sice_ICYC_reg[4]/NET0131 ,
		\sice_ICYC_reg[5]/NET0131 ,
		\sice_ICYC_reg[6]/NET0131 ,
		_w11931_,
		_w11932_
	);
	LUT2 #(
		.INIT('h6)
	) name7885 (
		\sice_ICYC_reg[7]/NET0131 ,
		_w11932_,
		_w11933_
	);
	LUT4 #(
		.INIT('h8000)
	) name7886 (
		\sice_IIRC_reg[0]/NET0131 ,
		\sice_IIRC_reg[1]/NET0131 ,
		\sice_IIRC_reg[2]/NET0131 ,
		\sice_IIRC_reg[3]/NET0131 ,
		_w11934_
	);
	LUT2 #(
		.INIT('h8)
	) name7887 (
		\sice_IIRC_reg[4]/NET0131 ,
		_w11934_,
		_w11935_
	);
	LUT4 #(
		.INIT('h8000)
	) name7888 (
		\sice_IIRC_reg[4]/NET0131 ,
		\sice_IIRC_reg[5]/NET0131 ,
		\sice_IIRC_reg[6]/NET0131 ,
		_w11934_,
		_w11936_
	);
	LUT2 #(
		.INIT('h6)
	) name7889 (
		\sice_IIRC_reg[7]/NET0131 ,
		_w11936_,
		_w11937_
	);
	LUT3 #(
		.INIT('ha8)
	) name7890 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w11938_
	);
	LUT3 #(
		.INIT('he2)
	) name7891 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001 ,
		_w11926_,
		_w11938_,
		_w11939_
	);
	LUT3 #(
		.INIT('ha8)
	) name7892 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w11940_
	);
	LUT3 #(
		.INIT('he2)
	) name7893 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		_w11926_,
		_w11940_,
		_w11941_
	);
	LUT4 #(
		.INIT('h4c08)
	) name7894 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11329_,
		_w11628_,
		_w11913_,
		_w11942_
	);
	LUT2 #(
		.INIT('h1)
	) name7895 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001 ,
		_w11329_,
		_w11943_
	);
	LUT2 #(
		.INIT('h1)
	) name7896 (
		_w11942_,
		_w11943_,
		_w11944_
	);
	LUT2 #(
		.INIT('h1)
	) name7897 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		\core_c_dec_updSR_E_reg/P0001 ,
		_w11945_
	);
	LUT3 #(
		.INIT('h04)
	) name7898 (
		_w9453_,
		_w9894_,
		_w11945_,
		_w11946_
	);
	LUT3 #(
		.INIT('ha8)
	) name7899 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w11626_,
		_w11627_,
		_w11947_
	);
	LUT2 #(
		.INIT('h4)
	) name7900 (
		_w11592_,
		_w11861_,
		_w11948_
	);
	LUT3 #(
		.INIT('he0)
	) name7901 (
		_w11393_,
		_w11589_,
		_w11852_,
		_w11949_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name7902 (
		_w11333_,
		_w11385_,
		_w11448_,
		_w11468_,
		_w11950_
	);
	LUT3 #(
		.INIT('h0e)
	) name7903 (
		_w11552_,
		_w11474_,
		_w11950_,
		_w11951_
	);
	LUT3 #(
		.INIT('h01)
	) name7904 (
		_w11949_,
		_w11951_,
		_w11948_,
		_w11952_
	);
	LUT4 #(
		.INIT('h00bf)
	) name7905 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11382_,
		_w11429_,
		_w11953_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name7906 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11434_,
		_w11445_,
		_w11954_
	);
	LUT4 #(
		.INIT('hfa32)
	) name7907 (
		_w11844_,
		_w11855_,
		_w11953_,
		_w11954_,
		_w11955_
	);
	LUT3 #(
		.INIT('he0)
	) name7908 (
		_w11393_,
		_w11589_,
		_w11873_,
		_w11956_
	);
	LUT4 #(
		.INIT('h37bf)
	) name7909 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11405_,
		_w11439_,
		_w11957_
	);
	LUT4 #(
		.INIT('hfd75)
	) name7910 (
		_w11333_,
		_w11385_,
		_w11514_,
		_w11464_,
		_w11958_
	);
	LUT2 #(
		.INIT('h1)
	) name7911 (
		_w11957_,
		_w11958_,
		_w11959_
	);
	LUT3 #(
		.INIT('h10)
	) name7912 (
		_w11956_,
		_w11959_,
		_w11955_,
		_w11960_
	);
	LUT3 #(
		.INIT('hc8)
	) name7913 (
		_w11397_,
		_w11532_,
		_w11519_,
		_w11961_
	);
	LUT2 #(
		.INIT('h2)
	) name7914 (
		_w11386_,
		_w11494_,
		_w11962_
	);
	LUT4 #(
		.INIT('ha820)
	) name7915 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001 ,
		_w11963_
	);
	LUT4 #(
		.INIT('h0045)
	) name7916 (
		_w11570_,
		_w11592_,
		_w11962_,
		_w11963_,
		_w11964_
	);
	LUT2 #(
		.INIT('h4)
	) name7917 (
		_w11961_,
		_w11964_,
		_w11965_
	);
	LUT3 #(
		.INIT('h80)
	) name7918 (
		_w11952_,
		_w11960_,
		_w11965_,
		_w11966_
	);
	LUT4 #(
		.INIT('h8000)
	) name7919 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11395_,
		_w11406_,
		_w11967_
	);
	LUT2 #(
		.INIT('h1)
	) name7920 (
		_w11438_,
		_w11885_,
		_w11968_
	);
	LUT4 #(
		.INIT('h0001)
	) name7921 (
		_w11403_,
		_w11438_,
		_w11885_,
		_w11967_,
		_w11969_
	);
	LUT3 #(
		.INIT('h40)
	) name7922 (
		_w11908_,
		_w11909_,
		_w11969_,
		_w11970_
	);
	LUT2 #(
		.INIT('h2)
	) name7923 (
		_w11402_,
		_w11593_,
		_w11971_
	);
	LUT4 #(
		.INIT('h0004)
	) name7924 (
		_w11426_,
		_w11568_,
		_w11832_,
		_w11971_,
		_w11972_
	);
	LUT4 #(
		.INIT('h1000)
	) name7925 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11395_,
		_w11973_
	);
	LUT2 #(
		.INIT('h4)
	) name7926 (
		_w11386_,
		_w11578_,
		_w11974_
	);
	LUT3 #(
		.INIT('ha8)
	) name7927 (
		_w11863_,
		_w11973_,
		_w11974_,
		_w11975_
	);
	LUT4 #(
		.INIT('h2000)
	) name7928 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11418_,
		_w11976_
	);
	LUT3 #(
		.INIT('hc8)
	) name7929 (
		_w11547_,
		_w11499_,
		_w11976_,
		_w11977_
	);
	LUT3 #(
		.INIT('h04)
	) name7930 (
		_w11536_,
		_w11386_,
		_w11954_,
		_w11978_
	);
	LUT3 #(
		.INIT('he0)
	) name7931 (
		_w11420_,
		_w11421_,
		_w11458_,
		_w11979_
	);
	LUT4 #(
		.INIT('h0001)
	) name7932 (
		_w11975_,
		_w11977_,
		_w11978_,
		_w11979_,
		_w11980_
	);
	LUT3 #(
		.INIT('h80)
	) name7933 (
		_w11972_,
		_w11970_,
		_w11980_,
		_w11981_
	);
	LUT4 #(
		.INIT('h2333)
	) name7934 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w11947_,
		_w11966_,
		_w11981_,
		_w11982_
	);
	LUT3 #(
		.INIT('he2)
	) name7935 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001 ,
		_w11946_,
		_w11982_,
		_w11983_
	);
	LUT4 #(
		.INIT('h4000)
	) name7936 (
		\memc_MMR_web_reg/NET0131 ,
		_w5672_,
		_w9431_,
		_w11604_,
		_w11984_
	);
	LUT2 #(
		.INIT('h2)
	) name7937 (
		\sport1_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w11984_,
		_w11985_
	);
	LUT3 #(
		.INIT('he0)
	) name7938 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w11986_
	);
	LUT4 #(
		.INIT('h4500)
	) name7939 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w11986_,
		_w11987_
	);
	LUT2 #(
		.INIT('he)
	) name7940 (
		_w11985_,
		_w11987_,
		_w11988_
	);
	LUT2 #(
		.INIT('h2)
	) name7941 (
		\sport1_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w11984_,
		_w11989_
	);
	LUT4 #(
		.INIT('h4500)
	) name7942 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w11986_,
		_w11990_
	);
	LUT2 #(
		.INIT('he)
	) name7943 (
		_w11989_,
		_w11990_,
		_w11991_
	);
	LUT2 #(
		.INIT('h2)
	) name7944 (
		\sport1_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w11984_,
		_w11992_
	);
	LUT4 #(
		.INIT('h4500)
	) name7945 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w11986_,
		_w11993_
	);
	LUT2 #(
		.INIT('he)
	) name7946 (
		_w11992_,
		_w11993_,
		_w11994_
	);
	LUT3 #(
		.INIT('hca)
	) name7947 (
		\sport1_regs_MWORDreg_DO_reg[8]/NET0131 ,
		_w5760_,
		_w11984_,
		_w11995_
	);
	LUT2 #(
		.INIT('h2)
	) name7948 (
		\sport1_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w11984_,
		_w11996_
	);
	LUT4 #(
		.INIT('h4500)
	) name7949 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w11986_,
		_w11997_
	);
	LUT2 #(
		.INIT('he)
	) name7950 (
		_w11996_,
		_w11997_,
		_w11998_
	);
	LUT2 #(
		.INIT('h2)
	) name7951 (
		\sport1_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w11984_,
		_w11999_
	);
	LUT4 #(
		.INIT('h4500)
	) name7952 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w11986_,
		_w12000_
	);
	LUT2 #(
		.INIT('he)
	) name7953 (
		_w11999_,
		_w12000_,
		_w12001_
	);
	LUT2 #(
		.INIT('h2)
	) name7954 (
		\sport1_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w11984_,
		_w12002_
	);
	LUT4 #(
		.INIT('h4500)
	) name7955 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w11986_,
		_w12003_
	);
	LUT2 #(
		.INIT('he)
	) name7956 (
		_w12002_,
		_w12003_,
		_w12004_
	);
	LUT3 #(
		.INIT('hca)
	) name7957 (
		\sport0_regs_MWORDreg_DO_reg[8]/NET0131 ,
		_w5760_,
		_w11609_,
		_w12005_
	);
	LUT4 #(
		.INIT('h4544)
	) name7958 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6774_,
		_w6894_,
		_w6896_,
		_w12006_
	);
	LUT2 #(
		.INIT('h2)
	) name7959 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8841_,
		_w12007_
	);
	LUT2 #(
		.INIT('h1)
	) name7960 (
		_w12006_,
		_w12007_,
		_w12008_
	);
	LUT3 #(
		.INIT('ha8)
	) name7961 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12006_,
		_w12007_,
		_w12009_
	);
	LUT3 #(
		.INIT('hc8)
	) name7962 (
		_w11572_,
		_w11854_,
		_w11831_,
		_w12010_
	);
	LUT3 #(
		.INIT('h0e)
	) name7963 (
		_w11420_,
		_w11421_,
		_w11452_,
		_w12011_
	);
	LUT3 #(
		.INIT('h02)
	) name7964 (
		_w11386_,
		_w11540_,
		_w11593_,
		_w12012_
	);
	LUT3 #(
		.INIT('hc8)
	) name7965 (
		_w11547_,
		_w11449_,
		_w11976_,
		_w12013_
	);
	LUT4 #(
		.INIT('h0001)
	) name7966 (
		_w12010_,
		_w12011_,
		_w12012_,
		_w12013_,
		_w12014_
	);
	LUT4 #(
		.INIT('ha820)
	) name7967 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001 ,
		_w12015_
	);
	LUT4 #(
		.INIT('h0001)
	) name7968 (
		_w11403_,
		_w11438_,
		_w11967_,
		_w12015_,
		_w12016_
	);
	LUT4 #(
		.INIT('hddd0)
	) name7969 (
		_w11538_,
		_w11593_,
		_w11512_,
		_w11957_,
		_w12017_
	);
	LUT4 #(
		.INIT('h1000)
	) name7970 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11392_,
		_w12018_
	);
	LUT3 #(
		.INIT('hc8)
	) name7971 (
		_w11557_,
		_w11532_,
		_w12018_,
		_w12019_
	);
	LUT4 #(
		.INIT('h2000)
	) name7972 (
		_w11571_,
		_w12019_,
		_w12016_,
		_w12017_,
		_w12020_
	);
	LUT4 #(
		.INIT('h0f08)
	) name7973 (
		_w11333_,
		_w11397_,
		_w11498_,
		_w11519_,
		_w12021_
	);
	LUT2 #(
		.INIT('h1)
	) name7974 (
		_w11592_,
		_w11471_,
		_w12022_
	);
	LUT3 #(
		.INIT('h32)
	) name7975 (
		_w11552_,
		_w11489_,
		_w11474_,
		_w12023_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name7976 (
		_w11333_,
		_w11385_,
		_w11514_,
		_w11457_,
		_w12024_
	);
	LUT4 #(
		.INIT('h7770)
	) name7977 (
		_w11424_,
		_w11495_,
		_w11954_,
		_w12024_,
		_w12025_
	);
	LUT4 #(
		.INIT('h0100)
	) name7978 (
		_w12022_,
		_w12021_,
		_w12023_,
		_w12025_,
		_w12026_
	);
	LUT3 #(
		.INIT('h80)
	) name7979 (
		_w12014_,
		_w12020_,
		_w12026_,
		_w12027_
	);
	LUT4 #(
		.INIT('h4000)
	) name7980 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12014_,
		_w12020_,
		_w12026_,
		_w12028_
	);
	LUT4 #(
		.INIT('h222e)
	) name7981 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001 ,
		_w11946_,
		_w12009_,
		_w12028_,
		_w12029_
	);
	LUT2 #(
		.INIT('h2)
	) name7982 (
		\sport0_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w11609_,
		_w12030_
	);
	LUT3 #(
		.INIT('he0)
	) name7983 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w12031_
	);
	LUT4 #(
		.INIT('h4500)
	) name7984 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w12031_,
		_w12032_
	);
	LUT2 #(
		.INIT('he)
	) name7985 (
		_w12030_,
		_w12032_,
		_w12033_
	);
	LUT2 #(
		.INIT('h2)
	) name7986 (
		\sport0_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w11609_,
		_w12034_
	);
	LUT4 #(
		.INIT('h4500)
	) name7987 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w12031_,
		_w12035_
	);
	LUT2 #(
		.INIT('he)
	) name7988 (
		_w12034_,
		_w12035_,
		_w12036_
	);
	LUT2 #(
		.INIT('h2)
	) name7989 (
		\sport0_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w11609_,
		_w12037_
	);
	LUT4 #(
		.INIT('h4500)
	) name7990 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w12031_,
		_w12038_
	);
	LUT2 #(
		.INIT('he)
	) name7991 (
		_w12037_,
		_w12038_,
		_w12039_
	);
	LUT4 #(
		.INIT('h0045)
	) name7992 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w11613_,
		_w12040_
	);
	LUT3 #(
		.INIT('he2)
	) name7993 (
		\sport0_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w11609_,
		_w12040_,
		_w12041_
	);
	LUT2 #(
		.INIT('h2)
	) name7994 (
		\sport0_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w11609_,
		_w12042_
	);
	LUT4 #(
		.INIT('h4500)
	) name7995 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w12031_,
		_w12043_
	);
	LUT2 #(
		.INIT('he)
	) name7996 (
		_w12042_,
		_w12043_,
		_w12044_
	);
	LUT2 #(
		.INIT('h2)
	) name7997 (
		\sport0_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w11609_,
		_w12045_
	);
	LUT4 #(
		.INIT('h4500)
	) name7998 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w12031_,
		_w12046_
	);
	LUT2 #(
		.INIT('he)
	) name7999 (
		_w12045_,
		_w12046_,
		_w12047_
	);
	LUT4 #(
		.INIT('h0004)
	) name8000 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9452_,
		_w9453_,
		_w11945_,
		_w12048_
	);
	LUT3 #(
		.INIT('hca)
	) name8001 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001 ,
		_w11982_,
		_w12048_,
		_w12049_
	);
	LUT4 #(
		.INIT('h00df)
	) name8002 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\memc_Dread_E_reg/NET0131 ,
		\memc_IOcmd_E_reg/NET0131 ,
		_w12050_
	);
	LUT3 #(
		.INIT('he0)
	) name8003 (
		PM_bdry_sel_pad,
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		_w12051_
	);
	LUT2 #(
		.INIT('h8)
	) name8004 (
		\core_c_dec_Double_E_reg/P0001 ,
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w12052_
	);
	LUT2 #(
		.INIT('h8)
	) name8005 (
		_w12051_,
		_w12052_,
		_w12053_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name8006 (
		_w4069_,
		_w4077_,
		_w4862_,
		_w4868_,
		_w12054_
	);
	LUT4 #(
		.INIT('hf4f5)
	) name8007 (
		_w4069_,
		_w4077_,
		_w4862_,
		_w4868_,
		_w12055_
	);
	LUT2 #(
		.INIT('h1)
	) name8008 (
		\core_c_psq_ECYC_reg/P0001 ,
		_w9936_,
		_w12056_
	);
	LUT4 #(
		.INIT('h2700)
	) name8009 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4069_,
		_w12054_,
		_w12056_,
		_w12057_
	);
	LUT2 #(
		.INIT('h4)
	) name8010 (
		_w12053_,
		_w12057_,
		_w12058_
	);
	LUT3 #(
		.INIT('h40)
	) name8011 (
		_w9936_,
		_w12051_,
		_w12052_,
		_w12059_
	);
	LUT4 #(
		.INIT('h4000)
	) name8012 (
		_w4747_,
		_w4768_,
		_w4798_,
		_w12059_,
		_w12060_
	);
	LUT4 #(
		.INIT('h00bf)
	) name8013 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w9936_,
		_w12061_
	);
	LUT2 #(
		.INIT('h2)
	) name8014 (
		\emc_DMDoe_reg/NET0131 ,
		_w12061_,
		_w12062_
	);
	LUT4 #(
		.INIT('h5754)
	) name8015 (
		_w12050_,
		_w12058_,
		_w12060_,
		_w12062_,
		_w12063_
	);
	LUT4 #(
		.INIT('h03aa)
	) name8016 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001 ,
		_w12009_,
		_w12028_,
		_w12048_,
		_w12064_
	);
	LUT4 #(
		.INIT('h03aa)
	) name8017 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w8757_,
		_w8760_,
		_w11984_,
		_w12065_
	);
	LUT4 #(
		.INIT('h03aa)
	) name8018 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w8757_,
		_w8760_,
		_w11609_,
		_w12066_
	);
	LUT4 #(
		.INIT('haf23)
	) name8019 (
		\sport1_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w12067_
	);
	LUT4 #(
		.INIT('haf23)
	) name8020 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w12068_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8021 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w12069_
	);
	LUT2 #(
		.INIT('h9)
	) name8022 (
		\sport1_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w12070_
	);
	LUT4 #(
		.INIT('h8000)
	) name8023 (
		_w12069_,
		_w12070_,
		_w12067_,
		_w12068_,
		_w12071_
	);
	LUT4 #(
		.INIT('h8421)
	) name8024 (
		\sport1_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w12072_
	);
	LUT4 #(
		.INIT('haf23)
	) name8025 (
		\sport1_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w12073_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8026 (
		\sport1_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w12074_
	);
	LUT3 #(
		.INIT('h80)
	) name8027 (
		_w12073_,
		_w12074_,
		_w12072_,
		_w12075_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8028 (
		\sport1_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w12076_
	);
	LUT4 #(
		.INIT('hf531)
	) name8029 (
		\sport1_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w12077_
	);
	LUT2 #(
		.INIT('h6)
	) name8030 (
		\sport1_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w12078_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8031 (
		\sport1_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w12079_
	);
	LUT4 #(
		.INIT('h4000)
	) name8032 (
		_w12078_,
		_w12079_,
		_w12076_,
		_w12077_,
		_w12080_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8033 (
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w12081_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8034 (
		\sport1_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w12082_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8035 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w12083_
	);
	LUT4 #(
		.INIT('haf23)
	) name8036 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w12084_
	);
	LUT4 #(
		.INIT('h8000)
	) name8037 (
		_w12083_,
		_w12084_,
		_w12081_,
		_w12082_,
		_w12085_
	);
	LUT4 #(
		.INIT('h8000)
	) name8038 (
		_w12080_,
		_w12085_,
		_w12071_,
		_w12075_,
		_w12086_
	);
	LUT2 #(
		.INIT('h2)
	) name8039 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12087_
	);
	LUT3 #(
		.INIT('h59)
	) name8040 (
		\sport1_cfg_SCLKi_h_reg/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12088_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8041 (
		\sport0_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w12089_
	);
	LUT4 #(
		.INIT('haf23)
	) name8042 (
		\sport0_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w12090_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8043 (
		\sport0_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w12091_
	);
	LUT2 #(
		.INIT('h9)
	) name8044 (
		\sport0_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w12092_
	);
	LUT4 #(
		.INIT('h8000)
	) name8045 (
		_w12091_,
		_w12092_,
		_w12089_,
		_w12090_,
		_w12093_
	);
	LUT4 #(
		.INIT('h8421)
	) name8046 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w12094_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8047 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w12095_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8048 (
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w12096_
	);
	LUT3 #(
		.INIT('h80)
	) name8049 (
		_w12095_,
		_w12096_,
		_w12094_,
		_w12097_
	);
	LUT4 #(
		.INIT('haf23)
	) name8050 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w12098_
	);
	LUT4 #(
		.INIT('hf531)
	) name8051 (
		\sport0_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w12099_
	);
	LUT2 #(
		.INIT('h6)
	) name8052 (
		\sport0_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w12100_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8053 (
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w12101_
	);
	LUT4 #(
		.INIT('h4000)
	) name8054 (
		_w12100_,
		_w12101_,
		_w12098_,
		_w12099_,
		_w12102_
	);
	LUT4 #(
		.INIT('haf23)
	) name8055 (
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w12103_
	);
	LUT4 #(
		.INIT('haf23)
	) name8056 (
		\sport0_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w12104_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8057 (
		\sport0_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w12105_
	);
	LUT4 #(
		.INIT('haf23)
	) name8058 (
		\sport0_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w12106_
	);
	LUT4 #(
		.INIT('h8000)
	) name8059 (
		_w12105_,
		_w12106_,
		_w12103_,
		_w12104_,
		_w12107_
	);
	LUT4 #(
		.INIT('h8000)
	) name8060 (
		_w12102_,
		_w12107_,
		_w12093_,
		_w12097_,
		_w12108_
	);
	LUT2 #(
		.INIT('h2)
	) name8061 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12109_
	);
	LUT3 #(
		.INIT('h59)
	) name8062 (
		\sport0_cfg_SCLKi_h_reg/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12110_
	);
	LUT4 #(
		.INIT('h4044)
	) name8063 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w12111_
	);
	LUT3 #(
		.INIT('h07)
	) name8064 (
		_w9910_,
		_w11802_,
		_w12111_,
		_w12112_
	);
	LUT4 #(
		.INIT('h0002)
	) name8065 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w4971_,
		_w9453_,
		_w12113_
	);
	LUT4 #(
		.INIT('h0007)
	) name8066 (
		_w9910_,
		_w11802_,
		_w12111_,
		_w12113_,
		_w12114_
	);
	LUT3 #(
		.INIT('h02)
	) name8067 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9453_,
		_w12115_
	);
	LUT4 #(
		.INIT('h0f04)
	) name8068 (
		_w9792_,
		_w9805_,
		_w9823_,
		_w9825_,
		_w12116_
	);
	LUT2 #(
		.INIT('h2)
	) name8069 (
		_w9794_,
		_w9803_,
		_w12117_
	);
	LUT4 #(
		.INIT('h0410)
	) name8070 (
		_w9456_,
		_w9794_,
		_w9803_,
		_w12116_,
		_w12118_
	);
	LUT4 #(
		.INIT('h50c5)
	) name8071 (
		_w9759_,
		_w9757_,
		_w9794_,
		_w9803_,
		_w12119_
	);
	LUT3 #(
		.INIT('h1e)
	) name8072 (
		_w9456_,
		_w12116_,
		_w12119_,
		_w12120_
	);
	LUT4 #(
		.INIT('h804c)
	) name8073 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12115_,
		_w12118_,
		_w12120_,
		_w12121_
	);
	LUT4 #(
		.INIT('h2022)
	) name8074 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w6774_,
		_w6894_,
		_w6896_,
		_w12122_
	);
	LUT4 #(
		.INIT('h4000)
	) name8075 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001 ,
		_w12123_
	);
	LUT4 #(
		.INIT('h0200)
	) name8076 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001 ,
		_w12124_
	);
	LUT4 #(
		.INIT('h2000)
	) name8077 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001 ,
		_w12125_
	);
	LUT3 #(
		.INIT('h01)
	) name8078 (
		_w12124_,
		_w12125_,
		_w12123_,
		_w12126_
	);
	LUT4 #(
		.INIT('h0400)
	) name8079 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001 ,
		_w12127_
	);
	LUT4 #(
		.INIT('h0100)
	) name8080 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001 ,
		_w12128_
	);
	LUT4 #(
		.INIT('h0800)
	) name8081 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001 ,
		_w12129_
	);
	LUT4 #(
		.INIT('h1000)
	) name8082 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001 ,
		_w12130_
	);
	LUT4 #(
		.INIT('h0001)
	) name8083 (
		_w12127_,
		_w12128_,
		_w12129_,
		_w12130_,
		_w12131_
	);
	LUT2 #(
		.INIT('h8)
	) name8084 (
		_w12126_,
		_w12131_,
		_w12132_
	);
	LUT2 #(
		.INIT('h2)
	) name8085 (
		_w9911_,
		_w12132_,
		_w12133_
	);
	LUT2 #(
		.INIT('h1)
	) name8086 (
		_w12122_,
		_w12133_,
		_w12134_
	);
	LUT2 #(
		.INIT('h8)
	) name8087 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w12135_
	);
	LUT4 #(
		.INIT('h2022)
	) name8088 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w6378_,
		_w6498_,
		_w6500_,
		_w12136_
	);
	LUT4 #(
		.INIT('h4000)
	) name8089 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001 ,
		_w12137_
	);
	LUT4 #(
		.INIT('h0200)
	) name8090 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001 ,
		_w12138_
	);
	LUT4 #(
		.INIT('h2000)
	) name8091 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001 ,
		_w12139_
	);
	LUT3 #(
		.INIT('h01)
	) name8092 (
		_w12138_,
		_w12139_,
		_w12137_,
		_w12140_
	);
	LUT4 #(
		.INIT('h0400)
	) name8093 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001 ,
		_w12141_
	);
	LUT4 #(
		.INIT('h0100)
	) name8094 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001 ,
		_w12142_
	);
	LUT4 #(
		.INIT('h0800)
	) name8095 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001 ,
		_w12143_
	);
	LUT4 #(
		.INIT('h1000)
	) name8096 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001 ,
		_w12144_
	);
	LUT4 #(
		.INIT('h0001)
	) name8097 (
		_w12141_,
		_w12142_,
		_w12143_,
		_w12144_,
		_w12145_
	);
	LUT2 #(
		.INIT('h8)
	) name8098 (
		_w12140_,
		_w12145_,
		_w12146_
	);
	LUT2 #(
		.INIT('h2)
	) name8099 (
		_w9911_,
		_w12146_,
		_w12147_
	);
	LUT2 #(
		.INIT('h1)
	) name8100 (
		_w12136_,
		_w12147_,
		_w12148_
	);
	LUT4 #(
		.INIT('h5700)
	) name8101 (
		_w12115_,
		_w12118_,
		_w12135_,
		_w12148_,
		_w12149_
	);
	LUT2 #(
		.INIT('h1)
	) name8102 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w12150_
	);
	LUT4 #(
		.INIT('h0010)
	) name8103 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12151_
	);
	LUT4 #(
		.INIT('hb400)
	) name8104 (
		_w12121_,
		_w12134_,
		_w12149_,
		_w12151_,
		_w12152_
	);
	LUT2 #(
		.INIT('h2)
	) name8105 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w12153_
	);
	LUT4 #(
		.INIT('h0020)
	) name8106 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12154_
	);
	LUT4 #(
		.INIT('h4b00)
	) name8107 (
		_w12121_,
		_w12134_,
		_w12149_,
		_w12154_,
		_w12155_
	);
	LUT2 #(
		.INIT('h8)
	) name8108 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w12156_
	);
	LUT4 #(
		.INIT('h0080)
	) name8109 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12157_
	);
	LUT2 #(
		.INIT('h4)
	) name8110 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w12158_
	);
	LUT4 #(
		.INIT('h0040)
	) name8111 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12159_
	);
	LUT4 #(
		.INIT('h0200)
	) name8112 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12160_
	);
	LUT4 #(
		.INIT('h0023)
	) name8113 (
		_w9792_,
		_w9804_,
		_w9805_,
		_w9825_,
		_w12161_
	);
	LUT3 #(
		.INIT('h0b)
	) name8114 (
		_w9790_,
		_w9823_,
		_w12117_,
		_w12162_
	);
	LUT3 #(
		.INIT('h45)
	) name8115 (
		_w9456_,
		_w12161_,
		_w12162_,
		_w12163_
	);
	LUT4 #(
		.INIT('h4044)
	) name8116 (
		_w9456_,
		_w12115_,
		_w12161_,
		_w12162_,
		_w12164_
	);
	LUT4 #(
		.INIT('h0400)
	) name8117 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001 ,
		_w12165_
	);
	LUT4 #(
		.INIT('h0200)
	) name8118 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001 ,
		_w12166_
	);
	LUT4 #(
		.INIT('h4000)
	) name8119 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001 ,
		_w12167_
	);
	LUT3 #(
		.INIT('h01)
	) name8120 (
		_w12166_,
		_w12167_,
		_w12165_,
		_w12168_
	);
	LUT4 #(
		.INIT('h2000)
	) name8121 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001 ,
		_w12169_
	);
	LUT4 #(
		.INIT('h0100)
	) name8122 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001 ,
		_w12170_
	);
	LUT4 #(
		.INIT('h0800)
	) name8123 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001 ,
		_w12171_
	);
	LUT4 #(
		.INIT('h1000)
	) name8124 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001 ,
		_w12172_
	);
	LUT4 #(
		.INIT('h0001)
	) name8125 (
		_w12169_,
		_w12170_,
		_w12171_,
		_w12172_,
		_w12173_
	);
	LUT2 #(
		.INIT('h8)
	) name8126 (
		_w12168_,
		_w12173_,
		_w12174_
	);
	LUT2 #(
		.INIT('h2)
	) name8127 (
		_w9911_,
		_w12174_,
		_w12175_
	);
	LUT4 #(
		.INIT('h2022)
	) name8128 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w6054_,
		_w6173_,
		_w6175_,
		_w12176_
	);
	LUT2 #(
		.INIT('h1)
	) name8129 (
		_w12175_,
		_w12176_,
		_w12177_
	);
	LUT4 #(
		.INIT('h0100)
	) name8130 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12178_
	);
	LUT4 #(
		.INIT('h10df)
	) name8131 (
		_w12160_,
		_w12164_,
		_w12177_,
		_w12178_,
		_w12179_
	);
	LUT4 #(
		.INIT('h1b00)
	) name8132 (
		_w12149_,
		_w12159_,
		_w12157_,
		_w12179_,
		_w12180_
	);
	LUT4 #(
		.INIT('h5455)
	) name8133 (
		_w12114_,
		_w12155_,
		_w12152_,
		_w12180_,
		_w12181_
	);
	LUT4 #(
		.INIT('h0020)
	) name8134 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[4]/NET0131 ,
		_w9453_,
		_w12182_
	);
	LUT3 #(
		.INIT('hb0)
	) name8135 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9458_,
		_w12183_
	);
	LUT2 #(
		.INIT('h8)
	) name8136 (
		_w12182_,
		_w12183_,
		_w12184_
	);
	LUT2 #(
		.INIT('h2)
	) name8137 (
		_w12112_,
		_w12184_,
		_w12185_
	);
	LUT3 #(
		.INIT('h48)
	) name8138 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w12186_
	);
	LUT3 #(
		.INIT('h20)
	) name8139 (
		_w12112_,
		_w12184_,
		_w12186_,
		_w12187_
	);
	LUT4 #(
		.INIT('h0200)
	) name8140 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001 ,
		_w12188_
	);
	LUT4 #(
		.INIT('h0400)
	) name8141 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001 ,
		_w12189_
	);
	LUT4 #(
		.INIT('h0800)
	) name8142 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001 ,
		_w12190_
	);
	LUT3 #(
		.INIT('h01)
	) name8143 (
		_w12189_,
		_w12190_,
		_w12188_,
		_w12191_
	);
	LUT4 #(
		.INIT('h2000)
	) name8144 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001 ,
		_w12192_
	);
	LUT4 #(
		.INIT('h0100)
	) name8145 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001 ,
		_w12193_
	);
	LUT4 #(
		.INIT('h4000)
	) name8146 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001 ,
		_w12194_
	);
	LUT4 #(
		.INIT('h1000)
	) name8147 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001 ,
		_w12195_
	);
	LUT4 #(
		.INIT('h0001)
	) name8148 (
		_w12192_,
		_w12193_,
		_w12194_,
		_w12195_,
		_w12196_
	);
	LUT2 #(
		.INIT('h8)
	) name8149 (
		_w12191_,
		_w12196_,
		_w12197_
	);
	LUT2 #(
		.INIT('h2)
	) name8150 (
		_w9911_,
		_w12197_,
		_w12198_
	);
	LUT2 #(
		.INIT('h8)
	) name8151 (
		_w9474_,
		_w12182_,
		_w12199_
	);
	LUT4 #(
		.INIT('h2022)
	) name8152 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w7257_,
		_w7375_,
		_w7377_,
		_w12200_
	);
	LUT4 #(
		.INIT('h0001)
	) name8153 (
		_w12156_,
		_w12199_,
		_w12200_,
		_w12198_,
		_w12201_
	);
	LUT4 #(
		.INIT('h5554)
	) name8154 (
		_w12158_,
		_w12199_,
		_w12200_,
		_w12198_,
		_w12202_
	);
	LUT4 #(
		.INIT('h3332)
	) name8155 (
		_w12185_,
		_w12187_,
		_w12202_,
		_w12201_,
		_w12203_
	);
	LUT4 #(
		.INIT('h45cf)
	) name8156 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w12157_,
		_w12178_,
		_w12204_
	);
	LUT4 #(
		.INIT('h236f)
	) name8157 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w12154_,
		_w12159_,
		_w12205_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name8158 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w4161_,
		_w12151_,
		_w12160_,
		_w12206_
	);
	LUT3 #(
		.INIT('h80)
	) name8159 (
		_w12204_,
		_w12205_,
		_w12206_,
		_w12207_
	);
	LUT4 #(
		.INIT('h8000)
	) name8160 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12208_
	);
	LUT4 #(
		.INIT('h00bf)
	) name8161 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12208_,
		_w12209_
	);
	LUT3 #(
		.INIT('hd0)
	) name8162 (
		_w12114_,
		_w12207_,
		_w12209_,
		_w12210_
	);
	LUT3 #(
		.INIT('hd0)
	) name8163 (
		_w5100_,
		_w12203_,
		_w12210_,
		_w12211_
	);
	LUT4 #(
		.INIT('h1000)
	) name8164 (
		\core_eu_ec_cun_condOK_CE_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12212_
	);
	LUT2 #(
		.INIT('h2)
	) name8165 (
		_w4140_,
		_w12212_,
		_w12213_
	);
	LUT3 #(
		.INIT('hb0)
	) name8166 (
		_w12181_,
		_w12211_,
		_w12213_,
		_w12214_
	);
	LUT4 #(
		.INIT('h9a55)
	) name8167 (
		_w10165_,
		_w11250_,
		_w11285_,
		_w11289_,
		_w12215_
	);
	LUT3 #(
		.INIT('h82)
	) name8168 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10132_,
		_w12215_,
		_w12216_
	);
	LUT2 #(
		.INIT('h9)
	) name8169 (
		_w11274_,
		_w11283_,
		_w12217_
	);
	LUT4 #(
		.INIT('h010f)
	) name8170 (
		_w11250_,
		_w11273_,
		_w11281_,
		_w11286_,
		_w12218_
	);
	LUT4 #(
		.INIT('h0514)
	) name8171 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11287_,
		_w12217_,
		_w12218_,
		_w12219_
	);
	LUT4 #(
		.INIT('h5040)
	) name8172 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w9893_,
		_w11305_,
		_w12220_
	);
	LUT2 #(
		.INIT('h2)
	) name8173 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 ,
		_w12220_,
		_w12221_
	);
	LUT2 #(
		.INIT('h2)
	) name8174 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w12222_
	);
	LUT3 #(
		.INIT('h80)
	) name8175 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 ,
		_w9894_,
		_w11305_,
		_w12223_
	);
	LUT3 #(
		.INIT('h80)
	) name8176 (
		_w9894_,
		_w11318_,
		_w11319_,
		_w12224_
	);
	LUT4 #(
		.INIT('h007f)
	) name8177 (
		_w9894_,
		_w11318_,
		_w11319_,
		_w12223_,
		_w12225_
	);
	LUT4 #(
		.INIT('h4454)
	) name8178 (
		_w11624_,
		_w12221_,
		_w12222_,
		_w12225_,
		_w12226_
	);
	LUT3 #(
		.INIT('hc4)
	) name8179 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 ,
		_w11308_,
		_w12227_
	);
	LUT2 #(
		.INIT('h1)
	) name8180 (
		_w12226_,
		_w12227_,
		_w12228_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name8181 (
		_w11624_,
		_w12216_,
		_w12219_,
		_w12228_,
		_w12229_
	);
	LUT2 #(
		.INIT('h2)
	) name8182 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 ,
		_w11310_,
		_w12230_
	);
	LUT2 #(
		.INIT('h1)
	) name8183 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w12231_
	);
	LUT4 #(
		.INIT('h007f)
	) name8184 (
		_w11300_,
		_w11318_,
		_w11319_,
		_w11324_,
		_w12232_
	);
	LUT4 #(
		.INIT('h4454)
	) name8185 (
		_w9946_,
		_w12230_,
		_w12231_,
		_w12232_,
		_w12233_
	);
	LUT3 #(
		.INIT('hc8)
	) name8186 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 ,
		_w11308_,
		_w12234_
	);
	LUT2 #(
		.INIT('h1)
	) name8187 (
		_w12233_,
		_w12234_,
		_w12235_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name8188 (
		_w9946_,
		_w12216_,
		_w12219_,
		_w12235_,
		_w12236_
	);
	LUT3 #(
		.INIT('h36)
	) name8189 (
		_w10131_,
		_w10133_,
		_w10166_,
		_w12237_
	);
	LUT4 #(
		.INIT('h5401)
	) name8190 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10132_,
		_w11290_,
		_w12237_,
		_w12238_
	);
	LUT4 #(
		.INIT('h007d)
	) name8191 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11293_,
		_w11295_,
		_w12238_,
		_w12239_
	);
	LUT4 #(
		.INIT('hff82)
	) name8192 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11293_,
		_w11295_,
		_w12238_,
		_w12240_
	);
	LUT2 #(
		.INIT('h6)
	) name8193 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		_w12241_
	);
	LUT3 #(
		.INIT('h20)
	) name8194 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12241_,
		_w12242_
	);
	LUT3 #(
		.INIT('h69)
	) name8195 (
		_w11250_,
		_w11268_,
		_w11272_,
		_w12243_
	);
	LUT4 #(
		.INIT('h8228)
	) name8196 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11250_,
		_w11268_,
		_w11272_,
		_w12244_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8197 (
		_w10433_,
		_w10640_,
		_w10645_,
		_w11231_,
		_w12245_
	);
	LUT4 #(
		.INIT('h50d0)
	) name8198 (
		_w11186_,
		_w11243_,
		_w11237_,
		_w12245_,
		_w12246_
	);
	LUT4 #(
		.INIT('h0c04)
	) name8199 (
		_w10923_,
		_w11245_,
		_w11246_,
		_w12246_,
		_w12247_
	);
	LUT4 #(
		.INIT('ha596)
	) name8200 (
		_w10964_,
		_w10970_,
		_w10972_,
		_w12247_,
		_w12248_
	);
	LUT3 #(
		.INIT('hdc)
	) name8201 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12244_,
		_w12248_,
		_w12249_
	);
	LUT2 #(
		.INIT('h6)
	) name8202 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		_w12250_
	);
	LUT3 #(
		.INIT('h20)
	) name8203 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12250_,
		_w12251_
	);
	LUT4 #(
		.INIT('h8000)
	) name8204 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_OUTcnt_reg[1]/NET0131 ,
		\clkc_OUTcnt_reg[2]/NET0131 ,
		\clkc_OUTcnt_reg[3]/NET0131 ,
		_w12252_
	);
	LUT4 #(
		.INIT('h8000)
	) name8205 (
		\clkc_OUTcnt_reg[4]/NET0131 ,
		\clkc_OUTcnt_reg[5]/NET0131 ,
		\clkc_OUTcnt_reg[6]/NET0131 ,
		_w12252_,
		_w12253_
	);
	LUT2 #(
		.INIT('h2)
	) name8206 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_ckr_reg_DO_reg[8]/NET0131 ,
		_w12254_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8207 (
		\clkc_OUTcnt_reg[2]/NET0131 ,
		\clkc_OUTcnt_reg[6]/NET0131 ,
		\clkc_ckr_reg_DO_reg[10]/NET0131 ,
		\clkc_ckr_reg_DO_reg[14]/NET0131 ,
		_w12255_
	);
	LUT4 #(
		.INIT('h8acf)
	) name8208 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_OUTcnt_reg[3]/NET0131 ,
		\clkc_ckr_reg_DO_reg[11]/NET0131 ,
		\clkc_ckr_reg_DO_reg[8]/NET0131 ,
		_w12256_
	);
	LUT4 #(
		.INIT('hf531)
	) name8209 (
		\clkc_OUTcnt_reg[2]/NET0131 ,
		\clkc_OUTcnt_reg[3]/NET0131 ,
		\clkc_ckr_reg_DO_reg[10]/NET0131 ,
		\clkc_ckr_reg_DO_reg[11]/NET0131 ,
		_w12257_
	);
	LUT3 #(
		.INIT('h80)
	) name8210 (
		_w12255_,
		_w12256_,
		_w12257_,
		_w12258_
	);
	LUT2 #(
		.INIT('h2)
	) name8211 (
		\clkc_OUTcnt_reg[6]/NET0131 ,
		\clkc_ckr_reg_DO_reg[14]/NET0131 ,
		_w12259_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name8212 (
		\clkc_OUTcnt_reg[4]/NET0131 ,
		\clkc_OUTcnt_reg[5]/NET0131 ,
		\clkc_ckr_reg_DO_reg[12]/NET0131 ,
		\clkc_ckr_reg_DO_reg[13]/NET0131 ,
		_w12260_
	);
	LUT4 #(
		.INIT('hcf45)
	) name8213 (
		\clkc_OUTcnt_reg[1]/NET0131 ,
		\clkc_OUTcnt_reg[4]/NET0131 ,
		\clkc_ckr_reg_DO_reg[12]/NET0131 ,
		\clkc_ckr_reg_DO_reg[9]/NET0131 ,
		_w12261_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name8214 (
		\clkc_OUTcnt_reg[1]/NET0131 ,
		\clkc_OUTcnt_reg[5]/NET0131 ,
		\clkc_ckr_reg_DO_reg[13]/NET0131 ,
		\clkc_ckr_reg_DO_reg[9]/NET0131 ,
		_w12262_
	);
	LUT4 #(
		.INIT('h4000)
	) name8215 (
		_w12259_,
		_w12261_,
		_w12262_,
		_w12260_,
		_w12263_
	);
	LUT4 #(
		.INIT('h070f)
	) name8216 (
		\clkc_OUTcnt_reg[4]/NET0131 ,
		\clkc_OUTcnt_reg[5]/NET0131 ,
		\clkc_OUTcnt_reg[6]/NET0131 ,
		_w12252_,
		_w12264_
	);
	LUT4 #(
		.INIT('h00bf)
	) name8217 (
		_w12254_,
		_w12258_,
		_w12263_,
		_w12264_,
		_w12265_
	);
	LUT2 #(
		.INIT('h4)
	) name8218 (
		_w12253_,
		_w12265_,
		_w12266_
	);
	LUT3 #(
		.INIT('h2a)
	) name8219 (
		\core_c_psq_INT_en_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12267_
	);
	LUT4 #(
		.INIT('hc444)
	) name8220 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		_w4073_,
		_w4084_,
		_w12268_
	);
	LUT3 #(
		.INIT('h13)
	) name8221 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_Iflag_reg[10]/NET0131 ,
		\core_c_psq_Iflag_reg[8]/NET0131 ,
		_w12269_
	);
	LUT4 #(
		.INIT('h00ec)
	) name8222 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_Iflag_reg[10]/NET0131 ,
		\core_c_psq_Iflag_reg[8]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w12270_
	);
	LUT4 #(
		.INIT('h002a)
	) name8223 (
		\core_c_psq_INT_en_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12270_,
		_w12271_
	);
	LUT3 #(
		.INIT('h08)
	) name8224 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		\core_c_psq_Iflag_reg[9]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w12272_
	);
	LUT3 #(
		.INIT('h08)
	) name8225 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_Iflag_reg[5]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w12273_
	);
	LUT2 #(
		.INIT('h8)
	) name8226 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_Iflag_reg[6]/NET0131 ,
		_w12274_
	);
	LUT3 #(
		.INIT('h08)
	) name8227 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_Iflag_reg[6]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w12275_
	);
	LUT3 #(
		.INIT('h08)
	) name8228 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_Iflag_reg[4]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w12276_
	);
	LUT3 #(
		.INIT('h08)
	) name8229 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		\core_c_psq_Iflag_reg[7]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w12277_
	);
	LUT2 #(
		.INIT('h1)
	) name8230 (
		_w12276_,
		_w12277_,
		_w12278_
	);
	LUT3 #(
		.INIT('h01)
	) name8231 (
		_w12275_,
		_w12276_,
		_w12277_,
		_w12279_
	);
	LUT4 #(
		.INIT('h0002)
	) name8232 (
		_w12273_,
		_w12275_,
		_w12276_,
		_w12277_,
		_w12280_
	);
	LUT4 #(
		.INIT('haeaa)
	) name8233 (
		_w12268_,
		_w12271_,
		_w12272_,
		_w12280_,
		_w12281_
	);
	LUT2 #(
		.INIT('h8)
	) name8234 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w9894_,
		_w12282_
	);
	LUT2 #(
		.INIT('h2)
	) name8235 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w9021_,
		_w12283_
	);
	LUT4 #(
		.INIT('h00ab)
	) name8236 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w7140_,
		_w7240_,
		_w12283_,
		_w12284_
	);
	LUT3 #(
		.INIT('h13)
	) name8237 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 ,
		_w9894_,
		_w12285_
	);
	LUT4 #(
		.INIT('h0002)
	) name8238 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w12285_,
		_w12286_
	);
	LUT4 #(
		.INIT('h313b)
	) name8239 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 ,
		_w11308_,
		_w11635_,
		_w12287_
	);
	LUT4 #(
		.INIT('h2f00)
	) name8240 (
		_w12282_,
		_w12284_,
		_w12286_,
		_w12287_,
		_w12288_
	);
	LUT2 #(
		.INIT('h1)
	) name8241 (
		_w11624_,
		_w12288_,
		_w12289_
	);
	LUT2 #(
		.INIT('h9)
	) name8242 (
		_w10967_,
		_w10969_,
		_w12290_
	);
	LUT4 #(
		.INIT('h3bc4)
	) name8243 (
		_w10923_,
		_w11245_,
		_w12246_,
		_w12290_,
		_w12291_
	);
	LUT2 #(
		.INIT('h6)
	) name8244 (
		_w10814_,
		_w10868_,
		_w12292_
	);
	LUT4 #(
		.INIT('h32cd)
	) name8245 (
		_w10922_,
		_w11244_,
		_w12246_,
		_w12292_,
		_w12293_
	);
	LUT4 #(
		.INIT('h4c08)
	) name8246 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w12291_,
		_w12293_,
		_w12294_
	);
	LUT2 #(
		.INIT('he)
	) name8247 (
		_w12289_,
		_w12294_,
		_w12295_
	);
	LUT3 #(
		.INIT('h80)
	) name8248 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12296_
	);
	LUT2 #(
		.INIT('h1)
	) name8249 (
		_w5047_,
		_w12296_,
		_w12297_
	);
	LUT4 #(
		.INIT('hbf00)
	) name8250 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12297_,
		_w12298_
	);
	LUT4 #(
		.INIT('h1000)
	) name8251 (
		\core_c_dec_SHTop_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12299_
	);
	LUT3 #(
		.INIT('h02)
	) name8252 (
		_w4102_,
		_w12299_,
		_w12298_,
		_w12300_
	);
	LUT4 #(
		.INIT('h8000)
	) name8253 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		_w12301_
	);
	LUT3 #(
		.INIT('h6c)
	) name8254 (
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		_w12301_,
		_w12302_
	);
	LUT3 #(
		.INIT('h20)
	) name8255 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12302_,
		_w12303_
	);
	LUT3 #(
		.INIT('h78)
	) name8256 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		_w12304_
	);
	LUT3 #(
		.INIT('h20)
	) name8257 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12304_,
		_w12305_
	);
	LUT4 #(
		.INIT('h8000)
	) name8258 (
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		_w12301_,
		_w12306_
	);
	LUT2 #(
		.INIT('h8)
	) name8259 (
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		_w12306_,
		_w12307_
	);
	LUT3 #(
		.INIT('h80)
	) name8260 (
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		_w12306_,
		_w12308_
	);
	LUT4 #(
		.INIT('h8000)
	) name8261 (
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		_w12306_,
		_w12309_
	);
	LUT2 #(
		.INIT('h8)
	) name8262 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		_w12309_,
		_w12310_
	);
	LUT3 #(
		.INIT('h80)
	) name8263 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		_w12309_,
		_w12311_
	);
	LUT4 #(
		.INIT('h8000)
	) name8264 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		_w12309_,
		_w12312_
	);
	LUT3 #(
		.INIT('h48)
	) name8265 (
		\sport0_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		_w12109_,
		_w12312_,
		_w12313_
	);
	LUT3 #(
		.INIT('h04)
	) name8266 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12314_
	);
	LUT4 #(
		.INIT('h4544)
	) name8267 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5784_,
		_w5911_,
		_w5913_,
		_w12315_
	);
	LUT2 #(
		.INIT('h2)
	) name8268 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8647_,
		_w12316_
	);
	LUT2 #(
		.INIT('h1)
	) name8269 (
		_w12315_,
		_w12316_,
		_w12317_
	);
	LUT3 #(
		.INIT('h13)
	) name8270 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 ,
		_w9894_,
		_w12318_
	);
	LUT4 #(
		.INIT('h0002)
	) name8271 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w12318_,
		_w12319_
	);
	LUT4 #(
		.INIT('h5700)
	) name8272 (
		_w12282_,
		_w12315_,
		_w12316_,
		_w12319_,
		_w12320_
	);
	LUT4 #(
		.INIT('h313b)
	) name8273 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 ,
		_w11308_,
		_w11635_,
		_w12321_
	);
	LUT3 #(
		.INIT('h45)
	) name8274 (
		_w11624_,
		_w12320_,
		_w12321_,
		_w12322_
	);
	LUT2 #(
		.INIT('h9)
	) name8275 (
		_w11226_,
		_w11228_,
		_w12323_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name8276 (
		_w10433_,
		_w10640_,
		_w10645_,
		_w12323_,
		_w12324_
	);
	LUT2 #(
		.INIT('h9)
	) name8277 (
		_w10626_,
		_w10628_,
		_w12325_
	);
	LUT4 #(
		.INIT('h80aa)
	) name8278 (
		_w10639_,
		_w10352_,
		_w10430_,
		_w10432_,
		_w12326_
	);
	LUT4 #(
		.INIT('h2232)
	) name8279 (
		_w10574_,
		_w10643_,
		_w10642_,
		_w12326_,
		_w12327_
	);
	LUT4 #(
		.INIT('h8dd8)
	) name8280 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12324_,
		_w12325_,
		_w12327_,
		_w12328_
	);
	LUT2 #(
		.INIT('h9)
	) name8281 (
		_w10563_,
		_w10573_,
		_w12329_
	);
	LUT4 #(
		.INIT('h0541)
	) name8282 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10642_,
		_w12329_,
		_w12326_,
		_w12330_
	);
	LUT4 #(
		.INIT('h1331)
	) name8283 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12330_,
		_w12325_,
		_w12327_,
		_w12331_
	);
	LUT2 #(
		.INIT('h9)
	) name8284 (
		_w10633_,
		_w10634_,
		_w12332_
	);
	LUT4 #(
		.INIT('h4055)
	) name8285 (
		_w10638_,
		_w10352_,
		_w10430_,
		_w10432_,
		_w12333_
	);
	LUT4 #(
		.INIT('h0514)
	) name8286 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10641_,
		_w12332_,
		_w12333_,
		_w12334_
	);
	LUT4 #(
		.INIT('h0a82)
	) name8287 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10642_,
		_w12329_,
		_w12326_,
		_w12335_
	);
	LUT2 #(
		.INIT('h1)
	) name8288 (
		_w12334_,
		_w12335_,
		_w12336_
	);
	LUT2 #(
		.INIT('h9)
	) name8289 (
		_w10636_,
		_w10637_,
		_w12337_
	);
	LUT4 #(
		.INIT('h708f)
	) name8290 (
		_w10352_,
		_w10430_,
		_w10432_,
		_w12337_,
		_w12338_
	);
	LUT2 #(
		.INIT('h1)
	) name8291 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12338_,
		_w12339_
	);
	LUT4 #(
		.INIT('ha082)
	) name8292 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10641_,
		_w12332_,
		_w12333_,
		_w12340_
	);
	LUT2 #(
		.INIT('h1)
	) name8293 (
		_w12339_,
		_w12340_,
		_w12341_
	);
	LUT2 #(
		.INIT('h9)
	) name8294 (
		_w10389_,
		_w10427_,
		_w12342_
	);
	LUT4 #(
		.INIT('h0df2)
	) name8295 (
		_w10352_,
		_w10429_,
		_w10431_,
		_w12342_,
		_w12343_
	);
	LUT3 #(
		.INIT('h36)
	) name8296 (
		_w10353_,
		_w10387_,
		_w10428_,
		_w12344_
	);
	LUT2 #(
		.INIT('h9)
	) name8297 (
		_w10352_,
		_w12344_,
		_w12345_
	);
	LUT3 #(
		.INIT('h41)
	) name8298 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10352_,
		_w12344_,
		_w12346_
	);
	LUT3 #(
		.INIT('h0d)
	) name8299 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12343_,
		_w12346_,
		_w12347_
	);
	LUT3 #(
		.INIT('h27)
	) name8300 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12338_,
		_w12343_,
		_w12348_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8301 (
		_w10253_,
		_w10254_,
		_w10319_,
		_w10351_,
		_w12349_
	);
	LUT4 #(
		.INIT('h349e)
	) name8302 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10320_,
		_w10351_,
		_w12344_,
		_w12350_
	);
	LUT2 #(
		.INIT('h9)
	) name8303 (
		_w10255_,
		_w10319_,
		_w12351_
	);
	LUT3 #(
		.INIT('h14)
	) name8304 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10255_,
		_w10319_,
		_w12352_
	);
	LUT3 #(
		.INIT('h0d)
	) name8305 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12349_,
		_w12352_,
		_w12353_
	);
	LUT4 #(
		.INIT('h0154)
	) name8306 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10289_,
		_w10318_,
		_w11639_,
		_w12354_
	);
	LUT4 #(
		.INIT('h007d)
	) name8307 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10255_,
		_w10319_,
		_w12354_,
		_w12355_
	);
	LUT2 #(
		.INIT('h9)
	) name8308 (
		_w10305_,
		_w10317_,
		_w12356_
	);
	LUT3 #(
		.INIT('h41)
	) name8309 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10305_,
		_w10317_,
		_w12357_
	);
	LUT3 #(
		.INIT('h07)
	) name8310 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11637_,
		_w12357_,
		_w12358_
	);
	LUT3 #(
		.INIT('h36)
	) name8311 (
		_w10300_,
		_w10301_,
		_w10314_,
		_w12359_
	);
	LUT3 #(
		.INIT('h14)
	) name8312 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10313_,
		_w12359_,
		_w12360_
	);
	LUT4 #(
		.INIT('h007d)
	) name8313 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10305_,
		_w10317_,
		_w12360_,
		_w12361_
	);
	LUT4 #(
		.INIT('hc16b)
	) name8314 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10311_,
		_w10312_,
		_w12359_,
		_w12362_
	);
	LUT3 #(
		.INIT('h41)
	) name8315 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10306_,
		_w10310_,
		_w12363_
	);
	LUT4 #(
		.INIT('h00d7)
	) name8316 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10311_,
		_w10312_,
		_w12363_,
		_w12364_
	);
	LUT2 #(
		.INIT('h8)
	) name8317 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		_w12365_
	);
	LUT4 #(
		.INIT('h0154)
	) name8318 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10308_,
		_w12365_,
		_w12366_
	);
	LUT4 #(
		.INIT('h00d7)
	) name8319 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10306_,
		_w10310_,
		_w12366_,
		_w12367_
	);
	LUT4 #(
		.INIT('ha802)
	) name8320 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10308_,
		_w12365_,
		_w12368_
	);
	LUT2 #(
		.INIT('h4)
	) name8321 (
		_w5869_,
		_w11083_,
		_w12369_
	);
	LUT2 #(
		.INIT('h1)
	) name8322 (
		_w12368_,
		_w12369_,
		_w12370_
	);
	LUT2 #(
		.INIT('h2)
	) name8323 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 ,
		\memc_usysr_DO_reg[10]/NET0131 ,
		_w12371_
	);
	LUT3 #(
		.INIT('h10)
	) name8324 (
		_w12368_,
		_w12369_,
		_w12371_,
		_w12372_
	);
	LUT2 #(
		.INIT('h4)
	) name8325 (
		_w12367_,
		_w12372_,
		_w12373_
	);
	LUT2 #(
		.INIT('h8)
	) name8326 (
		_w12364_,
		_w12373_,
		_w12374_
	);
	LUT2 #(
		.INIT('h8)
	) name8327 (
		_w12362_,
		_w12374_,
		_w12375_
	);
	LUT2 #(
		.INIT('h8)
	) name8328 (
		_w12361_,
		_w12375_,
		_w12376_
	);
	LUT4 #(
		.INIT('he000)
	) name8329 (
		_w11638_,
		_w11640_,
		_w12358_,
		_w12376_,
		_w12377_
	);
	LUT2 #(
		.INIT('h8)
	) name8330 (
		_w12355_,
		_w12377_,
		_w12378_
	);
	LUT3 #(
		.INIT('h40)
	) name8331 (
		_w12353_,
		_w12350_,
		_w12378_,
		_w12379_
	);
	LUT3 #(
		.INIT('h20)
	) name8332 (
		_w12348_,
		_w12347_,
		_w12379_,
		_w12380_
	);
	LUT4 #(
		.INIT('h2000)
	) name8333 (
		_w12331_,
		_w12341_,
		_w12336_,
		_w12380_,
		_w12381_
	);
	LUT2 #(
		.INIT('h4)
	) name8334 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12324_,
		_w12382_
	);
	LUT2 #(
		.INIT('h9)
	) name8335 (
		_w11219_,
		_w11225_,
		_w12383_
	);
	LUT4 #(
		.INIT('h004f)
	) name8336 (
		_w10433_,
		_w10640_,
		_w10645_,
		_w11229_,
		_w12384_
	);
	LUT4 #(
		.INIT('ha082)
	) name8337 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11239_,
		_w12383_,
		_w12384_,
		_w12385_
	);
	LUT2 #(
		.INIT('h1)
	) name8338 (
		_w12382_,
		_w12385_,
		_w12386_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8339 (
		_w11624_,
		_w12328_,
		_w12381_,
		_w12386_,
		_w12387_
	);
	LUT2 #(
		.INIT('he)
	) name8340 (
		_w12322_,
		_w12387_,
		_w12388_
	);
	LUT4 #(
		.INIT('h007f)
	) name8341 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w5045_,
		_w5046_,
		_w9323_,
		_w12389_
	);
	LUT2 #(
		.INIT('h4)
	) name8342 (
		_w4967_,
		_w12389_,
		_w12390_
	);
	LUT2 #(
		.INIT('hb)
	) name8343 (
		_w4967_,
		_w12389_,
		_w12391_
	);
	LUT2 #(
		.INIT('h4)
	) name8344 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w12392_
	);
	LUT2 #(
		.INIT('h4)
	) name8345 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w12393_
	);
	LUT2 #(
		.INIT('h8)
	) name8346 (
		_w5028_,
		_w12393_,
		_w12394_
	);
	LUT4 #(
		.INIT('h8000)
	) name8347 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w5028_,
		_w12392_,
		_w12393_,
		_w12395_
	);
	LUT3 #(
		.INIT('h01)
	) name8348 (
		_w5043_,
		_w5048_,
		_w12395_,
		_w12396_
	);
	LUT2 #(
		.INIT('h8)
	) name8349 (
		_w12390_,
		_w12396_,
		_w12397_
	);
	LUT2 #(
		.INIT('h1)
	) name8350 (
		_w4104_,
		_w12397_,
		_w12398_
	);
	LUT4 #(
		.INIT('h808c)
	) name8351 (
		\core_c_dec_Post2_E_reg/P0001 ,
		_w4102_,
		_w4104_,
		_w12397_,
		_w12399_
	);
	LUT3 #(
		.INIT('h80)
	) name8352 (
		_w11389_,
		_w11503_,
		_w11872_,
		_w12400_
	);
	LUT4 #(
		.INIT('h1000)
	) name8353 (
		_w11348_,
		_w11357_,
		_w11388_,
		_w11439_,
		_w12401_
	);
	LUT4 #(
		.INIT('h0f04)
	) name8354 (
		_w11444_,
		_w11405_,
		_w11487_,
		_w12401_,
		_w12402_
	);
	LUT2 #(
		.INIT('h1)
	) name8355 (
		_w12400_,
		_w12402_,
		_w12403_
	);
	LUT4 #(
		.INIT('hf400)
	) name8356 (
		_w11444_,
		_w11423_,
		_w11462_,
		_w11874_,
		_w12404_
	);
	LUT3 #(
		.INIT('h0b)
	) name8357 (
		_w11446_,
		_w11469_,
		_w12404_,
		_w12405_
	);
	LUT3 #(
		.INIT('h2a)
	) name8358 (
		_w11386_,
		_w12403_,
		_w12405_,
		_w12406_
	);
	LUT4 #(
		.INIT('h000d)
	) name8359 (
		_w11386_,
		_w11530_,
		_w11522_,
		_w11524_,
		_w12407_
	);
	LUT3 #(
		.INIT('h2a)
	) name8360 (
		_w11341_,
		_w11594_,
		_w12407_,
		_w12408_
	);
	LUT3 #(
		.INIT('h80)
	) name8361 (
		_w11580_,
		_w11437_,
		_w11479_,
		_w12409_
	);
	LUT3 #(
		.INIT('h04)
	) name8362 (
		_w12408_,
		_w12409_,
		_w12406_,
		_w12410_
	);
	LUT3 #(
		.INIT('h10)
	) name8363 (
		_w11586_,
		_w11590_,
		_w11441_,
		_w12411_
	);
	LUT3 #(
		.INIT('h02)
	) name8364 (
		_w11333_,
		_w11385_,
		_w11335_,
		_w12412_
	);
	LUT4 #(
		.INIT('hfd75)
	) name8365 (
		_w11333_,
		_w11385_,
		_w11335_,
		_w11528_,
		_w12413_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name8366 (
		_w11534_,
		_w11446_,
		_w11466_,
		_w12413_,
		_w12414_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name8367 (
		_w11406_,
		_w11530_,
		_w11504_,
		_w11450_,
		_w12415_
	);
	LUT3 #(
		.INIT('h02)
	) name8368 (
		_w11386_,
		_w11540_,
		_w11492_,
		_w12416_
	);
	LUT3 #(
		.INIT('h40)
	) name8369 (
		_w11444_,
		_w11476_,
		_w11453_,
		_w12417_
	);
	LUT4 #(
		.INIT('ha820)
	) name8370 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001 ,
		_w12418_
	);
	LUT4 #(
		.INIT('h007f)
	) name8371 (
		_w11389_,
		_w11538_,
		_w11491_,
		_w12418_,
		_w12419_
	);
	LUT3 #(
		.INIT('h10)
	) name8372 (
		_w11591_,
		_w12417_,
		_w12419_,
		_w12420_
	);
	LUT4 #(
		.INIT('h4000)
	) name8373 (
		_w12416_,
		_w12420_,
		_w12414_,
		_w12415_,
		_w12421_
	);
	LUT4 #(
		.INIT('hf040)
	) name8374 (
		_w11444_,
		_w11423_,
		_w11458_,
		_w11462_,
		_w12422_
	);
	LUT3 #(
		.INIT('h40)
	) name8375 (
		_w11444_,
		_w11537_,
		_w11392_,
		_w12423_
	);
	LUT3 #(
		.INIT('h54)
	) name8376 (
		_w11386_,
		_w12422_,
		_w12423_,
		_w12424_
	);
	LUT4 #(
		.INIT('h00f4)
	) name8377 (
		_w11444_,
		_w11414_,
		_w11481_,
		_w11512_,
		_w12425_
	);
	LUT4 #(
		.INIT('h0f04)
	) name8378 (
		_w11444_,
		_w11428_,
		_w11501_,
		_w11455_,
		_w12426_
	);
	LUT4 #(
		.INIT('hf040)
	) name8379 (
		_w11444_,
		_w11405_,
		_w11485_,
		_w12401_,
		_w12427_
	);
	LUT3 #(
		.INIT('h01)
	) name8380 (
		_w12426_,
		_w12427_,
		_w12425_,
		_w12428_
	);
	LUT2 #(
		.INIT('h4)
	) name8381 (
		_w12424_,
		_w12428_,
		_w12429_
	);
	LUT3 #(
		.INIT('h80)
	) name8382 (
		_w12411_,
		_w12421_,
		_w12429_,
		_w12430_
	);
	LUT2 #(
		.INIT('h4)
	) name8383 (
		_w11386_,
		_w11429_,
		_w12431_
	);
	LUT4 #(
		.INIT('hc480)
	) name8384 (
		_w11386_,
		_w11341_,
		_w11415_,
		_w11429_,
		_w12432_
	);
	LUT4 #(
		.INIT('h0004)
	) name8385 (
		_w11549_,
		_w11554_,
		_w11559_,
		_w12432_,
		_w12433_
	);
	LUT3 #(
		.INIT('h80)
	) name8386 (
		_w11910_,
		_w11834_,
		_w12433_,
		_w12434_
	);
	LUT4 #(
		.INIT('h8000)
	) name8387 (
		_w11433_,
		_w12434_,
		_w12410_,
		_w12430_,
		_w12435_
	);
	LUT4 #(
		.INIT('h7020)
	) name8388 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11318_,
		_w11830_,
		_w12435_,
		_w12436_
	);
	LUT4 #(
		.INIT('h5545)
	) name8389 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w12437_
	);
	LUT2 #(
		.INIT('h1)
	) name8390 (
		_w12436_,
		_w12437_,
		_w12438_
	);
	LUT4 #(
		.INIT('h80c4)
	) name8391 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w12291_,
		_w12293_,
		_w12439_
	);
	LUT4 #(
		.INIT('h0040)
	) name8392 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w9452_,
		_w11305_,
		_w12440_
	);
	LUT2 #(
		.INIT('h2)
	) name8393 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001 ,
		_w11310_,
		_w12441_
	);
	LUT3 #(
		.INIT('h10)
	) name8394 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11658_,
		_w12442_
	);
	LUT3 #(
		.INIT('h01)
	) name8395 (
		_w9946_,
		_w12441_,
		_w12442_,
		_w12443_
	);
	LUT3 #(
		.INIT('h70)
	) name8396 (
		_w12284_,
		_w12440_,
		_w12443_,
		_w12444_
	);
	LUT2 #(
		.INIT('h1)
	) name8397 (
		_w12439_,
		_w12444_,
		_w12445_
	);
	LUT4 #(
		.INIT('h4000)
	) name8398 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11406_,
		_w11476_,
		_w12446_
	);
	LUT2 #(
		.INIT('h1)
	) name8399 (
		_w11551_,
		_w12446_,
		_w12447_
	);
	LUT3 #(
		.INIT('h10)
	) name8400 (
		_w11549_,
		_w11595_,
		_w12447_,
		_w12448_
	);
	LUT4 #(
		.INIT('h1000)
	) name8401 (
		_w11549_,
		_w11595_,
		_w11968_,
		_w12447_,
		_w12449_
	);
	LUT3 #(
		.INIT('h80)
	) name8402 (
		_w11577_,
		_w11910_,
		_w11834_,
		_w12450_
	);
	LUT4 #(
		.INIT('h8000)
	) name8403 (
		_w11577_,
		_w11871_,
		_w11910_,
		_w11834_,
		_w12451_
	);
	LUT3 #(
		.INIT('hc8)
	) name8404 (
		_w11555_,
		_w11484_,
		_w11888_,
		_w12452_
	);
	LUT3 #(
		.INIT('h02)
	) name8405 (
		_w11386_,
		_w11528_,
		_w11957_,
		_w12453_
	);
	LUT3 #(
		.INIT('hc8)
	) name8406 (
		_w11587_,
		_w11872_,
		_w11880_,
		_w12454_
	);
	LUT3 #(
		.INIT('h20)
	) name8407 (
		_w11389_,
		_w11386_,
		_w11445_,
		_w12455_
	);
	LUT3 #(
		.INIT('hc8)
	) name8408 (
		_w11435_,
		_w11449_,
		_w12455_,
		_w12456_
	);
	LUT4 #(
		.INIT('h0001)
	) name8409 (
		_w12452_,
		_w12453_,
		_w12454_,
		_w12456_,
		_w12457_
	);
	LUT2 #(
		.INIT('h8)
	) name8410 (
		_w11588_,
		_w11507_,
		_w12458_
	);
	LUT4 #(
		.INIT('ha820)
	) name8411 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001 ,
		_w12459_
	);
	LUT3 #(
		.INIT('h0d)
	) name8412 (
		_w11578_,
		_w11471_,
		_w12459_,
		_w12460_
	);
	LUT3 #(
		.INIT('h08)
	) name8413 (
		_w11389_,
		_w11476_,
		_w11512_,
		_w12461_
	);
	LUT2 #(
		.INIT('h8)
	) name8414 (
		_w11415_,
		_w11488_,
		_w12462_
	);
	LUT3 #(
		.INIT('h10)
	) name8415 (
		_w12461_,
		_w12462_,
		_w12460_,
		_w12463_
	);
	LUT3 #(
		.INIT('h0e)
	) name8416 (
		_w11393_,
		_w11589_,
		_w11501_,
		_w12464_
	);
	LUT2 #(
		.INIT('h4)
	) name8417 (
		_w11957_,
		_w12412_,
		_w12465_
	);
	LUT4 #(
		.INIT('h0100)
	) name8418 (
		_w12458_,
		_w12464_,
		_w12465_,
		_w12463_,
		_w12466_
	);
	LUT4 #(
		.INIT('h2220)
	) name8419 (
		_w11386_,
		_w11540_,
		_w11552_,
		_w11474_,
		_w12467_
	);
	LUT4 #(
		.INIT('h1000)
	) name8420 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11385_,
		_w11358_,
		_w11382_,
		_w12468_
	);
	LUT3 #(
		.INIT('ha8)
	) name8421 (
		_w11458_,
		_w12431_,
		_w12468_,
		_w12469_
	);
	LUT2 #(
		.INIT('h1)
	) name8422 (
		_w12467_,
		_w12469_,
		_w12470_
	);
	LUT2 #(
		.INIT('h2)
	) name8423 (
		_w11515_,
		_w11953_,
		_w12471_
	);
	LUT4 #(
		.INIT('h8000)
	) name8424 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11341_,
		_w11358_,
		_w11395_,
		_w12472_
	);
	LUT2 #(
		.INIT('h1)
	) name8425 (
		_w11403_,
		_w12472_,
		_w12473_
	);
	LUT4 #(
		.INIT('h0015)
	) name8426 (
		_w11403_,
		_w11522_,
		_w11863_,
		_w12472_,
		_w12474_
	);
	LUT2 #(
		.INIT('h4)
	) name8427 (
		_w12471_,
		_w12474_,
		_w12475_
	);
	LUT4 #(
		.INIT('h135f)
	) name8428 (
		_w11409_,
		_w11558_,
		_w11469_,
		_w11841_,
		_w12476_
	);
	LUT3 #(
		.INIT('ha8)
	) name8429 (
		_w11538_,
		_w11552_,
		_w11474_,
		_w12477_
	);
	LUT2 #(
		.INIT('h8)
	) name8430 (
		_w11465_,
		_w11973_,
		_w12478_
	);
	LUT3 #(
		.INIT('h10)
	) name8431 (
		_w12477_,
		_w12478_,
		_w12476_,
		_w12479_
	);
	LUT4 #(
		.INIT('h8000)
	) name8432 (
		_w12475_,
		_w12479_,
		_w12466_,
		_w12470_,
		_w12480_
	);
	LUT4 #(
		.INIT('h8000)
	) name8433 (
		_w12449_,
		_w12451_,
		_w12457_,
		_w12480_,
		_w12481_
	);
	LUT4 #(
		.INIT('h7020)
	) name8434 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w11331_,
		_w11946_,
		_w12481_,
		_w12482_
	);
	LUT4 #(
		.INIT('h5545)
	) name8435 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001 ,
		_w9453_,
		_w9894_,
		_w11945_,
		_w12483_
	);
	LUT2 #(
		.INIT('h1)
	) name8436 (
		_w12482_,
		_w12483_,
		_w12484_
	);
	LUT2 #(
		.INIT('h2)
	) name8437 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8671_,
		_w12485_
	);
	LUT4 #(
		.INIT('h00ab)
	) name8438 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5937_,
		_w6038_,
		_w12485_,
		_w12486_
	);
	LUT2 #(
		.INIT('h2)
	) name8439 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12486_,
		_w12487_
	);
	LUT3 #(
		.INIT('h02)
	) name8440 (
		_w11386_,
		_w11335_,
		_w11592_,
		_w12488_
	);
	LUT3 #(
		.INIT('he0)
	) name8441 (
		_w11393_,
		_w11589_,
		_w11848_,
		_w12489_
	);
	LUT3 #(
		.INIT('h08)
	) name8442 (
		_w11389_,
		_w11445_,
		_w11844_,
		_w12490_
	);
	LUT4 #(
		.INIT('ha820)
	) name8443 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001 ,
		_w12491_
	);
	LUT3 #(
		.INIT('h07)
	) name8444 (
		_w11578_,
		_w11873_,
		_w12491_,
		_w12492_
	);
	LUT2 #(
		.INIT('h4)
	) name8445 (
		_w12490_,
		_w12492_,
		_w12493_
	);
	LUT3 #(
		.INIT('h10)
	) name8446 (
		_w12488_,
		_w12489_,
		_w12493_,
		_w12494_
	);
	LUT3 #(
		.INIT('ha8)
	) name8447 (
		_w11537_,
		_w11420_,
		_w11421_,
		_w12495_
	);
	LUT3 #(
		.INIT('h20)
	) name8448 (
		_w11389_,
		_w11386_,
		_w11476_,
		_w12496_
	);
	LUT3 #(
		.INIT('hc8)
	) name8449 (
		_w11588_,
		_w11863_,
		_w12496_,
		_w12497_
	);
	LUT2 #(
		.INIT('h1)
	) name8450 (
		_w12495_,
		_w12497_,
		_w12498_
	);
	LUT2 #(
		.INIT('h8)
	) name8451 (
		_w11435_,
		_w11841_,
		_w12499_
	);
	LUT4 #(
		.INIT('hfd75)
	) name8452 (
		_w11333_,
		_w11385_,
		_w11540_,
		_w11494_,
		_w12500_
	);
	LUT4 #(
		.INIT('h7770)
	) name8453 (
		_w11587_,
		_w11484_,
		_w11957_,
		_w12500_,
		_w12501_
	);
	LUT2 #(
		.INIT('h4)
	) name8454 (
		_w12499_,
		_w12501_,
		_w12502_
	);
	LUT2 #(
		.INIT('h8)
	) name8455 (
		_w11872_,
		_w11973_,
		_w12503_
	);
	LUT3 #(
		.INIT('h02)
	) name8456 (
		_w11333_,
		_w11385_,
		_w11498_,
		_w12504_
	);
	LUT2 #(
		.INIT('h2)
	) name8457 (
		_w11386_,
		_w11457_,
		_w12505_
	);
	LUT4 #(
		.INIT('hfd75)
	) name8458 (
		_w11333_,
		_w11385_,
		_w11498_,
		_w11457_,
		_w12506_
	);
	LUT3 #(
		.INIT('h0e)
	) name8459 (
		_w11552_,
		_w11474_,
		_w12506_,
		_w12507_
	);
	LUT2 #(
		.INIT('h1)
	) name8460 (
		_w11953_,
		_w11950_,
		_w12508_
	);
	LUT3 #(
		.INIT('he0)
	) name8461 (
		_w11393_,
		_w11589_,
		_w11875_,
		_w12509_
	);
	LUT4 #(
		.INIT('h0001)
	) name8462 (
		_w12503_,
		_w12507_,
		_w12508_,
		_w12509_,
		_w12510_
	);
	LUT4 #(
		.INIT('h8000)
	) name8463 (
		_w12502_,
		_w12510_,
		_w12494_,
		_w12498_,
		_w12511_
	);
	LUT4 #(
		.INIT('h0057)
	) name8464 (
		_w11341_,
		_w11396_,
		_w11548_,
		_w11438_,
		_w12512_
	);
	LUT3 #(
		.INIT('h10)
	) name8465 (
		_w11426_,
		_w11971_,
		_w12512_,
		_w12513_
	);
	LUT3 #(
		.INIT('hc8)
	) name8466 (
		_w11547_,
		_w11854_,
		_w11976_,
		_w12514_
	);
	LUT3 #(
		.INIT('hc8)
	) name8467 (
		_w11409_,
		_w11507_,
		_w11896_,
		_w12515_
	);
	LUT2 #(
		.INIT('h1)
	) name8468 (
		_w11403_,
		_w11885_,
		_w12516_
	);
	LUT4 #(
		.INIT('h0001)
	) name8469 (
		_w11403_,
		_w11551_,
		_w11885_,
		_w12446_,
		_w12517_
	);
	LUT3 #(
		.INIT('h04)
	) name8470 (
		_w12515_,
		_w12517_,
		_w12514_,
		_w12518_
	);
	LUT2 #(
		.INIT('h8)
	) name8471 (
		_w12513_,
		_w12518_,
		_w12519_
	);
	LUT4 #(
		.INIT('h4000)
	) name8472 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12450_,
		_w12511_,
		_w12519_,
		_w12520_
	);
	LUT4 #(
		.INIT('h222e)
	) name8473 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001 ,
		_w11946_,
		_w12487_,
		_w12520_,
		_w12521_
	);
	LUT4 #(
		.INIT('h7020)
	) name8474 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w11331_,
		_w12048_,
		_w12481_,
		_w12522_
	);
	LUT2 #(
		.INIT('h1)
	) name8475 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001 ,
		_w12048_,
		_w12523_
	);
	LUT2 #(
		.INIT('h1)
	) name8476 (
		_w12522_,
		_w12523_,
		_w12524_
	);
	LUT4 #(
		.INIT('h2000)
	) name8477 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12525_
	);
	LUT3 #(
		.INIT('ha8)
	) name8478 (
		_w4102_,
		_w11926_,
		_w12525_,
		_w12526_
	);
	LUT4 #(
		.INIT('h222e)
	) name8479 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001 ,
		_w12048_,
		_w12487_,
		_w12520_,
		_w12527_
	);
	LUT3 #(
		.INIT('h20)
	) name8480 (
		_w4884_,
		_w9412_,
		_w9413_,
		_w12528_
	);
	LUT4 #(
		.INIT('h0800)
	) name8481 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		_w4884_,
		_w9412_,
		_w9413_,
		_w12529_
	);
	LUT3 #(
		.INIT('h20)
	) name8482 (
		_w9076_,
		_w9412_,
		_w9413_,
		_w12530_
	);
	LUT4 #(
		.INIT('h3302)
	) name8483 (
		\bdma_CMcnt_reg[1]/NET0131 ,
		_w9414_,
		_w12529_,
		_w12530_,
		_w12531_
	);
	LUT3 #(
		.INIT('h12)
	) name8484 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		_w9414_,
		_w12528_,
		_w12532_
	);
	LUT3 #(
		.INIT('h01)
	) name8485 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w4762_,
		_w4763_,
		_w12533_
	);
	LUT4 #(
		.INIT('h8a00)
	) name8486 (
		_w4761_,
		_w5534_,
		_w9411_,
		_w12533_,
		_w12534_
	);
	LUT4 #(
		.INIT('h2223)
	) name8487 (
		\bdma_BMcyc_del_reg/P0001 ,
		\bdma_BSreq_reg/NET0131 ,
		_w5536_,
		_w9081_,
		_w12535_
	);
	LUT2 #(
		.INIT('hb)
	) name8488 (
		_w12534_,
		_w12535_,
		_w12536_
	);
	LUT4 #(
		.INIT('h7020)
	) name8489 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11318_,
		_w11329_,
		_w12435_,
		_w12537_
	);
	LUT2 #(
		.INIT('h1)
	) name8490 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001 ,
		_w11329_,
		_w12538_
	);
	LUT2 #(
		.INIT('h1)
	) name8491 (
		_w12537_,
		_w12538_,
		_w12539_
	);
	LUT2 #(
		.INIT('h1)
	) name8492 (
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w12540_
	);
	LUT4 #(
		.INIT('hb41e)
	) name8493 (
		\ITFS0_pad ,
		\T_TFS0_pad ,
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w9405_,
		_w12541_
	);
	LUT2 #(
		.INIT('h2)
	) name8494 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_cfg_TFSgi_d_reg/NET0131 ,
		_w12542_
	);
	LUT2 #(
		.INIT('h8)
	) name8495 (
		_w12541_,
		_w12542_,
		_w12543_
	);
	LUT4 #(
		.INIT('h3500)
	) name8496 (
		\sport0_cfg_TFSg_d2_reg/NET0131 ,
		\sport0_cfg_TFSg_d3_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w12544_
	);
	LUT4 #(
		.INIT('hfb00)
	) name8497 (
		\sport0_cfg_TFSg_d1_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		\sport0_txctl_TCS_reg[0]/NET0131 ,
		_w12545_
	);
	LUT2 #(
		.INIT('h4)
	) name8498 (
		_w12544_,
		_w12545_,
		_w12546_
	);
	LUT4 #(
		.INIT('hd500)
	) name8499 (
		_w12540_,
		_w12541_,
		_w12542_,
		_w12546_,
		_w12547_
	);
	LUT3 #(
		.INIT('h13)
	) name8500 (
		\sport0_txctl_TCS_reg[0]/NET0131 ,
		\sport0_txctl_TCS_reg[1]/NET0131 ,
		\sport0_txctl_TCS_reg[2]/NET0131 ,
		_w12548_
	);
	LUT3 #(
		.INIT('h04)
	) name8501 (
		\sport0_txctl_TCS_reg[0]/NET0131 ,
		\sport0_txctl_TCS_reg[1]/NET0131 ,
		\sport0_txctl_TCS_reg[2]/NET0131 ,
		_w12549_
	);
	LUT4 #(
		.INIT('h0001)
	) name8502 (
		\sport0_txctl_Bcnt_reg[0]/NET0131 ,
		\sport0_txctl_Bcnt_reg[1]/NET0131 ,
		\sport0_txctl_Bcnt_reg[2]/NET0131 ,
		\sport0_txctl_Bcnt_reg[3]/NET0131 ,
		_w12550_
	);
	LUT3 #(
		.INIT('h8c)
	) name8503 (
		\sport0_txctl_Bcnt_reg[4]/NET0131 ,
		_w12549_,
		_w12550_,
		_w12551_
	);
	LUT4 #(
		.INIT('h001f)
	) name8504 (
		\sport0_txctl_TCS_reg[2]/NET0131 ,
		_w12547_,
		_w12548_,
		_w12551_,
		_w12552_
	);
	LUT4 #(
		.INIT('hffe0)
	) name8505 (
		\sport0_txctl_TCS_reg[2]/NET0131 ,
		_w12547_,
		_w12548_,
		_w12551_,
		_w12553_
	);
	LUT3 #(
		.INIT('hca)
	) name8506 (
		\sport0_txctl_TXSHT_reg[14]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w12552_,
		_w12554_
	);
	LUT4 #(
		.INIT('h80aa)
	) name8507 (
		_w9946_,
		_w12328_,
		_w12381_,
		_w12386_,
		_w12555_
	);
	LUT2 #(
		.INIT('h2)
	) name8508 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001 ,
		_w11310_,
		_w12556_
	);
	LUT3 #(
		.INIT('h01)
	) name8509 (
		_w9946_,
		_w12442_,
		_w12556_,
		_w12557_
	);
	LUT4 #(
		.INIT('hef00)
	) name8510 (
		_w12315_,
		_w12316_,
		_w12440_,
		_w12557_,
		_w12558_
	);
	LUT2 #(
		.INIT('h1)
	) name8511 (
		_w12555_,
		_w12558_,
		_w12559_
	);
	LUT4 #(
		.INIT('h4544)
	) name8512 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w7793_,
		_w7903_,
		_w7905_,
		_w12560_
	);
	LUT2 #(
		.INIT('h2)
	) name8513 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8974_,
		_w12561_
	);
	LUT2 #(
		.INIT('h1)
	) name8514 (
		_w12560_,
		_w12561_,
		_w12562_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8515 (
		_w11410_,
		_w11558_,
		_w11894_,
		_w11860_,
		_w12563_
	);
	LUT4 #(
		.INIT('hf040)
	) name8516 (
		_w11444_,
		_w11423_,
		_w11485_,
		_w11462_,
		_w12564_
	);
	LUT3 #(
		.INIT('h0e)
	) name8517 (
		_w11530_,
		_w12024_,
		_w12564_,
		_w12565_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name8518 (
		_w11534_,
		_w11492_,
		_w11453_,
		_w11471_,
		_w12566_
	);
	LUT4 #(
		.INIT('h1000)
	) name8519 (
		_w11595_,
		_w12563_,
		_w12565_,
		_w12566_,
		_w12567_
	);
	LUT2 #(
		.INIT('h4)
	) name8520 (
		_w11386_,
		_w11415_,
		_w12568_
	);
	LUT3 #(
		.INIT('hc8)
	) name8521 (
		_w11555_,
		_w11495_,
		_w12568_,
		_w12569_
	);
	LUT3 #(
		.INIT('hc8)
	) name8522 (
		_w11587_,
		_w11854_,
		_w11880_,
		_w12570_
	);
	LUT3 #(
		.INIT('h0d)
	) name8523 (
		_w11406_,
		_w11585_,
		_w11901_,
		_w12571_
	);
	LUT3 #(
		.INIT('ha8)
	) name8524 (
		_w11499_,
		_w11522_,
		_w11523_,
		_w12572_
	);
	LUT4 #(
		.INIT('h0010)
	) name8525 (
		_w12569_,
		_w12570_,
		_w12571_,
		_w12572_,
		_w12573_
	);
	LUT4 #(
		.INIT('ha820)
	) name8526 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001 ,
		_w12574_
	);
	LUT3 #(
		.INIT('h07)
	) name8527 (
		_w11508_,
		_w11455_,
		_w12574_,
		_w12575_
	);
	LUT2 #(
		.INIT('h8)
	) name8528 (
		_w11488_,
		_w11462_,
		_w12576_
	);
	LUT3 #(
		.INIT('h80)
	) name8529 (
		_w11389_,
		_w11491_,
		_w11450_,
		_w12577_
	);
	LUT3 #(
		.INIT('h10)
	) name8530 (
		_w12576_,
		_w12577_,
		_w12575_,
		_w12578_
	);
	LUT2 #(
		.INIT('h1)
	) name8531 (
		_w11553_,
		_w11885_,
		_w12579_
	);
	LUT4 #(
		.INIT('hf040)
	) name8532 (
		_w11444_,
		_w11428_,
		_w11511_,
		_w11455_,
		_w12580_
	);
	LUT3 #(
		.INIT('h01)
	) name8533 (
		_w11575_,
		_w11576_,
		_w12580_,
		_w12581_
	);
	LUT3 #(
		.INIT('h80)
	) name8534 (
		_w12578_,
		_w12579_,
		_w12581_,
		_w12582_
	);
	LUT3 #(
		.INIT('h40)
	) name8535 (
		_w11444_,
		_w11428_,
		_w11508_,
		_w12583_
	);
	LUT3 #(
		.INIT('h40)
	) name8536 (
		_w11444_,
		_w11423_,
		_w11488_,
		_w12584_
	);
	LUT3 #(
		.INIT('h40)
	) name8537 (
		_w11444_,
		_w11392_,
		_w11450_,
		_w12585_
	);
	LUT3 #(
		.INIT('h01)
	) name8538 (
		_w12584_,
		_w12585_,
		_w12583_,
		_w12586_
	);
	LUT2 #(
		.INIT('h8)
	) name8539 (
		_w11903_,
		_w12586_,
		_w12587_
	);
	LUT4 #(
		.INIT('h8000)
	) name8540 (
		_w12582_,
		_w12587_,
		_w12573_,
		_w12567_,
		_w12588_
	);
	LUT4 #(
		.INIT('h0002)
	) name8541 (
		_w11568_,
		_w11570_,
		_w11582_,
		_w11832_,
		_w12589_
	);
	LUT3 #(
		.INIT('hd0)
	) name8542 (
		_w11341_,
		_w11398_,
		_w11479_,
		_w12590_
	);
	LUT2 #(
		.INIT('h8)
	) name8543 (
		_w12589_,
		_w12590_,
		_w12591_
	);
	LUT3 #(
		.INIT('h04)
	) name8544 (
		_w11549_,
		_w11441_,
		_w11869_,
		_w12592_
	);
	LUT4 #(
		.INIT('h0057)
	) name8545 (
		_w11341_,
		_w11419_,
		_w11425_,
		_w11430_,
		_w12593_
	);
	LUT2 #(
		.INIT('h8)
	) name8546 (
		_w11408_,
		_w12593_,
		_w12594_
	);
	LUT3 #(
		.INIT('ha8)
	) name8547 (
		_w11532_,
		_w11435_,
		_w12455_,
		_w12595_
	);
	LUT3 #(
		.INIT('ha8)
	) name8548 (
		_w11537_,
		_w11588_,
		_w12496_,
		_w12596_
	);
	LUT3 #(
		.INIT('ha8)
	) name8549 (
		_w11341_,
		_w11409_,
		_w11896_,
		_w12597_
	);
	LUT3 #(
		.INIT('h01)
	) name8550 (
		_w12596_,
		_w12597_,
		_w12595_,
		_w12598_
	);
	LUT3 #(
		.INIT('h80)
	) name8551 (
		_w12594_,
		_w12592_,
		_w12598_,
		_w12599_
	);
	LUT4 #(
		.INIT('h8000)
	) name8552 (
		_w11911_,
		_w12591_,
		_w12599_,
		_w12588_,
		_w12600_
	);
	LUT4 #(
		.INIT('h4c08)
	) name8553 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11830_,
		_w12562_,
		_w12600_,
		_w12601_
	);
	LUT4 #(
		.INIT('h5545)
	) name8554 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w12602_
	);
	LUT2 #(
		.INIT('h1)
	) name8555 (
		_w12601_,
		_w12602_,
		_w12603_
	);
	LUT2 #(
		.INIT('h8)
	) name8556 (
		\bdma_BWcnt_reg[0]/NET0131 ,
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w12604_
	);
	LUT4 #(
		.INIT('h4000)
	) name8557 (
		\bdma_BSreq_reg/NET0131 ,
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w4764_,
		_w12604_,
		_w12605_
	);
	LUT3 #(
		.INIT('h6c)
	) name8558 (
		\bdma_BWcnt_reg[3]/NET0131 ,
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w12605_,
		_w12606_
	);
	LUT2 #(
		.INIT('h4)
	) name8559 (
		_w9413_,
		_w12606_,
		_w12607_
	);
	LUT4 #(
		.INIT('hf600)
	) name8560 (
		_w9480_,
		_w9725_,
		_w9732_,
		_w9759_,
		_w12608_
	);
	LUT4 #(
		.INIT('h9f96)
	) name8561 (
		_w9480_,
		_w9725_,
		_w9732_,
		_w9757_,
		_w12609_
	);
	LUT2 #(
		.INIT('h4)
	) name8562 (
		_w12608_,
		_w12609_,
		_w12610_
	);
	LUT3 #(
		.INIT('h1e)
	) name8563 (
		_w9456_,
		_w9715_,
		_w12610_,
		_w12611_
	);
	LUT4 #(
		.INIT('h10b0)
	) name8564 (
		_w9455_,
		_w9768_,
		_w9895_,
		_w12611_,
		_w12612_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8565 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001 ,
		_w9451_,
		_w9453_,
		_w9894_,
		_w12613_
	);
	LUT2 #(
		.INIT('he)
	) name8566 (
		_w12612_,
		_w12613_,
		_w12614_
	);
	LUT4 #(
		.INIT('h028a)
	) name8567 (
		_w9454_,
		_w9455_,
		_w9768_,
		_w12611_,
		_w12615_
	);
	LUT2 #(
		.INIT('h2)
	) name8568 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001 ,
		_w9454_,
		_w12616_
	);
	LUT2 #(
		.INIT('he)
	) name8569 (
		_w12615_,
		_w12616_,
		_w12617_
	);
	LUT3 #(
		.INIT('h08)
	) name8570 (
		\idma_IADi_reg[15]/P0001 ,
		\idma_IAL_reg/P0001 ,
		\idma_ISn_reg/P0001 ,
		_w12618_
	);
	LUT4 #(
		.INIT('h007f)
	) name8571 (
		_w5804_,
		_w9431_,
		_w11604_,
		_w12618_,
		_w12619_
	);
	LUT3 #(
		.INIT('h04)
	) name8572 (
		\idma_IADi_reg[15]/P0001 ,
		\idma_IAL_reg/P0001 ,
		\idma_ISn_reg/P0001 ,
		_w12620_
	);
	LUT2 #(
		.INIT('h1)
	) name8573 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w12621_
	);
	LUT4 #(
		.INIT('h0001)
	) name8574 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w12622_
	);
	LUT4 #(
		.INIT('h070f)
	) name8575 (
		_w5658_,
		_w9431_,
		_w12620_,
		_w12622_,
		_w12623_
	);
	LUT4 #(
		.INIT('h3363)
	) name8576 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PCrd_1st_reg/NET0131 ,
		\idma_RDCMD_d1_reg/P0001 ,
		\idma_RDCMD_reg/P0001 ,
		_w12624_
	);
	LUT3 #(
		.INIT('h7f)
	) name8577 (
		_w12619_,
		_w12623_,
		_w12624_,
		_w12625_
	);
	LUT4 #(
		.INIT('h4544)
	) name8578 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w7257_,
		_w7375_,
		_w7377_,
		_w12626_
	);
	LUT2 #(
		.INIT('h2)
	) name8579 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8907_,
		_w12627_
	);
	LUT2 #(
		.INIT('h1)
	) name8580 (
		_w12626_,
		_w12627_,
		_w12628_
	);
	LUT4 #(
		.INIT('h0200)
	) name8581 (
		_w11577_,
		_w11907_,
		_w11908_,
		_w11909_,
		_w12629_
	);
	LUT2 #(
		.INIT('h8)
	) name8582 (
		_w11871_,
		_w12629_,
		_w12630_
	);
	LUT2 #(
		.INIT('h1)
	) name8583 (
		_w11530_,
		_w11950_,
		_w12631_
	);
	LUT4 #(
		.INIT('h153f)
	) name8584 (
		_w11555_,
		_w11558_,
		_w11458_,
		_w11874_,
		_w12632_
	);
	LUT2 #(
		.INIT('h4)
	) name8585 (
		_w12631_,
		_w12632_,
		_w12633_
	);
	LUT2 #(
		.INIT('h8)
	) name8586 (
		_w11537_,
		_w11409_,
		_w12634_
	);
	LUT3 #(
		.INIT('h80)
	) name8587 (
		_w11389_,
		_w11476_,
		_w12505_,
		_w12635_
	);
	LUT3 #(
		.INIT('h08)
	) name8588 (
		_w11389_,
		_w11491_,
		_w11844_,
		_w12636_
	);
	LUT4 #(
		.INIT('h153f)
	) name8589 (
		_w11415_,
		_w11455_,
		_w11864_,
		_w11848_,
		_w12637_
	);
	LUT3 #(
		.INIT('h10)
	) name8590 (
		_w12635_,
		_w12636_,
		_w12637_,
		_w12638_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name8591 (
		_w11333_,
		_w11385_,
		_w11506_,
		_w11452_,
		_w12639_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name8592 (
		_w11534_,
		_w11522_,
		_w11464_,
		_w12639_,
		_w12640_
	);
	LUT3 #(
		.INIT('h40)
	) name8593 (
		_w12634_,
		_w12638_,
		_w12640_,
		_w12641_
	);
	LUT2 #(
		.INIT('h1)
	) name8594 (
		_w11407_,
		_w11967_,
		_w12642_
	);
	LUT4 #(
		.INIT('h0001)
	) name8595 (
		_w11407_,
		_w11436_,
		_w11885_,
		_w11967_,
		_w12643_
	);
	LUT2 #(
		.INIT('h8)
	) name8596 (
		_w12571_,
		_w12643_,
		_w12644_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name8597 (
		_w11333_,
		_w11341_,
		_w11394_,
		_w11397_,
		_w12645_
	);
	LUT3 #(
		.INIT('h08)
	) name8598 (
		_w12571_,
		_w12643_,
		_w12645_,
		_w12646_
	);
	LUT3 #(
		.INIT('h80)
	) name8599 (
		_w12633_,
		_w12641_,
		_w12646_,
		_w12647_
	);
	LUT3 #(
		.INIT('h02)
	) name8600 (
		_w11386_,
		_w11335_,
		_w11953_,
		_w12648_
	);
	LUT3 #(
		.INIT('h01)
	) name8601 (
		_w11550_,
		_w11551_,
		_w12446_,
		_w12649_
	);
	LUT3 #(
		.INIT('hc8)
	) name8602 (
		_w11435_,
		_w11860_,
		_w12455_,
		_w12650_
	);
	LUT3 #(
		.INIT('ha8)
	) name8603 (
		_w11854_,
		_w11973_,
		_w11974_,
		_w12651_
	);
	LUT4 #(
		.INIT('h0004)
	) name8604 (
		_w12648_,
		_w12649_,
		_w12650_,
		_w12651_,
		_w12652_
	);
	LUT4 #(
		.INIT('h4000)
	) name8605 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11382_,
		_w11406_,
		_w12653_
	);
	LUT3 #(
		.INIT('h40)
	) name8606 (
		_w11385_,
		_w11415_,
		_w11874_,
		_w12654_
	);
	LUT3 #(
		.INIT('h40)
	) name8607 (
		_w11444_,
		_w11428_,
		_w11864_,
		_w12655_
	);
	LUT3 #(
		.INIT('h40)
	) name8608 (
		_w11536_,
		_w11386_,
		_w11578_,
		_w12656_
	);
	LUT4 #(
		.INIT('h0001)
	) name8609 (
		_w12653_,
		_w12654_,
		_w12655_,
		_w12656_,
		_w12657_
	);
	LUT4 #(
		.INIT('ha820)
	) name8610 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001 ,
		_w12658_
	);
	LUT4 #(
		.INIT('h007f)
	) name8611 (
		_w11473_,
		_w11389_,
		_w11341_,
		_w12658_,
		_w12659_
	);
	LUT3 #(
		.INIT('h04)
	) name8612 (
		_w11444_,
		_w11392_,
		_w11844_,
		_w12660_
	);
	LUT4 #(
		.INIT('h0100)
	) name8613 (
		_w11403_,
		_w11553_,
		_w12660_,
		_w12659_,
		_w12661_
	);
	LUT3 #(
		.INIT('hc8)
	) name8614 (
		_w11588_,
		_w11499_,
		_w12496_,
		_w12662_
	);
	LUT3 #(
		.INIT('hc8)
	) name8615 (
		_w11587_,
		_w11495_,
		_w11880_,
		_w12663_
	);
	LUT4 #(
		.INIT('h1000)
	) name8616 (
		_w12662_,
		_w12663_,
		_w12657_,
		_w12661_,
		_w12664_
	);
	LUT2 #(
		.INIT('h8)
	) name8617 (
		_w12652_,
		_w12664_,
		_w12665_
	);
	LUT3 #(
		.INIT('h10)
	) name8618 (
		_w11549_,
		_w11595_,
		_w11441_,
		_w12666_
	);
	LUT2 #(
		.INIT('h8)
	) name8619 (
		_w12589_,
		_w12666_,
		_w12667_
	);
	LUT4 #(
		.INIT('h8000)
	) name8620 (
		_w12630_,
		_w12647_,
		_w12665_,
		_w12667_,
		_w12668_
	);
	LUT4 #(
		.INIT('h4c08)
	) name8621 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11830_,
		_w12628_,
		_w12668_,
		_w12669_
	);
	LUT4 #(
		.INIT('h5545)
	) name8622 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w12670_
	);
	LUT2 #(
		.INIT('h1)
	) name8623 (
		_w12669_,
		_w12670_,
		_w12671_
	);
	LUT2 #(
		.INIT('h2)
	) name8624 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8781_,
		_w12672_
	);
	LUT4 #(
		.INIT('h00ab)
	) name8625 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8757_,
		_w8760_,
		_w12672_,
		_w12673_
	);
	LUT4 #(
		.INIT('ha820)
	) name8626 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001 ,
		_w12674_
	);
	LUT4 #(
		.INIT('h007f)
	) name8627 (
		_w11389_,
		_w11491_,
		_w11962_,
		_w12674_,
		_w12675_
	);
	LUT3 #(
		.INIT('hb0)
	) name8628 (
		_w11534_,
		_w11855_,
		_w12675_,
		_w12676_
	);
	LUT4 #(
		.INIT('haf8c)
	) name8629 (
		_w11504_,
		_w11446_,
		_w11873_,
		_w11950_,
		_w12677_
	);
	LUT3 #(
		.INIT('h02)
	) name8630 (
		_w11386_,
		_w11335_,
		_w11530_,
		_w12678_
	);
	LUT4 #(
		.INIT('h2000)
	) name8631 (
		_w11580_,
		_w12678_,
		_w12676_,
		_w12677_,
		_w12679_
	);
	LUT4 #(
		.INIT('h000e)
	) name8632 (
		_w11386_,
		_w11530_,
		_w11522_,
		_w11524_,
		_w12680_
	);
	LUT4 #(
		.INIT('h00f4)
	) name8633 (
		_w11444_,
		_w11414_,
		_w11481_,
		_w11844_,
		_w12681_
	);
	LUT4 #(
		.INIT('hf400)
	) name8634 (
		_w11444_,
		_w11428_,
		_w11455_,
		_w12504_,
		_w12682_
	);
	LUT4 #(
		.INIT('h000b)
	) name8635 (
		_w11492_,
		_w11861_,
		_w12681_,
		_w12682_,
		_w12683_
	);
	LUT3 #(
		.INIT('hd0)
	) name8636 (
		_w11341_,
		_w12680_,
		_w12683_,
		_w12684_
	);
	LUT4 #(
		.INIT('h8000)
	) name8637 (
		_w11417_,
		_w11432_,
		_w12679_,
		_w12684_,
		_w12685_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name8638 (
		_w11444_,
		_w11386_,
		_w11392_,
		_w11494_,
		_w12686_
	);
	LUT3 #(
		.INIT('he0)
	) name8639 (
		_w11534_,
		_w11536_,
		_w12686_,
		_w12687_
	);
	LUT4 #(
		.INIT('h00f4)
	) name8640 (
		_w11444_,
		_w11423_,
		_w11462_,
		_w11464_,
		_w12688_
	);
	LUT4 #(
		.INIT('h00f4)
	) name8641 (
		_w11444_,
		_w11428_,
		_w11455_,
		_w11457_,
		_w12689_
	);
	LUT4 #(
		.INIT('h000e)
	) name8642 (
		_w11504_,
		_w11506_,
		_w12689_,
		_w12688_,
		_w12690_
	);
	LUT4 #(
		.INIT('hf040)
	) name8643 (
		_w11444_,
		_w11405_,
		_w11863_,
		_w12401_,
		_w12691_
	);
	LUT3 #(
		.INIT('h01)
	) name8644 (
		_w11386_,
		_w12404_,
		_w12691_,
		_w12692_
	);
	LUT3 #(
		.INIT('h07)
	) name8645 (
		_w12687_,
		_w12690_,
		_w12692_,
		_w12693_
	);
	LUT2 #(
		.INIT('h2)
	) name8646 (
		_w11596_,
		_w12693_,
		_w12694_
	);
	LUT2 #(
		.INIT('h8)
	) name8647 (
		_w11442_,
		_w12590_,
		_w12695_
	);
	LUT4 #(
		.INIT('h8000)
	) name8648 (
		_w12434_,
		_w12695_,
		_w12685_,
		_w12694_,
		_w12696_
	);
	LUT4 #(
		.INIT('h4c08)
	) name8649 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11830_,
		_w12673_,
		_w12696_,
		_w12697_
	);
	LUT4 #(
		.INIT('h5545)
	) name8650 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w12698_
	);
	LUT2 #(
		.INIT('h1)
	) name8651 (
		_w12697_,
		_w12698_,
		_w12699_
	);
	LUT4 #(
		.INIT('h4c08)
	) name8652 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11329_,
		_w12562_,
		_w12600_,
		_w12700_
	);
	LUT2 #(
		.INIT('h1)
	) name8653 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001 ,
		_w11329_,
		_w12701_
	);
	LUT2 #(
		.INIT('h1)
	) name8654 (
		_w12700_,
		_w12701_,
		_w12702_
	);
	LUT4 #(
		.INIT('h0400)
	) name8655 (
		_w4747_,
		_w4768_,
		_w4781_,
		_w4796_,
		_w12703_
	);
	LUT3 #(
		.INIT('h10)
	) name8656 (
		_w4785_,
		_w4787_,
		_w12703_,
		_w12704_
	);
	LUT3 #(
		.INIT('h20)
	) name8657 (
		_w4787_,
		_w8595_,
		_w12703_,
		_w12705_
	);
	LUT4 #(
		.INIT('h4144)
	) name8658 (
		_w4750_,
		_w4781_,
		_w4784_,
		_w4786_,
		_w12706_
	);
	LUT4 #(
		.INIT('hb000)
	) name8659 (
		_w4747_,
		_w4768_,
		_w4796_,
		_w12706_,
		_w12707_
	);
	LUT2 #(
		.INIT('h1)
	) name8660 (
		_w9413_,
		_w12707_,
		_w12708_
	);
	LUT4 #(
		.INIT('hf8dd)
	) name8661 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w12709_
	);
	LUT4 #(
		.INIT('h0080)
	) name8662 (
		\emc_RWcnt_reg[0]/P0001 ,
		\emc_RWcnt_reg[1]/P0001 ,
		\emc_RWcnt_reg[2]/P0001 ,
		_w12709_,
		_w12710_
	);
	LUT4 #(
		.INIT('h78f0)
	) name8663 (
		\emc_RWcnt_reg[3]/P0001 ,
		\emc_RWcnt_reg[4]/P0001 ,
		\emc_RWcnt_reg[5]/P0001 ,
		_w12710_,
		_w12711_
	);
	LUT4 #(
		.INIT('h1000)
	) name8664 (
		_w12705_,
		_w12704_,
		_w12708_,
		_w12711_,
		_w12712_
	);
	LUT3 #(
		.INIT('h6c)
	) name8665 (
		\emc_RWcnt_reg[3]/P0001 ,
		\emc_RWcnt_reg[4]/P0001 ,
		_w12710_,
		_w12713_
	);
	LUT4 #(
		.INIT('h1000)
	) name8666 (
		_w12705_,
		_w12704_,
		_w12708_,
		_w12713_,
		_w12714_
	);
	LUT4 #(
		.INIT('h4c08)
	) name8667 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11329_,
		_w12628_,
		_w12668_,
		_w12715_
	);
	LUT2 #(
		.INIT('h1)
	) name8668 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001 ,
		_w11329_,
		_w12716_
	);
	LUT2 #(
		.INIT('h1)
	) name8669 (
		_w12715_,
		_w12716_,
		_w12717_
	);
	LUT4 #(
		.INIT('h4c08)
	) name8670 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11329_,
		_w12673_,
		_w12696_,
		_w12718_
	);
	LUT2 #(
		.INIT('h1)
	) name8671 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001 ,
		_w11329_,
		_w12719_
	);
	LUT2 #(
		.INIT('h1)
	) name8672 (
		_w12718_,
		_w12719_,
		_w12720_
	);
	LUT4 #(
		.INIT('h8000)
	) name8673 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		_w12721_
	);
	LUT4 #(
		.INIT('h8000)
	) name8674 (
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		_w12721_,
		_w12722_
	);
	LUT2 #(
		.INIT('h8)
	) name8675 (
		\sport1_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		_w12722_,
		_w12723_
	);
	LUT3 #(
		.INIT('h80)
	) name8676 (
		\sport1_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		_w12722_,
		_w12724_
	);
	LUT4 #(
		.INIT('h8000)
	) name8677 (
		\sport1_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		_w12722_,
		_w12725_
	);
	LUT4 #(
		.INIT('h0408)
	) name8678 (
		\sport1_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12724_,
		_w12726_
	);
	LUT3 #(
		.INIT('h6c)
	) name8679 (
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		_w12721_,
		_w12727_
	);
	LUT3 #(
		.INIT('h20)
	) name8680 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12727_,
		_w12728_
	);
	LUT3 #(
		.INIT('h78)
	) name8681 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		_w12729_
	);
	LUT3 #(
		.INIT('h20)
	) name8682 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12729_,
		_w12730_
	);
	LUT2 #(
		.INIT('h8)
	) name8683 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		_w12725_,
		_w12731_
	);
	LUT3 #(
		.INIT('h80)
	) name8684 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		_w12725_,
		_w12732_
	);
	LUT4 #(
		.INIT('h8000)
	) name8685 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		_w12725_,
		_w12733_
	);
	LUT3 #(
		.INIT('h48)
	) name8686 (
		\sport1_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		_w12087_,
		_w12733_,
		_w12734_
	);
	LUT3 #(
		.INIT('h04)
	) name8687 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12735_
	);
	LUT4 #(
		.INIT('h4544)
	) name8688 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w7592_,
		_w7707_,
		_w7709_,
		_w12736_
	);
	LUT2 #(
		.INIT('h2)
	) name8689 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8929_,
		_w12737_
	);
	LUT2 #(
		.INIT('h1)
	) name8690 (
		_w12736_,
		_w12737_,
		_w12738_
	);
	LUT3 #(
		.INIT('ha8)
	) name8691 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12736_,
		_w12737_,
		_w12739_
	);
	LUT2 #(
		.INIT('h8)
	) name8692 (
		_w11834_,
		_w11970_,
		_w12740_
	);
	LUT3 #(
		.INIT('h02)
	) name8693 (
		_w11386_,
		_w11540_,
		_w11954_,
		_w12741_
	);
	LUT3 #(
		.INIT('he0)
	) name8694 (
		_w11420_,
		_w11421_,
		_w11874_,
		_w12742_
	);
	LUT3 #(
		.INIT('hc8)
	) name8695 (
		_w11547_,
		_w11458_,
		_w11976_,
		_w12743_
	);
	LUT3 #(
		.INIT('h01)
	) name8696 (
		_w12742_,
		_w12743_,
		_w12741_,
		_w12744_
	);
	LUT3 #(
		.INIT('h0e)
	) name8697 (
		_w11393_,
		_w11589_,
		_w11512_,
		_w12745_
	);
	LUT4 #(
		.INIT('h7770)
	) name8698 (
		_w11424_,
		_w11532_,
		_w11489_,
		_w11953_,
		_w12746_
	);
	LUT2 #(
		.INIT('h4)
	) name8699 (
		_w12745_,
		_w12746_,
		_w12747_
	);
	LUT3 #(
		.INIT('h32)
	) name8700 (
		_w11552_,
		_w11454_,
		_w11474_,
		_w12748_
	);
	LUT2 #(
		.INIT('h2)
	) name8701 (
		_w11538_,
		_w11954_,
		_w12749_
	);
	LUT4 #(
		.INIT('heee0)
	) name8702 (
		_w11592_,
		_w11501_,
		_w11471_,
		_w11957_,
		_w12750_
	);
	LUT3 #(
		.INIT('h10)
	) name8703 (
		_w12748_,
		_w12749_,
		_w12750_,
		_w12751_
	);
	LUT3 #(
		.INIT('he0)
	) name8704 (
		_w11397_,
		_w11519_,
		_w11854_,
		_w12752_
	);
	LUT4 #(
		.INIT('ha820)
	) name8705 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001 ,
		_w12753_
	);
	LUT4 #(
		.INIT('h8000)
	) name8706 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11382_,
		_w11406_,
		_w12754_
	);
	LUT4 #(
		.INIT('h000d)
	) name8707 (
		_w11402_,
		_w11593_,
		_w12753_,
		_w12754_,
		_w12755_
	);
	LUT2 #(
		.INIT('h4)
	) name8708 (
		_w12752_,
		_w12755_,
		_w12756_
	);
	LUT4 #(
		.INIT('h8000)
	) name8709 (
		_w12747_,
		_w12751_,
		_w12756_,
		_w12744_,
		_w12757_
	);
	LUT4 #(
		.INIT('h2333)
	) name8710 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12739_,
		_w12740_,
		_w12757_,
		_w12758_
	);
	LUT3 #(
		.INIT('he2)
	) name8711 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001 ,
		_w11946_,
		_w12758_,
		_w12759_
	);
	LUT3 #(
		.INIT('hc8)
	) name8712 (
		_w11557_,
		_w11854_,
		_w12018_,
		_w12760_
	);
	LUT3 #(
		.INIT('ha8)
	) name8713 (
		_w11537_,
		_w11572_,
		_w11831_,
		_w12761_
	);
	LUT3 #(
		.INIT('he0)
	) name8714 (
		_w11397_,
		_w11519_,
		_w11458_,
		_w12762_
	);
	LUT3 #(
		.INIT('he0)
	) name8715 (
		_w11420_,
		_w11421_,
		_w11507_,
		_w12763_
	);
	LUT4 #(
		.INIT('h0001)
	) name8716 (
		_w12760_,
		_w12761_,
		_w12762_,
		_w12763_,
		_w12764_
	);
	LUT4 #(
		.INIT('h7707)
	) name8717 (
		_w11424_,
		_w11499_,
		_w11848_,
		_w11954_,
		_w12765_
	);
	LUT3 #(
		.INIT('he0)
	) name8718 (
		_w11552_,
		_w11474_,
		_w11864_,
		_w12766_
	);
	LUT3 #(
		.INIT('h08)
	) name8719 (
		_w11333_,
		_w11385_,
		_w11335_,
		_w12767_
	);
	LUT3 #(
		.INIT('h0b)
	) name8720 (
		_w11385_,
		_w11341_,
		_w12767_,
		_w12768_
	);
	LUT4 #(
		.INIT('h1bff)
	) name8721 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11473_,
		_w11401_,
		_w11358_,
		_w12769_
	);
	LUT2 #(
		.INIT('h1)
	) name8722 (
		_w12768_,
		_w12769_,
		_w12770_
	);
	LUT3 #(
		.INIT('h10)
	) name8723 (
		_w12766_,
		_w12770_,
		_w12765_,
		_w12771_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name8724 (
		_w11593_,
		_w11875_,
		_w11954_,
		_w12500_,
		_w12772_
	);
	LUT4 #(
		.INIT('hfca8)
	) name8725 (
		_w11592_,
		_w11844_,
		_w11957_,
		_w11950_,
		_w12773_
	);
	LUT2 #(
		.INIT('h8)
	) name8726 (
		_w12772_,
		_w12773_,
		_w12774_
	);
	LUT3 #(
		.INIT('hc8)
	) name8727 (
		_w11547_,
		_w11872_,
		_w11976_,
		_w12775_
	);
	LUT4 #(
		.INIT('ha820)
	) name8728 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001 ,
		_w12776_
	);
	LUT2 #(
		.INIT('h1)
	) name8729 (
		_w11967_,
		_w12776_,
		_w12777_
	);
	LUT3 #(
		.INIT('h20)
	) name8730 (
		_w11569_,
		_w12775_,
		_w12777_,
		_w12778_
	);
	LUT4 #(
		.INIT('h8000)
	) name8731 (
		_w12771_,
		_w12774_,
		_w12778_,
		_w12764_,
		_w12779_
	);
	LUT4 #(
		.INIT('h4c08)
	) name8732 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w11946_,
		_w12317_,
		_w12779_,
		_w12780_
	);
	LUT4 #(
		.INIT('h5545)
	) name8733 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001 ,
		_w9453_,
		_w9894_,
		_w11945_,
		_w12781_
	);
	LUT2 #(
		.INIT('h1)
	) name8734 (
		_w12780_,
		_w12781_,
		_w12782_
	);
	LUT3 #(
		.INIT('he2)
	) name8735 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001 ,
		_w12048_,
		_w12758_,
		_w12783_
	);
	LUT4 #(
		.INIT('h4c08)
	) name8736 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12048_,
		_w12317_,
		_w12779_,
		_w12784_
	);
	LUT2 #(
		.INIT('h1)
	) name8737 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001 ,
		_w12048_,
		_w12785_
	);
	LUT2 #(
		.INIT('h1)
	) name8738 (
		_w12784_,
		_w12785_,
		_w12786_
	);
	LUT4 #(
		.INIT('h0408)
	) name8739 (
		\sport0_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12308_,
		_w12787_
	);
	LUT2 #(
		.INIT('h8)
	) name8740 (
		\emc_PMcst_reg/NET0131 ,
		_w9936_,
		_w12788_
	);
	LUT4 #(
		.INIT('ha820)
	) name8741 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		_w12789_
	);
	LUT3 #(
		.INIT('h80)
	) name8742 (
		\memc_Pread_E_reg/NET0131 ,
		_w12051_,
		_w12789_,
		_w12790_
	);
	LUT3 #(
		.INIT('h13)
	) name8743 (
		_w12057_,
		_w12788_,
		_w12790_,
		_w12791_
	);
	LUT3 #(
		.INIT('h80)
	) name8744 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12051_,
		_w12789_,
		_w12792_
	);
	LUT3 #(
		.INIT('h02)
	) name8745 (
		\emc_PMcst_reg/NET0131 ,
		_w4794_,
		_w4804_,
		_w12793_
	);
	LUT3 #(
		.INIT('h27)
	) name8746 (
		_w12057_,
		_w12792_,
		_w12793_,
		_w12794_
	);
	LUT2 #(
		.INIT('h7)
	) name8747 (
		_w12791_,
		_w12794_,
		_w12795_
	);
	LUT3 #(
		.INIT('h01)
	) name8748 (
		\tm_TCR_TMP_reg[1]/NET0131 ,
		\tm_TCR_TMP_reg[2]/NET0131 ,
		\tm_TCR_TMP_reg[3]/NET0131 ,
		_w12796_
	);
	LUT4 #(
		.INIT('h0001)
	) name8749 (
		\tm_TCR_TMP_reg[0]/NET0131 ,
		\tm_TCR_TMP_reg[1]/NET0131 ,
		\tm_TCR_TMP_reg[2]/NET0131 ,
		\tm_TCR_TMP_reg[3]/NET0131 ,
		_w12797_
	);
	LUT4 #(
		.INIT('h0001)
	) name8750 (
		\tm_TCR_TMP_reg[4]/NET0131 ,
		\tm_TCR_TMP_reg[5]/NET0131 ,
		\tm_TCR_TMP_reg[6]/NET0131 ,
		\tm_TCR_TMP_reg[7]/NET0131 ,
		_w12798_
	);
	LUT4 #(
		.INIT('h0001)
	) name8751 (
		\tm_TCR_TMP_reg[14]/NET0131 ,
		\tm_TCR_TMP_reg[15]/NET0131 ,
		\tm_TCR_TMP_reg[8]/NET0131 ,
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w12799_
	);
	LUT4 #(
		.INIT('h0001)
	) name8752 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		\tm_TCR_TMP_reg[11]/NET0131 ,
		\tm_TCR_TMP_reg[12]/NET0131 ,
		\tm_TCR_TMP_reg[13]/NET0131 ,
		_w12800_
	);
	LUT4 #(
		.INIT('h8000)
	) name8753 (
		_w12797_,
		_w12798_,
		_w12799_,
		_w12800_,
		_w12801_
	);
	LUT3 #(
		.INIT('h04)
	) name8754 (
		\T_TMODE[0]_pad ,
		\tm_WR_TSR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TSR_TMP_GEN2_reg/P0001 ,
		_w12802_
	);
	LUT3 #(
		.INIT('h04)
	) name8755 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		_w12803_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name8756 (
		\T_TMODE[0]_pad ,
		\tm_MSTAT5_syn_reg/NET0131 ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		_w12804_
	);
	LUT2 #(
		.INIT('h4)
	) name8757 (
		_w12802_,
		_w12804_,
		_w12805_
	);
	LUT2 #(
		.INIT('h8)
	) name8758 (
		_w12801_,
		_w12805_,
		_w12806_
	);
	LUT2 #(
		.INIT('h8)
	) name8759 (
		\core_c_dec_updAF_E_reg/P0001 ,
		_w4106_,
		_w12807_
	);
	LUT4 #(
		.INIT('h0400)
	) name8760 (
		_w4094_,
		_w4097_,
		_w4101_,
		_w11927_,
		_w12808_
	);
	LUT3 #(
		.INIT('h20)
	) name8761 (
		_w4834_,
		_w11921_,
		_w12808_,
		_w12809_
	);
	LUT2 #(
		.INIT('he)
	) name8762 (
		_w12807_,
		_w12809_,
		_w12810_
	);
	LUT2 #(
		.INIT('h1)
	) name8763 (
		\idma_WRcnt_reg[0]/NET0131 ,
		\idma_WRcnt_reg[1]/NET0131 ,
		_w12811_
	);
	LUT3 #(
		.INIT('h01)
	) name8764 (
		\idma_WRcnt_reg[0]/NET0131 ,
		\idma_WRcnt_reg[1]/NET0131 ,
		\idma_WRcnt_reg[2]/NET0131 ,
		_w12812_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8765 (
		\idma_WRcnt_reg[0]/NET0131 ,
		\idma_WRcnt_reg[1]/NET0131 ,
		\idma_WRcnt_reg[2]/NET0131 ,
		\idma_WRtrue_reg/NET0131 ,
		_w12813_
	);
	LUT2 #(
		.INIT('h4)
	) name8766 (
		\idma_WRCMD_d1_reg/P0001 ,
		\idma_WRCMD_reg/P0001 ,
		_w12814_
	);
	LUT2 #(
		.INIT('he)
	) name8767 (
		_w12813_,
		_w12814_,
		_w12815_
	);
	LUT2 #(
		.INIT('h1)
	) name8768 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12816_
	);
	LUT3 #(
		.INIT('h10)
	) name8769 (
		\idma_ISn_reg/P0001 ,
		\idma_IWRn_reg/P0001 ,
		\idma_WRtrue_reg/NET0131 ,
		_w12817_
	);
	LUT3 #(
		.INIT('ha8)
	) name8770 (
		\auctl_DSack_reg/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12818_
	);
	LUT2 #(
		.INIT('h1)
	) name8771 (
		\idma_RDcnt_reg[0]/NET0131 ,
		\idma_RDcnt_reg[1]/NET0131 ,
		_w12819_
	);
	LUT3 #(
		.INIT('h01)
	) name8772 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		\idma_RDcnt_reg[2]/NET0131 ,
		_w12820_
	);
	LUT4 #(
		.INIT('ha888)
	) name8773 (
		\idma_RDcyc_reg/NET0131 ,
		_w12818_,
		_w12819_,
		_w12820_,
		_w12821_
	);
	LUT3 #(
		.INIT('h54)
	) name8774 (
		_w12816_,
		_w12817_,
		_w12821_,
		_w12822_
	);
	LUT3 #(
		.INIT('hca)
	) name8775 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 ,
		_w11922_,
		_w11926_,
		_w12823_
	);
	LUT4 #(
		.INIT('h0008)
	) name8776 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w12824_
	);
	LUT3 #(
		.INIT('h80)
	) name8777 (
		_w9431_,
		_w11604_,
		_w12824_,
		_w12825_
	);
	LUT4 #(
		.INIT('h4000)
	) name8778 (
		\memc_MMR_web_reg/NET0131 ,
		_w9431_,
		_w11604_,
		_w12824_,
		_w12826_
	);
	LUT4 #(
		.INIT('h03aa)
	) name8779 (
		\sport0_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w7140_,
		_w7240_,
		_w12826_,
		_w12827_
	);
	LUT3 #(
		.INIT('h01)
	) name8780 (
		\sport1_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[5]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[6]/NET0131 ,
		_w12828_
	);
	LUT4 #(
		.INIT('h0001)
	) name8781 (
		\sport1_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[5]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[6]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[7]/NET0131 ,
		_w12829_
	);
	LUT4 #(
		.INIT('h0800)
	) name8782 (
		\sport1_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[1]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[2]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		_w12830_
	);
	LUT4 #(
		.INIT('h0002)
	) name8783 (
		\sport1_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[2]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[3]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[4]/NET0131 ,
		_w12831_
	);
	LUT4 #(
		.INIT('h4000)
	) name8784 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		_w12829_,
		_w12830_,
		_w12831_,
		_w12832_
	);
	LUT4 #(
		.INIT('h1d00)
	) name8785 (
		\T_RD1_pad ,
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w9403_,
		_w12832_,
		_w12833_
	);
	LUT2 #(
		.INIT('h1)
	) name8786 (
		\sport1_rxctl_SLOT1_EXT_reg[2]/NET0131 ,
		_w12832_,
		_w12834_
	);
	LUT2 #(
		.INIT('h1)
	) name8787 (
		_w12833_,
		_w12834_,
		_w12835_
	);
	LUT4 #(
		.INIT('h8000)
	) name8788 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		_w12829_,
		_w12830_,
		_w12831_,
		_w12836_
	);
	LUT4 #(
		.INIT('h1d00)
	) name8789 (
		\T_RD1_pad ,
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w9403_,
		_w12836_,
		_w12837_
	);
	LUT2 #(
		.INIT('h1)
	) name8790 (
		\sport1_rxctl_SLOT1_EXT_reg[3]/NET0131 ,
		_w12836_,
		_w12838_
	);
	LUT2 #(
		.INIT('h1)
	) name8791 (
		_w12837_,
		_w12838_,
		_w12839_
	);
	LUT3 #(
		.INIT('h01)
	) name8792 (
		\sport0_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[5]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[6]/NET0131 ,
		_w12840_
	);
	LUT4 #(
		.INIT('h0001)
	) name8793 (
		\sport0_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[5]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[6]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[7]/NET0131 ,
		_w12841_
	);
	LUT4 #(
		.INIT('h0800)
	) name8794 (
		\sport0_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[1]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[2]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		_w12842_
	);
	LUT4 #(
		.INIT('h0002)
	) name8795 (
		\sport0_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[2]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[3]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[4]/NET0131 ,
		_w12843_
	);
	LUT4 #(
		.INIT('h4000)
	) name8796 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		_w12841_,
		_w12842_,
		_w12843_,
		_w12844_
	);
	LUT4 #(
		.INIT('h1d00)
	) name8797 (
		\T_RD0_pad ,
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w9377_,
		_w12844_,
		_w12845_
	);
	LUT2 #(
		.INIT('h1)
	) name8798 (
		\sport0_rxctl_SLOT1_EXT_reg[2]/NET0131 ,
		_w12844_,
		_w12846_
	);
	LUT2 #(
		.INIT('h1)
	) name8799 (
		_w12845_,
		_w12846_,
		_w12847_
	);
	LUT4 #(
		.INIT('h8000)
	) name8800 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		_w12841_,
		_w12842_,
		_w12843_,
		_w12848_
	);
	LUT4 #(
		.INIT('h1d00)
	) name8801 (
		\T_RD0_pad ,
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w9377_,
		_w12848_,
		_w12849_
	);
	LUT2 #(
		.INIT('h1)
	) name8802 (
		\sport0_rxctl_SLOT1_EXT_reg[3]/NET0131 ,
		_w12848_,
		_w12850_
	);
	LUT2 #(
		.INIT('h1)
	) name8803 (
		_w12849_,
		_w12850_,
		_w12851_
	);
	LUT4 #(
		.INIT('h03aa)
	) name8804 (
		\sport0_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w7465_,
		_w7565_,
		_w12826_,
		_w12852_
	);
	LUT3 #(
		.INIT('h40)
	) name8805 (
		IACKn_pad,
		\idma_IRDn_reg/P0001 ,
		\idma_IWRn_reg/P0001 ,
		_w12853_
	);
	LUT4 #(
		.INIT('hbf00)
	) name8806 (
		IACKn_pad,
		\idma_IRDn_reg/P0001 ,
		\idma_IWRn_reg/P0001 ,
		\idma_WRtrue_reg/NET0131 ,
		_w12854_
	);
	LUT3 #(
		.INIT('h8c)
	) name8807 (
		\idma_WRcnt_reg[0]/NET0131 ,
		\idma_WRcnt_reg[1]/NET0131 ,
		_w12854_,
		_w12855_
	);
	LUT2 #(
		.INIT('h2)
	) name8808 (
		_w12814_,
		_w12853_,
		_w12856_
	);
	LUT4 #(
		.INIT('hff07)
	) name8809 (
		\idma_WRtrue_reg/NET0131 ,
		_w12811_,
		_w12814_,
		_w12853_,
		_w12857_
	);
	LUT3 #(
		.INIT('h04)
	) name8810 (
		\memc_usysr_DO_reg[8]/NET0131 ,
		_w12814_,
		_w12853_,
		_w12858_
	);
	LUT3 #(
		.INIT('h0b)
	) name8811 (
		_w12855_,
		_w12857_,
		_w12858_,
		_w12859_
	);
	LUT4 #(
		.INIT('h0001)
	) name8812 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w12860_
	);
	LUT3 #(
		.INIT('h04)
	) name8813 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w9931_,
		_w12860_,
		_w12861_
	);
	LUT3 #(
		.INIT('h04)
	) name8814 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w12862_
	);
	LUT4 #(
		.INIT('hd777)
	) name8815 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12862_,
		_w12863_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8816 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001 ,
		_w4834_,
		_w12861_,
		_w12863_,
		_w12864_
	);
	LUT4 #(
		.INIT('h7d77)
	) name8817 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12862_,
		_w12865_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8818 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001 ,
		_w4834_,
		_w12861_,
		_w12865_,
		_w12866_
	);
	LUT3 #(
		.INIT('h20)
	) name8819 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w12867_
	);
	LUT4 #(
		.INIT('hd777)
	) name8820 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12867_,
		_w12868_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8821 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001 ,
		_w4834_,
		_w12861_,
		_w12868_,
		_w12869_
	);
	LUT4 #(
		.INIT('h7d77)
	) name8822 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12867_,
		_w12870_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8823 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001 ,
		_w4834_,
		_w12861_,
		_w12870_,
		_w12871_
	);
	LUT3 #(
		.INIT('h02)
	) name8824 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w12872_
	);
	LUT4 #(
		.INIT('hd777)
	) name8825 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12872_,
		_w12873_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8826 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001 ,
		_w4834_,
		_w12861_,
		_w12873_,
		_w12874_
	);
	LUT4 #(
		.INIT('h7d77)
	) name8827 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12872_,
		_w12875_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8828 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001 ,
		_w4834_,
		_w12861_,
		_w12875_,
		_w12876_
	);
	LUT3 #(
		.INIT('h10)
	) name8829 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w12877_
	);
	LUT4 #(
		.INIT('hd777)
	) name8830 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12877_,
		_w12878_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8831 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001 ,
		_w4834_,
		_w12861_,
		_w12878_,
		_w12879_
	);
	LUT4 #(
		.INIT('h7d77)
	) name8832 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12877_,
		_w12880_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8833 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001 ,
		_w4834_,
		_w12861_,
		_w12880_,
		_w12881_
	);
	LUT3 #(
		.INIT('h01)
	) name8834 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w12882_
	);
	LUT4 #(
		.INIT('hd777)
	) name8835 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12882_,
		_w12883_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8836 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001 ,
		_w4834_,
		_w12861_,
		_w12883_,
		_w12884_
	);
	LUT3 #(
		.INIT('h40)
	) name8837 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w12885_
	);
	LUT4 #(
		.INIT('hd777)
	) name8838 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12885_,
		_w12886_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8839 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001 ,
		_w4834_,
		_w12861_,
		_w12886_,
		_w12887_
	);
	LUT4 #(
		.INIT('h7d77)
	) name8840 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12885_,
		_w12888_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8841 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001 ,
		_w4834_,
		_w12861_,
		_w12888_,
		_w12889_
	);
	LUT4 #(
		.INIT('h7d77)
	) name8842 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w12882_,
		_w12890_
	);
	LUT4 #(
		.INIT('h2aea)
	) name8843 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001 ,
		_w4834_,
		_w12861_,
		_w12890_,
		_w12891_
	);
	LUT4 #(
		.INIT('h03aa)
	) name8844 (
		\sport0_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w12826_,
		_w12892_
	);
	LUT4 #(
		.INIT('h03aa)
	) name8845 (
		\sport0_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w12826_,
		_w12893_
	);
	LUT3 #(
		.INIT('h01)
	) name8846 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		\core_c_dec_MpopLP_Eg_reg/P0001 ,
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		_w12894_
	);
	LUT3 #(
		.INIT('h08)
	) name8847 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[2]/NET0131 ,
		_w12895_
	);
	LUT3 #(
		.INIT('h8a)
	) name8848 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w12896_
	);
	LUT4 #(
		.INIT('h008a)
	) name8849 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w12895_,
		_w12897_
	);
	LUT2 #(
		.INIT('h4)
	) name8850 (
		_w12894_,
		_w12897_,
		_w12898_
	);
	LUT4 #(
		.INIT('h5551)
	) name8851 (
		\core_c_dec_MpopLP_Eg_reg/P0001 ,
		_w4169_,
		_w4430_,
		_w4178_,
		_w12899_
	);
	LUT4 #(
		.INIT('h0001)
	) name8852 (
		\core_c_psq_lpstk_ptr_reg[2]/NET0131 ,
		_w4971_,
		_w12894_,
		_w12899_,
		_w12900_
	);
	LUT2 #(
		.INIT('h9)
	) name8853 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w12901_
	);
	LUT4 #(
		.INIT('h008a)
	) name8854 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w12901_,
		_w12902_
	);
	LUT3 #(
		.INIT('h0b)
	) name8855 (
		_w12897_,
		_w12901_,
		_w12902_,
		_w12903_
	);
	LUT4 #(
		.INIT('h02fe)
	) name8856 (
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w12898_,
		_w12900_,
		_w12903_,
		_w12904_
	);
	LUT3 #(
		.INIT('h56)
	) name8857 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		_w12898_,
		_w12900_,
		_w12905_
	);
	LUT4 #(
		.INIT('hc444)
	) name8858 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[7]/NET0131 ,
		_w4073_,
		_w4084_,
		_w12906_
	);
	LUT4 #(
		.INIT('hff20)
	) name8859 (
		_w12271_,
		_w12272_,
		_w12275_,
		_w12906_,
		_w12907_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name8860 (
		\core_c_psq_lpstk_ptr_reg[2]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12896_,
		_w12908_
	);
	LUT2 #(
		.INIT('h2)
	) name8861 (
		_w4434_,
		_w12894_,
		_w12909_
	);
	LUT2 #(
		.INIT('h4)
	) name8862 (
		_w12897_,
		_w12909_,
		_w12910_
	);
	LUT4 #(
		.INIT('hf1f0)
	) name8863 (
		_w4971_,
		_w12899_,
		_w12908_,
		_w12910_,
		_w12911_
	);
	LUT3 #(
		.INIT('ha8)
	) name8864 (
		_w5327_,
		_w7465_,
		_w7565_,
		_w12912_
	);
	LUT4 #(
		.INIT('h00ef)
	) name8865 (
		_w5327_,
		_w8118_,
		_w8121_,
		_w12912_,
		_w12913_
	);
	LUT3 #(
		.INIT('h73)
	) name8866 (
		_w5041_,
		_w8093_,
		_w12913_,
		_w12914_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8867 (
		_w5029_,
		_w5041_,
		_w8093_,
		_w12913_,
		_w12915_
	);
	LUT2 #(
		.INIT('h2)
	) name8868 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w12916_
	);
	LUT2 #(
		.INIT('h8)
	) name8869 (
		_w5046_,
		_w12916_,
		_w12917_
	);
	LUT3 #(
		.INIT('h80)
	) name8870 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12918_
	);
	LUT3 #(
		.INIT('h07)
	) name8871 (
		_w4073_,
		_w4084_,
		_w12918_,
		_w12919_
	);
	LUT3 #(
		.INIT('h40)
	) name8872 (
		\core_c_psq_Taddr_Eb_reg[8]/P0001 ,
		_w4073_,
		_w4084_,
		_w12920_
	);
	LUT3 #(
		.INIT('h0b)
	) name8873 (
		_w12915_,
		_w12919_,
		_w12920_,
		_w12921_
	);
	LUT4 #(
		.INIT('h8a88)
	) name8874 (
		_w5327_,
		_w7793_,
		_w7903_,
		_w7905_,
		_w12922_
	);
	LUT4 #(
		.INIT('h00ef)
	) name8875 (
		_w5327_,
		_w8052_,
		_w8055_,
		_w12922_,
		_w12923_
	);
	LUT3 #(
		.INIT('h73)
	) name8876 (
		_w5041_,
		_w8061_,
		_w12923_,
		_w12924_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8877 (
		_w5029_,
		_w5041_,
		_w8061_,
		_w12923_,
		_w12925_
	);
	LUT3 #(
		.INIT('h80)
	) name8878 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12926_
	);
	LUT3 #(
		.INIT('h07)
	) name8879 (
		_w4073_,
		_w4084_,
		_w12926_,
		_w12927_
	);
	LUT3 #(
		.INIT('h40)
	) name8880 (
		\core_c_psq_Taddr_Eb_reg[7]/P0001 ,
		_w4073_,
		_w4084_,
		_w12928_
	);
	LUT3 #(
		.INIT('h0b)
	) name8881 (
		_w12925_,
		_w12927_,
		_w12928_,
		_w12929_
	);
	LUT4 #(
		.INIT('h8a88)
	) name8882 (
		_w5327_,
		_w7927_,
		_w8040_,
		_w8042_,
		_w12930_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8883 (
		_w5327_,
		_w7715_,
		_w7720_,
		_w12930_,
		_w12931_
	);
	LUT3 #(
		.INIT('h73)
	) name8884 (
		_w5041_,
		_w7748_,
		_w12931_,
		_w12932_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8885 (
		_w5029_,
		_w5041_,
		_w7748_,
		_w12931_,
		_w12933_
	);
	LUT3 #(
		.INIT('h80)
	) name8886 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12934_
	);
	LUT3 #(
		.INIT('h07)
	) name8887 (
		_w4073_,
		_w4084_,
		_w12934_,
		_w12935_
	);
	LUT3 #(
		.INIT('h40)
	) name8888 (
		\core_c_psq_Taddr_Eb_reg[6]/P0001 ,
		_w4073_,
		_w4084_,
		_w12936_
	);
	LUT3 #(
		.INIT('h0b)
	) name8889 (
		_w12933_,
		_w12935_,
		_w12936_,
		_w12937_
	);
	LUT4 #(
		.INIT('h8a88)
	) name8890 (
		_w5327_,
		_w7592_,
		_w7707_,
		_w7709_,
		_w12938_
	);
	LUT4 #(
		.INIT('h00ef)
	) name8891 (
		_w5327_,
		_w7386_,
		_w7390_,
		_w12938_,
		_w12939_
	);
	LUT3 #(
		.INIT('h73)
	) name8892 (
		_w5041_,
		_w7419_,
		_w12939_,
		_w12940_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8893 (
		_w5029_,
		_w5041_,
		_w7419_,
		_w12939_,
		_w12941_
	);
	LUT3 #(
		.INIT('h80)
	) name8894 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12942_
	);
	LUT3 #(
		.INIT('h07)
	) name8895 (
		_w4073_,
		_w4084_,
		_w12942_,
		_w12943_
	);
	LUT3 #(
		.INIT('h40)
	) name8896 (
		\core_c_psq_Taddr_Eb_reg[5]/P0001 ,
		_w4073_,
		_w4084_,
		_w12944_
	);
	LUT3 #(
		.INIT('h0b)
	) name8897 (
		_w12941_,
		_w12943_,
		_w12944_,
		_w12945_
	);
	LUT4 #(
		.INIT('h8a88)
	) name8898 (
		_w5327_,
		_w7257_,
		_w7375_,
		_w7377_,
		_w12946_
	);
	LUT4 #(
		.INIT('h00ef)
	) name8899 (
		_w5327_,
		_w7083_,
		_w7086_,
		_w12946_,
		_w12947_
	);
	LUT3 #(
		.INIT('h73)
	) name8900 (
		_w5041_,
		_w7096_,
		_w12947_,
		_w12948_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8901 (
		_w5029_,
		_w5041_,
		_w7096_,
		_w12947_,
		_w12949_
	);
	LUT3 #(
		.INIT('h80)
	) name8902 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12950_
	);
	LUT3 #(
		.INIT('h07)
	) name8903 (
		_w4073_,
		_w4084_,
		_w12950_,
		_w12951_
	);
	LUT3 #(
		.INIT('h40)
	) name8904 (
		\core_c_psq_Taddr_Eb_reg[4]/P0001 ,
		_w4073_,
		_w4084_,
		_w12952_
	);
	LUT3 #(
		.INIT('h0b)
	) name8905 (
		_w12949_,
		_w12951_,
		_w12952_,
		_w12953_
	);
	LUT3 #(
		.INIT('h73)
	) name8906 (
		_w5041_,
		_w7034_,
		_w9156_,
		_w12954_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8907 (
		_w5029_,
		_w5041_,
		_w7034_,
		_w9156_,
		_w12955_
	);
	LUT3 #(
		.INIT('h80)
	) name8908 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12956_
	);
	LUT3 #(
		.INIT('h07)
	) name8909 (
		_w4073_,
		_w4084_,
		_w12956_,
		_w12957_
	);
	LUT3 #(
		.INIT('h40)
	) name8910 (
		\core_c_psq_Taddr_Eb_reg[3]/P0001 ,
		_w4073_,
		_w4084_,
		_w12958_
	);
	LUT3 #(
		.INIT('h0b)
	) name8911 (
		_w12955_,
		_w12957_,
		_w12958_,
		_w12959_
	);
	LUT4 #(
		.INIT('h2022)
	) name8912 (
		_w5327_,
		_w6378_,
		_w6498_,
		_w6500_,
		_w12960_
	);
	LUT4 #(
		.INIT('h00ba)
	) name8913 (
		_w5327_,
		_w7004_,
		_w7008_,
		_w12960_,
		_w12961_
	);
	LUT3 #(
		.INIT('h37)
	) name8914 (
		_w5041_,
		_w6996_,
		_w12961_,
		_w12962_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name8915 (
		_w5029_,
		_w5041_,
		_w6996_,
		_w12961_,
		_w12963_
	);
	LUT3 #(
		.INIT('h80)
	) name8916 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12964_
	);
	LUT3 #(
		.INIT('h07)
	) name8917 (
		_w4073_,
		_w4084_,
		_w12964_,
		_w12965_
	);
	LUT3 #(
		.INIT('h40)
	) name8918 (
		\core_c_psq_Taddr_Eb_reg[2]/P0001 ,
		_w4073_,
		_w4084_,
		_w12966_
	);
	LUT3 #(
		.INIT('h0b)
	) name8919 (
		_w12963_,
		_w12965_,
		_w12966_,
		_w12967_
	);
	LUT4 #(
		.INIT('h2022)
	) name8920 (
		_w5327_,
		_w6774_,
		_w6894_,
		_w6896_,
		_w12968_
	);
	LUT4 #(
		.INIT('h00ba)
	) name8921 (
		_w5327_,
		_w6965_,
		_w6970_,
		_w12968_,
		_w12969_
	);
	LUT3 #(
		.INIT('h37)
	) name8922 (
		_w5041_,
		_w6955_,
		_w12969_,
		_w12970_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name8923 (
		_w5029_,
		_w5041_,
		_w6955_,
		_w12969_,
		_w12971_
	);
	LUT3 #(
		.INIT('h80)
	) name8924 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12972_
	);
	LUT3 #(
		.INIT('h07)
	) name8925 (
		_w4073_,
		_w4084_,
		_w12972_,
		_w12973_
	);
	LUT3 #(
		.INIT('h40)
	) name8926 (
		\core_c_psq_Taddr_Eb_reg[1]/P0001 ,
		_w4073_,
		_w4084_,
		_w12974_
	);
	LUT3 #(
		.INIT('h0b)
	) name8927 (
		_w12971_,
		_w12973_,
		_w12974_,
		_w12975_
	);
	LUT4 #(
		.INIT('h5554)
	) name8928 (
		_w5327_,
		_w6909_,
		_w6910_,
		_w6911_,
		_w12976_
	);
	LUT2 #(
		.INIT('h8)
	) name8929 (
		_w5327_,
		_w5760_,
		_w12977_
	);
	LUT4 #(
		.INIT('h888c)
	) name8930 (
		_w5041_,
		_w6918_,
		_w12976_,
		_w12977_,
		_w12978_
	);
	LUT3 #(
		.INIT('h80)
	) name8931 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12979_
	);
	LUT3 #(
		.INIT('h07)
	) name8932 (
		_w4073_,
		_w4084_,
		_w12979_,
		_w12980_
	);
	LUT3 #(
		.INIT('h40)
	) name8933 (
		\core_c_psq_Taddr_Eb_reg[13]/P0001 ,
		_w4073_,
		_w4084_,
		_w12981_
	);
	LUT4 #(
		.INIT('h002f)
	) name8934 (
		_w5029_,
		_w12978_,
		_w12980_,
		_w12981_,
		_w12982_
	);
	LUT2 #(
		.INIT('h8)
	) name8935 (
		_w5327_,
		_w6758_,
		_w12983_
	);
	LUT4 #(
		.INIT('h00ba)
	) name8936 (
		_w5327_,
		_w6576_,
		_w6580_,
		_w12983_,
		_w12984_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name8937 (
		_w5029_,
		_w5041_,
		_w6608_,
		_w12984_,
		_w12985_
	);
	LUT3 #(
		.INIT('h80)
	) name8938 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12986_
	);
	LUT3 #(
		.INIT('h07)
	) name8939 (
		_w4073_,
		_w4084_,
		_w12986_,
		_w12987_
	);
	LUT3 #(
		.INIT('h40)
	) name8940 (
		\core_c_psq_Taddr_Eb_reg[12]/P0001 ,
		_w4073_,
		_w4084_,
		_w12988_
	);
	LUT3 #(
		.INIT('h0b)
	) name8941 (
		_w12985_,
		_w12987_,
		_w12988_,
		_w12989_
	);
	LUT3 #(
		.INIT('h02)
	) name8942 (
		_w5327_,
		_w6263_,
		_w6362_,
		_w12990_
	);
	LUT4 #(
		.INIT('h00ba)
	) name8943 (
		_w5327_,
		_w6529_,
		_w6533_,
		_w12990_,
		_w12991_
	);
	LUT4 #(
		.INIT('hff45)
	) name8944 (
		_w5327_,
		_w6529_,
		_w6533_,
		_w12990_,
		_w12992_
	);
	LUT3 #(
		.INIT('h37)
	) name8945 (
		_w5041_,
		_w6506_,
		_w12991_,
		_w12993_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name8946 (
		_w5029_,
		_w5041_,
		_w6506_,
		_w12991_,
		_w12994_
	);
	LUT3 #(
		.INIT('h80)
	) name8947 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w5046_,
		_w12916_,
		_w12995_
	);
	LUT3 #(
		.INIT('h07)
	) name8948 (
		_w4073_,
		_w4084_,
		_w12995_,
		_w12996_
	);
	LUT3 #(
		.INIT('h40)
	) name8949 (
		\core_c_psq_Taddr_Eb_reg[11]/P0001 ,
		_w4073_,
		_w4084_,
		_w12997_
	);
	LUT3 #(
		.INIT('h0b)
	) name8950 (
		_w12994_,
		_w12996_,
		_w12997_,
		_w12998_
	);
	LUT3 #(
		.INIT('ha8)
	) name8951 (
		_w5327_,
		_w5937_,
		_w6038_,
		_w12999_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8952 (
		_w5327_,
		_w6209_,
		_w6215_,
		_w12999_,
		_w13000_
	);
	LUT3 #(
		.INIT('h73)
	) name8953 (
		_w5041_,
		_w6181_,
		_w13000_,
		_w13001_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8954 (
		_w5029_,
		_w5041_,
		_w6181_,
		_w13000_,
		_w13002_
	);
	LUT3 #(
		.INIT('h80)
	) name8955 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w5046_,
		_w12916_,
		_w13003_
	);
	LUT3 #(
		.INIT('h07)
	) name8956 (
		_w4073_,
		_w4084_,
		_w13003_,
		_w13004_
	);
	LUT3 #(
		.INIT('h40)
	) name8957 (
		\core_c_psq_Taddr_Eb_reg[10]/P0001 ,
		_w4073_,
		_w4084_,
		_w13005_
	);
	LUT3 #(
		.INIT('h0b)
	) name8958 (
		_w13002_,
		_w13004_,
		_w13005_,
		_w13006_
	);
	LUT4 #(
		.INIT('h2022)
	) name8959 (
		_w5327_,
		_w5784_,
		_w5911_,
		_w5913_,
		_w13007_
	);
	LUT4 #(
		.INIT('h00ba)
	) name8960 (
		_w5327_,
		_w5439_,
		_w5529_,
		_w13007_,
		_w13008_
	);
	LUT3 #(
		.INIT('h37)
	) name8961 (
		_w5041_,
		_w5549_,
		_w13008_,
		_w13009_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name8962 (
		_w5029_,
		_w5041_,
		_w5549_,
		_w13008_,
		_w13010_
	);
	LUT3 #(
		.INIT('h80)
	) name8963 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w5046_,
		_w12916_,
		_w13011_
	);
	LUT3 #(
		.INIT('h07)
	) name8964 (
		_w4073_,
		_w4084_,
		_w13011_,
		_w13012_
	);
	LUT3 #(
		.INIT('h40)
	) name8965 (
		\core_c_psq_Taddr_Eb_reg[0]/P0001 ,
		_w4073_,
		_w4084_,
		_w13013_
	);
	LUT3 #(
		.INIT('h0b)
	) name8966 (
		_w13010_,
		_w13012_,
		_w13013_,
		_w13014_
	);
	LUT4 #(
		.INIT('h8000)
	) name8967 (
		\sice_ICYC_reg[7]/NET0131 ,
		\sice_ICYC_reg[8]/NET0131 ,
		\sice_ICYC_reg[9]/NET0131 ,
		_w11932_,
		_w13015_
	);
	LUT4 #(
		.INIT('h8000)
	) name8968 (
		\sice_ICYC_reg[10]/NET0131 ,
		\sice_ICYC_reg[11]/NET0131 ,
		\sice_ICYC_reg[12]/NET0131 ,
		_w13015_,
		_w13016_
	);
	LUT4 #(
		.INIT('h8000)
	) name8969 (
		\sice_ICYC_reg[13]/NET0131 ,
		\sice_ICYC_reg[14]/NET0131 ,
		\sice_ICYC_reg[15]/NET0131 ,
		_w13016_,
		_w13017_
	);
	LUT4 #(
		.INIT('h8000)
	) name8970 (
		\sice_ICYC_reg[16]/NET0131 ,
		\sice_ICYC_reg[17]/NET0131 ,
		\sice_ICYC_reg[18]/NET0131 ,
		_w13017_,
		_w13018_
	);
	LUT4 #(
		.INIT('h8000)
	) name8971 (
		\sice_ICYC_reg[19]/NET0131 ,
		\sice_ICYC_reg[20]/NET0131 ,
		\sice_ICYC_reg[21]/NET0131 ,
		_w13018_,
		_w13019_
	);
	LUT4 #(
		.INIT('h78f0)
	) name8972 (
		\sice_ICYC_reg[19]/NET0131 ,
		\sice_ICYC_reg[20]/NET0131 ,
		\sice_ICYC_reg[21]/NET0131 ,
		_w13018_,
		_w13020_
	);
	LUT3 #(
		.INIT('ha8)
	) name8973 (
		_w5327_,
		_w7140_,
		_w7240_,
		_w13021_
	);
	LUT4 #(
		.INIT('h00ef)
	) name8974 (
		_w5327_,
		_w8157_,
		_w8162_,
		_w13021_,
		_w13022_
	);
	LUT3 #(
		.INIT('h73)
	) name8975 (
		_w5041_,
		_w8132_,
		_w13022_,
		_w13023_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8976 (
		_w5029_,
		_w5041_,
		_w8132_,
		_w13022_,
		_w13024_
	);
	LUT3 #(
		.INIT('h80)
	) name8977 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		_w5046_,
		_w12916_,
		_w13025_
	);
	LUT3 #(
		.INIT('h07)
	) name8978 (
		_w4073_,
		_w4084_,
		_w13025_,
		_w13026_
	);
	LUT3 #(
		.INIT('h40)
	) name8979 (
		\core_c_psq_Taddr_Eb_reg[9]/P0001 ,
		_w4073_,
		_w4084_,
		_w13027_
	);
	LUT3 #(
		.INIT('h0b)
	) name8980 (
		_w13024_,
		_w13026_,
		_w13027_,
		_w13028_
	);
	LUT4 #(
		.INIT('h1555)
	) name8981 (
		\bdma_BEAD_reg[0]/NET0131 ,
		_w4885_,
		_w4884_,
		_w9075_,
		_w13029_
	);
	LUT3 #(
		.INIT('h04)
	) name8982 (
		_w9412_,
		_w9413_,
		_w13029_,
		_w13030_
	);
	LUT4 #(
		.INIT('h0020)
	) name8983 (
		\bdma_BEAD_reg[1]/NET0131 ,
		_w9412_,
		_w9413_,
		_w13029_,
		_w13031_
	);
	LUT4 #(
		.INIT('h8000)
	) name8984 (
		_w5643_,
		_w5658_,
		_w9431_,
		_w12621_,
		_w13032_
	);
	LUT3 #(
		.INIT('h12)
	) name8985 (
		\bdma_BEAD_reg[1]/NET0131 ,
		_w13032_,
		_w13030_,
		_w13033_
	);
	LUT4 #(
		.INIT('h4500)
	) name8986 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13032_,
		_w13034_
	);
	LUT2 #(
		.INIT('he)
	) name8987 (
		_w13033_,
		_w13034_,
		_w13035_
	);
	LUT4 #(
		.INIT('h5655)
	) name8988 (
		\bdma_BEAD_reg[0]/NET0131 ,
		_w9077_,
		_w9412_,
		_w9413_,
		_w13036_
	);
	LUT2 #(
		.INIT('h1)
	) name8989 (
		_w13032_,
		_w13036_,
		_w13037_
	);
	LUT4 #(
		.INIT('h4500)
	) name8990 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13032_,
		_w13038_
	);
	LUT2 #(
		.INIT('he)
	) name8991 (
		_w13037_,
		_w13038_,
		_w13039_
	);
	LUT4 #(
		.INIT('h9aaa)
	) name8992 (
		\clkc_CLKOUT_reg/NET0131 ,
		_w12254_,
		_w12258_,
		_w12263_,
		_w13040_
	);
	LUT2 #(
		.INIT('h6)
	) name8993 (
		\sice_ICYC_reg[22]/NET0131 ,
		_w13019_,
		_w13041_
	);
	LUT3 #(
		.INIT('h80)
	) name8994 (
		_w5790_,
		_w9431_,
		_w11604_,
		_w13042_
	);
	LUT4 #(
		.INIT('h4000)
	) name8995 (
		\memc_MMR_web_reg/NET0131 ,
		_w5790_,
		_w9431_,
		_w11604_,
		_w13043_
	);
	LUT4 #(
		.INIT('hba00)
	) name8996 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13043_,
		_w13044_
	);
	LUT2 #(
		.INIT('h1)
	) name8997 (
		\tm_tsr_reg_DO_reg[7]/NET0131 ,
		_w13043_,
		_w13045_
	);
	LUT2 #(
		.INIT('h1)
	) name8998 (
		_w13044_,
		_w13045_,
		_w13046_
	);
	LUT4 #(
		.INIT('hba00)
	) name8999 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13043_,
		_w13047_
	);
	LUT2 #(
		.INIT('h1)
	) name9000 (
		\tm_tsr_reg_DO_reg[6]/NET0131 ,
		_w13043_,
		_w13048_
	);
	LUT2 #(
		.INIT('h1)
	) name9001 (
		_w13047_,
		_w13048_,
		_w13049_
	);
	LUT4 #(
		.INIT('hba00)
	) name9002 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13043_,
		_w13050_
	);
	LUT2 #(
		.INIT('h1)
	) name9003 (
		\tm_tsr_reg_DO_reg[5]/NET0131 ,
		_w13043_,
		_w13051_
	);
	LUT2 #(
		.INIT('h1)
	) name9004 (
		_w13050_,
		_w13051_,
		_w13052_
	);
	LUT4 #(
		.INIT('hba00)
	) name9005 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13043_,
		_w13053_
	);
	LUT2 #(
		.INIT('h1)
	) name9006 (
		\tm_tsr_reg_DO_reg[3]/NET0131 ,
		_w13043_,
		_w13054_
	);
	LUT2 #(
		.INIT('h1)
	) name9007 (
		_w13053_,
		_w13054_,
		_w13055_
	);
	LUT4 #(
		.INIT('hba00)
	) name9008 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13043_,
		_w13056_
	);
	LUT2 #(
		.INIT('h1)
	) name9009 (
		\tm_tsr_reg_DO_reg[2]/NET0131 ,
		_w13043_,
		_w13057_
	);
	LUT2 #(
		.INIT('h1)
	) name9010 (
		_w13056_,
		_w13057_,
		_w13058_
	);
	LUT4 #(
		.INIT('hba00)
	) name9011 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13043_,
		_w13059_
	);
	LUT2 #(
		.INIT('h1)
	) name9012 (
		\tm_tsr_reg_DO_reg[4]/NET0131 ,
		_w13043_,
		_w13060_
	);
	LUT2 #(
		.INIT('h1)
	) name9013 (
		_w13059_,
		_w13060_,
		_w13061_
	);
	LUT4 #(
		.INIT('hba00)
	) name9014 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13043_,
		_w13062_
	);
	LUT2 #(
		.INIT('h1)
	) name9015 (
		\tm_tsr_reg_DO_reg[1]/NET0131 ,
		_w13043_,
		_w13063_
	);
	LUT2 #(
		.INIT('h1)
	) name9016 (
		_w13062_,
		_w13063_,
		_w13064_
	);
	LUT4 #(
		.INIT('hba00)
	) name9017 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13043_,
		_w13065_
	);
	LUT2 #(
		.INIT('h1)
	) name9018 (
		\tm_tsr_reg_DO_reg[0]/NET0131 ,
		_w13043_,
		_w13066_
	);
	LUT2 #(
		.INIT('h1)
	) name9019 (
		_w13065_,
		_w13066_,
		_w13067_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9020 (
		\tm_tsr_reg_DO_reg[8]/NET0131 ,
		_w8798_,
		_w8801_,
		_w13043_,
		_w13068_
	);
	LUT3 #(
		.INIT('h04)
	) name9021 (
		\memc_usysr_DO_reg[7]/NET0131 ,
		_w12814_,
		_w12853_,
		_w13069_
	);
	LUT4 #(
		.INIT('h5509)
	) name9022 (
		\idma_WRcnt_reg[0]/NET0131 ,
		\idma_WRtrue_reg/NET0131 ,
		_w12814_,
		_w12853_,
		_w13070_
	);
	LUT2 #(
		.INIT('h1)
	) name9023 (
		_w13069_,
		_w13070_,
		_w13071_
	);
	LUT4 #(
		.INIT('h2333)
	) name9024 (
		IACKn_pad,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_IRDn_reg/P0001 ,
		\idma_IWRn_reg/P0001 ,
		_w13072_
	);
	LUT3 #(
		.INIT('h40)
	) name9025 (
		\idma_PM_1st_reg/NET0131 ,
		\idma_RDcyc_reg/NET0131 ,
		_w13072_,
		_w13073_
	);
	LUT2 #(
		.INIT('h4)
	) name9026 (
		\idma_RDCMD_d1_reg/P0001 ,
		\idma_RDCMD_reg/P0001 ,
		_w13074_
	);
	LUT3 #(
		.INIT('h40)
	) name9027 (
		\idma_PM_1st_reg/NET0131 ,
		_w13074_,
		_w13072_,
		_w13075_
	);
	LUT4 #(
		.INIT('h4000)
	) name9028 (
		\idma_PM_1st_reg/NET0131 ,
		\idma_RDcyc_reg/NET0131 ,
		_w12819_,
		_w13072_,
		_w13076_
	);
	LUT4 #(
		.INIT('h0603)
	) name9029 (
		\idma_RDcnt_reg[0]/NET0131 ,
		\idma_RDcnt_reg[1]/NET0131 ,
		_w13075_,
		_w13073_,
		_w13077_
	);
	LUT4 #(
		.INIT('h1000)
	) name9030 (
		\idma_PM_1st_reg/NET0131 ,
		\memc_usysr_DO_reg[5]/NET0131 ,
		_w13074_,
		_w13072_,
		_w13078_
	);
	LUT2 #(
		.INIT('h1)
	) name9031 (
		_w13077_,
		_w13078_,
		_w13079_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name9032 (
		\idma_RDcnt_reg[0]/NET0131 ,
		\memc_usysr_DO_reg[4]/NET0131 ,
		_w13075_,
		_w13073_,
		_w13080_
	);
	LUT2 #(
		.INIT('h8)
	) name9033 (
		\core_c_dec_updAR_E_reg/P0001 ,
		_w4106_,
		_w13081_
	);
	LUT3 #(
		.INIT('h20)
	) name9034 (
		_w4834_,
		_w11921_,
		_w11928_,
		_w13082_
	);
	LUT2 #(
		.INIT('he)
	) name9035 (
		_w13081_,
		_w13082_,
		_w13083_
	);
	LUT4 #(
		.INIT('h7f80)
	) name9036 (
		\sice_ICYC_reg[0]/NET0131 ,
		\sice_ICYC_reg[1]/NET0131 ,
		\sice_ICYC_reg[2]/NET0131 ,
		\sice_ICYC_reg[3]/NET0131 ,
		_w13084_
	);
	LUT4 #(
		.INIT('h7f80)
	) name9037 (
		\sice_IIRC_reg[0]/NET0131 ,
		\sice_IIRC_reg[1]/NET0131 ,
		\sice_IIRC_reg[2]/NET0131 ,
		\sice_IIRC_reg[3]/NET0131 ,
		_w13085_
	);
	LUT4 #(
		.INIT('h7f80)
	) name9038 (
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[1]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[2]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[3]/NET0131 ,
		_w13086_
	);
	LUT4 #(
		.INIT('h8000)
	) name9039 (
		\sice_IIRC_reg[7]/NET0131 ,
		\sice_IIRC_reg[8]/NET0131 ,
		\sice_IIRC_reg[9]/NET0131 ,
		_w11936_,
		_w13087_
	);
	LUT4 #(
		.INIT('h8000)
	) name9040 (
		\sice_IIRC_reg[10]/NET0131 ,
		\sice_IIRC_reg[11]/NET0131 ,
		\sice_IIRC_reg[12]/NET0131 ,
		_w13087_,
		_w13088_
	);
	LUT3 #(
		.INIT('h6c)
	) name9041 (
		\sice_IIRC_reg[13]/NET0131 ,
		\sice_IIRC_reg[14]/NET0131 ,
		_w13088_,
		_w13089_
	);
	LUT3 #(
		.INIT('h6c)
	) name9042 (
		\sice_ICYC_reg[13]/NET0131 ,
		\sice_ICYC_reg[14]/NET0131 ,
		_w13016_,
		_w13090_
	);
	LUT3 #(
		.INIT('h20)
	) name9043 (
		\core_c_dec_updMF_E_reg/P0001 ,
		_w9453_,
		_w9894_,
		_w13091_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name9044 (
		\core_c_dec_updMF_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001 ,
		_w9453_,
		_w9894_,
		_w13092_
	);
	LUT4 #(
		.INIT('h7200)
	) name9045 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12291_,
		_w12293_,
		_w13091_,
		_w13093_
	);
	LUT2 #(
		.INIT('he)
	) name9046 (
		_w13092_,
		_w13093_,
		_w13094_
	);
	LUT3 #(
		.INIT('h60)
	) name9047 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13095_
	);
	LUT3 #(
		.INIT('h15)
	) name9048 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13096_
	);
	LUT4 #(
		.INIT('h4800)
	) name9049 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13097_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9050 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13098_
	);
	LUT2 #(
		.INIT('h9)
	) name9051 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		_w13099_
	);
	LUT3 #(
		.INIT('h09)
	) name9052 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w13100_
	);
	LUT4 #(
		.INIT('h458a)
	) name9053 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13101_
	);
	LUT2 #(
		.INIT('h8)
	) name9054 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w13102_
	);
	LUT4 #(
		.INIT('h8040)
	) name9055 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13103_
	);
	LUT4 #(
		.INIT('h2022)
	) name9056 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13103_,
		_w13100_,
		_w13101_,
		_w13104_
	);
	LUT4 #(
		.INIT('h0e0d)
	) name9057 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13105_
	);
	LUT4 #(
		.INIT('h4020)
	) name9058 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13106_
	);
	LUT3 #(
		.INIT('h02)
	) name9059 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13106_,
		_w13105_,
		_w13107_
	);
	LUT4 #(
		.INIT('h3331)
	) name9060 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13098_,
		_w13106_,
		_w13105_,
		_w13108_
	);
	LUT4 #(
		.INIT('h082a)
	) name9061 (
		_w13096_,
		_w13098_,
		_w13104_,
		_w13107_,
		_w13109_
	);
	LUT4 #(
		.INIT('h8010)
	) name9062 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13110_
	);
	LUT3 #(
		.INIT('h84)
	) name9063 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13111_
	);
	LUT4 #(
		.INIT('h0b07)
	) name9064 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13112_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9065 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13110_,
		_w13111_,
		_w13112_,
		_w13113_
	);
	LUT3 #(
		.INIT('h60)
	) name9066 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13114_
	);
	LUT3 #(
		.INIT('h48)
	) name9067 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13115_
	);
	LUT2 #(
		.INIT('h4)
	) name9068 (
		_w13114_,
		_w13115_,
		_w13116_
	);
	LUT4 #(
		.INIT('h111b)
	) name9069 (
		_w13098_,
		_w13104_,
		_w13113_,
		_w13116_,
		_w13117_
	);
	LUT3 #(
		.INIT('h24)
	) name9070 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13118_
	);
	LUT4 #(
		.INIT('h4200)
	) name9071 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13119_
	);
	LUT3 #(
		.INIT('h54)
	) name9072 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w13118_,
		_w13119_,
		_w13120_
	);
	LUT4 #(
		.INIT('h152a)
	) name9073 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13121_
	);
	LUT3 #(
		.INIT('h84)
	) name9074 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13122_
	);
	LUT4 #(
		.INIT('h8040)
	) name9075 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13123_
	);
	LUT3 #(
		.INIT('h0e)
	) name9076 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13121_,
		_w13123_,
		_w13124_
	);
	LUT3 #(
		.INIT('h8a)
	) name9077 (
		_w13098_,
		_w13120_,
		_w13124_,
		_w13125_
	);
	LUT3 #(
		.INIT('h01)
	) name9078 (
		_w13098_,
		_w13113_,
		_w13116_,
		_w13126_
	);
	LUT2 #(
		.INIT('h1)
	) name9079 (
		_w13125_,
		_w13126_,
		_w13127_
	);
	LUT4 #(
		.INIT('h0007)
	) name9080 (
		_w13109_,
		_w13117_,
		_w13125_,
		_w13126_,
		_w13128_
	);
	LUT4 #(
		.INIT('h0008)
	) name9081 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13098_,
		_w13106_,
		_w13105_,
		_w13129_
	);
	LUT3 #(
		.INIT('h02)
	) name9082 (
		_w13095_,
		_w13098_,
		_w13102_,
		_w13130_
	);
	LUT2 #(
		.INIT('h1)
	) name9083 (
		_w13129_,
		_w13130_,
		_w13131_
	);
	LUT4 #(
		.INIT('h1555)
	) name9084 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13132_
	);
	LUT4 #(
		.INIT('h4a00)
	) name9085 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13133_
	);
	LUT4 #(
		.INIT('h0027)
	) name9086 (
		_w13098_,
		_w13104_,
		_w13107_,
		_w13133_,
		_w13134_
	);
	LUT3 #(
		.INIT('h80)
	) name9087 (
		_w13117_,
		_w13131_,
		_w13134_,
		_w13135_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name9088 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w13127_,
		_w13128_,
		_w13135_,
		_w13136_
	);
	LUT4 #(
		.INIT('h55a6)
	) name9089 (
		_w13096_,
		_w13098_,
		_w13104_,
		_w13108_,
		_w13137_
	);
	LUT4 #(
		.INIT('he0aa)
	) name9090 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13138_
	);
	LUT3 #(
		.INIT('h10)
	) name9091 (
		_w13129_,
		_w13130_,
		_w13138_,
		_w13139_
	);
	LUT3 #(
		.INIT('h80)
	) name9092 (
		_w13117_,
		_w13137_,
		_w13139_,
		_w13140_
	);
	LUT3 #(
		.INIT('h15)
	) name9093 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w13136_,
		_w13140_,
		_w13141_
	);
	LUT4 #(
		.INIT('h00bd)
	) name9094 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13142_
	);
	LUT4 #(
		.INIT('h70e0)
	) name9095 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w13143_
	);
	LUT2 #(
		.INIT('h4)
	) name9096 (
		_w13142_,
		_w13143_,
		_w13144_
	);
	LUT4 #(
		.INIT('h00ed)
	) name9097 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13145_
	);
	LUT3 #(
		.INIT('h54)
	) name9098 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w13122_,
		_w13145_,
		_w13146_
	);
	LUT2 #(
		.INIT('h1)
	) name9099 (
		_w13144_,
		_w13146_,
		_w13147_
	);
	LUT3 #(
		.INIT('h02)
	) name9100 (
		_w13098_,
		_w13144_,
		_w13146_,
		_w13148_
	);
	LUT3 #(
		.INIT('h10)
	) name9101 (
		_w13098_,
		_w13120_,
		_w13124_,
		_w13149_
	);
	LUT4 #(
		.INIT('h0800)
	) name9102 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13150_
	);
	LUT3 #(
		.INIT('h0e)
	) name9103 (
		_w13148_,
		_w13149_,
		_w13150_,
		_w13151_
	);
	LUT4 #(
		.INIT('h1055)
	) name9104 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w13127_,
		_w13135_,
		_w13151_,
		_w13152_
	);
	LUT4 #(
		.INIT('h1045)
	) name9105 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w13127_,
		_w13135_,
		_w13151_,
		_w13153_
	);
	LUT2 #(
		.INIT('h1)
	) name9106 (
		_w13148_,
		_w13153_,
		_w13154_
	);
	LUT2 #(
		.INIT('h8)
	) name9107 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13155_
	);
	LUT3 #(
		.INIT('h82)
	) name9108 (
		_w13155_,
		_w13141_,
		_w13154_,
		_w13156_
	);
	LUT4 #(
		.INIT('h1011)
	) name9109 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w7592_,
		_w7707_,
		_w7709_,
		_w13157_
	);
	LUT2 #(
		.INIT('h2)
	) name9110 (
		\sport0_rxctl_a_sync1_reg/P0001 ,
		\sport0_rxctl_a_sync2_reg/P0001 ,
		_w13158_
	);
	LUT3 #(
		.INIT('h40)
	) name9111 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13159_
	);
	LUT2 #(
		.INIT('h1)
	) name9112 (
		_w13158_,
		_w13159_,
		_w13160_
	);
	LUT4 #(
		.INIT('h4044)
	) name9113 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTRX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w13161_
	);
	LUT2 #(
		.INIT('he)
	) name9114 (
		_w13158_,
		_w13161_,
		_w13162_
	);
	LUT4 #(
		.INIT('hafac)
	) name9115 (
		\sport0_rxctl_RXSHT_reg[5]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w13163_
	);
	LUT4 #(
		.INIT('hef00)
	) name9116 (
		_w13156_,
		_w13157_,
		_w13160_,
		_w13163_,
		_w13164_
	);
	LUT4 #(
		.INIT('h0002)
	) name9117 (
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w13165_
	);
	LUT2 #(
		.INIT('he)
	) name9118 (
		_w13164_,
		_w13165_,
		_w13166_
	);
	LUT3 #(
		.INIT('h15)
	) name9119 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		_w12258_,
		_w12263_,
		_w13167_
	);
	LUT4 #(
		.INIT('h0040)
	) name9120 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_updMF_E_reg/P0001 ,
		_w9452_,
		_w9453_,
		_w13168_
	);
	LUT2 #(
		.INIT('h2)
	) name9121 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001 ,
		_w13168_,
		_w13169_
	);
	LUT4 #(
		.INIT('h7200)
	) name9122 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12291_,
		_w12293_,
		_w13168_,
		_w13170_
	);
	LUT2 #(
		.INIT('he)
	) name9123 (
		_w13169_,
		_w13170_,
		_w13171_
	);
	LUT4 #(
		.INIT('h135f)
	) name9124 (
		_w11555_,
		_w11435_,
		_w11449_,
		_w11458_,
		_w13172_
	);
	LUT4 #(
		.INIT('h0777)
	) name9125 (
		_w11341_,
		_w11397_,
		_w11558_,
		_w11469_,
		_w13173_
	);
	LUT2 #(
		.INIT('h8)
	) name9126 (
		_w13172_,
		_w13173_,
		_w13174_
	);
	LUT4 #(
		.INIT('hfa32)
	) name9127 (
		_w11534_,
		_w11538_,
		_w11489_,
		_w11953_,
		_w13175_
	);
	LUT2 #(
		.INIT('h4)
	) name9128 (
		_w11530_,
		_w11508_,
		_w13176_
	);
	LUT3 #(
		.INIT('he0)
	) name9129 (
		_w11393_,
		_w11589_,
		_w12412_,
		_w13177_
	);
	LUT3 #(
		.INIT('h10)
	) name9130 (
		_w13176_,
		_w13177_,
		_w13175_,
		_w13178_
	);
	LUT4 #(
		.INIT('h1311)
	) name9131 (
		_w11406_,
		_w11403_,
		_w11556_,
		_w11585_,
		_w13179_
	);
	LUT2 #(
		.INIT('h8)
	) name9132 (
		_w12642_,
		_w13179_,
		_w13180_
	);
	LUT2 #(
		.INIT('h8)
	) name9133 (
		_w11495_,
		_w11973_,
		_w13181_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name9134 (
		_w11588_,
		_w11510_,
		_w11465_,
		_w11839_,
		_w13182_
	);
	LUT4 #(
		.INIT('h0800)
	) name9135 (
		_w12642_,
		_w13179_,
		_w13181_,
		_w13182_,
		_w13183_
	);
	LUT3 #(
		.INIT('h80)
	) name9136 (
		_w13174_,
		_w13178_,
		_w13183_,
		_w13184_
	);
	LUT3 #(
		.INIT('hc8)
	) name9137 (
		_w11409_,
		_w11499_,
		_w11896_,
		_w13185_
	);
	LUT3 #(
		.INIT('h02)
	) name9138 (
		_w11386_,
		_w11540_,
		_w11953_,
		_w13186_
	);
	LUT3 #(
		.INIT('hc8)
	) name9139 (
		_w11587_,
		_w11874_,
		_w11880_,
		_w13187_
	);
	LUT3 #(
		.INIT('h01)
	) name9140 (
		_w13186_,
		_w13187_,
		_w13185_,
		_w13188_
	);
	LUT4 #(
		.INIT('ha820)
	) name9141 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001 ,
		_w13189_
	);
	LUT4 #(
		.INIT('h007f)
	) name9142 (
		_w11473_,
		_w11389_,
		_w11341_,
		_w13189_,
		_w13190_
	);
	LUT3 #(
		.INIT('h08)
	) name9143 (
		_w11389_,
		_w11476_,
		_w11471_,
		_w13191_
	);
	LUT3 #(
		.INIT('h80)
	) name9144 (
		_w11389_,
		_w11445_,
		_w11459_,
		_w13192_
	);
	LUT4 #(
		.INIT('h0100)
	) name9145 (
		_w11553_,
		_w13191_,
		_w13192_,
		_w13190_,
		_w13193_
	);
	LUT2 #(
		.INIT('h2)
	) name9146 (
		_w11415_,
		_w11454_,
		_w13194_
	);
	LUT4 #(
		.INIT('h135f)
	) name9147 (
		_w11578_,
		_w11529_,
		_w11496_,
		_w11511_,
		_w13195_
	);
	LUT4 #(
		.INIT('h0700)
	) name9148 (
		_w11522_,
		_w11872_,
		_w13194_,
		_w13195_,
		_w13196_
	);
	LUT4 #(
		.INIT('h00a8)
	) name9149 (
		_w11386_,
		_w11393_,
		_w11589_,
		_w11528_,
		_w13197_
	);
	LUT4 #(
		.INIT('h2000)
	) name9150 (
		_w12649_,
		_w13197_,
		_w13193_,
		_w13196_,
		_w13198_
	);
	LUT2 #(
		.INIT('h8)
	) name9151 (
		_w13188_,
		_w13198_,
		_w13199_
	);
	LUT4 #(
		.INIT('h8000)
	) name9152 (
		_w12451_,
		_w12666_,
		_w13184_,
		_w13199_,
		_w13200_
	);
	LUT4 #(
		.INIT('h4c08)
	) name9153 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11830_,
		_w12008_,
		_w13200_,
		_w13201_
	);
	LUT4 #(
		.INIT('h5545)
	) name9154 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w13202_
	);
	LUT2 #(
		.INIT('h1)
	) name9155 (
		_w13201_,
		_w13202_,
		_w13203_
	);
	LUT3 #(
		.INIT('h6c)
	) name9156 (
		\clkc_OUTcnt_reg[4]/NET0131 ,
		\clkc_OUTcnt_reg[5]/NET0131 ,
		_w12252_,
		_w13204_
	);
	LUT4 #(
		.INIT('hbf00)
	) name9157 (
		_w12254_,
		_w12258_,
		_w12263_,
		_w13204_,
		_w13205_
	);
	LUT4 #(
		.INIT('h4c08)
	) name9158 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11329_,
		_w12008_,
		_w13200_,
		_w13206_
	);
	LUT2 #(
		.INIT('h1)
	) name9159 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001 ,
		_w11329_,
		_w13207_
	);
	LUT2 #(
		.INIT('h1)
	) name9160 (
		_w13206_,
		_w13207_,
		_w13208_
	);
	LUT3 #(
		.INIT('h78)
	) name9161 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_OUTcnt_reg[1]/NET0131 ,
		\clkc_OUTcnt_reg[2]/NET0131 ,
		_w13209_
	);
	LUT4 #(
		.INIT('hbf00)
	) name9162 (
		_w12254_,
		_w12258_,
		_w12263_,
		_w13209_,
		_w13210_
	);
	LUT3 #(
		.INIT('h13)
	) name9163 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001 ,
		_w9894_,
		_w13211_
	);
	LUT4 #(
		.INIT('h0002)
	) name9164 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w13211_,
		_w13212_
	);
	LUT4 #(
		.INIT('h5700)
	) name9165 (
		_w11625_,
		_w12736_,
		_w12737_,
		_w13212_,
		_w13213_
	);
	LUT4 #(
		.INIT('h313b)
	) name9166 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001 ,
		_w11631_,
		_w11635_,
		_w13214_
	);
	LUT4 #(
		.INIT('hc480)
	) name9167 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w11637_,
		_w12356_,
		_w13215_
	);
	LUT4 #(
		.INIT('hff45)
	) name9168 (
		_w11624_,
		_w13213_,
		_w13214_,
		_w13215_,
		_w13216_
	);
	LUT4 #(
		.INIT('h084c)
	) name9169 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w11637_,
		_w12356_,
		_w13217_
	);
	LUT2 #(
		.INIT('h2)
	) name9170 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001 ,
		_w11656_,
		_w13218_
	);
	LUT3 #(
		.INIT('h01)
	) name9171 (
		_w9946_,
		_w11659_,
		_w13218_,
		_w13219_
	);
	LUT4 #(
		.INIT('hfd00)
	) name9172 (
		_w11655_,
		_w12736_,
		_w12737_,
		_w13219_,
		_w13220_
	);
	LUT2 #(
		.INIT('h1)
	) name9173 (
		_w13217_,
		_w13220_,
		_w13221_
	);
	LUT3 #(
		.INIT('h01)
	) name9174 (
		_w11550_,
		_w11553_,
		_w11475_,
		_w13222_
	);
	LUT3 #(
		.INIT('h20)
	) name9175 (
		_w11441_,
		_w12645_,
		_w13222_,
		_w13223_
	);
	LUT2 #(
		.INIT('h8)
	) name9176 (
		_w12448_,
		_w13223_,
		_w13224_
	);
	LUT4 #(
		.INIT('h7707)
	) name9177 (
		_w11522_,
		_w11449_,
		_w11855_,
		_w11953_,
		_w13225_
	);
	LUT3 #(
		.INIT('he0)
	) name9178 (
		_w11393_,
		_w11589_,
		_w12767_,
		_w13226_
	);
	LUT2 #(
		.INIT('h4)
	) name9179 (
		_w11492_,
		_w11864_,
		_w13227_
	);
	LUT3 #(
		.INIT('h10)
	) name9180 (
		_w13226_,
		_w13227_,
		_w13225_,
		_w13228_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name9181 (
		_w11587_,
		_w11530_,
		_w11458_,
		_w12639_,
		_w13229_
	);
	LUT4 #(
		.INIT('h3f2a)
	) name9182 (
		_w11534_,
		_w11409_,
		_w11495_,
		_w11844_,
		_w13230_
	);
	LUT2 #(
		.INIT('h8)
	) name9183 (
		_w13229_,
		_w13230_,
		_w13231_
	);
	LUT3 #(
		.INIT('h80)
	) name9184 (
		_w13180_,
		_w13228_,
		_w13231_,
		_w13232_
	);
	LUT3 #(
		.INIT('h04)
	) name9185 (
		_w11536_,
		_w11386_,
		_w11953_,
		_w13233_
	);
	LUT3 #(
		.INIT('hc8)
	) name9186 (
		_w11555_,
		_w11469_,
		_w11888_,
		_w13234_
	);
	LUT3 #(
		.INIT('ha8)
	) name9187 (
		_w11499_,
		_w11435_,
		_w12455_,
		_w13235_
	);
	LUT3 #(
		.INIT('h01)
	) name9188 (
		_w13234_,
		_w13235_,
		_w13233_,
		_w13236_
	);
	LUT4 #(
		.INIT('h0080)
	) name9189 (
		_w11389_,
		_w11386_,
		_w11476_,
		_w11464_,
		_w13237_
	);
	LUT4 #(
		.INIT('h8000)
	) name9190 (
		_w11389_,
		_w11385_,
		_w11445_,
		_w11458_,
		_w13238_
	);
	LUT4 #(
		.INIT('h4000)
	) name9191 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11406_,
		_w11491_,
		_w13239_
	);
	LUT3 #(
		.INIT('h01)
	) name9192 (
		_w13238_,
		_w13239_,
		_w13237_,
		_w13240_
	);
	LUT2 #(
		.INIT('h8)
	) name9193 (
		_w11415_,
		_w11838_,
		_w13241_
	);
	LUT4 #(
		.INIT('ha820)
	) name9194 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001 ,
		_w13242_
	);
	LUT3 #(
		.INIT('h07)
	) name9195 (
		_w11578_,
		_w11962_,
		_w13242_,
		_w13243_
	);
	LUT4 #(
		.INIT('h0700)
	) name9196 (
		_w11558_,
		_w11465_,
		_w13241_,
		_w13243_,
		_w13244_
	);
	LUT3 #(
		.INIT('hc8)
	) name9197 (
		_w11588_,
		_w11874_,
		_w12496_,
		_w13245_
	);
	LUT3 #(
		.INIT('ha8)
	) name9198 (
		_w11860_,
		_w11973_,
		_w11974_,
		_w13246_
	);
	LUT4 #(
		.INIT('h1000)
	) name9199 (
		_w13245_,
		_w13246_,
		_w13240_,
		_w13244_,
		_w13247_
	);
	LUT2 #(
		.INIT('h8)
	) name9200 (
		_w13236_,
		_w13247_,
		_w13248_
	);
	LUT4 #(
		.INIT('h8000)
	) name9201 (
		_w12451_,
		_w13224_,
		_w13232_,
		_w13248_,
		_w13249_
	);
	LUT4 #(
		.INIT('h7020)
	) name9202 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11315_,
		_w11830_,
		_w13249_,
		_w13250_
	);
	LUT4 #(
		.INIT('h5545)
	) name9203 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w13251_
	);
	LUT2 #(
		.INIT('h1)
	) name9204 (
		_w13250_,
		_w13251_,
		_w13252_
	);
	LUT4 #(
		.INIT('h7020)
	) name9205 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11315_,
		_w11329_,
		_w13249_,
		_w13253_
	);
	LUT2 #(
		.INIT('h1)
	) name9206 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001 ,
		_w11329_,
		_w13254_
	);
	LUT2 #(
		.INIT('h1)
	) name9207 (
		_w13253_,
		_w13254_,
		_w13255_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9208 (
		\core_c_dec_Call_Ed_reg/P0001 ,
		_w4160_,
		_w4158_,
		_w4167_,
		_w13256_
	);
	LUT2 #(
		.INIT('h1)
	) name9209 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w13257_
	);
	LUT4 #(
		.INIT('h2322)
	) name9210 (
		_w4971_,
		_w11600_,
		_w13256_,
		_w13257_,
		_w13258_
	);
	LUT2 #(
		.INIT('h4)
	) name9211 (
		\core_c_psq_pcstk_ptr_reg[4]/NET0131 ,
		_w4114_,
		_w13259_
	);
	LUT3 #(
		.INIT('hba)
	) name9212 (
		\core_c_psq_SSTAT_reg[1]/NET0131 ,
		_w13258_,
		_w13259_,
		_w13260_
	);
	LUT3 #(
		.INIT('ha8)
	) name9213 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w11313_,
		_w11314_,
		_w13261_
	);
	LUT4 #(
		.INIT('h0f08)
	) name9214 (
		_w11333_,
		_w11397_,
		_w11494_,
		_w11519_,
		_w13262_
	);
	LUT4 #(
		.INIT('hfac8)
	) name9215 (
		_w11592_,
		_w11954_,
		_w11958_,
		_w12506_,
		_w13263_
	);
	LUT2 #(
		.INIT('h8)
	) name9216 (
		_w11424_,
		_w11860_,
		_w13264_
	);
	LUT3 #(
		.INIT('he0)
	) name9217 (
		_w11393_,
		_w11589_,
		_w11864_,
		_w13265_
	);
	LUT3 #(
		.INIT('h10)
	) name9218 (
		_w13264_,
		_w13265_,
		_w13263_,
		_w13266_
	);
	LUT4 #(
		.INIT('ha820)
	) name9219 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001 ,
		_w13267_
	);
	LUT3 #(
		.INIT('h0b)
	) name9220 (
		_w11593_,
		_w11855_,
		_w13267_,
		_w13268_
	);
	LUT2 #(
		.INIT('h8)
	) name9221 (
		_w11571_,
		_w13268_,
		_w13269_
	);
	LUT3 #(
		.INIT('h40)
	) name9222 (
		_w13262_,
		_w13266_,
		_w13269_,
		_w13270_
	);
	LUT2 #(
		.INIT('h2)
	) name9223 (
		_w11872_,
		_w11957_,
		_w13271_
	);
	LUT3 #(
		.INIT('he0)
	) name9224 (
		_w11552_,
		_w11474_,
		_w11841_,
		_w13272_
	);
	LUT4 #(
		.INIT('h5554)
	) name9225 (
		_w11386_,
		_w11581_,
		_w13271_,
		_w13272_,
		_w13273_
	);
	LUT3 #(
		.INIT('hc8)
	) name9226 (
		_w11572_,
		_w11532_,
		_w11831_,
		_w13274_
	);
	LUT3 #(
		.INIT('h02)
	) name9227 (
		_w11386_,
		_w11506_,
		_w11957_,
		_w13275_
	);
	LUT3 #(
		.INIT('h04)
	) name9228 (
		_w11536_,
		_w11386_,
		_w11593_,
		_w13276_
	);
	LUT3 #(
		.INIT('h01)
	) name9229 (
		_w13275_,
		_w13276_,
		_w13274_,
		_w13277_
	);
	LUT3 #(
		.INIT('hc8)
	) name9230 (
		_w11547_,
		_w11469_,
		_w11976_,
		_w13278_
	);
	LUT4 #(
		.INIT('h0a08)
	) name9231 (
		_w11386_,
		_w11552_,
		_w11483_,
		_w11474_,
		_w13279_
	);
	LUT3 #(
		.INIT('he0)
	) name9232 (
		_w11420_,
		_w11421_,
		_w11449_,
		_w13280_
	);
	LUT4 #(
		.INIT('h0002)
	) name9233 (
		_w11969_,
		_w13278_,
		_w13279_,
		_w13280_,
		_w13281_
	);
	LUT3 #(
		.INIT('h40)
	) name9234 (
		_w13273_,
		_w13277_,
		_w13281_,
		_w13282_
	);
	LUT4 #(
		.INIT('h2333)
	) name9235 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w13261_,
		_w13270_,
		_w13282_,
		_w13283_
	);
	LUT3 #(
		.INIT('he2)
	) name9236 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001 ,
		_w11946_,
		_w13283_,
		_w13284_
	);
	LUT3 #(
		.INIT('hc8)
	) name9237 (
		_w11555_,
		_w11841_,
		_w11888_,
		_w13285_
	);
	LUT3 #(
		.INIT('ha8)
	) name9238 (
		_w11484_,
		_w11522_,
		_w11523_,
		_w13286_
	);
	LUT3 #(
		.INIT('hc8)
	) name9239 (
		_w11409_,
		_w11465_,
		_w11896_,
		_w13287_
	);
	LUT4 #(
		.INIT('h4440)
	) name9240 (
		_w11536_,
		_w11386_,
		_w11552_,
		_w11474_,
		_w13288_
	);
	LUT4 #(
		.INIT('h0001)
	) name9241 (
		_w13285_,
		_w13286_,
		_w13287_,
		_w13288_,
		_w13289_
	);
	LUT4 #(
		.INIT('h4000)
	) name9242 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11382_,
		_w12504_,
		_w13290_
	);
	LUT4 #(
		.INIT('h4000)
	) name9243 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11382_,
		_w12505_,
		_w13291_
	);
	LUT4 #(
		.INIT('h4000)
	) name9244 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11401_,
		_w11358_,
		_w11855_,
		_w13292_
	);
	LUT4 #(
		.INIT('h8000)
	) name9245 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11406_,
		_w11439_,
		_w13293_
	);
	LUT4 #(
		.INIT('h0001)
	) name9246 (
		_w13290_,
		_w13291_,
		_w13292_,
		_w13293_,
		_w13294_
	);
	LUT3 #(
		.INIT('h80)
	) name9247 (
		_w11473_,
		_w11389_,
		_w11855_,
		_w13295_
	);
	LUT3 #(
		.INIT('h80)
	) name9248 (
		_w11389_,
		_w11445_,
		_w11838_,
		_w13296_
	);
	LUT3 #(
		.INIT('h08)
	) name9249 (
		_w11389_,
		_w11476_,
		_w12639_,
		_w13297_
	);
	LUT3 #(
		.INIT('h01)
	) name9250 (
		_w13296_,
		_w13297_,
		_w13295_,
		_w13298_
	);
	LUT4 #(
		.INIT('ha820)
	) name9251 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001 ,
		_w13299_
	);
	LUT3 #(
		.INIT('h0d)
	) name9252 (
		_w11429_,
		_w12506_,
		_w13299_,
		_w13300_
	);
	LUT2 #(
		.INIT('h4)
	) name9253 (
		_w12472_,
		_w13300_,
		_w13301_
	);
	LUT3 #(
		.INIT('h80)
	) name9254 (
		_w13298_,
		_w13301_,
		_w13294_,
		_w13302_
	);
	LUT3 #(
		.INIT('hc8)
	) name9255 (
		_w11435_,
		_w11469_,
		_w12455_,
		_w13303_
	);
	LUT3 #(
		.INIT('ha8)
	) name9256 (
		_w11874_,
		_w11973_,
		_w11974_,
		_w13304_
	);
	LUT2 #(
		.INIT('h1)
	) name9257 (
		_w13303_,
		_w13304_,
		_w13305_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9258 (
		_w11530_,
		_w11864_,
		_w11957_,
		_w12767_,
		_w13306_
	);
	LUT4 #(
		.INIT('h153f)
	) name9259 (
		_w11588_,
		_w11587_,
		_w11449_,
		_w11872_,
		_w13307_
	);
	LUT2 #(
		.INIT('h8)
	) name9260 (
		_w13306_,
		_w13307_,
		_w13308_
	);
	LUT3 #(
		.INIT('he0)
	) name9261 (
		_w11393_,
		_w11589_,
		_w11962_,
		_w13309_
	);
	LUT3 #(
		.INIT('he0)
	) name9262 (
		_w11393_,
		_w11589_,
		_w11861_,
		_w13310_
	);
	LUT2 #(
		.INIT('h8)
	) name9263 (
		_w11558_,
		_w11507_,
		_w13311_
	);
	LUT4 #(
		.INIT('h0002)
	) name9264 (
		_w11408_,
		_w13309_,
		_w13310_,
		_w13311_,
		_w13312_
	);
	LUT4 #(
		.INIT('h8000)
	) name9265 (
		_w13308_,
		_w13312_,
		_w13302_,
		_w13305_,
		_w13313_
	);
	LUT4 #(
		.INIT('h8000)
	) name9266 (
		_w12449_,
		_w12451_,
		_w13289_,
		_w13313_,
		_w13314_
	);
	LUT4 #(
		.INIT('h4c08)
	) name9267 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w11946_,
		_w12673_,
		_w13314_,
		_w13315_
	);
	LUT4 #(
		.INIT('h5545)
	) name9268 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001 ,
		_w9453_,
		_w9894_,
		_w11945_,
		_w13316_
	);
	LUT2 #(
		.INIT('h1)
	) name9269 (
		_w13315_,
		_w13316_,
		_w13317_
	);
	LUT3 #(
		.INIT('he2)
	) name9270 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001 ,
		_w12048_,
		_w13283_,
		_w13318_
	);
	LUT4 #(
		.INIT('h4c08)
	) name9271 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12048_,
		_w12673_,
		_w13314_,
		_w13319_
	);
	LUT2 #(
		.INIT('h1)
	) name9272 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001 ,
		_w12048_,
		_w13320_
	);
	LUT2 #(
		.INIT('h1)
	) name9273 (
		_w13319_,
		_w13320_,
		_w13321_
	);
	LUT2 #(
		.INIT('h8)
	) name9274 (
		\core_c_psq_PCS_reg[14]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w13322_
	);
	LUT4 #(
		.INIT('h028a)
	) name9275 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		_w13323_
	);
	LUT4 #(
		.INIT('h4000)
	) name9276 (
		\core_c_psq_SRST_reg/P0001 ,
		_w4065_,
		_w4066_,
		_w13323_,
		_w13324_
	);
	LUT2 #(
		.INIT('h1)
	) name9277 (
		_w13322_,
		_w13324_,
		_w13325_
	);
	LUT2 #(
		.INIT('he)
	) name9278 (
		_w13322_,
		_w13324_,
		_w13326_
	);
	LUT3 #(
		.INIT('h80)
	) name9279 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w13327_
	);
	LUT3 #(
		.INIT('h07)
	) name9280 (
		_w4461_,
		_w4498_,
		_w13327_,
		_w13328_
	);
	LUT4 #(
		.INIT('h4000)
	) name9281 (
		\core_c_psq_Eqend_D_reg/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w13329_
	);
	LUT2 #(
		.INIT('h2)
	) name9282 (
		_w4102_,
		_w13329_,
		_w13330_
	);
	LUT2 #(
		.INIT('h4)
	) name9283 (
		_w13328_,
		_w13330_,
		_w13331_
	);
	LUT4 #(
		.INIT('h2000)
	) name9284 (
		\core_c_dec_MpopLP_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w13332_
	);
	LUT2 #(
		.INIT('h8)
	) name9285 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w13333_
	);
	LUT3 #(
		.INIT('h80)
	) name9286 (
		_w5028_,
		_w5045_,
		_w13333_,
		_w13334_
	);
	LUT4 #(
		.INIT('h070f)
	) name9287 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w8174_,
		_w13332_,
		_w13334_,
		_w13335_
	);
	LUT2 #(
		.INIT('h2)
	) name9288 (
		_w4102_,
		_w13335_,
		_w13336_
	);
	LUT4 #(
		.INIT('h2000)
	) name9289 (
		\core_c_dec_Call_Ed_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w13337_
	);
	LUT2 #(
		.INIT('h1)
	) name9290 (
		_w5029_,
		_w12917_,
		_w13338_
	);
	LUT3 #(
		.INIT('h15)
	) name9291 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w5046_,
		_w12916_,
		_w13339_
	);
	LUT4 #(
		.INIT('h3331)
	) name9292 (
		_w8174_,
		_w13337_,
		_w13338_,
		_w13339_,
		_w13340_
	);
	LUT2 #(
		.INIT('h2)
	) name9293 (
		_w4102_,
		_w13340_,
		_w13341_
	);
	LUT4 #(
		.INIT('h2000)
	) name9294 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w13342_
	);
	LUT4 #(
		.INIT('haa08)
	) name9295 (
		_w4102_,
		_w4834_,
		_w11921_,
		_w13342_,
		_w13343_
	);
	LUT2 #(
		.INIT('h6)
	) name9296 (
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w12605_,
		_w13344_
	);
	LUT2 #(
		.INIT('h4)
	) name9297 (
		_w9413_,
		_w13344_,
		_w13345_
	);
	LUT3 #(
		.INIT('h80)
	) name9298 (
		_w5658_,
		_w9431_,
		_w12824_,
		_w13346_
	);
	LUT4 #(
		.INIT('hba00)
	) name9299 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13346_,
		_w13347_
	);
	LUT4 #(
		.INIT('h0100)
	) name9300 (
		_w7710_,
		_w7906_,
		_w8043_,
		_w13347_,
		_w13348_
	);
	LUT4 #(
		.INIT('h4500)
	) name9301 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13346_,
		_w13349_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name9302 (
		\bdma_BCTL_reg[7]/NET0131 ,
		_w5658_,
		_w9431_,
		_w12824_,
		_w13350_
	);
	LUT2 #(
		.INIT('h1)
	) name9303 (
		_w13349_,
		_w13350_,
		_w13351_
	);
	LUT2 #(
		.INIT('hb)
	) name9304 (
		_w13348_,
		_w13351_,
		_w13352_
	);
	LUT4 #(
		.INIT('h4500)
	) name9305 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13346_,
		_w13353_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name9306 (
		\bdma_BCTL_reg[6]/NET0131 ,
		_w5658_,
		_w9431_,
		_w12824_,
		_w13354_
	);
	LUT2 #(
		.INIT('h1)
	) name9307 (
		_w13353_,
		_w13354_,
		_w13355_
	);
	LUT2 #(
		.INIT('hb)
	) name9308 (
		_w13348_,
		_w13355_,
		_w13356_
	);
	LUT4 #(
		.INIT('h4500)
	) name9309 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13346_,
		_w13357_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name9310 (
		\bdma_BCTL_reg[5]/NET0131 ,
		_w5658_,
		_w9431_,
		_w12824_,
		_w13358_
	);
	LUT2 #(
		.INIT('h1)
	) name9311 (
		_w13357_,
		_w13358_,
		_w13359_
	);
	LUT2 #(
		.INIT('hb)
	) name9312 (
		_w13348_,
		_w13359_,
		_w13360_
	);
	LUT4 #(
		.INIT('h1555)
	) name9313 (
		\bdma_BCTL_reg[4]/NET0131 ,
		_w5658_,
		_w9431_,
		_w12824_,
		_w13361_
	);
	LUT2 #(
		.INIT('h1)
	) name9314 (
		_w13347_,
		_w13361_,
		_w13362_
	);
	LUT2 #(
		.INIT('he)
	) name9315 (
		_w13348_,
		_w13362_,
		_w13363_
	);
	LUT2 #(
		.INIT('h6)
	) name9316 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_OUTcnt_reg[1]/NET0131 ,
		_w13364_
	);
	LUT4 #(
		.INIT('hbf00)
	) name9317 (
		_w12254_,
		_w12258_,
		_w12263_,
		_w13364_,
		_w13365_
	);
	LUT3 #(
		.INIT('h80)
	) name9318 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13366_
	);
	LUT4 #(
		.INIT('h1400)
	) name9319 (
		\PIO_oe[8]_pad ,
		\pio_PIO_RES_OUT_reg[8]/P0001 ,
		\pio_PIO_RES_reg[8]/NET0131 ,
		\pio_pmask_reg_DO_reg[8]/NET0131 ,
		_w13367_
	);
	LUT2 #(
		.INIT('h1)
	) name9320 (
		\pio_PINT_reg[8]/NET0131 ,
		_w13367_,
		_w13368_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9321 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13368_,
		_w13369_
	);
	LUT3 #(
		.INIT('h0b)
	) name9322 (
		_w6758_,
		_w13366_,
		_w13369_,
		_w13370_
	);
	LUT2 #(
		.INIT('he)
	) name9323 (
		\tm_WR_TSR_KEEP_TO_TMCLK_p_reg/NET0131 ,
		\tm_WR_TSR_p_reg/P0001 ,
		_w13371_
	);
	LUT2 #(
		.INIT('h6)
	) name9324 (
		\emc_RWcnt_reg[3]/P0001 ,
		_w12710_,
		_w13372_
	);
	LUT4 #(
		.INIT('h1000)
	) name9325 (
		_w12705_,
		_w12704_,
		_w12708_,
		_w13372_,
		_w13373_
	);
	LUT4 #(
		.INIT('hf078)
	) name9326 (
		\emc_RWcnt_reg[0]/P0001 ,
		\emc_RWcnt_reg[1]/P0001 ,
		\emc_RWcnt_reg[2]/P0001 ,
		_w12709_,
		_w13374_
	);
	LUT4 #(
		.INIT('h1000)
	) name9327 (
		_w12705_,
		_w12704_,
		_w12708_,
		_w13374_,
		_w13375_
	);
	LUT3 #(
		.INIT('hc6)
	) name9328 (
		\emc_RWcnt_reg[0]/P0001 ,
		\emc_RWcnt_reg[1]/P0001 ,
		_w12709_,
		_w13376_
	);
	LUT4 #(
		.INIT('h1000)
	) name9329 (
		_w12705_,
		_w12704_,
		_w12708_,
		_w13376_,
		_w13377_
	);
	LUT2 #(
		.INIT('h9)
	) name9330 (
		\emc_RWcnt_reg[0]/P0001 ,
		_w12709_,
		_w13378_
	);
	LUT4 #(
		.INIT('h1000)
	) name9331 (
		_w12705_,
		_w12704_,
		_w12708_,
		_w13378_,
		_w13379_
	);
	LUT4 #(
		.INIT('h0004)
	) name9332 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MACop_E_reg/P0001 ,
		_w4971_,
		_w9453_,
		_w13380_
	);
	LUT4 #(
		.INIT('hfff8)
	) name9333 (
		_w9910_,
		_w11802_,
		_w12111_,
		_w13380_,
		_w13381_
	);
	LUT3 #(
		.INIT('h32)
	) name9334 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13382_
	);
	LUT3 #(
		.INIT('h01)
	) name9335 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13383_
	);
	LUT4 #(
		.INIT('h0004)
	) name9336 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[9]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13384_
	);
	LUT2 #(
		.INIT('h4)
	) name9337 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w13385_
	);
	LUT2 #(
		.INIT('h1)
	) name9338 (
		_w13384_,
		_w13385_,
		_w13386_
	);
	LUT4 #(
		.INIT('h10ff)
	) name9339 (
		_w7140_,
		_w7240_,
		_w13382_,
		_w13386_,
		_w13387_
	);
	LUT4 #(
		.INIT('h0004)
	) name9340 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[8]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13388_
	);
	LUT2 #(
		.INIT('h1)
	) name9341 (
		_w13385_,
		_w13388_,
		_w13389_
	);
	LUT4 #(
		.INIT('h10ff)
	) name9342 (
		_w7465_,
		_w7565_,
		_w13382_,
		_w13389_,
		_w13390_
	);
	LUT4 #(
		.INIT('h4500)
	) name9343 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13382_,
		_w13391_
	);
	LUT4 #(
		.INIT('h0004)
	) name9344 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[7]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13392_
	);
	LUT2 #(
		.INIT('h1)
	) name9345 (
		_w13385_,
		_w13392_,
		_w13393_
	);
	LUT2 #(
		.INIT('hb)
	) name9346 (
		_w13391_,
		_w13393_,
		_w13394_
	);
	LUT4 #(
		.INIT('h1400)
	) name9347 (
		\PIO_oe[9]_pad ,
		\pio_PIO_RES_OUT_reg[9]/P0001 ,
		\pio_PIO_RES_reg[9]/NET0131 ,
		\pio_pmask_reg_DO_reg[9]/NET0131 ,
		_w13395_
	);
	LUT2 #(
		.INIT('h1)
	) name9348 (
		\pio_PINT_reg[9]/NET0131 ,
		_w13395_,
		_w13396_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9349 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13396_,
		_w13397_
	);
	LUT3 #(
		.INIT('h0b)
	) name9350 (
		_w5760_,
		_w13366_,
		_w13397_,
		_w13398_
	);
	LUT4 #(
		.INIT('hcfcb)
	) name9351 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13399_
	);
	LUT4 #(
		.INIT('h10ff)
	) name9352 (
		_w8798_,
		_w8801_,
		_w13382_,
		_w13399_,
		_w13400_
	);
	LUT4 #(
		.INIT('h0004)
	) name9353 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[13]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13401_
	);
	LUT2 #(
		.INIT('h1)
	) name9354 (
		_w13385_,
		_w13401_,
		_w13402_
	);
	LUT3 #(
		.INIT('h8f)
	) name9355 (
		_w5760_,
		_w13382_,
		_w13402_,
		_w13403_
	);
	LUT4 #(
		.INIT('h0004)
	) name9356 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[14]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13404_
	);
	LUT2 #(
		.INIT('h1)
	) name9357 (
		_w13385_,
		_w13404_,
		_w13405_
	);
	LUT4 #(
		.INIT('h10ff)
	) name9358 (
		_w8757_,
		_w8760_,
		_w13382_,
		_w13405_,
		_w13406_
	);
	LUT4 #(
		.INIT('h0004)
	) name9359 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[12]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13407_
	);
	LUT2 #(
		.INIT('h1)
	) name9360 (
		_w13385_,
		_w13407_,
		_w13408_
	);
	LUT3 #(
		.INIT('h8f)
	) name9361 (
		_w6758_,
		_w13382_,
		_w13408_,
		_w13409_
	);
	LUT4 #(
		.INIT('h0004)
	) name9362 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[11]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13410_
	);
	LUT2 #(
		.INIT('h1)
	) name9363 (
		_w13385_,
		_w13410_,
		_w13411_
	);
	LUT4 #(
		.INIT('h10ff)
	) name9364 (
		_w6263_,
		_w6362_,
		_w13382_,
		_w13411_,
		_w13412_
	);
	LUT4 #(
		.INIT('h0004)
	) name9365 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[10]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w13413_
	);
	LUT2 #(
		.INIT('h1)
	) name9366 (
		_w13385_,
		_w13413_,
		_w13414_
	);
	LUT4 #(
		.INIT('h10ff)
	) name9367 (
		_w5937_,
		_w6038_,
		_w13382_,
		_w13414_,
		_w13415_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name9368 (
		\core_c_dec_updMF_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001 ,
		_w9453_,
		_w9894_,
		_w13416_
	);
	LUT4 #(
		.INIT('h7000)
	) name9369 (
		_w12328_,
		_w12381_,
		_w12386_,
		_w13091_,
		_w13417_
	);
	LUT2 #(
		.INIT('he)
	) name9370 (
		_w13416_,
		_w13417_,
		_w13418_
	);
	LUT4 #(
		.INIT('h2227)
	) name9371 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w13419_
	);
	LUT2 #(
		.INIT('h8)
	) name9372 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w13420_
	);
	LUT3 #(
		.INIT('hba)
	) name9373 (
		\sport0_rxctl_RSreq_reg/NET0131 ,
		_w13419_,
		_w13420_,
		_w13421_
	);
	LUT2 #(
		.INIT('h2)
	) name9374 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001 ,
		_w13168_,
		_w13422_
	);
	LUT4 #(
		.INIT('h7000)
	) name9375 (
		_w12328_,
		_w12381_,
		_w12386_,
		_w13168_,
		_w13423_
	);
	LUT2 #(
		.INIT('he)
	) name9376 (
		_w13422_,
		_w13423_,
		_w13424_
	);
	LUT4 #(
		.INIT('hb41e)
	) name9377 (
		\IRFS1_pad ,
		\T_RFS1_pad ,
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w9352_,
		_w13425_
	);
	LUT2 #(
		.INIT('h4)
	) name9378 (
		\sport1_cfg_RFSgi_d_reg/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w13426_
	);
	LUT2 #(
		.INIT('h8)
	) name9379 (
		_w13425_,
		_w13426_,
		_w13427_
	);
	LUT4 #(
		.INIT('hb41e)
	) name9380 (
		\IRFS0_pad ,
		\T_RFS0_pad ,
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w9350_,
		_w13428_
	);
	LUT2 #(
		.INIT('h4)
	) name9381 (
		\sport0_cfg_RFSgi_d_reg/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w13429_
	);
	LUT2 #(
		.INIT('h8)
	) name9382 (
		_w13428_,
		_w13429_,
		_w13430_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9383 (
		\core_c_psq_Iact_E_reg[9]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w13431_
	);
	LUT3 #(
		.INIT('h70)
	) name9384 (
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_T_IRQ2_s1_reg/P0001 ,
		\core_c_psq_irq2_de_OUT_reg/P0001 ,
		_w13432_
	);
	LUT3 #(
		.INIT('ha8)
	) name9385 (
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_IFC_reg[15]/NET0131 ,
		\core_c_psq_Iflag_reg[9]/NET0131 ,
		_w13433_
	);
	LUT2 #(
		.INIT('h1)
	) name9386 (
		_w13432_,
		_w13433_,
		_w13434_
	);
	LUT4 #(
		.INIT('h0057)
	) name9387 (
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_IFC_reg[7]/NET0131 ,
		_w13431_,
		_w13434_,
		_w13435_
	);
	LUT2 #(
		.INIT('h4)
	) name9388 (
		\core_c_psq_ICNTL_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_irq1_de_OUT_reg/P0001 ,
		_w13436_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9389 (
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w13437_
	);
	LUT4 #(
		.INIT('h00ba)
	) name9390 (
		\core_c_psq_IFC_reg[10]/NET0131 ,
		\core_c_psq_T_IRQ1_s1_reg/P0001 ,
		\core_c_psq_irq1_de_OUT_reg/P0001 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w13438_
	);
	LUT3 #(
		.INIT('ha8)
	) name9391 (
		\core_c_psq_ICNTL_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_Iflag_reg[12]/NET0131 ,
		_w13438_,
		_w13439_
	);
	LUT4 #(
		.INIT('hcdcc)
	) name9392 (
		\core_c_psq_IFC_reg[2]/NET0131 ,
		_w13436_,
		_w13437_,
		_w13439_,
		_w13440_
	);
	LUT2 #(
		.INIT('h4)
	) name9393 (
		\core_c_psq_ICNTL_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_irq0_de_OUT_reg/P0001 ,
		_w13441_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9394 (
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w13442_
	);
	LUT4 #(
		.INIT('h00ba)
	) name9395 (
		\core_c_psq_IFC_reg[9]/NET0131 ,
		\core_c_psq_T_IRQ0_s1_reg/P0001 ,
		\core_c_psq_irq0_de_OUT_reg/P0001 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w13443_
	);
	LUT3 #(
		.INIT('ha8)
	) name9396 (
		\core_c_psq_ICNTL_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_Iflag_reg[11]/NET0131 ,
		_w13443_,
		_w13444_
	);
	LUT4 #(
		.INIT('hcdcc)
	) name9397 (
		\core_c_psq_IFC_reg[1]/NET0131 ,
		_w13441_,
		_w13442_,
		_w13444_,
		_w13445_
	);
	LUT4 #(
		.INIT('hbf00)
	) name9398 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4102_,
		_w13446_
	);
	LUT2 #(
		.INIT('h8)
	) name9399 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w13447_
	);
	LUT3 #(
		.INIT('h0e)
	) name9400 (
		_w5047_,
		_w12296_,
		_w13447_,
		_w13448_
	);
	LUT4 #(
		.INIT('h8c80)
	) name9401 (
		\core_c_dec_updSR_E_reg/P0001 ,
		_w4102_,
		_w4104_,
		_w13448_,
		_w13449_
	);
	LUT4 #(
		.INIT('h4000)
	) name9402 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w5028_,
		_w5044_,
		_w12393_,
		_w13450_
	);
	LUT4 #(
		.INIT('h2000)
	) name9403 (
		\core_c_dec_Nseq_Ed_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w13451_
	);
	LUT4 #(
		.INIT('h050d)
	) name9404 (
		_w8174_,
		_w13338_,
		_w13451_,
		_w13450_,
		_w13452_
	);
	LUT2 #(
		.INIT('h2)
	) name9405 (
		_w4102_,
		_w13452_,
		_w13453_
	);
	LUT3 #(
		.INIT('h40)
	) name9406 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w8174_,
		_w13450_,
		_w13454_
	);
	LUT4 #(
		.INIT('h2000)
	) name9407 (
		\core_c_dec_Nrti_Ed_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w13455_
	);
	LUT3 #(
		.INIT('h0d)
	) name9408 (
		_w8174_,
		_w13338_,
		_w13455_,
		_w13456_
	);
	LUT3 #(
		.INIT('h8a)
	) name9409 (
		_w4102_,
		_w13454_,
		_w13456_,
		_w13457_
	);
	LUT4 #(
		.INIT('h1400)
	) name9410 (
		\PIO_oe[5]_pad ,
		\pio_PIO_RES_OUT_reg[5]/P0001 ,
		\pio_PIO_RES_reg[5]/NET0131 ,
		\pio_pmask_reg_DO_reg[5]/NET0131 ,
		_w13458_
	);
	LUT2 #(
		.INIT('h1)
	) name9411 (
		\pio_PINT_reg[5]/NET0131 ,
		_w13458_,
		_w13459_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9412 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13459_,
		_w13460_
	);
	LUT4 #(
		.INIT('hba00)
	) name9413 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13366_,
		_w13461_
	);
	LUT2 #(
		.INIT('h1)
	) name9414 (
		_w13460_,
		_w13461_,
		_w13462_
	);
	LUT4 #(
		.INIT('h1400)
	) name9415 (
		\PIO_oe[4]_pad ,
		\pio_PIO_RES_OUT_reg[4]/P0001 ,
		\pio_PIO_RES_reg[4]/NET0131 ,
		\pio_pmask_reg_DO_reg[4]/NET0131 ,
		_w13463_
	);
	LUT2 #(
		.INIT('h1)
	) name9416 (
		\pio_PINT_reg[4]/NET0131 ,
		_w13463_,
		_w13464_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9417 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13464_,
		_w13465_
	);
	LUT4 #(
		.INIT('hba00)
	) name9418 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13366_,
		_w13466_
	);
	LUT2 #(
		.INIT('h1)
	) name9419 (
		_w13465_,
		_w13466_,
		_w13467_
	);
	LUT4 #(
		.INIT('h1400)
	) name9420 (
		\PIO_oe[11]_pad ,
		\pio_PIO_RES_OUT_reg[11]/P0001 ,
		\pio_PIO_RES_reg[11]/NET0131 ,
		\pio_pmask_reg_DO_reg[11]/NET0131 ,
		_w13468_
	);
	LUT2 #(
		.INIT('h1)
	) name9421 (
		\pio_PINT_reg[11]/NET0131 ,
		_w13468_,
		_w13469_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9422 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13469_,
		_w13470_
	);
	LUT4 #(
		.INIT('h001f)
	) name9423 (
		_w8798_,
		_w8801_,
		_w13366_,
		_w13470_,
		_w13471_
	);
	LUT4 #(
		.INIT('h1400)
	) name9424 (
		\PIO_oe[2]_pad ,
		\pio_PIO_RES_OUT_reg[2]/P0001 ,
		\pio_PIO_RES_reg[2]/NET0131 ,
		\pio_pmask_reg_DO_reg[2]/NET0131 ,
		_w13472_
	);
	LUT2 #(
		.INIT('h1)
	) name9425 (
		\pio_PINT_reg[2]/NET0131 ,
		_w13472_,
		_w13473_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9426 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13473_,
		_w13474_
	);
	LUT4 #(
		.INIT('hba00)
	) name9427 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13366_,
		_w13475_
	);
	LUT2 #(
		.INIT('h1)
	) name9428 (
		_w13474_,
		_w13475_,
		_w13476_
	);
	LUT4 #(
		.INIT('h1400)
	) name9429 (
		\PIO_oe[10]_pad ,
		\pio_PIO_RES_OUT_reg[10]/P0001 ,
		\pio_PIO_RES_reg[10]/NET0131 ,
		\pio_pmask_reg_DO_reg[10]/NET0131 ,
		_w13477_
	);
	LUT2 #(
		.INIT('h1)
	) name9430 (
		\pio_PINT_reg[10]/NET0131 ,
		_w13477_,
		_w13478_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9431 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13478_,
		_w13479_
	);
	LUT4 #(
		.INIT('h001f)
	) name9432 (
		_w8757_,
		_w8760_,
		_w13366_,
		_w13479_,
		_w13480_
	);
	LUT4 #(
		.INIT('h1400)
	) name9433 (
		\PIO_oe[0]_pad ,
		\pio_PIO_RES_OUT_reg[0]/P0001 ,
		\pio_PIO_RES_reg[0]/NET0131 ,
		\pio_pmask_reg_DO_reg[0]/NET0131 ,
		_w13481_
	);
	LUT2 #(
		.INIT('h1)
	) name9434 (
		\pio_PINT_reg[0]/NET0131 ,
		_w13481_,
		_w13482_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9435 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13482_,
		_w13483_
	);
	LUT4 #(
		.INIT('hba00)
	) name9436 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13366_,
		_w13484_
	);
	LUT2 #(
		.INIT('h1)
	) name9437 (
		_w13483_,
		_w13484_,
		_w13485_
	);
	LUT4 #(
		.INIT('hc444)
	) name9438 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		_w4073_,
		_w4084_,
		_w13486_
	);
	LUT3 #(
		.INIT('h04)
	) name9439 (
		_w12274_,
		_w12276_,
		_w12277_,
		_w13487_
	);
	LUT4 #(
		.INIT('hf2f0)
	) name9440 (
		_w12271_,
		_w12272_,
		_w13486_,
		_w13487_,
		_w13488_
	);
	LUT4 #(
		.INIT('h1400)
	) name9441 (
		\PIO_oe[1]_pad ,
		\pio_PIO_RES_OUT_reg[1]/P0001 ,
		\pio_PIO_RES_reg[1]/NET0131 ,
		\pio_pmask_reg_DO_reg[1]/NET0131 ,
		_w13489_
	);
	LUT2 #(
		.INIT('h1)
	) name9442 (
		\pio_PINT_reg[1]/NET0131 ,
		_w13489_,
		_w13490_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9443 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13490_,
		_w13491_
	);
	LUT4 #(
		.INIT('hba00)
	) name9444 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13366_,
		_w13492_
	);
	LUT2 #(
		.INIT('h1)
	) name9445 (
		_w13491_,
		_w13492_,
		_w13493_
	);
	LUT4 #(
		.INIT('h1400)
	) name9446 (
		\PIO_oe[3]_pad ,
		\pio_PIO_RES_OUT_reg[3]/P0001 ,
		\pio_PIO_RES_reg[3]/NET0131 ,
		\pio_pmask_reg_DO_reg[3]/NET0131 ,
		_w13494_
	);
	LUT2 #(
		.INIT('h1)
	) name9447 (
		\pio_PINT_reg[3]/NET0131 ,
		_w13494_,
		_w13495_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9448 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13495_,
		_w13496_
	);
	LUT4 #(
		.INIT('hba00)
	) name9449 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13366_,
		_w13497_
	);
	LUT2 #(
		.INIT('h1)
	) name9450 (
		_w13496_,
		_w13497_,
		_w13498_
	);
	LUT4 #(
		.INIT('h1400)
	) name9451 (
		\PIO_oe[6]_pad ,
		\pio_PIO_RES_OUT_reg[6]/P0001 ,
		\pio_PIO_RES_reg[6]/NET0131 ,
		\pio_pmask_reg_DO_reg[6]/NET0131 ,
		_w13499_
	);
	LUT2 #(
		.INIT('h1)
	) name9452 (
		\pio_PINT_reg[6]/NET0131 ,
		_w13499_,
		_w13500_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9453 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13500_,
		_w13501_
	);
	LUT4 #(
		.INIT('hba00)
	) name9454 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13366_,
		_w13502_
	);
	LUT2 #(
		.INIT('h1)
	) name9455 (
		_w13501_,
		_w13502_,
		_w13503_
	);
	LUT3 #(
		.INIT('h2a)
	) name9456 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001 ,
		_w4834_,
		_w12861_,
		_w13504_
	);
	LUT3 #(
		.INIT('h40)
	) name9457 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w9931_,
		_w13505_
	);
	LUT3 #(
		.INIT('h80)
	) name9458 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w13506_
	);
	LUT3 #(
		.INIT('h95)
	) name9459 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w13506_,
		_w13507_
	);
	LUT3 #(
		.INIT('h08)
	) name9460 (
		_w4834_,
		_w13505_,
		_w13507_,
		_w13508_
	);
	LUT2 #(
		.INIT('he)
	) name9461 (
		_w13504_,
		_w13508_,
		_w13509_
	);
	LUT3 #(
		.INIT('h2a)
	) name9462 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001 ,
		_w4834_,
		_w12861_,
		_w13510_
	);
	LUT3 #(
		.INIT('h65)
	) name9463 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w13506_,
		_w13511_
	);
	LUT3 #(
		.INIT('h08)
	) name9464 (
		_w4834_,
		_w13505_,
		_w13511_,
		_w13512_
	);
	LUT2 #(
		.INIT('he)
	) name9465 (
		_w13510_,
		_w13512_,
		_w13513_
	);
	LUT3 #(
		.INIT('h2a)
	) name9466 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001 ,
		_w4834_,
		_w12861_,
		_w13514_
	);
	LUT3 #(
		.INIT('h08)
	) name9467 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w13515_
	);
	LUT3 #(
		.INIT('h95)
	) name9468 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w13515_,
		_w13516_
	);
	LUT3 #(
		.INIT('h08)
	) name9469 (
		_w4834_,
		_w13505_,
		_w13516_,
		_w13517_
	);
	LUT2 #(
		.INIT('he)
	) name9470 (
		_w13514_,
		_w13517_,
		_w13518_
	);
	LUT3 #(
		.INIT('h2a)
	) name9471 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001 ,
		_w4834_,
		_w12861_,
		_w13519_
	);
	LUT3 #(
		.INIT('h65)
	) name9472 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w13515_,
		_w13520_
	);
	LUT3 #(
		.INIT('h08)
	) name9473 (
		_w4834_,
		_w13505_,
		_w13520_,
		_w13521_
	);
	LUT2 #(
		.INIT('he)
	) name9474 (
		_w13519_,
		_w13521_,
		_w13522_
	);
	LUT3 #(
		.INIT('h40)
	) name9475 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w4818_,
		_w12394_,
		_w13523_
	);
	LUT2 #(
		.INIT('h8)
	) name9476 (
		_w5028_,
		_w12916_,
		_w13524_
	);
	LUT4 #(
		.INIT('hbf00)
	) name9477 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w13524_,
		_w13525_
	);
	LUT4 #(
		.INIT('h31f5)
	) name9478 (
		_w4834_,
		_w5044_,
		_w11921_,
		_w13525_,
		_w13526_
	);
	LUT2 #(
		.INIT('hb)
	) name9479 (
		_w13523_,
		_w13526_,
		_w13527_
	);
	LUT4 #(
		.INIT('h1011)
	) name9480 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w7257_,
		_w7375_,
		_w7377_,
		_w13528_
	);
	LUT4 #(
		.INIT('h1555)
	) name9481 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w13117_,
		_w13137_,
		_w13139_,
		_w13529_
	);
	LUT3 #(
		.INIT('h40)
	) name9482 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13530_
	);
	LUT2 #(
		.INIT('h1)
	) name9483 (
		_w13158_,
		_w13530_,
		_w13531_
	);
	LUT4 #(
		.INIT('h7d00)
	) name9484 (
		_w13155_,
		_w13136_,
		_w13529_,
		_w13531_,
		_w13532_
	);
	LUT4 #(
		.INIT('hafac)
	) name9485 (
		\sport0_rxctl_RXSHT_reg[4]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w13533_
	);
	LUT4 #(
		.INIT('h0002)
	) name9486 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w13534_
	);
	LUT4 #(
		.INIT('hffb0)
	) name9487 (
		_w13528_,
		_w13532_,
		_w13533_,
		_w13534_,
		_w13535_
	);
	LUT3 #(
		.INIT('hc8)
	) name9488 (
		_w4063_,
		_w4857_,
		_w4845_,
		_w13536_
	);
	LUT2 #(
		.INIT('hb)
	) name9489 (
		_w12398_,
		_w13536_,
		_w13537_
	);
	LUT4 #(
		.INIT('h1400)
	) name9490 (
		\PIO_oe[7]_pad ,
		\pio_PIO_RES_OUT_reg[7]/P0001 ,
		\pio_PIO_RES_reg[7]/NET0131 ,
		\pio_pmask_reg_DO_reg[7]/NET0131 ,
		_w13538_
	);
	LUT2 #(
		.INIT('h1)
	) name9491 (
		\pio_PINT_reg[7]/NET0131 ,
		_w13538_,
		_w13539_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9492 (
		_w5672_,
		_w5658_,
		_w9431_,
		_w13539_,
		_w13540_
	);
	LUT4 #(
		.INIT('hba00)
	) name9493 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13366_,
		_w13541_
	);
	LUT2 #(
		.INIT('h1)
	) name9494 (
		_w13540_,
		_w13541_,
		_w13542_
	);
	LUT4 #(
		.INIT('h4000)
	) name9495 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w5028_,
		_w12392_,
		_w12393_,
		_w13543_
	);
	LUT3 #(
		.INIT('h01)
	) name9496 (
		_w4967_,
		_w4969_,
		_w13543_,
		_w13544_
	);
	LUT4 #(
		.INIT('h00bf)
	) name9497 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w13544_,
		_w13545_
	);
	LUT4 #(
		.INIT('h00c8)
	) name9498 (
		_w4063_,
		_w4857_,
		_w4845_,
		_w13545_,
		_w13546_
	);
	LUT4 #(
		.INIT('hff37)
	) name9499 (
		_w4063_,
		_w4857_,
		_w4845_,
		_w13545_,
		_w13547_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9500 (
		\core_c_psq_SSTAT_reg[4]/NET0131 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4094_,
		_w4097_,
		_w13548_
	);
	LUT4 #(
		.INIT('hab00)
	) name9501 (
		_w4971_,
		_w9906_,
		_w9907_,
		_w13548_,
		_w13549_
	);
	LUT3 #(
		.INIT('h7e)
	) name9502 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w13550_
	);
	LUT3 #(
		.INIT('h0e)
	) name9503 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w9906_,
		_w13550_,
		_w13551_
	);
	LUT3 #(
		.INIT('hec)
	) name9504 (
		_w11802_,
		_w13549_,
		_w13551_,
		_w13552_
	);
	LUT4 #(
		.INIT('hce02)
	) name9505 (
		\emc_PMDoe_reg/NET0131 ,
		_w12057_,
		_w12061_,
		_w12790_,
		_w13553_
	);
	LUT2 #(
		.INIT('h9)
	) name9506 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		_w13554_
	);
	LUT3 #(
		.INIT('hc1)
	) name9507 (
		_w9916_,
		_w11602_,
		_w13554_,
		_w13555_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9508 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13556_
	);
	LUT4 #(
		.INIT('h0800)
	) name9509 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13557_
	);
	LUT2 #(
		.INIT('he)
	) name9510 (
		_w13556_,
		_w13557_,
		_w13558_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9511 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13559_
	);
	LUT4 #(
		.INIT('h0800)
	) name9512 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13560_
	);
	LUT2 #(
		.INIT('he)
	) name9513 (
		_w13559_,
		_w13560_,
		_w13561_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9514 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13562_
	);
	LUT4 #(
		.INIT('h0800)
	) name9515 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13563_
	);
	LUT2 #(
		.INIT('he)
	) name9516 (
		_w13562_,
		_w13563_,
		_w13564_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9517 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13565_
	);
	LUT4 #(
		.INIT('h0800)
	) name9518 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13566_
	);
	LUT2 #(
		.INIT('he)
	) name9519 (
		_w13565_,
		_w13566_,
		_w13567_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9520 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13568_
	);
	LUT4 #(
		.INIT('h0800)
	) name9521 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13569_
	);
	LUT2 #(
		.INIT('he)
	) name9522 (
		_w13568_,
		_w13569_,
		_w13570_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9523 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13571_
	);
	LUT4 #(
		.INIT('h0800)
	) name9524 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13572_
	);
	LUT2 #(
		.INIT('he)
	) name9525 (
		_w13571_,
		_w13572_,
		_w13573_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9526 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13574_
	);
	LUT4 #(
		.INIT('h0800)
	) name9527 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13575_
	);
	LUT2 #(
		.INIT('he)
	) name9528 (
		_w13574_,
		_w13575_,
		_w13576_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9529 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13577_
	);
	LUT4 #(
		.INIT('h0800)
	) name9530 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13578_
	);
	LUT2 #(
		.INIT('he)
	) name9531 (
		_w13577_,
		_w13578_,
		_w13579_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9532 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13580_
	);
	LUT4 #(
		.INIT('h0800)
	) name9533 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13581_
	);
	LUT2 #(
		.INIT('he)
	) name9534 (
		_w13580_,
		_w13581_,
		_w13582_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9535 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13583_
	);
	LUT4 #(
		.INIT('h0800)
	) name9536 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13584_
	);
	LUT2 #(
		.INIT('he)
	) name9537 (
		_w13583_,
		_w13584_,
		_w13585_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9538 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13586_
	);
	LUT4 #(
		.INIT('h0800)
	) name9539 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13587_
	);
	LUT2 #(
		.INIT('he)
	) name9540 (
		_w13586_,
		_w13587_,
		_w13588_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9541 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13589_
	);
	LUT4 #(
		.INIT('h0800)
	) name9542 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13590_
	);
	LUT2 #(
		.INIT('he)
	) name9543 (
		_w13589_,
		_w13590_,
		_w13591_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9544 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13592_
	);
	LUT4 #(
		.INIT('h0800)
	) name9545 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13593_
	);
	LUT2 #(
		.INIT('he)
	) name9546 (
		_w13592_,
		_w13593_,
		_w13594_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9547 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13595_
	);
	LUT4 #(
		.INIT('h0800)
	) name9548 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13596_
	);
	LUT2 #(
		.INIT('he)
	) name9549 (
		_w13595_,
		_w13596_,
		_w13597_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9550 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13598_
	);
	LUT4 #(
		.INIT('h0800)
	) name9551 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13599_
	);
	LUT2 #(
		.INIT('he)
	) name9552 (
		_w13598_,
		_w13599_,
		_w13600_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9553 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13601_
	);
	LUT4 #(
		.INIT('h0800)
	) name9554 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13602_
	);
	LUT2 #(
		.INIT('he)
	) name9555 (
		_w13601_,
		_w13602_,
		_w13603_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9556 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13604_
	);
	LUT4 #(
		.INIT('h0800)
	) name9557 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13605_
	);
	LUT2 #(
		.INIT('he)
	) name9558 (
		_w13604_,
		_w13605_,
		_w13606_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9559 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13607_
	);
	LUT4 #(
		.INIT('h0800)
	) name9560 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w4438_,
		_w12894_,
		_w12897_,
		_w13608_
	);
	LUT2 #(
		.INIT('he)
	) name9561 (
		_w13607_,
		_w13608_,
		_w13609_
	);
	LUT4 #(
		.INIT('h4544)
	) name9562 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6054_,
		_w6173_,
		_w6175_,
		_w13610_
	);
	LUT2 #(
		.INIT('h2)
	) name9563 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8885_,
		_w13611_
	);
	LUT3 #(
		.INIT('ha8)
	) name9564 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w13610_,
		_w13611_,
		_w13612_
	);
	LUT2 #(
		.INIT('h8)
	) name9565 (
		_w11555_,
		_w11465_,
		_w13613_
	);
	LUT4 #(
		.INIT('hfca8)
	) name9566 (
		_w11530_,
		_w11489_,
		_w11492_,
		_w11454_,
		_w13614_
	);
	LUT4 #(
		.INIT('h135f)
	) name9567 (
		_w11558_,
		_w11532_,
		_w11874_,
		_w12468_,
		_w13615_
	);
	LUT4 #(
		.INIT('h0eee)
	) name9568 (
		_w11534_,
		_w11512_,
		_w11522_,
		_w11469_,
		_w13616_
	);
	LUT4 #(
		.INIT('h4000)
	) name9569 (
		_w13613_,
		_w13615_,
		_w13616_,
		_w13614_,
		_w13617_
	);
	LUT3 #(
		.INIT('h54)
	) name9570 (
		_w11540_,
		_w11409_,
		_w11896_,
		_w13618_
	);
	LUT3 #(
		.INIT('ha8)
	) name9571 (
		_w11537_,
		_w11973_,
		_w11974_,
		_w13619_
	);
	LUT3 #(
		.INIT('h02)
	) name9572 (
		_w11386_,
		_w11528_,
		_w11953_,
		_w13620_
	);
	LUT3 #(
		.INIT('h01)
	) name9573 (
		_w13619_,
		_w13620_,
		_w13618_,
		_w13621_
	);
	LUT3 #(
		.INIT('ha8)
	) name9574 (
		_w11495_,
		_w11435_,
		_w12455_,
		_w13622_
	);
	LUT4 #(
		.INIT('ha820)
	) name9575 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001 ,
		_w13623_
	);
	LUT3 #(
		.INIT('h07)
	) name9576 (
		_w11429_,
		_w12412_,
		_w13623_,
		_w13624_
	);
	LUT2 #(
		.INIT('h2)
	) name9577 (
		_w11415_,
		_w11471_,
		_w13625_
	);
	LUT3 #(
		.INIT('h80)
	) name9578 (
		_w11389_,
		_w11476_,
		_w11515_,
		_w13626_
	);
	LUT4 #(
		.INIT('h0100)
	) name9579 (
		_w11403_,
		_w13625_,
		_w13626_,
		_w13624_,
		_w13627_
	);
	LUT3 #(
		.INIT('hc8)
	) name9580 (
		_w11588_,
		_w11458_,
		_w12496_,
		_w13628_
	);
	LUT3 #(
		.INIT('hc8)
	) name9581 (
		_w11587_,
		_w11499_,
		_w11880_,
		_w13629_
	);
	LUT4 #(
		.INIT('h0100)
	) name9582 (
		_w13622_,
		_w13628_,
		_w13629_,
		_w13627_,
		_w13630_
	);
	LUT4 #(
		.INIT('h8000)
	) name9583 (
		_w12644_,
		_w13621_,
		_w13630_,
		_w13617_,
		_w13631_
	);
	LUT4 #(
		.INIT('h4000)
	) name9584 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w12451_,
		_w13224_,
		_w13631_,
		_w13632_
	);
	LUT4 #(
		.INIT('h222e)
	) name9585 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001 ,
		_w11830_,
		_w13612_,
		_w13632_,
		_w13633_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9586 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13634_
	);
	LUT4 #(
		.INIT('h0800)
	) name9587 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13635_
	);
	LUT2 #(
		.INIT('he)
	) name9588 (
		_w13634_,
		_w13635_,
		_w13636_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9589 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13637_
	);
	LUT4 #(
		.INIT('h0800)
	) name9590 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13638_
	);
	LUT2 #(
		.INIT('he)
	) name9591 (
		_w13637_,
		_w13638_,
		_w13639_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9592 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13640_
	);
	LUT4 #(
		.INIT('h0800)
	) name9593 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13641_
	);
	LUT2 #(
		.INIT('he)
	) name9594 (
		_w13640_,
		_w13641_,
		_w13642_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9595 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13643_
	);
	LUT4 #(
		.INIT('h0800)
	) name9596 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13644_
	);
	LUT2 #(
		.INIT('he)
	) name9597 (
		_w13643_,
		_w13644_,
		_w13645_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9598 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13646_
	);
	LUT4 #(
		.INIT('h0800)
	) name9599 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13647_
	);
	LUT2 #(
		.INIT('he)
	) name9600 (
		_w13646_,
		_w13647_,
		_w13648_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9601 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13649_
	);
	LUT4 #(
		.INIT('h0800)
	) name9602 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13650_
	);
	LUT2 #(
		.INIT('he)
	) name9603 (
		_w13649_,
		_w13650_,
		_w13651_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9604 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13652_
	);
	LUT4 #(
		.INIT('h0800)
	) name9605 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13653_
	);
	LUT2 #(
		.INIT('he)
	) name9606 (
		_w13652_,
		_w13653_,
		_w13654_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9607 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13655_
	);
	LUT4 #(
		.INIT('h0800)
	) name9608 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13656_
	);
	LUT2 #(
		.INIT('he)
	) name9609 (
		_w13655_,
		_w13656_,
		_w13657_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9610 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13658_
	);
	LUT4 #(
		.INIT('h0800)
	) name9611 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13659_
	);
	LUT2 #(
		.INIT('he)
	) name9612 (
		_w13658_,
		_w13659_,
		_w13660_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9613 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13661_
	);
	LUT4 #(
		.INIT('h0800)
	) name9614 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13662_
	);
	LUT2 #(
		.INIT('he)
	) name9615 (
		_w13661_,
		_w13662_,
		_w13663_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9616 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13664_
	);
	LUT4 #(
		.INIT('h0800)
	) name9617 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13665_
	);
	LUT2 #(
		.INIT('he)
	) name9618 (
		_w13664_,
		_w13665_,
		_w13666_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9619 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13667_
	);
	LUT4 #(
		.INIT('h0800)
	) name9620 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13668_
	);
	LUT2 #(
		.INIT('he)
	) name9621 (
		_w13667_,
		_w13668_,
		_w13669_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9622 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13670_
	);
	LUT4 #(
		.INIT('h0800)
	) name9623 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13671_
	);
	LUT2 #(
		.INIT('he)
	) name9624 (
		_w13670_,
		_w13671_,
		_w13672_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9625 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13673_
	);
	LUT4 #(
		.INIT('h0800)
	) name9626 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13674_
	);
	LUT2 #(
		.INIT('he)
	) name9627 (
		_w13673_,
		_w13674_,
		_w13675_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9628 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13676_
	);
	LUT4 #(
		.INIT('h0800)
	) name9629 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13677_
	);
	LUT2 #(
		.INIT('he)
	) name9630 (
		_w13676_,
		_w13677_,
		_w13678_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9631 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13679_
	);
	LUT4 #(
		.INIT('h0800)
	) name9632 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13680_
	);
	LUT2 #(
		.INIT('he)
	) name9633 (
		_w13679_,
		_w13680_,
		_w13681_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9634 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13682_
	);
	LUT4 #(
		.INIT('h0800)
	) name9635 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13683_
	);
	LUT2 #(
		.INIT('he)
	) name9636 (
		_w13682_,
		_w13683_,
		_w13684_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9637 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13685_
	);
	LUT4 #(
		.INIT('h0800)
	) name9638 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w4435_,
		_w12894_,
		_w12897_,
		_w13686_
	);
	LUT2 #(
		.INIT('he)
	) name9639 (
		_w13685_,
		_w13686_,
		_w13687_
	);
	LUT4 #(
		.INIT('haccc)
	) name9640 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001 ,
		_w12897_,
		_w12909_,
		_w13688_
	);
	LUT4 #(
		.INIT('haccc)
	) name9641 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001 ,
		_w12897_,
		_w12909_,
		_w13689_
	);
	LUT4 #(
		.INIT('haccc)
	) name9642 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001 ,
		_w12897_,
		_w12909_,
		_w13690_
	);
	LUT4 #(
		.INIT('haccc)
	) name9643 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001 ,
		_w12897_,
		_w12909_,
		_w13691_
	);
	LUT4 #(
		.INIT('haccc)
	) name9644 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001 ,
		_w12897_,
		_w12909_,
		_w13692_
	);
	LUT4 #(
		.INIT('haccc)
	) name9645 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001 ,
		_w12897_,
		_w12909_,
		_w13693_
	);
	LUT4 #(
		.INIT('haccc)
	) name9646 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001 ,
		_w12897_,
		_w12909_,
		_w13694_
	);
	LUT4 #(
		.INIT('haccc)
	) name9647 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001 ,
		_w12897_,
		_w12909_,
		_w13695_
	);
	LUT4 #(
		.INIT('haccc)
	) name9648 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001 ,
		_w12897_,
		_w12909_,
		_w13696_
	);
	LUT4 #(
		.INIT('haccc)
	) name9649 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001 ,
		_w12897_,
		_w12909_,
		_w13697_
	);
	LUT4 #(
		.INIT('haccc)
	) name9650 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001 ,
		_w12897_,
		_w12909_,
		_w13698_
	);
	LUT4 #(
		.INIT('haccc)
	) name9651 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001 ,
		_w12897_,
		_w12909_,
		_w13699_
	);
	LUT3 #(
		.INIT('h28)
	) name9652 (
		_w9455_,
		_w9883_,
		_w9885_,
		_w13700_
	);
	LUT4 #(
		.INIT('h5401)
	) name9653 (
		_w9455_,
		_w9456_,
		_w9715_,
		_w12610_,
		_w13701_
	);
	LUT4 #(
		.INIT('heee2)
	) name9654 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001 ,
		_w9895_,
		_w13700_,
		_w13701_,
		_w13702_
	);
	LUT4 #(
		.INIT('haccc)
	) name9655 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001 ,
		_w12897_,
		_w12909_,
		_w13703_
	);
	LUT4 #(
		.INIT('haccc)
	) name9656 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001 ,
		_w12897_,
		_w12909_,
		_w13704_
	);
	LUT4 #(
		.INIT('haccc)
	) name9657 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001 ,
		_w12897_,
		_w12909_,
		_w13705_
	);
	LUT4 #(
		.INIT('haccc)
	) name9658 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001 ,
		_w12897_,
		_w12909_,
		_w13706_
	);
	LUT4 #(
		.INIT('haccc)
	) name9659 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001 ,
		_w12897_,
		_w12909_,
		_w13707_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9660 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13708_
	);
	LUT4 #(
		.INIT('h0800)
	) name9661 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13709_
	);
	LUT2 #(
		.INIT('he)
	) name9662 (
		_w13708_,
		_w13709_,
		_w13710_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9663 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13711_
	);
	LUT4 #(
		.INIT('h0800)
	) name9664 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13712_
	);
	LUT2 #(
		.INIT('he)
	) name9665 (
		_w13711_,
		_w13712_,
		_w13713_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9666 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13714_
	);
	LUT4 #(
		.INIT('h0800)
	) name9667 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13715_
	);
	LUT2 #(
		.INIT('he)
	) name9668 (
		_w13714_,
		_w13715_,
		_w13716_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9669 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13717_
	);
	LUT4 #(
		.INIT('h0800)
	) name9670 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13718_
	);
	LUT2 #(
		.INIT('he)
	) name9671 (
		_w13717_,
		_w13718_,
		_w13719_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9672 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13720_
	);
	LUT4 #(
		.INIT('h0800)
	) name9673 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13721_
	);
	LUT2 #(
		.INIT('he)
	) name9674 (
		_w13720_,
		_w13721_,
		_w13722_
	);
	LUT4 #(
		.INIT('heee2)
	) name9675 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001 ,
		_w9454_,
		_w13700_,
		_w13701_,
		_w13723_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9676 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13724_
	);
	LUT4 #(
		.INIT('h0800)
	) name9677 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13725_
	);
	LUT2 #(
		.INIT('he)
	) name9678 (
		_w13724_,
		_w13725_,
		_w13726_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9679 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13727_
	);
	LUT4 #(
		.INIT('h0800)
	) name9680 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13728_
	);
	LUT2 #(
		.INIT('he)
	) name9681 (
		_w13727_,
		_w13728_,
		_w13729_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9682 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13730_
	);
	LUT4 #(
		.INIT('h0800)
	) name9683 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13731_
	);
	LUT2 #(
		.INIT('he)
	) name9684 (
		_w13730_,
		_w13731_,
		_w13732_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9685 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13733_
	);
	LUT4 #(
		.INIT('h0800)
	) name9686 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13734_
	);
	LUT2 #(
		.INIT('he)
	) name9687 (
		_w13733_,
		_w13734_,
		_w13735_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9688 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13736_
	);
	LUT4 #(
		.INIT('h0800)
	) name9689 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13737_
	);
	LUT2 #(
		.INIT('he)
	) name9690 (
		_w13736_,
		_w13737_,
		_w13738_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9691 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13739_
	);
	LUT4 #(
		.INIT('h0800)
	) name9692 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13740_
	);
	LUT2 #(
		.INIT('he)
	) name9693 (
		_w13739_,
		_w13740_,
		_w13741_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9694 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13742_
	);
	LUT4 #(
		.INIT('h0800)
	) name9695 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13743_
	);
	LUT2 #(
		.INIT('he)
	) name9696 (
		_w13742_,
		_w13743_,
		_w13744_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9697 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13745_
	);
	LUT4 #(
		.INIT('h0800)
	) name9698 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13746_
	);
	LUT2 #(
		.INIT('he)
	) name9699 (
		_w13745_,
		_w13746_,
		_w13747_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9700 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13748_
	);
	LUT4 #(
		.INIT('h0800)
	) name9701 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13749_
	);
	LUT2 #(
		.INIT('he)
	) name9702 (
		_w13748_,
		_w13749_,
		_w13750_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9703 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13751_
	);
	LUT4 #(
		.INIT('h0800)
	) name9704 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13752_
	);
	LUT2 #(
		.INIT('he)
	) name9705 (
		_w13751_,
		_w13752_,
		_w13753_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9706 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13754_
	);
	LUT4 #(
		.INIT('h0800)
	) name9707 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13755_
	);
	LUT2 #(
		.INIT('he)
	) name9708 (
		_w13754_,
		_w13755_,
		_w13756_
	);
	LUT2 #(
		.INIT('h9)
	) name9709 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w13757_
	);
	LUT3 #(
		.INIT('hbc)
	) name9710 (
		_w9437_,
		_w9439_,
		_w13757_,
		_w13758_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9711 (
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w13759_
	);
	LUT4 #(
		.INIT('h1101)
	) name9712 (
		\core_c_psq_IFC_reg[12]/NET0131 ,
		\core_c_psq_Iflag_reg[4]/NET0131 ,
		\core_c_psq_T_IRQE1_reg/P0001 ,
		\core_c_psq_T_IRQE1_s1_reg/P0001 ,
		_w13760_
	);
	LUT2 #(
		.INIT('h1)
	) name9713 (
		\core_c_psq_IFC_reg[4]/NET0131 ,
		_w13760_,
		_w13761_
	);
	LUT2 #(
		.INIT('h4)
	) name9714 (
		_w13759_,
		_w13761_,
		_w13762_
	);
	LUT3 #(
		.INIT('hae)
	) name9715 (
		\core_c_psq_SSTAT_reg[5]/NET0131 ,
		_w9916_,
		_w11602_,
		_w13763_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9716 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13764_
	);
	LUT4 #(
		.INIT('h0800)
	) name9717 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13765_
	);
	LUT2 #(
		.INIT('he)
	) name9718 (
		_w13764_,
		_w13765_,
		_w13766_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name9719 (
		\bdma_DM_2nd_reg/NET0131 ,
		_w5531_,
		_w9412_,
		_w9413_,
		_w13767_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name9720 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13768_
	);
	LUT4 #(
		.INIT('h0800)
	) name9721 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w4437_,
		_w12894_,
		_w12897_,
		_w13769_
	);
	LUT2 #(
		.INIT('he)
	) name9722 (
		_w13768_,
		_w13769_,
		_w13770_
	);
	LUT4 #(
		.INIT('h4000)
	) name9723 (
		\memc_MMR_web_reg/NET0131 ,
		_w5658_,
		_w9431_,
		_w11608_,
		_w13771_
	);
	LUT3 #(
		.INIT('hca)
	) name9724 (
		\pio_pmask_reg_DO_reg[9]/NET0131 ,
		_w5760_,
		_w13771_,
		_w13772_
	);
	LUT4 #(
		.INIT('h4000)
	) name9725 (
		\memc_MMR_web_reg/NET0131 ,
		_w5658_,
		_w9431_,
		_w11606_,
		_w13773_
	);
	LUT3 #(
		.INIT('hca)
	) name9726 (
		\PIO_oe[8]_pad ,
		_w6758_,
		_w13773_,
		_w13774_
	);
	LUT4 #(
		.INIT('h222e)
	) name9727 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001 ,
		_w11329_,
		_w13612_,
		_w13632_,
		_w13775_
	);
	LUT4 #(
		.INIT('haccc)
	) name9728 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001 ,
		_w12897_,
		_w12909_,
		_w13776_
	);
	LUT4 #(
		.INIT('h4000)
	) name9729 (
		\memc_MMR_web_reg/NET0131 ,
		_w5810_,
		_w9431_,
		_w11604_,
		_w13777_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9730 (
		\memc_usysr_DO_reg[9]/NET0131 ,
		_w7140_,
		_w7240_,
		_w13777_,
		_w13778_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9731 (
		\memc_usysr_DO_reg[8]/NET0131 ,
		_w7465_,
		_w7565_,
		_w13777_,
		_w13779_
	);
	LUT3 #(
		.INIT('hca)
	) name9732 (
		\memc_usysr_DO_reg[13]/NET0131 ,
		_w5760_,
		_w13777_,
		_w13780_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9733 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w13777_,
		_w13781_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9734 (
		\memc_usysr_DO_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w13777_,
		_w13782_
	);
	LUT4 #(
		.INIT('h4000)
	) name9735 (
		\memc_MMR_web_reg/NET0131 ,
		_w5647_,
		_w9431_,
		_w11604_,
		_w13783_
	);
	LUT2 #(
		.INIT('h8)
	) name9736 (
		_w12621_,
		_w13783_,
		_w13784_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9737 (
		\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w7140_,
		_w7240_,
		_w13784_,
		_w13785_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9738 (
		\sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w7465_,
		_w7565_,
		_w13784_,
		_w13786_
	);
	LUT3 #(
		.INIT('ha8)
	) name9739 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w13610_,
		_w13611_,
		_w13787_
	);
	LUT3 #(
		.INIT('ha8)
	) name9740 (
		_w11386_,
		_w13271_,
		_w13272_,
		_w13788_
	);
	LUT2 #(
		.INIT('h8)
	) name9741 (
		_w11537_,
		_w11424_,
		_w13789_
	);
	LUT3 #(
		.INIT('hc8)
	) name9742 (
		_w11552_,
		_w11508_,
		_w11474_,
		_w13790_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name9743 (
		_w11593_,
		_w11450_,
		_w11957_,
		_w12412_,
		_w13791_
	);
	LUT3 #(
		.INIT('h10)
	) name9744 (
		_w13789_,
		_w13790_,
		_w13791_,
		_w13792_
	);
	LUT3 #(
		.INIT('h20)
	) name9745 (
		_w11574_,
		_w13788_,
		_w13792_,
		_w13793_
	);
	LUT3 #(
		.INIT('hc8)
	) name9746 (
		_w11547_,
		_w11465_,
		_w11976_,
		_w13794_
	);
	LUT3 #(
		.INIT('he0)
	) name9747 (
		_w11397_,
		_w11519_,
		_w11860_,
		_w13795_
	);
	LUT3 #(
		.INIT('he0)
	) name9748 (
		_w11420_,
		_w11421_,
		_w11469_,
		_w13796_
	);
	LUT3 #(
		.INIT('h01)
	) name9749 (
		_w13795_,
		_w13796_,
		_w13794_,
		_w13797_
	);
	LUT4 #(
		.INIT('ha820)
	) name9750 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001 ,
		_w13798_
	);
	LUT4 #(
		.INIT('h0054)
	) name9751 (
		_w11581_,
		_w11501_,
		_w11954_,
		_w13798_,
		_w13799_
	);
	LUT2 #(
		.INIT('h1)
	) name9752 (
		_w11592_,
		_w12024_,
		_w13800_
	);
	LUT3 #(
		.INIT('h0e)
	) name9753 (
		_w11393_,
		_w11589_,
		_w11489_,
		_w13801_
	);
	LUT3 #(
		.INIT('h10)
	) name9754 (
		_w13800_,
		_w13801_,
		_w13799_,
		_w13802_
	);
	LUT3 #(
		.INIT('h02)
	) name9755 (
		_w11386_,
		_w11593_,
		_w11528_,
		_w13803_
	);
	LUT2 #(
		.INIT('h2)
	) name9756 (
		_w11969_,
		_w13803_,
		_w13804_
	);
	LUT3 #(
		.INIT('h80)
	) name9757 (
		_w13802_,
		_w13804_,
		_w13797_,
		_w13805_
	);
	LUT4 #(
		.INIT('h2333)
	) name9758 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w13787_,
		_w13793_,
		_w13805_,
		_w13806_
	);
	LUT3 #(
		.INIT('he2)
	) name9759 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001 ,
		_w11946_,
		_w13806_,
		_w13807_
	);
	LUT3 #(
		.INIT('hca)
	) name9760 (
		\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w5760_,
		_w13784_,
		_w13808_
	);
	LUT3 #(
		.INIT('hca)
	) name9761 (
		\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w6758_,
		_w13784_,
		_w13809_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9762 (
		\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w13784_,
		_w13810_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9763 (
		\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w13784_,
		_w13811_
	);
	LUT4 #(
		.INIT('h4000)
	) name9764 (
		\memc_MMR_web_reg/NET0131 ,
		_w5658_,
		_w5810_,
		_w9431_,
		_w13812_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9765 (
		\sport1_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w7465_,
		_w7565_,
		_w13812_,
		_w13813_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9766 (
		\sport1_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w7140_,
		_w7240_,
		_w13812_,
		_w13814_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9767 (
		\sport1_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w13812_,
		_w13815_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9768 (
		\sport1_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w13812_,
		_w13816_
	);
	LUT3 #(
		.INIT('h01)
	) name9769 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_c_dec_DIVS_E_reg/P0001 ,
		\core_c_dec_MTAY0_E_reg/P0001 ,
		_w13817_
	);
	LUT2 #(
		.INIT('h2)
	) name9770 (
		_w9894_,
		_w13817_,
		_w13818_
	);
	LUT2 #(
		.INIT('h1)
	) name9771 (
		\core_c_dec_Double_E_reg/P0001 ,
		\core_c_dec_accPM_E_reg/P0001 ,
		_w13819_
	);
	LUT2 #(
		.INIT('h1)
	) name9772 (
		_w9021_,
		_w13819_,
		_w13820_
	);
	LUT4 #(
		.INIT('h001f)
	) name9773 (
		_w7140_,
		_w7240_,
		_w13819_,
		_w13820_,
		_w13821_
	);
	LUT4 #(
		.INIT('h80b0)
	) name9774 (
		_w7540_,
		_w9455_,
		_w13818_,
		_w13821_,
		_w13822_
	);
	LUT3 #(
		.INIT('h51)
	) name9775 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001 ,
		_w9894_,
		_w13817_,
		_w13823_
	);
	LUT2 #(
		.INIT('h1)
	) name9776 (
		_w13822_,
		_w13823_,
		_w13824_
	);
	LUT2 #(
		.INIT('h2)
	) name9777 (
		_w8998_,
		_w13819_,
		_w13825_
	);
	LUT4 #(
		.INIT('h00ef)
	) name9778 (
		_w7465_,
		_w7565_,
		_w13819_,
		_w13825_,
		_w13826_
	);
	LUT4 #(
		.INIT('hb080)
	) name9779 (
		_w7872_,
		_w9455_,
		_w13818_,
		_w13826_,
		_w13827_
	);
	LUT3 #(
		.INIT('h51)
	) name9780 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001 ,
		_w9894_,
		_w13817_,
		_w13828_
	);
	LUT2 #(
		.INIT('h1)
	) name9781 (
		_w13827_,
		_w13828_,
		_w13829_
	);
	LUT4 #(
		.INIT('hba00)
	) name9782 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13819_,
		_w13830_
	);
	LUT2 #(
		.INIT('h1)
	) name9783 (
		_w8974_,
		_w13819_,
		_w13831_
	);
	LUT2 #(
		.INIT('h8)
	) name9784 (
		_w7931_,
		_w9455_,
		_w13832_
	);
	LUT4 #(
		.INIT('h00ab)
	) name9785 (
		_w9455_,
		_w13830_,
		_w13831_,
		_w13832_,
		_w13833_
	);
	LUT3 #(
		.INIT('he2)
	) name9786 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001 ,
		_w13818_,
		_w13833_,
		_w13834_
	);
	LUT4 #(
		.INIT('hba00)
	) name9787 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13819_,
		_w13835_
	);
	LUT2 #(
		.INIT('h1)
	) name9788 (
		_w8952_,
		_w13819_,
		_w13836_
	);
	LUT2 #(
		.INIT('h8)
	) name9789 (
		_w7681_,
		_w9455_,
		_w13837_
	);
	LUT4 #(
		.INIT('h00ab)
	) name9790 (
		_w9455_,
		_w13835_,
		_w13836_,
		_w13837_,
		_w13838_
	);
	LUT3 #(
		.INIT('he2)
	) name9791 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001 ,
		_w13818_,
		_w13838_,
		_w13839_
	);
	LUT4 #(
		.INIT('hba00)
	) name9792 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13819_,
		_w13840_
	);
	LUT2 #(
		.INIT('h1)
	) name9793 (
		_w8929_,
		_w13819_,
		_w13841_
	);
	LUT2 #(
		.INIT('h8)
	) name9794 (
		_w7359_,
		_w9455_,
		_w13842_
	);
	LUT4 #(
		.INIT('h00ab)
	) name9795 (
		_w9455_,
		_w13840_,
		_w13841_,
		_w13842_,
		_w13843_
	);
	LUT3 #(
		.INIT('he2)
	) name9796 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001 ,
		_w13818_,
		_w13843_,
		_w13844_
	);
	LUT4 #(
		.INIT('hba00)
	) name9797 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13819_,
		_w13845_
	);
	LUT2 #(
		.INIT('h1)
	) name9798 (
		_w8907_,
		_w13819_,
		_w13846_
	);
	LUT2 #(
		.INIT('h8)
	) name9799 (
		_w6158_,
		_w9455_,
		_w13847_
	);
	LUT4 #(
		.INIT('h00ab)
	) name9800 (
		_w9455_,
		_w13845_,
		_w13846_,
		_w13847_,
		_w13848_
	);
	LUT3 #(
		.INIT('he2)
	) name9801 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001 ,
		_w13818_,
		_w13848_,
		_w13849_
	);
	LUT4 #(
		.INIT('hba00)
	) name9802 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13819_,
		_w13850_
	);
	LUT2 #(
		.INIT('h1)
	) name9803 (
		_w8885_,
		_w13819_,
		_w13851_
	);
	LUT2 #(
		.INIT('h8)
	) name9804 (
		_w6452_,
		_w9455_,
		_w13852_
	);
	LUT4 #(
		.INIT('h00ab)
	) name9805 (
		_w9455_,
		_w13850_,
		_w13851_,
		_w13852_,
		_w13853_
	);
	LUT3 #(
		.INIT('he2)
	) name9806 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001 ,
		_w13818_,
		_w13853_,
		_w13854_
	);
	LUT4 #(
		.INIT('hba00)
	) name9807 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13819_,
		_w13855_
	);
	LUT2 #(
		.INIT('h1)
	) name9808 (
		_w8863_,
		_w13819_,
		_w13856_
	);
	LUT2 #(
		.INIT('h8)
	) name9809 (
		_w6854_,
		_w9455_,
		_w13857_
	);
	LUT4 #(
		.INIT('h00ab)
	) name9810 (
		_w9455_,
		_w13855_,
		_w13856_,
		_w13857_,
		_w13858_
	);
	LUT3 #(
		.INIT('he2)
	) name9811 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001 ,
		_w13818_,
		_w13858_,
		_w13859_
	);
	LUT2 #(
		.INIT('h1)
	) name9812 (
		_w8821_,
		_w13819_,
		_w13860_
	);
	LUT4 #(
		.INIT('h001f)
	) name9813 (
		_w8798_,
		_w8801_,
		_w13819_,
		_w13860_,
		_w13861_
	);
	LUT4 #(
		.INIT('h80b0)
	) name9814 (
		_w8269_,
		_w9455_,
		_w13818_,
		_w13861_,
		_w13862_
	);
	LUT3 #(
		.INIT('h51)
	) name9815 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001 ,
		_w9894_,
		_w13817_,
		_w13863_
	);
	LUT2 #(
		.INIT('h1)
	) name9816 (
		_w13862_,
		_w13863_,
		_w13864_
	);
	LUT2 #(
		.INIT('h1)
	) name9817 (
		_w8781_,
		_w13819_,
		_w13865_
	);
	LUT4 #(
		.INIT('h001f)
	) name9818 (
		_w8757_,
		_w8760_,
		_w13819_,
		_w13865_,
		_w13866_
	);
	LUT4 #(
		.INIT('h80b0)
	) name9819 (
		_w5736_,
		_w9455_,
		_w13818_,
		_w13866_,
		_w13867_
	);
	LUT3 #(
		.INIT('h51)
	) name9820 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001 ,
		_w9894_,
		_w13817_,
		_w13868_
	);
	LUT2 #(
		.INIT('h1)
	) name9821 (
		_w13867_,
		_w13868_,
		_w13869_
	);
	LUT4 #(
		.INIT('h0503)
	) name9822 (
		_w5760_,
		_w8740_,
		_w9455_,
		_w13819_,
		_w13870_
	);
	LUT2 #(
		.INIT('h8)
	) name9823 (
		_w6748_,
		_w9455_,
		_w13871_
	);
	LUT4 #(
		.INIT('h222e)
	) name9824 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001 ,
		_w13818_,
		_w13870_,
		_w13871_,
		_w13872_
	);
	LUT4 #(
		.INIT('h0503)
	) name9825 (
		_w6758_,
		_w8717_,
		_w9455_,
		_w13819_,
		_w13873_
	);
	LUT2 #(
		.INIT('h8)
	) name9826 (
		_w6351_,
		_w9455_,
		_w13874_
	);
	LUT4 #(
		.INIT('h222e)
	) name9827 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001 ,
		_w13818_,
		_w13873_,
		_w13874_,
		_w13875_
	);
	LUT3 #(
		.INIT('he2)
	) name9828 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001 ,
		_w12048_,
		_w13806_,
		_w13876_
	);
	LUT2 #(
		.INIT('h2)
	) name9829 (
		_w8694_,
		_w13819_,
		_w13877_
	);
	LUT4 #(
		.INIT('h00ef)
	) name9830 (
		_w6263_,
		_w6362_,
		_w13819_,
		_w13877_,
		_w13878_
	);
	LUT4 #(
		.INIT('hb080)
	) name9831 (
		_w6028_,
		_w9455_,
		_w13818_,
		_w13878_,
		_w13879_
	);
	LUT3 #(
		.INIT('h51)
	) name9832 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001 ,
		_w9894_,
		_w13817_,
		_w13880_
	);
	LUT2 #(
		.INIT('h1)
	) name9833 (
		_w13879_,
		_w13880_,
		_w13881_
	);
	LUT2 #(
		.INIT('h1)
	) name9834 (
		_w8671_,
		_w13819_,
		_w13882_
	);
	LUT4 #(
		.INIT('h001f)
	) name9835 (
		_w5937_,
		_w6038_,
		_w13819_,
		_w13882_,
		_w13883_
	);
	LUT4 #(
		.INIT('h80b0)
	) name9836 (
		_w7230_,
		_w9455_,
		_w13818_,
		_w13883_,
		_w13884_
	);
	LUT3 #(
		.INIT('h51)
	) name9837 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001 ,
		_w9894_,
		_w13817_,
		_w13885_
	);
	LUT2 #(
		.INIT('h1)
	) name9838 (
		_w13884_,
		_w13885_,
		_w13886_
	);
	LUT3 #(
		.INIT('hca)
	) name9839 (
		\PIO_oe[9]_pad ,
		_w5760_,
		_w13773_,
		_w13887_
	);
	LUT2 #(
		.INIT('h8)
	) name9840 (
		_w5656_,
		_w13783_,
		_w13888_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9841 (
		\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w7140_,
		_w7240_,
		_w13888_,
		_w13889_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9842 (
		\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w7465_,
		_w7565_,
		_w13888_,
		_w13890_
	);
	LUT3 #(
		.INIT('hca)
	) name9843 (
		\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w5760_,
		_w13888_,
		_w13891_
	);
	LUT3 #(
		.INIT('hca)
	) name9844 (
		\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w6758_,
		_w13888_,
		_w13892_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9845 (
		\sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w13888_,
		_w13893_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9846 (
		\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w13888_,
		_w13894_
	);
	LUT3 #(
		.INIT('hca)
	) name9847 (
		\pio_pmask_reg_DO_reg[8]/NET0131 ,
		_w6758_,
		_w13771_,
		_w13895_
	);
	LUT3 #(
		.INIT('hca)
	) name9848 (
		\sport0_regs_AUTO_a_reg[12]/NET0131 ,
		_w6758_,
		_w12825_,
		_w13896_
	);
	LUT4 #(
		.INIT('hba00)
	) name9849 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13819_,
		_w13897_
	);
	LUT2 #(
		.INIT('h1)
	) name9850 (
		_w8841_,
		_w13819_,
		_w13898_
	);
	LUT2 #(
		.INIT('h4)
	) name9851 (
		_w5895_,
		_w9455_,
		_w13899_
	);
	LUT4 #(
		.INIT('h00fe)
	) name9852 (
		_w9455_,
		_w13897_,
		_w13898_,
		_w13899_,
		_w13900_
	);
	LUT3 #(
		.INIT('h2e)
	) name9853 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001 ,
		_w13818_,
		_w13900_,
		_w13901_
	);
	LUT2 #(
		.INIT('h2)
	) name9854 (
		_w11300_,
		_w13817_,
		_w13902_
	);
	LUT4 #(
		.INIT('h8b00)
	) name9855 (
		_w7540_,
		_w9455_,
		_w13821_,
		_w13902_,
		_w13903_
	);
	LUT3 #(
		.INIT('h51)
	) name9856 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001 ,
		_w11300_,
		_w13817_,
		_w13904_
	);
	LUT2 #(
		.INIT('h1)
	) name9857 (
		_w13903_,
		_w13904_,
		_w13905_
	);
	LUT4 #(
		.INIT('hb800)
	) name9858 (
		_w7872_,
		_w9455_,
		_w13826_,
		_w13902_,
		_w13906_
	);
	LUT3 #(
		.INIT('h51)
	) name9859 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001 ,
		_w11300_,
		_w13817_,
		_w13907_
	);
	LUT2 #(
		.INIT('h1)
	) name9860 (
		_w13906_,
		_w13907_,
		_w13908_
	);
	LUT3 #(
		.INIT('hca)
	) name9861 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001 ,
		_w13833_,
		_w13902_,
		_w13909_
	);
	LUT3 #(
		.INIT('hca)
	) name9862 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001 ,
		_w13838_,
		_w13902_,
		_w13910_
	);
	LUT3 #(
		.INIT('hca)
	) name9863 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001 ,
		_w13843_,
		_w13902_,
		_w13911_
	);
	LUT3 #(
		.INIT('hca)
	) name9864 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001 ,
		_w13848_,
		_w13902_,
		_w13912_
	);
	LUT3 #(
		.INIT('hca)
	) name9865 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001 ,
		_w13853_,
		_w13902_,
		_w13913_
	);
	LUT3 #(
		.INIT('hca)
	) name9866 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001 ,
		_w13858_,
		_w13902_,
		_w13914_
	);
	LUT3 #(
		.INIT('h3a)
	) name9867 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001 ,
		_w13900_,
		_w13902_,
		_w13915_
	);
	LUT4 #(
		.INIT('h8b00)
	) name9868 (
		_w8269_,
		_w9455_,
		_w13861_,
		_w13902_,
		_w13916_
	);
	LUT3 #(
		.INIT('h51)
	) name9869 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001 ,
		_w11300_,
		_w13817_,
		_w13917_
	);
	LUT2 #(
		.INIT('h1)
	) name9870 (
		_w13916_,
		_w13917_,
		_w13918_
	);
	LUT4 #(
		.INIT('h8b00)
	) name9871 (
		_w5736_,
		_w9455_,
		_w13866_,
		_w13902_,
		_w13919_
	);
	LUT3 #(
		.INIT('h51)
	) name9872 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001 ,
		_w11300_,
		_w13817_,
		_w13920_
	);
	LUT2 #(
		.INIT('h1)
	) name9873 (
		_w13919_,
		_w13920_,
		_w13921_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9874 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001 ,
		_w13870_,
		_w13871_,
		_w13902_,
		_w13922_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9875 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001 ,
		_w13873_,
		_w13874_,
		_w13902_,
		_w13923_
	);
	LUT4 #(
		.INIT('hb800)
	) name9876 (
		_w6028_,
		_w9455_,
		_w13878_,
		_w13902_,
		_w13924_
	);
	LUT3 #(
		.INIT('h51)
	) name9877 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001 ,
		_w11300_,
		_w13817_,
		_w13925_
	);
	LUT2 #(
		.INIT('h1)
	) name9878 (
		_w13924_,
		_w13925_,
		_w13926_
	);
	LUT4 #(
		.INIT('h8b00)
	) name9879 (
		_w7230_,
		_w9455_,
		_w13883_,
		_w13902_,
		_w13927_
	);
	LUT3 #(
		.INIT('h51)
	) name9880 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001 ,
		_w11300_,
		_w13817_,
		_w13928_
	);
	LUT2 #(
		.INIT('h1)
	) name9881 (
		_w13927_,
		_w13928_,
		_w13929_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9882 (
		\sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w8798_,
		_w8801_,
		_w13888_,
		_w13930_
	);
	LUT4 #(
		.INIT('hba00)
	) name9883 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13888_,
		_w13931_
	);
	LUT3 #(
		.INIT('h15)
	) name9884 (
		\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w5656_,
		_w13783_,
		_w13932_
	);
	LUT2 #(
		.INIT('h1)
	) name9885 (
		_w13931_,
		_w13932_,
		_w13933_
	);
	LUT4 #(
		.INIT('hba00)
	) name9886 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13888_,
		_w13934_
	);
	LUT3 #(
		.INIT('h15)
	) name9887 (
		\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w5656_,
		_w13783_,
		_w13935_
	);
	LUT2 #(
		.INIT('h1)
	) name9888 (
		_w13934_,
		_w13935_,
		_w13936_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9889 (
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w8798_,
		_w8801_,
		_w12825_,
		_w13937_
	);
	LUT4 #(
		.INIT('hba00)
	) name9890 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13771_,
		_w13938_
	);
	LUT2 #(
		.INIT('h1)
	) name9891 (
		\pio_pmask_reg_DO_reg[7]/NET0131 ,
		_w13771_,
		_w13939_
	);
	LUT2 #(
		.INIT('h1)
	) name9892 (
		_w13938_,
		_w13939_,
		_w13940_
	);
	LUT4 #(
		.INIT('hba00)
	) name9893 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13771_,
		_w13941_
	);
	LUT2 #(
		.INIT('h1)
	) name9894 (
		\pio_pmask_reg_DO_reg[6]/NET0131 ,
		_w13771_,
		_w13942_
	);
	LUT2 #(
		.INIT('h1)
	) name9895 (
		_w13941_,
		_w13942_,
		_w13943_
	);
	LUT4 #(
		.INIT('hba00)
	) name9896 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13771_,
		_w13944_
	);
	LUT2 #(
		.INIT('h1)
	) name9897 (
		\pio_pmask_reg_DO_reg[3]/NET0131 ,
		_w13771_,
		_w13945_
	);
	LUT2 #(
		.INIT('h1)
	) name9898 (
		_w13944_,
		_w13945_,
		_w13946_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9899 (
		\pio_pmask_reg_DO_reg[11]/NET0131 ,
		_w8798_,
		_w8801_,
		_w13771_,
		_w13947_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9900 (
		\sice_ICYC_reg[16]/NET0131 ,
		\sice_ICYC_reg[17]/NET0131 ,
		\sice_ICYC_reg[18]/NET0131 ,
		_w13017_,
		_w13948_
	);
	LUT4 #(
		.INIT('hba00)
	) name9901 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13771_,
		_w13949_
	);
	LUT2 #(
		.INIT('h1)
	) name9902 (
		\pio_pmask_reg_DO_reg[2]/NET0131 ,
		_w13771_,
		_w13950_
	);
	LUT2 #(
		.INIT('h1)
	) name9903 (
		_w13949_,
		_w13950_,
		_w13951_
	);
	LUT4 #(
		.INIT('hba00)
	) name9904 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13771_,
		_w13952_
	);
	LUT2 #(
		.INIT('h1)
	) name9905 (
		\pio_pmask_reg_DO_reg[0]/NET0131 ,
		_w13771_,
		_w13953_
	);
	LUT2 #(
		.INIT('h1)
	) name9906 (
		_w13952_,
		_w13953_,
		_w13954_
	);
	LUT4 #(
		.INIT('hba00)
	) name9907 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13773_,
		_w13955_
	);
	LUT2 #(
		.INIT('h1)
	) name9908 (
		\PIO_oe[7]_pad ,
		_w13773_,
		_w13956_
	);
	LUT2 #(
		.INIT('h1)
	) name9909 (
		_w13955_,
		_w13956_,
		_w13957_
	);
	LUT4 #(
		.INIT('hba00)
	) name9910 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13773_,
		_w13958_
	);
	LUT2 #(
		.INIT('h1)
	) name9911 (
		\PIO_oe[6]_pad ,
		_w13773_,
		_w13959_
	);
	LUT2 #(
		.INIT('h1)
	) name9912 (
		_w13958_,
		_w13959_,
		_w13960_
	);
	LUT4 #(
		.INIT('hba00)
	) name9913 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13773_,
		_w13961_
	);
	LUT2 #(
		.INIT('h1)
	) name9914 (
		\PIO_oe[4]_pad ,
		_w13773_,
		_w13962_
	);
	LUT2 #(
		.INIT('h1)
	) name9915 (
		_w13961_,
		_w13962_,
		_w13963_
	);
	LUT4 #(
		.INIT('hba00)
	) name9916 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13773_,
		_w13964_
	);
	LUT2 #(
		.INIT('h1)
	) name9917 (
		\PIO_oe[2]_pad ,
		_w13773_,
		_w13965_
	);
	LUT2 #(
		.INIT('h1)
	) name9918 (
		_w13964_,
		_w13965_,
		_w13966_
	);
	LUT4 #(
		.INIT('hba00)
	) name9919 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13773_,
		_w13967_
	);
	LUT2 #(
		.INIT('h1)
	) name9920 (
		\PIO_oe[1]_pad ,
		_w13773_,
		_w13968_
	);
	LUT2 #(
		.INIT('h1)
	) name9921 (
		_w13967_,
		_w13968_,
		_w13969_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9922 (
		\PIO_oe[11]_pad ,
		_w8798_,
		_w8801_,
		_w13773_,
		_w13970_
	);
	LUT4 #(
		.INIT('hba00)
	) name9923 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13777_,
		_w13971_
	);
	LUT2 #(
		.INIT('h1)
	) name9924 (
		\memc_usysr_DO_reg[7]/NET0131 ,
		_w13777_,
		_w13972_
	);
	LUT2 #(
		.INIT('h1)
	) name9925 (
		_w13971_,
		_w13972_,
		_w13973_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9926 (
		\pio_pmask_reg_DO_reg[10]/NET0131 ,
		_w8757_,
		_w8760_,
		_w13771_,
		_w13974_
	);
	LUT4 #(
		.INIT('hba00)
	) name9927 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13771_,
		_w13975_
	);
	LUT2 #(
		.INIT('h1)
	) name9928 (
		\pio_pmask_reg_DO_reg[5]/NET0131 ,
		_w13771_,
		_w13976_
	);
	LUT2 #(
		.INIT('h1)
	) name9929 (
		_w13975_,
		_w13976_,
		_w13977_
	);
	LUT4 #(
		.INIT('hba00)
	) name9930 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13777_,
		_w13978_
	);
	LUT2 #(
		.INIT('h1)
	) name9931 (
		\memc_usysr_DO_reg[5]/NET0131 ,
		_w13777_,
		_w13979_
	);
	LUT2 #(
		.INIT('h1)
	) name9932 (
		_w13978_,
		_w13979_,
		_w13980_
	);
	LUT4 #(
		.INIT('hba00)
	) name9933 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13777_,
		_w13981_
	);
	LUT2 #(
		.INIT('h1)
	) name9934 (
		\memc_usysr_DO_reg[6]/NET0131 ,
		_w13777_,
		_w13982_
	);
	LUT2 #(
		.INIT('h1)
	) name9935 (
		_w13981_,
		_w13982_,
		_w13983_
	);
	LUT4 #(
		.INIT('hba00)
	) name9936 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13777_,
		_w13984_
	);
	LUT2 #(
		.INIT('h1)
	) name9937 (
		\memc_usysr_DO_reg[4]/NET0131 ,
		_w13777_,
		_w13985_
	);
	LUT2 #(
		.INIT('h1)
	) name9938 (
		_w13984_,
		_w13985_,
		_w13986_
	);
	LUT4 #(
		.INIT('hba00)
	) name9939 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13777_,
		_w13987_
	);
	LUT2 #(
		.INIT('h1)
	) name9940 (
		\memc_usysr_DO_reg[2]/NET0131 ,
		_w13777_,
		_w13988_
	);
	LUT2 #(
		.INIT('h1)
	) name9941 (
		_w13987_,
		_w13988_,
		_w13989_
	);
	LUT4 #(
		.INIT('hba00)
	) name9942 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13777_,
		_w13990_
	);
	LUT2 #(
		.INIT('h1)
	) name9943 (
		\memc_usysr_DO_reg[1]/NET0131 ,
		_w13777_,
		_w13991_
	);
	LUT2 #(
		.INIT('h1)
	) name9944 (
		_w13990_,
		_w13991_,
		_w13992_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9945 (
		\memc_usysr_DO_reg[15]/NET0131 ,
		_w8798_,
		_w8801_,
		_w13777_,
		_w13993_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9946 (
		\memc_usysr_DO_reg[14]/NET0131 ,
		_w8757_,
		_w8760_,
		_w13777_,
		_w13994_
	);
	LUT4 #(
		.INIT('hba00)
	) name9947 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13777_,
		_w13995_
	);
	LUT2 #(
		.INIT('h1)
	) name9948 (
		\memc_usysr_DO_reg[0]/NET0131 ,
		_w13777_,
		_w13996_
	);
	LUT2 #(
		.INIT('h1)
	) name9949 (
		_w13995_,
		_w13996_,
		_w13997_
	);
	LUT4 #(
		.INIT('h0222)
	) name9950 (
		\idma_RDcyc_reg/NET0131 ,
		_w12818_,
		_w12819_,
		_w12820_,
		_w13998_
	);
	LUT2 #(
		.INIT('he)
	) name9951 (
		_w13074_,
		_w13998_,
		_w13999_
	);
	LUT4 #(
		.INIT('h1000)
	) name9952 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w14000_
	);
	LUT3 #(
		.INIT('h80)
	) name9953 (
		_w9431_,
		_w11604_,
		_w14000_,
		_w14001_
	);
	LUT4 #(
		.INIT('h4000)
	) name9954 (
		\memc_MMR_web_reg/NET0131 ,
		_w9431_,
		_w11604_,
		_w14000_,
		_w14002_
	);
	LUT4 #(
		.INIT('h03aa)
	) name9955 (
		\tm_tcr_reg_DO_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w14002_,
		_w14003_
	);
	LUT4 #(
		.INIT('hba00)
	) name9956 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13773_,
		_w14004_
	);
	LUT2 #(
		.INIT('h1)
	) name9957 (
		\PIO_oe[3]_pad ,
		_w13773_,
		_w14005_
	);
	LUT2 #(
		.INIT('h1)
	) name9958 (
		_w14004_,
		_w14005_,
		_w14006_
	);
	LUT4 #(
		.INIT('h4000)
	) name9959 (
		\memc_MMR_web_reg/NET0131 ,
		_w5658_,
		_w5790_,
		_w9431_,
		_w14007_
	);
	LUT4 #(
		.INIT('hba00)
	) name9960 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w14007_,
		_w14008_
	);
	LUT2 #(
		.INIT('h1)
	) name9961 (
		\emc_WSCRext_reg_DO_reg[7]/NET0131 ,
		_w14007_,
		_w14009_
	);
	LUT2 #(
		.INIT('h1)
	) name9962 (
		_w14008_,
		_w14009_,
		_w14010_
	);
	LUT4 #(
		.INIT('hba00)
	) name9963 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w14007_,
		_w14011_
	);
	LUT2 #(
		.INIT('h1)
	) name9964 (
		\emc_WSCRext_reg_DO_reg[6]/NET0131 ,
		_w14007_,
		_w14012_
	);
	LUT2 #(
		.INIT('h1)
	) name9965 (
		_w14011_,
		_w14012_,
		_w14013_
	);
	LUT4 #(
		.INIT('hba00)
	) name9966 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w14007_,
		_w14014_
	);
	LUT2 #(
		.INIT('h1)
	) name9967 (
		\emc_WSCRext_reg_DO_reg[5]/NET0131 ,
		_w14007_,
		_w14015_
	);
	LUT2 #(
		.INIT('h1)
	) name9968 (
		_w14014_,
		_w14015_,
		_w14016_
	);
	LUT4 #(
		.INIT('hba00)
	) name9969 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w14007_,
		_w14017_
	);
	LUT2 #(
		.INIT('h1)
	) name9970 (
		\emc_WSCRext_reg_DO_reg[4]/NET0131 ,
		_w14007_,
		_w14018_
	);
	LUT2 #(
		.INIT('h1)
	) name9971 (
		_w14017_,
		_w14018_,
		_w14019_
	);
	LUT4 #(
		.INIT('hba00)
	) name9972 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w14007_,
		_w14020_
	);
	LUT2 #(
		.INIT('h1)
	) name9973 (
		\emc_WSCRext_reg_DO_reg[3]/NET0131 ,
		_w14007_,
		_w14021_
	);
	LUT2 #(
		.INIT('h1)
	) name9974 (
		_w14020_,
		_w14021_,
		_w14022_
	);
	LUT4 #(
		.INIT('hba00)
	) name9975 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w14007_,
		_w14023_
	);
	LUT2 #(
		.INIT('h1)
	) name9976 (
		\emc_WSCRext_reg_DO_reg[2]/NET0131 ,
		_w14007_,
		_w14024_
	);
	LUT2 #(
		.INIT('h1)
	) name9977 (
		_w14023_,
		_w14024_,
		_w14025_
	);
	LUT4 #(
		.INIT('hba00)
	) name9978 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w14007_,
		_w14026_
	);
	LUT2 #(
		.INIT('h1)
	) name9979 (
		\emc_WSCRext_reg_DO_reg[1]/NET0131 ,
		_w14007_,
		_w14027_
	);
	LUT2 #(
		.INIT('h1)
	) name9980 (
		_w14026_,
		_w14027_,
		_w14028_
	);
	LUT4 #(
		.INIT('hba00)
	) name9981 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w14007_,
		_w14029_
	);
	LUT2 #(
		.INIT('h1)
	) name9982 (
		\emc_WSCRext_reg_DO_reg[0]/NET0131 ,
		_w14007_,
		_w14030_
	);
	LUT2 #(
		.INIT('h1)
	) name9983 (
		_w14029_,
		_w14030_,
		_w14031_
	);
	LUT4 #(
		.INIT('hba00)
	) name9984 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13784_,
		_w14032_
	);
	LUT3 #(
		.INIT('h15)
	) name9985 (
		\sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w12621_,
		_w13783_,
		_w14033_
	);
	LUT2 #(
		.INIT('h1)
	) name9986 (
		_w14032_,
		_w14033_,
		_w14034_
	);
	LUT4 #(
		.INIT('hba00)
	) name9987 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13784_,
		_w14035_
	);
	LUT3 #(
		.INIT('h15)
	) name9988 (
		\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w12621_,
		_w13783_,
		_w14036_
	);
	LUT2 #(
		.INIT('h1)
	) name9989 (
		_w14035_,
		_w14036_,
		_w14037_
	);
	LUT4 #(
		.INIT('hba00)
	) name9990 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13784_,
		_w14038_
	);
	LUT3 #(
		.INIT('h15)
	) name9991 (
		\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w12621_,
		_w13783_,
		_w14039_
	);
	LUT2 #(
		.INIT('h1)
	) name9992 (
		_w14038_,
		_w14039_,
		_w14040_
	);
	LUT4 #(
		.INIT('hba00)
	) name9993 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13784_,
		_w14041_
	);
	LUT3 #(
		.INIT('h15)
	) name9994 (
		\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w12621_,
		_w13783_,
		_w14042_
	);
	LUT2 #(
		.INIT('h1)
	) name9995 (
		_w14041_,
		_w14042_,
		_w14043_
	);
	LUT4 #(
		.INIT('hba00)
	) name9996 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13784_,
		_w14044_
	);
	LUT3 #(
		.INIT('h15)
	) name9997 (
		\sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w12621_,
		_w13783_,
		_w14045_
	);
	LUT2 #(
		.INIT('h1)
	) name9998 (
		_w14044_,
		_w14045_,
		_w14046_
	);
	LUT4 #(
		.INIT('hba00)
	) name9999 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13784_,
		_w14047_
	);
	LUT3 #(
		.INIT('h15)
	) name10000 (
		\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w12621_,
		_w13783_,
		_w14048_
	);
	LUT2 #(
		.INIT('h1)
	) name10001 (
		_w14047_,
		_w14048_,
		_w14049_
	);
	LUT4 #(
		.INIT('hba00)
	) name10002 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13784_,
		_w14050_
	);
	LUT3 #(
		.INIT('h15)
	) name10003 (
		\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w12621_,
		_w13783_,
		_w14051_
	);
	LUT2 #(
		.INIT('h1)
	) name10004 (
		_w14050_,
		_w14051_,
		_w14052_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10005 (
		\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w8798_,
		_w8801_,
		_w13784_,
		_w14053_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10006 (
		\sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w8757_,
		_w8760_,
		_w13784_,
		_w14054_
	);
	LUT4 #(
		.INIT('hba00)
	) name10007 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13784_,
		_w14055_
	);
	LUT3 #(
		.INIT('h15)
	) name10008 (
		\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w12621_,
		_w13783_,
		_w14056_
	);
	LUT2 #(
		.INIT('h1)
	) name10009 (
		_w14055_,
		_w14056_,
		_w14057_
	);
	LUT4 #(
		.INIT('hba00)
	) name10010 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13812_,
		_w14058_
	);
	LUT2 #(
		.INIT('h1)
	) name10011 (
		\sport1_regs_AUTOreg_DO_reg[7]/NET0131 ,
		_w13812_,
		_w14059_
	);
	LUT2 #(
		.INIT('h1)
	) name10012 (
		_w14058_,
		_w14059_,
		_w14060_
	);
	LUT4 #(
		.INIT('hba00)
	) name10013 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13812_,
		_w14061_
	);
	LUT2 #(
		.INIT('h1)
	) name10014 (
		\sport1_regs_AUTOreg_DO_reg[6]/NET0131 ,
		_w13812_,
		_w14062_
	);
	LUT2 #(
		.INIT('h1)
	) name10015 (
		_w14061_,
		_w14062_,
		_w14063_
	);
	LUT4 #(
		.INIT('hba00)
	) name10016 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13812_,
		_w14064_
	);
	LUT2 #(
		.INIT('h1)
	) name10017 (
		\sport1_regs_AUTOreg_DO_reg[5]/NET0131 ,
		_w13812_,
		_w14065_
	);
	LUT2 #(
		.INIT('h1)
	) name10018 (
		_w14064_,
		_w14065_,
		_w14066_
	);
	LUT4 #(
		.INIT('hba00)
	) name10019 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13812_,
		_w14067_
	);
	LUT2 #(
		.INIT('h1)
	) name10020 (
		\sport1_regs_AUTOreg_DO_reg[4]/NET0131 ,
		_w13812_,
		_w14068_
	);
	LUT2 #(
		.INIT('h1)
	) name10021 (
		_w14067_,
		_w14068_,
		_w14069_
	);
	LUT4 #(
		.INIT('hba00)
	) name10022 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13812_,
		_w14070_
	);
	LUT2 #(
		.INIT('h1)
	) name10023 (
		\sport1_regs_AUTOreg_DO_reg[3]/NET0131 ,
		_w13812_,
		_w14071_
	);
	LUT2 #(
		.INIT('h1)
	) name10024 (
		_w14070_,
		_w14071_,
		_w14072_
	);
	LUT4 #(
		.INIT('hba00)
	) name10025 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13812_,
		_w14073_
	);
	LUT2 #(
		.INIT('h1)
	) name10026 (
		\sport1_regs_AUTOreg_DO_reg[2]/NET0131 ,
		_w13812_,
		_w14074_
	);
	LUT2 #(
		.INIT('h1)
	) name10027 (
		_w14073_,
		_w14074_,
		_w14075_
	);
	LUT4 #(
		.INIT('hba00)
	) name10028 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13812_,
		_w14076_
	);
	LUT2 #(
		.INIT('h1)
	) name10029 (
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w13812_,
		_w14077_
	);
	LUT2 #(
		.INIT('h1)
	) name10030 (
		_w14076_,
		_w14077_,
		_w14078_
	);
	LUT4 #(
		.INIT('hba00)
	) name10031 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13812_,
		_w14079_
	);
	LUT2 #(
		.INIT('h1)
	) name10032 (
		\sport1_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w13812_,
		_w14080_
	);
	LUT2 #(
		.INIT('h1)
	) name10033 (
		_w14079_,
		_w14080_,
		_w14081_
	);
	LUT4 #(
		.INIT('hba00)
	) name10034 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13773_,
		_w14082_
	);
	LUT2 #(
		.INIT('h1)
	) name10035 (
		\PIO_oe[5]_pad ,
		_w13773_,
		_w14083_
	);
	LUT2 #(
		.INIT('h1)
	) name10036 (
		_w14082_,
		_w14083_,
		_w14084_
	);
	LUT4 #(
		.INIT('hba00)
	) name10037 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13771_,
		_w14085_
	);
	LUT2 #(
		.INIT('h1)
	) name10038 (
		\pio_pmask_reg_DO_reg[4]/NET0131 ,
		_w13771_,
		_w14086_
	);
	LUT2 #(
		.INIT('h1)
	) name10039 (
		_w14085_,
		_w14086_,
		_w14087_
	);
	LUT4 #(
		.INIT('hba00)
	) name10040 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13773_,
		_w14088_
	);
	LUT2 #(
		.INIT('h1)
	) name10041 (
		\PIO_oe[0]_pad ,
		_w13773_,
		_w14089_
	);
	LUT2 #(
		.INIT('h1)
	) name10042 (
		_w14088_,
		_w14089_,
		_w14090_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10043 (
		\sport0_regs_AUTO_a_reg[14]/NET0131 ,
		_w9431_,
		_w11604_,
		_w12824_,
		_w14091_
	);
	LUT4 #(
		.INIT('h1000)
	) name10044 (
		_w8757_,
		_w8760_,
		_w11605_,
		_w12824_,
		_w14092_
	);
	LUT2 #(
		.INIT('he)
	) name10045 (
		_w14091_,
		_w14092_,
		_w14093_
	);
	LUT4 #(
		.INIT('hba00)
	) name10046 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13771_,
		_w14094_
	);
	LUT2 #(
		.INIT('h1)
	) name10047 (
		\pio_pmask_reg_DO_reg[1]/NET0131 ,
		_w13771_,
		_w14095_
	);
	LUT2 #(
		.INIT('h1)
	) name10048 (
		_w14094_,
		_w14095_,
		_w14096_
	);
	LUT4 #(
		.INIT('hba00)
	) name10049 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13777_,
		_w14097_
	);
	LUT2 #(
		.INIT('h1)
	) name10050 (
		\memc_usysr_DO_reg[3]/NET0131 ,
		_w13777_,
		_w14098_
	);
	LUT2 #(
		.INIT('h1)
	) name10051 (
		_w14097_,
		_w14098_,
		_w14099_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10052 (
		\PIO_oe[10]_pad ,
		_w8757_,
		_w8760_,
		_w13773_,
		_w14100_
	);
	LUT4 #(
		.INIT('h0400)
	) name10053 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[10]/NET0131 ,
		_w14101_
	);
	LUT2 #(
		.INIT('h4)
	) name10054 (
		\T_TMODE[0]_pad ,
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w14102_
	);
	LUT2 #(
		.INIT('h8)
	) name10055 (
		_w12801_,
		_w14102_,
		_w14103_
	);
	LUT2 #(
		.INIT('h1)
	) name10056 (
		\tm_TSR_TMP_reg[1]/NET0131 ,
		\tm_TSR_TMP_reg[2]/NET0131 ,
		_w14104_
	);
	LUT4 #(
		.INIT('h0001)
	) name10057 (
		\tm_TSR_TMP_reg[0]/NET0131 ,
		\tm_TSR_TMP_reg[1]/NET0131 ,
		\tm_TSR_TMP_reg[2]/NET0131 ,
		\tm_TSR_TMP_reg[3]/NET0131 ,
		_w14105_
	);
	LUT4 #(
		.INIT('h0001)
	) name10058 (
		\tm_TSR_TMP_reg[4]/NET0131 ,
		\tm_TSR_TMP_reg[5]/NET0131 ,
		\tm_TSR_TMP_reg[6]/NET0131 ,
		\tm_TSR_TMP_reg[7]/NET0131 ,
		_w14106_
	);
	LUT4 #(
		.INIT('h1555)
	) name10059 (
		\T_TMODE[0]_pad ,
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w14105_,
		_w14106_,
		_w14107_
	);
	LUT2 #(
		.INIT('h1)
	) name10060 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w14107_,
		_w14108_
	);
	LUT3 #(
		.INIT('h15)
	) name10061 (
		\T_TMODE[0]_pad ,
		_w12797_,
		_w12798_,
		_w14109_
	);
	LUT4 #(
		.INIT('h0444)
	) name10062 (
		\T_TMODE[0]_pad ,
		\tm_TCR_TMP_reg[8]/NET0131 ,
		_w12797_,
		_w12798_,
		_w14110_
	);
	LUT2 #(
		.INIT('h8)
	) name10063 (
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w14110_,
		_w14111_
	);
	LUT3 #(
		.INIT('h80)
	) name10064 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w14110_,
		_w14112_
	);
	LUT4 #(
		.INIT('hc999)
	) name10065 (
		\T_TMODE[0]_pad ,
		\tm_TCR_TMP_reg[8]/NET0131 ,
		_w12797_,
		_w12798_,
		_w14113_
	);
	LUT3 #(
		.INIT('h81)
	) name10066 (
		\tm_TCR_TMP_reg[8]/NET0131 ,
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w14109_,
		_w14114_
	);
	LUT4 #(
		.INIT('h8001)
	) name10067 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		\tm_TCR_TMP_reg[8]/NET0131 ,
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w14109_,
		_w14115_
	);
	LUT4 #(
		.INIT('ha66a)
	) name10068 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		_w14108_,
		_w14111_,
		_w14114_,
		_w14116_
	);
	LUT4 #(
		.INIT('h2333)
	) name10069 (
		\tm_tpr_reg_DO_reg[10]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w14117_
	);
	LUT4 #(
		.INIT('hfeaa)
	) name10070 (
		_w14101_,
		_w14103_,
		_w14116_,
		_w14117_,
		_w14118_
	);
	LUT4 #(
		.INIT('hba00)
	) name10071 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13888_,
		_w14119_
	);
	LUT3 #(
		.INIT('h15)
	) name10072 (
		\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w5656_,
		_w13783_,
		_w14120_
	);
	LUT2 #(
		.INIT('h1)
	) name10073 (
		_w14119_,
		_w14120_,
		_w14121_
	);
	LUT4 #(
		.INIT('hba00)
	) name10074 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13888_,
		_w14122_
	);
	LUT3 #(
		.INIT('h15)
	) name10075 (
		\sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w5656_,
		_w13783_,
		_w14123_
	);
	LUT2 #(
		.INIT('h1)
	) name10076 (
		_w14122_,
		_w14123_,
		_w14124_
	);
	LUT4 #(
		.INIT('hba00)
	) name10077 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13888_,
		_w14125_
	);
	LUT3 #(
		.INIT('h15)
	) name10078 (
		\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w5656_,
		_w13783_,
		_w14126_
	);
	LUT2 #(
		.INIT('h1)
	) name10079 (
		_w14125_,
		_w14126_,
		_w14127_
	);
	LUT4 #(
		.INIT('hba00)
	) name10080 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13888_,
		_w14128_
	);
	LUT3 #(
		.INIT('h15)
	) name10081 (
		\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w5656_,
		_w13783_,
		_w14129_
	);
	LUT2 #(
		.INIT('h1)
	) name10082 (
		_w14128_,
		_w14129_,
		_w14130_
	);
	LUT4 #(
		.INIT('hba00)
	) name10083 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13888_,
		_w14131_
	);
	LUT3 #(
		.INIT('h15)
	) name10084 (
		\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w5656_,
		_w13783_,
		_w14132_
	);
	LUT2 #(
		.INIT('h1)
	) name10085 (
		_w14131_,
		_w14132_,
		_w14133_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10086 (
		\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w8757_,
		_w8760_,
		_w13888_,
		_w14134_
	);
	LUT4 #(
		.INIT('hba00)
	) name10087 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13888_,
		_w14135_
	);
	LUT3 #(
		.INIT('h15)
	) name10088 (
		\sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w5656_,
		_w13783_,
		_w14136_
	);
	LUT2 #(
		.INIT('h1)
	) name10089 (
		_w14135_,
		_w14136_,
		_w14137_
	);
	LUT4 #(
		.INIT('hc444)
	) name10090 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[8]/NET0131 ,
		_w4073_,
		_w4084_,
		_w14138_
	);
	LUT3 #(
		.INIT('hf8)
	) name10091 (
		_w12271_,
		_w12272_,
		_w14138_,
		_w14139_
	);
	LUT4 #(
		.INIT('h4000)
	) name10092 (
		\memc_MMR_web_reg/NET0131 ,
		_w5643_,
		_w9431_,
		_w11604_,
		_w14140_
	);
	LUT2 #(
		.INIT('h8)
	) name10093 (
		_w5671_,
		_w14140_,
		_w14141_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10094 (
		\clkc_ckr_reg_DO_reg[9]/NET0131 ,
		_w7140_,
		_w7240_,
		_w14141_,
		_w14142_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10095 (
		\clkc_ckr_reg_DO_reg[8]/NET0131 ,
		_w7465_,
		_w7565_,
		_w14141_,
		_w14143_
	);
	LUT3 #(
		.INIT('hca)
	) name10096 (
		\clkc_ckr_reg_DO_reg[13]/NET0131 ,
		_w5760_,
		_w14141_,
		_w14144_
	);
	LUT3 #(
		.INIT('hca)
	) name10097 (
		\clkc_ckr_reg_DO_reg[12]/NET0131 ,
		_w6758_,
		_w14141_,
		_w14145_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10098 (
		\clkc_ckr_reg_DO_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w14141_,
		_w14146_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10099 (
		\clkc_ckr_reg_DO_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w14141_,
		_w14147_
	);
	LUT2 #(
		.INIT('h8)
	) name10100 (
		_w5809_,
		_w13783_,
		_w14148_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10101 (
		\tm_tpr_reg_DO_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w14148_,
		_w14149_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10102 (
		\tm_tpr_reg_DO_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w14148_,
		_w14150_
	);
	LUT2 #(
		.INIT('h8)
	) name10103 (
		_w5809_,
		_w14140_,
		_w14151_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10104 (
		\emc_WSCRreg_DO_reg[9]/NET0131 ,
		_w7140_,
		_w7240_,
		_w14151_,
		_w14152_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10105 (
		\emc_WSCRreg_DO_reg[8]/NET0131 ,
		_w7465_,
		_w7565_,
		_w14151_,
		_w14153_
	);
	LUT3 #(
		.INIT('hca)
	) name10106 (
		\emc_WSCRreg_DO_reg[13]/NET0131 ,
		_w5760_,
		_w14151_,
		_w14154_
	);
	LUT3 #(
		.INIT('hca)
	) name10107 (
		\emc_WSCRreg_DO_reg[12]/NET0131 ,
		_w6758_,
		_w14151_,
		_w14155_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10108 (
		\emc_WSCRreg_DO_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w14151_,
		_w14156_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10109 (
		\emc_WSCRreg_DO_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w14151_,
		_w14157_
	);
	LUT2 #(
		.INIT('h6)
	) name10110 (
		\sice_ICYC_reg[10]/NET0131 ,
		_w13015_,
		_w14158_
	);
	LUT2 #(
		.INIT('h6)
	) name10111 (
		\sice_IIRC_reg[10]/NET0131 ,
		_w13087_,
		_w14159_
	);
	LUT4 #(
		.INIT('haccc)
	) name10112 (
		\T_ED[7]_pad ,
		\emc_PMDreg_reg[7]/P0001 ,
		_w9937_,
		_w9943_,
		_w14160_
	);
	LUT4 #(
		.INIT('haccc)
	) name10113 (
		\T_ED[6]_pad ,
		\emc_PMDreg_reg[6]/P0001 ,
		_w9937_,
		_w9943_,
		_w14161_
	);
	LUT4 #(
		.INIT('haccc)
	) name10114 (
		\T_ED[5]_pad ,
		\emc_PMDreg_reg[5]/P0001 ,
		_w9937_,
		_w9943_,
		_w14162_
	);
	LUT4 #(
		.INIT('haccc)
	) name10115 (
		\T_ED[4]_pad ,
		\emc_PMDreg_reg[4]/P0001 ,
		_w9937_,
		_w9943_,
		_w14163_
	);
	LUT4 #(
		.INIT('haccc)
	) name10116 (
		\T_ED[3]_pad ,
		\emc_PMDreg_reg[3]/P0001 ,
		_w9937_,
		_w9943_,
		_w14164_
	);
	LUT4 #(
		.INIT('haccc)
	) name10117 (
		\T_ED[2]_pad ,
		\emc_PMDreg_reg[2]/P0001 ,
		_w9937_,
		_w9943_,
		_w14165_
	);
	LUT4 #(
		.INIT('haccc)
	) name10118 (
		\T_ED[1]_pad ,
		\emc_PMDreg_reg[1]/P0001 ,
		_w9937_,
		_w9943_,
		_w14166_
	);
	LUT4 #(
		.INIT('haccc)
	) name10119 (
		\T_ED[15]_pad ,
		\emc_PMDreg_reg[15]/P0001 ,
		_w9937_,
		_w9943_,
		_w14167_
	);
	LUT4 #(
		.INIT('haccc)
	) name10120 (
		\T_ED[14]_pad ,
		\emc_PMDreg_reg[14]/P0001 ,
		_w9937_,
		_w9943_,
		_w14168_
	);
	LUT4 #(
		.INIT('haccc)
	) name10121 (
		\T_ED[13]_pad ,
		\emc_PMDreg_reg[13]/P0001 ,
		_w9937_,
		_w9943_,
		_w14169_
	);
	LUT4 #(
		.INIT('haccc)
	) name10122 (
		\T_ED[12]_pad ,
		\emc_PMDreg_reg[12]/P0001 ,
		_w9937_,
		_w9943_,
		_w14170_
	);
	LUT4 #(
		.INIT('haccc)
	) name10123 (
		\T_ED[11]_pad ,
		\emc_PMDreg_reg[11]/P0001 ,
		_w9937_,
		_w9943_,
		_w14171_
	);
	LUT4 #(
		.INIT('haccc)
	) name10124 (
		\T_ED[10]_pad ,
		\emc_PMDreg_reg[10]/P0001 ,
		_w9937_,
		_w9943_,
		_w14172_
	);
	LUT4 #(
		.INIT('haccc)
	) name10125 (
		\T_ED[0]_pad ,
		\emc_PMDreg_reg[0]/P0001 ,
		_w9937_,
		_w9943_,
		_w14173_
	);
	LUT4 #(
		.INIT('hba00)
	) name10126 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w14141_,
		_w14174_
	);
	LUT3 #(
		.INIT('h15)
	) name10127 (
		\clkc_ckr_reg_DO_reg[7]/NET0131 ,
		_w5671_,
		_w14140_,
		_w14175_
	);
	LUT2 #(
		.INIT('h1)
	) name10128 (
		_w14174_,
		_w14175_,
		_w14176_
	);
	LUT4 #(
		.INIT('hba00)
	) name10129 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w14141_,
		_w14177_
	);
	LUT3 #(
		.INIT('h15)
	) name10130 (
		\clkc_ckr_reg_DO_reg[6]/NET0131 ,
		_w5671_,
		_w14140_,
		_w14178_
	);
	LUT2 #(
		.INIT('h1)
	) name10131 (
		_w14177_,
		_w14178_,
		_w14179_
	);
	LUT4 #(
		.INIT('hba00)
	) name10132 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w14141_,
		_w14180_
	);
	LUT3 #(
		.INIT('h15)
	) name10133 (
		\clkc_ckr_reg_DO_reg[5]/NET0131 ,
		_w5671_,
		_w14140_,
		_w14181_
	);
	LUT2 #(
		.INIT('h1)
	) name10134 (
		_w14180_,
		_w14181_,
		_w14182_
	);
	LUT4 #(
		.INIT('hba00)
	) name10135 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w14141_,
		_w14183_
	);
	LUT3 #(
		.INIT('h15)
	) name10136 (
		\clkc_ckr_reg_DO_reg[4]/NET0131 ,
		_w5671_,
		_w14140_,
		_w14184_
	);
	LUT2 #(
		.INIT('h1)
	) name10137 (
		_w14183_,
		_w14184_,
		_w14185_
	);
	LUT4 #(
		.INIT('hba00)
	) name10138 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w14141_,
		_w14186_
	);
	LUT3 #(
		.INIT('h15)
	) name10139 (
		\clkc_ckr_reg_DO_reg[3]/NET0131 ,
		_w5671_,
		_w14140_,
		_w14187_
	);
	LUT2 #(
		.INIT('h1)
	) name10140 (
		_w14186_,
		_w14187_,
		_w14188_
	);
	LUT4 #(
		.INIT('hba00)
	) name10141 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w14141_,
		_w14189_
	);
	LUT3 #(
		.INIT('h15)
	) name10142 (
		\clkc_ckr_reg_DO_reg[2]/NET0131 ,
		_w5671_,
		_w14140_,
		_w14190_
	);
	LUT2 #(
		.INIT('h1)
	) name10143 (
		_w14189_,
		_w14190_,
		_w14191_
	);
	LUT4 #(
		.INIT('hba00)
	) name10144 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w14141_,
		_w14192_
	);
	LUT3 #(
		.INIT('h15)
	) name10145 (
		\clkc_ckr_reg_DO_reg[1]/NET0131 ,
		_w5671_,
		_w14140_,
		_w14193_
	);
	LUT2 #(
		.INIT('h1)
	) name10146 (
		_w14192_,
		_w14193_,
		_w14194_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10147 (
		\clkc_ckr_reg_DO_reg[15]/NET0131 ,
		_w8798_,
		_w8801_,
		_w14141_,
		_w14195_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10148 (
		\clkc_ckr_reg_DO_reg[14]/NET0131 ,
		_w8757_,
		_w8760_,
		_w14141_,
		_w14196_
	);
	LUT4 #(
		.INIT('hba00)
	) name10149 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w14141_,
		_w14197_
	);
	LUT3 #(
		.INIT('h15)
	) name10150 (
		\clkc_ckr_reg_DO_reg[0]/NET0131 ,
		_w5671_,
		_w14140_,
		_w14198_
	);
	LUT2 #(
		.INIT('h1)
	) name10151 (
		_w14197_,
		_w14198_,
		_w14199_
	);
	LUT3 #(
		.INIT('h6c)
	) name10152 (
		\sice_ICYC_reg[16]/NET0131 ,
		\sice_ICYC_reg[17]/NET0131 ,
		_w13017_,
		_w14200_
	);
	LUT4 #(
		.INIT('h8000)
	) name10153 (
		\sice_IIRC_reg[13]/NET0131 ,
		\sice_IIRC_reg[14]/NET0131 ,
		\sice_IIRC_reg[15]/NET0131 ,
		_w13088_,
		_w14201_
	);
	LUT3 #(
		.INIT('h80)
	) name10154 (
		\sice_IIRC_reg[16]/NET0131 ,
		\sice_IIRC_reg[17]/NET0131 ,
		_w14201_,
		_w14202_
	);
	LUT3 #(
		.INIT('h6c)
	) name10155 (
		\sice_IIRC_reg[16]/NET0131 ,
		\sice_IIRC_reg[17]/NET0131 ,
		_w14201_,
		_w14203_
	);
	LUT2 #(
		.INIT('h6)
	) name10156 (
		\sice_IIRC_reg[13]/NET0131 ,
		_w13088_,
		_w14204_
	);
	LUT2 #(
		.INIT('h6)
	) name10157 (
		\sice_ICYC_reg[13]/NET0131 ,
		_w13016_,
		_w14205_
	);
	LUT4 #(
		.INIT('hba00)
	) name10158 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w14148_,
		_w14206_
	);
	LUT3 #(
		.INIT('h15)
	) name10159 (
		\tm_tpr_reg_DO_reg[7]/NET0131 ,
		_w5809_,
		_w13783_,
		_w14207_
	);
	LUT2 #(
		.INIT('h1)
	) name10160 (
		_w14206_,
		_w14207_,
		_w14208_
	);
	LUT4 #(
		.INIT('hba00)
	) name10161 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w14148_,
		_w14209_
	);
	LUT3 #(
		.INIT('h15)
	) name10162 (
		\tm_tpr_reg_DO_reg[6]/NET0131 ,
		_w5809_,
		_w13783_,
		_w14210_
	);
	LUT2 #(
		.INIT('h1)
	) name10163 (
		_w14209_,
		_w14210_,
		_w14211_
	);
	LUT4 #(
		.INIT('hba00)
	) name10164 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w14148_,
		_w14212_
	);
	LUT3 #(
		.INIT('h15)
	) name10165 (
		\tm_tpr_reg_DO_reg[5]/NET0131 ,
		_w5809_,
		_w13783_,
		_w14213_
	);
	LUT2 #(
		.INIT('h1)
	) name10166 (
		_w14212_,
		_w14213_,
		_w14214_
	);
	LUT4 #(
		.INIT('hba00)
	) name10167 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w14148_,
		_w14215_
	);
	LUT3 #(
		.INIT('h15)
	) name10168 (
		\tm_tpr_reg_DO_reg[3]/NET0131 ,
		_w5809_,
		_w13783_,
		_w14216_
	);
	LUT2 #(
		.INIT('h1)
	) name10169 (
		_w14215_,
		_w14216_,
		_w14217_
	);
	LUT4 #(
		.INIT('hba00)
	) name10170 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w14148_,
		_w14218_
	);
	LUT3 #(
		.INIT('h15)
	) name10171 (
		\tm_tpr_reg_DO_reg[2]/NET0131 ,
		_w5809_,
		_w13783_,
		_w14219_
	);
	LUT2 #(
		.INIT('h1)
	) name10172 (
		_w14218_,
		_w14219_,
		_w14220_
	);
	LUT4 #(
		.INIT('hba00)
	) name10173 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w14148_,
		_w14221_
	);
	LUT3 #(
		.INIT('h15)
	) name10174 (
		\tm_tpr_reg_DO_reg[1]/NET0131 ,
		_w5809_,
		_w13783_,
		_w14222_
	);
	LUT2 #(
		.INIT('h1)
	) name10175 (
		_w14221_,
		_w14222_,
		_w14223_
	);
	LUT4 #(
		.INIT('hba00)
	) name10176 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w14148_,
		_w14224_
	);
	LUT3 #(
		.INIT('h15)
	) name10177 (
		\tm_tpr_reg_DO_reg[4]/NET0131 ,
		_w5809_,
		_w13783_,
		_w14225_
	);
	LUT2 #(
		.INIT('h1)
	) name10178 (
		_w14224_,
		_w14225_,
		_w14226_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10179 (
		\tm_tpr_reg_DO_reg[15]/NET0131 ,
		_w8798_,
		_w8801_,
		_w14148_,
		_w14227_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10180 (
		\tm_tpr_reg_DO_reg[14]/NET0131 ,
		_w8757_,
		_w8760_,
		_w14148_,
		_w14228_
	);
	LUT4 #(
		.INIT('hba00)
	) name10181 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w14148_,
		_w14229_
	);
	LUT3 #(
		.INIT('h15)
	) name10182 (
		\tm_tpr_reg_DO_reg[0]/NET0131 ,
		_w5809_,
		_w13783_,
		_w14230_
	);
	LUT2 #(
		.INIT('h1)
	) name10183 (
		_w14229_,
		_w14230_,
		_w14231_
	);
	LUT4 #(
		.INIT('hba00)
	) name10184 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w14151_,
		_w14232_
	);
	LUT3 #(
		.INIT('h15)
	) name10185 (
		\emc_WSCRreg_DO_reg[7]/NET0131 ,
		_w5809_,
		_w14140_,
		_w14233_
	);
	LUT2 #(
		.INIT('h1)
	) name10186 (
		_w14232_,
		_w14233_,
		_w14234_
	);
	LUT4 #(
		.INIT('hba00)
	) name10187 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w14151_,
		_w14235_
	);
	LUT3 #(
		.INIT('h15)
	) name10188 (
		\emc_WSCRreg_DO_reg[6]/NET0131 ,
		_w5809_,
		_w14140_,
		_w14236_
	);
	LUT2 #(
		.INIT('h1)
	) name10189 (
		_w14235_,
		_w14236_,
		_w14237_
	);
	LUT4 #(
		.INIT('hba00)
	) name10190 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w14151_,
		_w14238_
	);
	LUT3 #(
		.INIT('h15)
	) name10191 (
		\emc_WSCRreg_DO_reg[5]/NET0131 ,
		_w5809_,
		_w14140_,
		_w14239_
	);
	LUT2 #(
		.INIT('h1)
	) name10192 (
		_w14238_,
		_w14239_,
		_w14240_
	);
	LUT4 #(
		.INIT('hba00)
	) name10193 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w14151_,
		_w14241_
	);
	LUT3 #(
		.INIT('h15)
	) name10194 (
		\emc_WSCRreg_DO_reg[4]/NET0131 ,
		_w5809_,
		_w14140_,
		_w14242_
	);
	LUT2 #(
		.INIT('h1)
	) name10195 (
		_w14241_,
		_w14242_,
		_w14243_
	);
	LUT4 #(
		.INIT('hba00)
	) name10196 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w14151_,
		_w14244_
	);
	LUT3 #(
		.INIT('h15)
	) name10197 (
		\emc_WSCRreg_DO_reg[3]/NET0131 ,
		_w5809_,
		_w14140_,
		_w14245_
	);
	LUT2 #(
		.INIT('h1)
	) name10198 (
		_w14244_,
		_w14245_,
		_w14246_
	);
	LUT4 #(
		.INIT('hba00)
	) name10199 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w14151_,
		_w14247_
	);
	LUT3 #(
		.INIT('h15)
	) name10200 (
		\emc_WSCRreg_DO_reg[2]/NET0131 ,
		_w5809_,
		_w14140_,
		_w14248_
	);
	LUT2 #(
		.INIT('h1)
	) name10201 (
		_w14247_,
		_w14248_,
		_w14249_
	);
	LUT4 #(
		.INIT('hba00)
	) name10202 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w14151_,
		_w14250_
	);
	LUT3 #(
		.INIT('h15)
	) name10203 (
		\emc_WSCRreg_DO_reg[1]/NET0131 ,
		_w5809_,
		_w14140_,
		_w14251_
	);
	LUT2 #(
		.INIT('h1)
	) name10204 (
		_w14250_,
		_w14251_,
		_w14252_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10205 (
		\emc_WSCRreg_DO_reg[14]/NET0131 ,
		_w8757_,
		_w8760_,
		_w14151_,
		_w14253_
	);
	LUT4 #(
		.INIT('hba00)
	) name10206 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w14151_,
		_w14254_
	);
	LUT3 #(
		.INIT('h15)
	) name10207 (
		\emc_WSCRreg_DO_reg[0]/NET0131 ,
		_w5809_,
		_w14140_,
		_w14255_
	);
	LUT2 #(
		.INIT('h1)
	) name10208 (
		_w14254_,
		_w14255_,
		_w14256_
	);
	LUT2 #(
		.INIT('h1)
	) name10209 (
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w14257_
	);
	LUT4 #(
		.INIT('hb41e)
	) name10210 (
		\ITFS1_pad ,
		\T_TFS1_pad ,
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w9407_,
		_w14258_
	);
	LUT2 #(
		.INIT('h2)
	) name10211 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_cfg_TFSgi_d_reg/NET0131 ,
		_w14259_
	);
	LUT2 #(
		.INIT('h8)
	) name10212 (
		_w14258_,
		_w14259_,
		_w14260_
	);
	LUT4 #(
		.INIT('h3500)
	) name10213 (
		\sport1_cfg_TFSg_d2_reg/NET0131 ,
		\sport1_cfg_TFSg_d3_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w14261_
	);
	LUT4 #(
		.INIT('hfb00)
	) name10214 (
		\sport1_cfg_TFSg_d1_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		\sport1_txctl_TCS_reg[0]/NET0131 ,
		_w14262_
	);
	LUT2 #(
		.INIT('h4)
	) name10215 (
		_w14261_,
		_w14262_,
		_w14263_
	);
	LUT4 #(
		.INIT('hd500)
	) name10216 (
		_w14257_,
		_w14258_,
		_w14259_,
		_w14263_,
		_w14264_
	);
	LUT3 #(
		.INIT('h13)
	) name10217 (
		\sport1_txctl_TCS_reg[0]/NET0131 ,
		\sport1_txctl_TCS_reg[1]/NET0131 ,
		\sport1_txctl_TCS_reg[2]/NET0131 ,
		_w14265_
	);
	LUT3 #(
		.INIT('h04)
	) name10218 (
		\sport1_txctl_TCS_reg[0]/NET0131 ,
		\sport1_txctl_TCS_reg[1]/NET0131 ,
		\sport1_txctl_TCS_reg[2]/NET0131 ,
		_w14266_
	);
	LUT4 #(
		.INIT('h0001)
	) name10219 (
		\sport1_txctl_Bcnt_reg[0]/NET0131 ,
		\sport1_txctl_Bcnt_reg[1]/NET0131 ,
		\sport1_txctl_Bcnt_reg[2]/NET0131 ,
		\sport1_txctl_Bcnt_reg[3]/NET0131 ,
		_w14267_
	);
	LUT3 #(
		.INIT('h8c)
	) name10220 (
		\sport1_txctl_Bcnt_reg[4]/NET0131 ,
		_w14266_,
		_w14267_,
		_w14268_
	);
	LUT4 #(
		.INIT('h001f)
	) name10221 (
		\sport1_txctl_TCS_reg[2]/NET0131 ,
		_w14264_,
		_w14265_,
		_w14268_,
		_w14269_
	);
	LUT4 #(
		.INIT('hffe0)
	) name10222 (
		\sport1_txctl_TCS_reg[2]/NET0131 ,
		_w14264_,
		_w14265_,
		_w14268_,
		_w14270_
	);
	LUT3 #(
		.INIT('hca)
	) name10223 (
		\sport1_txctl_TXSHT_reg[9]/P0001 ,
		\sport1_txctl_TX_reg[10]/P0001 ,
		_w14269_,
		_w14271_
	);
	LUT3 #(
		.INIT('h13)
	) name10224 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001 ,
		_w9894_,
		_w14272_
	);
	LUT4 #(
		.INIT('h0002)
	) name10225 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w14272_,
		_w14273_
	);
	LUT4 #(
		.INIT('h5700)
	) name10226 (
		_w11625_,
		_w12626_,
		_w12627_,
		_w14273_,
		_w14274_
	);
	LUT4 #(
		.INIT('h313b)
	) name10227 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001 ,
		_w11631_,
		_w11635_,
		_w14275_
	);
	LUT2 #(
		.INIT('h2)
	) name10228 (
		_w11624_,
		_w12361_,
		_w14276_
	);
	LUT4 #(
		.INIT('hff45)
	) name10229 (
		_w11624_,
		_w14274_,
		_w14275_,
		_w14276_,
		_w14277_
	);
	LUT2 #(
		.INIT('h8)
	) name10230 (
		_w9946_,
		_w12361_,
		_w14278_
	);
	LUT2 #(
		.INIT('h2)
	) name10231 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001 ,
		_w11656_,
		_w14279_
	);
	LUT3 #(
		.INIT('h01)
	) name10232 (
		_w9946_,
		_w11659_,
		_w14279_,
		_w14280_
	);
	LUT4 #(
		.INIT('hfd00)
	) name10233 (
		_w11655_,
		_w12626_,
		_w12627_,
		_w14280_,
		_w14281_
	);
	LUT2 #(
		.INIT('h1)
	) name10234 (
		_w14278_,
		_w14281_,
		_w14282_
	);
	LUT4 #(
		.INIT('h8000)
	) name10235 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11710_,
		_w11713_,
		_w11735_,
		_w14283_
	);
	LUT4 #(
		.INIT('h0004)
	) name10236 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[6]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w14284_
	);
	LUT4 #(
		.INIT('h4500)
	) name10237 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13382_,
		_w14285_
	);
	LUT3 #(
		.INIT('hfe)
	) name10238 (
		_w14284_,
		_w14283_,
		_w14285_,
		_w14286_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name10239 (
		_w10049_,
		_w10072_,
		_w10101_,
		_w10102_,
		_w14287_
	);
	LUT4 #(
		.INIT('hae00)
	) name10240 (
		_w10134_,
		_w10165_,
		_w10167_,
		_w14287_,
		_w14288_
	);
	LUT4 #(
		.INIT('h4f00)
	) name10241 (
		_w11250_,
		_w11285_,
		_w11289_,
		_w14288_,
		_w14289_
	);
	LUT4 #(
		.INIT('hf800)
	) name10242 (
		_w10134_,
		_w10165_,
		_w11291_,
		_w14287_,
		_w14290_
	);
	LUT4 #(
		.INIT('hbb2b)
	) name10243 (
		_w10049_,
		_w10072_,
		_w10101_,
		_w10102_,
		_w14291_
	);
	LUT2 #(
		.INIT('h4)
	) name10244 (
		_w14290_,
		_w14291_,
		_w14292_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name10245 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w6145_,
		_w7346_,
		_w14293_
	);
	LUT2 #(
		.INIT('h1)
	) name10246 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w14293_,
		_w14294_
	);
	LUT3 #(
		.INIT('h1a)
	) name10247 (
		_w10010_,
		_w10039_,
		_w14294_,
		_w14295_
	);
	LUT3 #(
		.INIT('h40)
	) name10248 (
		_w10010_,
		_w10039_,
		_w14293_,
		_w14296_
	);
	LUT4 #(
		.INIT('h0376)
	) name10249 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10010_,
		_w10039_,
		_w14293_,
		_w14297_
	);
	LUT4 #(
		.INIT('h32c8)
	) name10250 (
		_w9997_,
		_w10020_,
		_w10040_,
		_w14297_,
		_w14298_
	);
	LUT4 #(
		.INIT('hc936)
	) name10251 (
		_w9997_,
		_w10020_,
		_w10040_,
		_w14297_,
		_w14299_
	);
	LUT4 #(
		.INIT('h0014)
	) name10252 (
		_w10019_,
		_w10020_,
		_w10040_,
		_w10041_,
		_w14300_
	);
	LUT3 #(
		.INIT('hc8)
	) name10253 (
		_w10043_,
		_w14299_,
		_w14300_,
		_w14301_
	);
	LUT4 #(
		.INIT('h0515)
	) name10254 (
		_w9974_,
		_w10043_,
		_w14299_,
		_w14300_,
		_w14302_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name10255 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w7346_,
		_w7664_,
		_w14303_
	);
	LUT2 #(
		.INIT('h1)
	) name10256 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w14303_,
		_w14304_
	);
	LUT3 #(
		.INIT('h1a)
	) name10257 (
		_w10010_,
		_w14294_,
		_w14304_,
		_w14305_
	);
	LUT3 #(
		.INIT('h40)
	) name10258 (
		_w10010_,
		_w14294_,
		_w14303_,
		_w14306_
	);
	LUT4 #(
		.INIT('h0376)
	) name10259 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10010_,
		_w14294_,
		_w14303_,
		_w14307_
	);
	LUT4 #(
		.INIT('h0104)
	) name10260 (
		_w9997_,
		_w10020_,
		_w14295_,
		_w14307_,
		_w14308_
	);
	LUT4 #(
		.INIT('h36c9)
	) name10261 (
		_w9997_,
		_w10020_,
		_w14295_,
		_w14307_,
		_w14309_
	);
	LUT4 #(
		.INIT('h0014)
	) name10262 (
		_w10019_,
		_w10020_,
		_w14295_,
		_w14296_,
		_w14310_
	);
	LUT3 #(
		.INIT('h32)
	) name10263 (
		_w14298_,
		_w14309_,
		_w14310_,
		_w14311_
	);
	LUT3 #(
		.INIT('hc9)
	) name10264 (
		_w14298_,
		_w14309_,
		_w14310_,
		_w14312_
	);
	LUT4 #(
		.INIT('h5a69)
	) name10265 (
		_w9974_,
		_w14298_,
		_w14309_,
		_w14310_,
		_w14313_
	);
	LUT3 #(
		.INIT('h4b)
	) name10266 (
		_w9974_,
		_w14301_,
		_w14312_,
		_w14314_
	);
	LUT3 #(
		.INIT('h04)
	) name10267 (
		_w9974_,
		_w10044_,
		_w10046_,
		_w14315_
	);
	LUT3 #(
		.INIT('h36)
	) name10268 (
		_w10043_,
		_w14299_,
		_w14300_,
		_w14316_
	);
	LUT2 #(
		.INIT('h6)
	) name10269 (
		_w14315_,
		_w14316_,
		_w14317_
	);
	LUT3 #(
		.INIT('ha8)
	) name10270 (
		_w9974_,
		_w10043_,
		_w14300_,
		_w14318_
	);
	LUT3 #(
		.INIT('h01)
	) name10271 (
		_w14315_,
		_w14316_,
		_w14318_,
		_w14319_
	);
	LUT3 #(
		.INIT('h49)
	) name10272 (
		_w9974_,
		_w10044_,
		_w10046_,
		_w14320_
	);
	LUT3 #(
		.INIT('h0b)
	) name10273 (
		_w10037_,
		_w10048_,
		_w14320_,
		_w14321_
	);
	LUT4 #(
		.INIT('h0abb)
	) name10274 (
		_w14314_,
		_w14317_,
		_w14319_,
		_w14321_,
		_w14322_
	);
	LUT4 #(
		.INIT('habaf)
	) name10275 (
		_w14314_,
		_w14317_,
		_w14319_,
		_w14321_,
		_w14323_
	);
	LUT4 #(
		.INIT('hf400)
	) name10276 (
		_w14289_,
		_w14292_,
		_w14322_,
		_w14323_,
		_w14324_
	);
	LUT4 #(
		.INIT('h5051)
	) name10277 (
		_w9974_,
		_w14298_,
		_w14309_,
		_w14310_,
		_w14325_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name10278 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w7664_,
		_w8026_,
		_w14326_
	);
	LUT2 #(
		.INIT('h1)
	) name10279 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w14326_,
		_w14327_
	);
	LUT3 #(
		.INIT('h1a)
	) name10280 (
		_w10010_,
		_w14304_,
		_w14327_,
		_w14328_
	);
	LUT3 #(
		.INIT('h40)
	) name10281 (
		_w10010_,
		_w14304_,
		_w14326_,
		_w14329_
	);
	LUT4 #(
		.INIT('h0376)
	) name10282 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w10010_,
		_w14304_,
		_w14326_,
		_w14330_
	);
	LUT4 #(
		.INIT('h0104)
	) name10283 (
		_w9997_,
		_w10020_,
		_w14305_,
		_w14330_,
		_w14331_
	);
	LUT4 #(
		.INIT('h36c9)
	) name10284 (
		_w9997_,
		_w10020_,
		_w14305_,
		_w14330_,
		_w14332_
	);
	LUT4 #(
		.INIT('h3328)
	) name10285 (
		_w10019_,
		_w10020_,
		_w14305_,
		_w14306_,
		_w14333_
	);
	LUT3 #(
		.INIT('h36)
	) name10286 (
		_w14308_,
		_w14332_,
		_w14333_,
		_w14334_
	);
	LUT4 #(
		.INIT('ha596)
	) name10287 (
		_w9974_,
		_w14308_,
		_w14332_,
		_w14333_,
		_w14335_
	);
	LUT4 #(
		.INIT('h0516)
	) name10288 (
		_w9974_,
		_w14308_,
		_w14332_,
		_w14333_,
		_w14336_
	);
	LUT3 #(
		.INIT('h0e)
	) name10289 (
		_w14325_,
		_w14335_,
		_w14336_,
		_w14337_
	);
	LUT4 #(
		.INIT('hfd75)
	) name10290 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w5713_,
		_w8026_,
		_w14338_
	);
	LUT2 #(
		.INIT('h1)
	) name10291 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w14338_,
		_w14339_
	);
	LUT2 #(
		.INIT('h1)
	) name10292 (
		_w10010_,
		_w14339_,
		_w14340_
	);
	LUT3 #(
		.INIT('h1a)
	) name10293 (
		_w10010_,
		_w14327_,
		_w14339_,
		_w14341_
	);
	LUT3 #(
		.INIT('h04)
	) name10294 (
		_w10010_,
		_w14327_,
		_w14339_,
		_w14342_
	);
	LUT3 #(
		.INIT('he1)
	) name10295 (
		_w10010_,
		_w14327_,
		_w14339_,
		_w14343_
	);
	LUT4 #(
		.INIT('h0104)
	) name10296 (
		_w9997_,
		_w10020_,
		_w14328_,
		_w14343_,
		_w14344_
	);
	LUT4 #(
		.INIT('h36c9)
	) name10297 (
		_w9997_,
		_w10020_,
		_w14328_,
		_w14343_,
		_w14345_
	);
	LUT4 #(
		.INIT('h3328)
	) name10298 (
		_w10019_,
		_w10020_,
		_w14328_,
		_w14329_,
		_w14346_
	);
	LUT3 #(
		.INIT('h01)
	) name10299 (
		_w14331_,
		_w14345_,
		_w14346_,
		_w14347_
	);
	LUT3 #(
		.INIT('hc8)
	) name10300 (
		_w14331_,
		_w14345_,
		_w14346_,
		_w14348_
	);
	LUT3 #(
		.INIT('h36)
	) name10301 (
		_w14331_,
		_w14345_,
		_w14346_,
		_w14349_
	);
	LUT4 #(
		.INIT('h0001)
	) name10302 (
		_w9974_,
		_w14308_,
		_w14332_,
		_w14333_,
		_w14350_
	);
	LUT2 #(
		.INIT('h9)
	) name10303 (
		_w14349_,
		_w14350_,
		_w14351_
	);
	LUT4 #(
		.INIT('h5a49)
	) name10304 (
		_w9974_,
		_w14298_,
		_w14309_,
		_w14310_,
		_w14352_
	);
	LUT3 #(
		.INIT('h0e)
	) name10305 (
		_w14302_,
		_w14313_,
		_w14352_,
		_w14353_
	);
	LUT3 #(
		.INIT('h4b)
	) name10306 (
		_w9974_,
		_w14311_,
		_w14334_,
		_w14354_
	);
	LUT2 #(
		.INIT('h4)
	) name10307 (
		_w14353_,
		_w14354_,
		_w14355_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name10308 (
		_w14337_,
		_w14351_,
		_w14353_,
		_w14354_,
		_w14356_
	);
	LUT2 #(
		.INIT('h2)
	) name10309 (
		_w14353_,
		_w14354_,
		_w14357_
	);
	LUT4 #(
		.INIT('hdd4d)
	) name10310 (
		_w14337_,
		_w14351_,
		_w14353_,
		_w14354_,
		_w14358_
	);
	LUT2 #(
		.INIT('h4)
	) name10311 (
		_w5713_,
		_w11131_,
		_w14359_
	);
	LUT4 #(
		.INIT('h3328)
	) name10312 (
		_w10019_,
		_w10020_,
		_w14341_,
		_w14342_,
		_w14360_
	);
	LUT4 #(
		.INIT('ha596)
	) name10313 (
		_w14340_,
		_w14344_,
		_w14359_,
		_w14360_,
		_w14361_
	);
	LUT4 #(
		.INIT('hac53)
	) name10314 (
		_w14347_,
		_w14348_,
		_w14350_,
		_w14361_,
		_w14362_
	);
	LUT3 #(
		.INIT('hca)
	) name10315 (
		_w10019_,
		_w10020_,
		_w14341_,
		_w14363_
	);
	LUT2 #(
		.INIT('h9)
	) name10316 (
		_w14362_,
		_w14363_,
		_w14364_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name10317 (
		_w14324_,
		_w14356_,
		_w14358_,
		_w14364_,
		_w14365_
	);
	LUT2 #(
		.INIT('h9)
	) name10318 (
		_w14337_,
		_w14351_,
		_w14366_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name10319 (
		_w14324_,
		_w14355_,
		_w14357_,
		_w14366_,
		_w14367_
	);
	LUT3 #(
		.INIT('h72)
	) name10320 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14365_,
		_w14367_,
		_w14368_
	);
	LUT3 #(
		.INIT('ha8)
	) name10321 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12626_,
		_w12627_,
		_w14369_
	);
	LUT3 #(
		.INIT('he0)
	) name10322 (
		_w11420_,
		_w11421_,
		_w11465_,
		_w14370_
	);
	LUT3 #(
		.INIT('ha8)
	) name10323 (
		_w11537_,
		_w11397_,
		_w11519_,
		_w14371_
	);
	LUT3 #(
		.INIT('h02)
	) name10324 (
		_w11386_,
		_w11335_,
		_w11593_,
		_w14372_
	);
	LUT3 #(
		.INIT('h01)
	) name10325 (
		_w14371_,
		_w14372_,
		_w14370_,
		_w14373_
	);
	LUT2 #(
		.INIT('h8)
	) name10326 (
		_w11424_,
		_w11854_,
		_w14374_
	);
	LUT3 #(
		.INIT('he0)
	) name10327 (
		_w11552_,
		_w11474_,
		_w11873_,
		_w14375_
	);
	LUT3 #(
		.INIT('h0e)
	) name10328 (
		_w11393_,
		_w11589_,
		_w11844_,
		_w14376_
	);
	LUT3 #(
		.INIT('h01)
	) name10329 (
		_w14375_,
		_w14376_,
		_w14374_,
		_w14377_
	);
	LUT4 #(
		.INIT('hddd0)
	) name10330 (
		_w11864_,
		_w11953_,
		_w11957_,
		_w11950_,
		_w14378_
	);
	LUT3 #(
		.INIT('he0)
	) name10331 (
		_w11552_,
		_w11474_,
		_w11852_,
		_w14379_
	);
	LUT2 #(
		.INIT('h1)
	) name10332 (
		_w11592_,
		_w12506_,
		_w14380_
	);
	LUT3 #(
		.INIT('h10)
	) name10333 (
		_w14379_,
		_w14380_,
		_w14378_,
		_w14381_
	);
	LUT3 #(
		.INIT('hc8)
	) name10334 (
		_w11547_,
		_w11874_,
		_w11976_,
		_w14382_
	);
	LUT4 #(
		.INIT('ha820)
	) name10335 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001 ,
		_w14383_
	);
	LUT4 #(
		.INIT('h000e)
	) name10336 (
		_w11954_,
		_w12500_,
		_w12754_,
		_w14383_,
		_w14384_
	);
	LUT2 #(
		.INIT('h4)
	) name10337 (
		_w14382_,
		_w14384_,
		_w14385_
	);
	LUT4 #(
		.INIT('h8000)
	) name10338 (
		_w14377_,
		_w14381_,
		_w14385_,
		_w14373_,
		_w14386_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name10339 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12740_,
		_w14369_,
		_w14386_,
		_w14387_
	);
	LUT3 #(
		.INIT('he2)
	) name10340 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001 ,
		_w11946_,
		_w14387_,
		_w14388_
	);
	LUT3 #(
		.INIT('he2)
	) name10341 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001 ,
		_w12048_,
		_w14387_,
		_w14389_
	);
	LUT2 #(
		.INIT('h9)
	) name10342 (
		_w14353_,
		_w14354_,
		_w14390_
	);
	LUT2 #(
		.INIT('h9)
	) name10343 (
		_w14324_,
		_w14390_,
		_w14391_
	);
	LUT3 #(
		.INIT('h41)
	) name10344 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14324_,
		_w14390_,
		_w14392_
	);
	LUT3 #(
		.INIT('hf8)
	) name10345 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14367_,
		_w14392_,
		_w14393_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name10346 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001 ,
		_w12216_,
		_w12219_,
		_w13380_,
		_w14394_
	);
	LUT4 #(
		.INIT('h2000)
	) name10347 (
		\core_c_dec_satMR_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14395_
	);
	LUT4 #(
		.INIT('haa80)
	) name10348 (
		_w4102_,
		_w12392_,
		_w13525_,
		_w14395_,
		_w14396_
	);
	LUT4 #(
		.INIT('h2000)
	) name10349 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14397_
	);
	LUT4 #(
		.INIT('haa80)
	) name10350 (
		_w4102_,
		_w5044_,
		_w13525_,
		_w14397_,
		_w14398_
	);
	LUT3 #(
		.INIT('h13)
	) name10351 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 ,
		_w9894_,
		_w14399_
	);
	LUT4 #(
		.INIT('h0002)
	) name10352 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w14399_,
		_w14400_
	);
	LUT4 #(
		.INIT('h5700)
	) name10353 (
		_w12282_,
		_w12560_,
		_w12561_,
		_w14400_,
		_w14401_
	);
	LUT4 #(
		.INIT('h313b)
	) name10354 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 ,
		_w11308_,
		_w11635_,
		_w14402_
	);
	LUT3 #(
		.INIT('h45)
	) name10355 (
		_w11624_,
		_w14401_,
		_w14402_,
		_w14403_
	);
	LUT2 #(
		.INIT('h6)
	) name10356 (
		_w10869_,
		_w10921_,
		_w14404_
	);
	LUT2 #(
		.INIT('h9)
	) name10357 (
		_w12246_,
		_w14404_,
		_w14405_
	);
	LUT3 #(
		.INIT('h28)
	) name10358 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12246_,
		_w14404_,
		_w14406_
	);
	LUT4 #(
		.INIT('h050d)
	) name10359 (
		_w11175_,
		_w11243_,
		_w11234_,
		_w12245_,
		_w14407_
	);
	LUT2 #(
		.INIT('h6)
	) name10360 (
		_w11183_,
		_w11184_,
		_w14408_
	);
	LUT4 #(
		.INIT('hcd32)
	) name10361 (
		_w11181_,
		_w11235_,
		_w14407_,
		_w14408_,
		_w14409_
	);
	LUT3 #(
		.INIT('h23)
	) name10362 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14406_,
		_w14409_,
		_w14410_
	);
	LUT4 #(
		.INIT('h80c4)
	) name10363 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w14405_,
		_w14409_,
		_w14411_
	);
	LUT2 #(
		.INIT('he)
	) name10364 (
		_w14403_,
		_w14411_,
		_w14412_
	);
	LUT2 #(
		.INIT('h8)
	) name10365 (
		_w5760_,
		_w12825_,
		_w14413_
	);
	LUT4 #(
		.INIT('hff35)
	) name10366 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w14414_
	);
	LUT4 #(
		.INIT('h35ff)
	) name10367 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w14415_
	);
	LUT2 #(
		.INIT('h8)
	) name10368 (
		_w14414_,
		_w14415_,
		_w14416_
	);
	LUT4 #(
		.INIT('hbf00)
	) name10369 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14416_,
		_w14417_
	);
	LUT4 #(
		.INIT('h1000)
	) name10370 (
		\core_eu_ec_cun_TERM_E_reg[3]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14418_
	);
	LUT3 #(
		.INIT('h02)
	) name10371 (
		_w4142_,
		_w14418_,
		_w14417_,
		_w14419_
	);
	LUT4 #(
		.INIT('hff35)
	) name10372 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w14420_
	);
	LUT4 #(
		.INIT('h35ff)
	) name10373 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w14421_
	);
	LUT2 #(
		.INIT('h8)
	) name10374 (
		_w14420_,
		_w14421_,
		_w14422_
	);
	LUT4 #(
		.INIT('hbf00)
	) name10375 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14422_,
		_w14423_
	);
	LUT4 #(
		.INIT('h1000)
	) name10376 (
		\core_eu_ec_cun_TERM_E_reg[2]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14424_
	);
	LUT3 #(
		.INIT('h02)
	) name10377 (
		_w4142_,
		_w14424_,
		_w14423_,
		_w14425_
	);
	LUT3 #(
		.INIT('h13)
	) name10378 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 ,
		_w9894_,
		_w14426_
	);
	LUT4 #(
		.INIT('h0002)
	) name10379 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w14426_,
		_w14427_
	);
	LUT4 #(
		.INIT('h313b)
	) name10380 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 ,
		_w11308_,
		_w11635_,
		_w14428_
	);
	LUT4 #(
		.INIT('h2f00)
	) name10381 (
		_w12282_,
		_w12673_,
		_w14427_,
		_w14428_,
		_w14429_
	);
	LUT2 #(
		.INIT('h1)
	) name10382 (
		_w11624_,
		_w14429_,
		_w14430_
	);
	LUT2 #(
		.INIT('h9)
	) name10383 (
		_w11276_,
		_w11280_,
		_w14431_
	);
	LUT4 #(
		.INIT('he01f)
	) name10384 (
		_w11250_,
		_w11273_,
		_w11286_,
		_w14431_,
		_w14432_
	);
	LUT2 #(
		.INIT('h4)
	) name10385 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14432_,
		_w14433_
	);
	LUT4 #(
		.INIT('h0a28)
	) name10386 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11287_,
		_w12217_,
		_w12218_,
		_w14434_
	);
	LUT2 #(
		.INIT('he)
	) name10387 (
		_w14433_,
		_w14434_,
		_w14435_
	);
	LUT4 #(
		.INIT('heeec)
	) name10388 (
		_w11624_,
		_w14430_,
		_w14433_,
		_w14434_,
		_w14436_
	);
	LUT4 #(
		.INIT('h2000)
	) name10389 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14437_
	);
	LUT4 #(
		.INIT('haa08)
	) name10390 (
		_w4102_,
		_w8174_,
		_w13338_,
		_w14437_,
		_w14438_
	);
	LUT4 #(
		.INIT('h2000)
	) name10391 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14439_
	);
	LUT4 #(
		.INIT('h00bf)
	) name10392 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w4818_,
		_w5047_,
		_w14439_,
		_w14440_
	);
	LUT2 #(
		.INIT('h2)
	) name10393 (
		_w4102_,
		_w14440_,
		_w14441_
	);
	LUT4 #(
		.INIT('h2000)
	) name10394 (
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14442_
	);
	LUT4 #(
		.INIT('haa80)
	) name10395 (
		_w4102_,
		_w8174_,
		_w13334_,
		_w14442_,
		_w14443_
	);
	LUT4 #(
		.INIT('h4c08)
	) name10396 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w14405_,
		_w14409_,
		_w14444_
	);
	LUT2 #(
		.INIT('h2)
	) name10397 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001 ,
		_w11310_,
		_w14445_
	);
	LUT3 #(
		.INIT('h01)
	) name10398 (
		_w9946_,
		_w12442_,
		_w14445_,
		_w14446_
	);
	LUT4 #(
		.INIT('hfd00)
	) name10399 (
		_w12440_,
		_w12560_,
		_w12561_,
		_w14446_,
		_w14447_
	);
	LUT2 #(
		.INIT('h1)
	) name10400 (
		_w14444_,
		_w14447_,
		_w14448_
	);
	LUT2 #(
		.INIT('h8)
	) name10401 (
		\clkc_CTR_cnt_reg[0]/NET0131 ,
		\clkc_CTR_cnt_reg[1]/NET0131 ,
		_w14449_
	);
	LUT2 #(
		.INIT('h7)
	) name10402 (
		\clkc_CTR_cnt_reg[0]/NET0131 ,
		\clkc_CTR_cnt_reg[1]/NET0131 ,
		_w14450_
	);
	LUT3 #(
		.INIT('h08)
	) name10403 (
		\clkc_CTR_cnt_reg[0]/NET0131 ,
		\clkc_CTR_cnt_reg[1]/NET0131 ,
		\clkc_RSTtext_reg/P0001 ,
		_w14451_
	);
	LUT3 #(
		.INIT('hf7)
	) name10404 (
		\clkc_CTR_cnt_reg[0]/NET0131 ,
		\clkc_CTR_cnt_reg[1]/NET0131 ,
		\clkc_RSTtext_reg/P0001 ,
		_w14452_
	);
	LUT2 #(
		.INIT('h1)
	) name10405 (
		\sice_GOICE_1_reg/NET0131 ,
		\sice_GOICE_2_reg/NET0131 ,
		_w14453_
	);
	LUT2 #(
		.INIT('he)
	) name10406 (
		\sice_GOICE_1_reg/NET0131 ,
		\sice_GOICE_2_reg/NET0131 ,
		_w14454_
	);
	LUT3 #(
		.INIT('h0e)
	) name10407 (
		\sice_GOICE_1_reg/NET0131 ,
		\sice_GOICE_2_reg/NET0131 ,
		\sice_GOICE_s1_reg/NET0131 ,
		_w14455_
	);
	LUT3 #(
		.INIT('h20)
	) name10408 (
		_w4140_,
		_w14455_,
		_w14451_,
		_w14456_
	);
	LUT4 #(
		.INIT('h9ccc)
	) name10409 (
		\bdma_BSreq_reg/NET0131 ,
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w4764_,
		_w12604_,
		_w14457_
	);
	LUT2 #(
		.INIT('h4)
	) name10410 (
		_w9413_,
		_w14457_,
		_w14458_
	);
	LUT4 #(
		.INIT('h0002)
	) name10411 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w14459_
	);
	LUT4 #(
		.INIT('h0800)
	) name10412 (
		T_IMS_pad,
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w14460_
	);
	LUT2 #(
		.INIT('h8)
	) name10413 (
		_w14459_,
		_w14460_,
		_w14461_
	);
	LUT2 #(
		.INIT('h4)
	) name10414 (
		\sice_IRST_reg/NET0131 ,
		\sice_SPC_reg[18]/P0001 ,
		_w14462_
	);
	LUT3 #(
		.INIT('h80)
	) name10415 (
		_w14459_,
		_w14460_,
		_w14462_,
		_w14463_
	);
	LUT2 #(
		.INIT('h4)
	) name10416 (
		\sice_CLR_I_reg/NET0131 ,
		\sice_SPC_reg[21]/P0001 ,
		_w14464_
	);
	LUT3 #(
		.INIT('h80)
	) name10417 (
		_w14459_,
		_w14460_,
		_w14464_,
		_w14465_
	);
	LUT4 #(
		.INIT('h4000)
	) name10418 (
		_w11698_,
		_w11705_,
		_w11724_,
		_w11728_,
		_w14466_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name10419 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11697_,
		_w11705_,
		_w11720_,
		_w14467_
	);
	LUT2 #(
		.INIT('h8)
	) name10420 (
		_w14466_,
		_w14467_,
		_w14468_
	);
	LUT2 #(
		.INIT('h8)
	) name10421 (
		_w11736_,
		_w14468_,
		_w14469_
	);
	LUT4 #(
		.INIT('h4000)
	) name10422 (
		_w11698_,
		_w11705_,
		_w11724_,
		_w11733_,
		_w14470_
	);
	LUT2 #(
		.INIT('h1)
	) name10423 (
		_w11729_,
		_w14470_,
		_w14471_
	);
	LUT4 #(
		.INIT('h8000)
	) name10424 (
		_w11710_,
		_w11713_,
		_w11729_,
		_w11735_,
		_w14472_
	);
	LUT2 #(
		.INIT('h4)
	) name10425 (
		_w11725_,
		_w14472_,
		_w14473_
	);
	LUT4 #(
		.INIT('ha251)
	) name10426 (
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w11679_,
		_w11680_,
		_w11681_,
		_w14474_
	);
	LUT4 #(
		.INIT('h59a6)
	) name10427 (
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w11679_,
		_w11680_,
		_w11681_,
		_w14475_
	);
	LUT4 #(
		.INIT('hbe9c)
	) name10428 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11682_,
		_w11683_,
		_w14474_,
		_w14476_
	);
	LUT3 #(
		.INIT('h04)
	) name10429 (
		_w11698_,
		_w11705_,
		_w14476_,
		_w14477_
	);
	LUT4 #(
		.INIT('h4f00)
	) name10430 (
		_w11721_,
		_w11725_,
		_w14472_,
		_w14477_,
		_w14478_
	);
	LUT4 #(
		.INIT('h4eb4)
	) name10431 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11677_,
		_w11682_,
		_w11683_,
		_w14479_
	);
	LUT4 #(
		.INIT('h4000)
	) name10432 (
		_w11698_,
		_w11705_,
		_w11724_,
		_w14479_,
		_w14480_
	);
	LUT2 #(
		.INIT('h2)
	) name10433 (
		_w11721_,
		_w14480_,
		_w14481_
	);
	LUT2 #(
		.INIT('h8)
	) name10434 (
		_w14472_,
		_w14481_,
		_w14482_
	);
	LUT4 #(
		.INIT('h0080)
	) name10435 (
		_w11710_,
		_w11713_,
		_w11718_,
		_w11734_,
		_w14483_
	);
	LUT4 #(
		.INIT('h0800)
	) name10436 (
		_w11710_,
		_w11713_,
		_w11729_,
		_w11735_,
		_w14484_
	);
	LUT2 #(
		.INIT('h1)
	) name10437 (
		_w14483_,
		_w14484_,
		_w14485_
	);
	LUT4 #(
		.INIT('h0155)
	) name10438 (
		_w14471_,
		_w14478_,
		_w14482_,
		_w14485_,
		_w14486_
	);
	LUT4 #(
		.INIT('hc040)
	) name10439 (
		_w11710_,
		_w11713_,
		_w11718_,
		_w14486_,
		_w14487_
	);
	LUT4 #(
		.INIT('ha020)
	) name10440 (
		_w11714_,
		_w11718_,
		_w11734_,
		_w14486_,
		_w14488_
	);
	LUT3 #(
		.INIT('h04)
	) name10441 (
		_w11698_,
		_w11705_,
		_w14479_,
		_w14489_
	);
	LUT2 #(
		.INIT('h2)
	) name10442 (
		_w11710_,
		_w11713_,
		_w14490_
	);
	LUT4 #(
		.INIT('h00df)
	) name10443 (
		_w11736_,
		_w14489_,
		_w14468_,
		_w14490_,
		_w14491_
	);
	LUT4 #(
		.INIT('hab00)
	) name10444 (
		_w14469_,
		_w14487_,
		_w14488_,
		_w14491_,
		_w14492_
	);
	LUT4 #(
		.INIT('h1011)
	) name10445 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w6054_,
		_w6173_,
		_w6175_,
		_w14493_
	);
	LUT4 #(
		.INIT('h007b)
	) name10446 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w14492_,
		_w14493_,
		_w14494_
	);
	LUT3 #(
		.INIT('h8b)
	) name10447 (
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w13383_,
		_w14494_,
		_w14495_
	);
	LUT2 #(
		.INIT('h4)
	) name10448 (
		\sice_CLR_M_reg/NET0131 ,
		\sice_SPC_reg[22]/P0001 ,
		_w14496_
	);
	LUT3 #(
		.INIT('h80)
	) name10449 (
		_w14459_,
		_w14460_,
		_w14496_,
		_w14497_
	);
	LUT3 #(
		.INIT('hea)
	) name10450 (
		\clkc_OSCoff_reg/NET0131 ,
		\clkc_OSCoff_set_reg/P0001 ,
		\clkc_SLEEP_reg/NET0131 ,
		_w14498_
	);
	LUT4 #(
		.INIT('h135f)
	) name10451 (
		\pio_PINT_reg[11]/NET0131 ,
		\pio_PINT_reg[5]/NET0131 ,
		\pio_pmask_reg_DO_reg[11]/NET0131 ,
		\pio_pmask_reg_DO_reg[5]/NET0131 ,
		_w14499_
	);
	LUT4 #(
		.INIT('h135f)
	) name10452 (
		\pio_PINT_reg[2]/NET0131 ,
		\pio_PINT_reg[9]/NET0131 ,
		\pio_pmask_reg_DO_reg[2]/NET0131 ,
		\pio_pmask_reg_DO_reg[9]/NET0131 ,
		_w14500_
	);
	LUT2 #(
		.INIT('h8)
	) name10453 (
		_w14499_,
		_w14500_,
		_w14501_
	);
	LUT4 #(
		.INIT('h135f)
	) name10454 (
		\pio_PINT_reg[10]/NET0131 ,
		\pio_PINT_reg[6]/NET0131 ,
		\pio_pmask_reg_DO_reg[10]/NET0131 ,
		\pio_pmask_reg_DO_reg[6]/NET0131 ,
		_w14502_
	);
	LUT4 #(
		.INIT('h135f)
	) name10455 (
		\pio_PINT_reg[0]/NET0131 ,
		\pio_PINT_reg[4]/NET0131 ,
		\pio_pmask_reg_DO_reg[0]/NET0131 ,
		\pio_pmask_reg_DO_reg[4]/NET0131 ,
		_w14503_
	);
	LUT4 #(
		.INIT('h135f)
	) name10456 (
		\pio_PINT_reg[3]/NET0131 ,
		\pio_PINT_reg[8]/NET0131 ,
		\pio_pmask_reg_DO_reg[3]/NET0131 ,
		\pio_pmask_reg_DO_reg[8]/NET0131 ,
		_w14504_
	);
	LUT4 #(
		.INIT('h135f)
	) name10457 (
		\pio_PINT_reg[1]/NET0131 ,
		\pio_PINT_reg[7]/NET0131 ,
		\pio_pmask_reg_DO_reg[1]/NET0131 ,
		\pio_pmask_reg_DO_reg[7]/NET0131 ,
		_w14505_
	);
	LUT4 #(
		.INIT('h8000)
	) name10458 (
		_w14504_,
		_w14505_,
		_w14502_,
		_w14503_,
		_w14506_
	);
	LUT2 #(
		.INIT('h7)
	) name10459 (
		_w14501_,
		_w14506_,
		_w14507_
	);
	LUT2 #(
		.INIT('hd)
	) name10460 (
		_w4140_,
		_w12802_,
		_w14508_
	);
	LUT2 #(
		.INIT('he)
	) name10461 (
		\tm_WR_TCR_KEEP_TO_TMCLK_p_reg/NET0131 ,
		\tm_WR_TCR_p_reg/P0001 ,
		_w14509_
	);
	LUT2 #(
		.INIT('h2)
	) name10462 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001 ,
		_w11310_,
		_w14510_
	);
	LUT3 #(
		.INIT('h01)
	) name10463 (
		_w9946_,
		_w12442_,
		_w14510_,
		_w14511_
	);
	LUT3 #(
		.INIT('h70)
	) name10464 (
		_w12440_,
		_w12673_,
		_w14511_,
		_w14512_
	);
	LUT4 #(
		.INIT('h00fd)
	) name10465 (
		_w9946_,
		_w14433_,
		_w14434_,
		_w14512_,
		_w14513_
	);
	LUT4 #(
		.INIT('h35ff)
	) name10466 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w14514_
	);
	LUT4 #(
		.INIT('hff35)
	) name10467 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w14515_
	);
	LUT2 #(
		.INIT('h8)
	) name10468 (
		_w14514_,
		_w14515_,
		_w14516_
	);
	LUT4 #(
		.INIT('hbf00)
	) name10469 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14516_,
		_w14517_
	);
	LUT4 #(
		.INIT('h1000)
	) name10470 (
		\core_eu_ec_cun_TERM_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14518_
	);
	LUT3 #(
		.INIT('h02)
	) name10471 (
		_w4142_,
		_w14518_,
		_w14517_,
		_w14519_
	);
	LUT4 #(
		.INIT('hff35)
	) name10472 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w14520_
	);
	LUT4 #(
		.INIT('h35ff)
	) name10473 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w14521_
	);
	LUT2 #(
		.INIT('h8)
	) name10474 (
		_w14520_,
		_w14521_,
		_w14522_
	);
	LUT4 #(
		.INIT('hbf00)
	) name10475 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14522_,
		_w14523_
	);
	LUT4 #(
		.INIT('h1000)
	) name10476 (
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14524_
	);
	LUT3 #(
		.INIT('h02)
	) name10477 (
		_w4142_,
		_w14524_,
		_w14523_,
		_w14525_
	);
	LUT3 #(
		.INIT('h40)
	) name10478 (
		_w11710_,
		_w11713_,
		_w11729_,
		_w14526_
	);
	LUT4 #(
		.INIT('h0e5b)
	) name10479 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_txctl_TX_reg[0]/P0001 ,
		_w11678_,
		_w11680_,
		_w14527_
	);
	LUT3 #(
		.INIT('h40)
	) name10480 (
		_w11698_,
		_w11705_,
		_w14527_,
		_w14528_
	);
	LUT2 #(
		.INIT('h2)
	) name10481 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w11680_,
		_w14529_
	);
	LUT3 #(
		.INIT('h0b)
	) name10482 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w14475_,
		_w14529_,
		_w14530_
	);
	LUT3 #(
		.INIT('h04)
	) name10483 (
		_w11698_,
		_w11705_,
		_w14530_,
		_w14531_
	);
	LUT4 #(
		.INIT('hf780)
	) name10484 (
		_w11726_,
		_w14472_,
		_w14531_,
		_w14528_,
		_w14532_
	);
	LUT4 #(
		.INIT('h3323)
	) name10485 (
		_w11725_,
		_w14484_,
		_w14472_,
		_w14477_,
		_w14533_
	);
	LUT3 #(
		.INIT('h13)
	) name10486 (
		_w14489_,
		_w14483_,
		_w14484_,
		_w14534_
	);
	LUT4 #(
		.INIT('h1f00)
	) name10487 (
		_w14473_,
		_w14532_,
		_w14533_,
		_w14534_,
		_w14535_
	);
	LUT3 #(
		.INIT('h8a)
	) name10488 (
		_w11718_,
		_w11721_,
		_w14483_,
		_w14536_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name10489 (
		_w11698_,
		_w11705_,
		_w11717_,
		_w11724_,
		_w14537_
	);
	LUT3 #(
		.INIT('h08)
	) name10490 (
		_w11710_,
		_w11713_,
		_w14537_,
		_w14538_
	);
	LUT4 #(
		.INIT('h1055)
	) name10491 (
		_w14526_,
		_w14535_,
		_w14536_,
		_w14538_,
		_w14539_
	);
	LUT2 #(
		.INIT('h4)
	) name10492 (
		_w11713_,
		_w11734_,
		_w14540_
	);
	LUT4 #(
		.INIT('h00f7)
	) name10493 (
		_w11736_,
		_w14468_,
		_w14531_,
		_w14540_,
		_w14541_
	);
	LUT4 #(
		.INIT('h56aa)
	) name10494 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w14469_,
		_w14539_,
		_w14541_,
		_w14542_
	);
	LUT4 #(
		.INIT('h040e)
	) name10495 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w6897_,
		_w13383_,
		_w14542_,
		_w14543_
	);
	LUT4 #(
		.INIT('h0004)
	) name10496 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w14544_
	);
	LUT2 #(
		.INIT('he)
	) name10497 (
		_w14543_,
		_w14544_,
		_w14545_
	);
	LUT4 #(
		.INIT('h1011)
	) name10498 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w6054_,
		_w6173_,
		_w6175_,
		_w14546_
	);
	LUT2 #(
		.INIT('h6)
	) name10499 (
		_w13109_,
		_w13117_,
		_w14547_
	);
	LUT3 #(
		.INIT('h15)
	) name10500 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w13137_,
		_w13139_,
		_w14548_
	);
	LUT3 #(
		.INIT('h40)
	) name10501 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w14549_
	);
	LUT2 #(
		.INIT('h1)
	) name10502 (
		_w13158_,
		_w14549_,
		_w14550_
	);
	LUT4 #(
		.INIT('h7d00)
	) name10503 (
		_w13155_,
		_w14547_,
		_w14548_,
		_w14550_,
		_w14551_
	);
	LUT4 #(
		.INIT('hafac)
	) name10504 (
		\sport0_rxctl_RXSHT_reg[3]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w14552_
	);
	LUT4 #(
		.INIT('h0002)
	) name10505 (
		\sport0_rxctl_RX_reg[3]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w14553_
	);
	LUT4 #(
		.INIT('hffb0)
	) name10506 (
		_w14546_,
		_w14551_,
		_w14552_,
		_w14553_,
		_w14554_
	);
	LUT3 #(
		.INIT('h13)
	) name10507 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 ,
		_w9894_,
		_w14555_
	);
	LUT4 #(
		.INIT('h0002)
	) name10508 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w14555_,
		_w14556_
	);
	LUT4 #(
		.INIT('h1f00)
	) name10509 (
		_w11626_,
		_w11627_,
		_w12282_,
		_w14556_,
		_w14557_
	);
	LUT4 #(
		.INIT('h313b)
	) name10510 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 ,
		_w11308_,
		_w11635_,
		_w14558_
	);
	LUT3 #(
		.INIT('h45)
	) name10511 (
		_w11624_,
		_w14557_,
		_w14558_,
		_w14559_
	);
	LUT2 #(
		.INIT('h9)
	) name10512 (
		_w11178_,
		_w11180_,
		_w14560_
	);
	LUT2 #(
		.INIT('h9)
	) name10513 (
		_w14407_,
		_w14560_,
		_w14561_
	);
	LUT4 #(
		.INIT('h4c08)
	) name10514 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w14409_,
		_w14561_,
		_w14562_
	);
	LUT2 #(
		.INIT('he)
	) name10515 (
		_w14559_,
		_w14562_,
		_w14563_
	);
	LUT4 #(
		.INIT('h80c4)
	) name10516 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w14409_,
		_w14561_,
		_w14564_
	);
	LUT2 #(
		.INIT('h2)
	) name10517 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001 ,
		_w11310_,
		_w14565_
	);
	LUT3 #(
		.INIT('h01)
	) name10518 (
		_w9946_,
		_w12442_,
		_w14565_,
		_w14566_
	);
	LUT4 #(
		.INIT('hef00)
	) name10519 (
		_w11626_,
		_w11627_,
		_w12440_,
		_w14566_,
		_w14567_
	);
	LUT2 #(
		.INIT('h1)
	) name10520 (
		_w14564_,
		_w14567_,
		_w14568_
	);
	LUT2 #(
		.INIT('h8)
	) name10521 (
		\core_c_dec_IDLE_Eg_reg/P0001 ,
		_w4106_,
		_w14569_
	);
	LUT4 #(
		.INIT('h1000)
	) name10522 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4428_,
		_w8172_,
		_w13446_,
		_w14570_
	);
	LUT4 #(
		.INIT('h4000)
	) name10523 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w5026_,
		_w5028_,
		_w5045_,
		_w14571_
	);
	LUT3 #(
		.INIT('hea)
	) name10524 (
		_w14569_,
		_w14570_,
		_w14571_,
		_w14572_
	);
	LUT4 #(
		.INIT('h4000)
	) name10525 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4861_,
		_w14573_
	);
	LUT2 #(
		.INIT('h2)
	) name10526 (
		_w8181_,
		_w8183_,
		_w14574_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name10527 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w8170_,
		_w14573_,
		_w14574_,
		_w14575_
	);
	LUT2 #(
		.INIT('h1)
	) name10528 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w14576_
	);
	LUT3 #(
		.INIT('h45)
	) name10529 (
		_w4971_,
		_w9911_,
		_w14576_,
		_w14577_
	);
	LUT4 #(
		.INIT('h6f00)
	) name10530 (
		_w9480_,
		_w9625_,
		_w9632_,
		_w9759_,
		_w14578_
	);
	LUT4 #(
		.INIT('hf969)
	) name10531 (
		_w9480_,
		_w9625_,
		_w9632_,
		_w9757_,
		_w14579_
	);
	LUT2 #(
		.INIT('h4)
	) name10532 (
		_w14578_,
		_w14579_,
		_w14580_
	);
	LUT4 #(
		.INIT('h00b0)
	) name10533 (
		_w9593_,
		_w9612_,
		_w9615_,
		_w9655_,
		_w14581_
	);
	LUT4 #(
		.INIT('h5541)
	) name10534 (
		_w9456_,
		_w9480_,
		_w9643_,
		_w9650_,
		_w14582_
	);
	LUT3 #(
		.INIT('h65)
	) name10535 (
		_w14580_,
		_w14581_,
		_w14582_,
		_w14583_
	);
	LUT4 #(
		.INIT('h10b0)
	) name10536 (
		_w9455_,
		_w9890_,
		_w9895_,
		_w14583_,
		_w14584_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10537 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001 ,
		_w9451_,
		_w9453_,
		_w9894_,
		_w14585_
	);
	LUT2 #(
		.INIT('he)
	) name10538 (
		_w14584_,
		_w14585_,
		_w14586_
	);
	LUT4 #(
		.INIT('h028a)
	) name10539 (
		_w9454_,
		_w9455_,
		_w9890_,
		_w14583_,
		_w14587_
	);
	LUT2 #(
		.INIT('h2)
	) name10540 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001 ,
		_w9454_,
		_w14588_
	);
	LUT2 #(
		.INIT('he)
	) name10541 (
		_w14587_,
		_w14588_,
		_w14589_
	);
	LUT4 #(
		.INIT('he8eb)
	) name10542 (
		\sport1_txctl_TCS_reg[0]/NET0131 ,
		\sport1_txctl_TCS_reg[1]/NET0131 ,
		\sport1_txctl_TCS_reg[2]/NET0131 ,
		_w14264_,
		_w14590_
	);
	LUT3 #(
		.INIT('h40)
	) name10543 (
		\sport1_txctl_Bcnt_reg[4]/NET0131 ,
		_w14266_,
		_w14267_,
		_w14591_
	);
	LUT4 #(
		.INIT('h0001)
	) name10544 (
		\sport1_txctl_Wcnt_reg[4]/NET0131 ,
		\sport1_txctl_Wcnt_reg[5]/NET0131 ,
		\sport1_txctl_Wcnt_reg[6]/NET0131 ,
		\sport1_txctl_Wcnt_reg[7]/NET0131 ,
		_w14592_
	);
	LUT4 #(
		.INIT('h0001)
	) name10545 (
		\sport1_txctl_Wcnt_reg[0]/NET0131 ,
		\sport1_txctl_Wcnt_reg[1]/NET0131 ,
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		\sport1_txctl_Wcnt_reg[3]/NET0131 ,
		_w14593_
	);
	LUT2 #(
		.INIT('h8)
	) name10546 (
		_w14592_,
		_w14593_,
		_w14594_
	);
	LUT3 #(
		.INIT('hea)
	) name10547 (
		_w14590_,
		_w14591_,
		_w14594_,
		_w14595_
	);
	LUT4 #(
		.INIT('he8eb)
	) name10548 (
		\sport0_txctl_TCS_reg[0]/NET0131 ,
		\sport0_txctl_TCS_reg[1]/NET0131 ,
		\sport0_txctl_TCS_reg[2]/NET0131 ,
		_w12547_,
		_w14596_
	);
	LUT3 #(
		.INIT('h40)
	) name10549 (
		\sport0_txctl_Bcnt_reg[4]/NET0131 ,
		_w12549_,
		_w12550_,
		_w14597_
	);
	LUT4 #(
		.INIT('h0001)
	) name10550 (
		\sport0_txctl_Wcnt_reg[4]/NET0131 ,
		\sport0_txctl_Wcnt_reg[5]/NET0131 ,
		\sport0_txctl_Wcnt_reg[6]/NET0131 ,
		\sport0_txctl_Wcnt_reg[7]/NET0131 ,
		_w14598_
	);
	LUT4 #(
		.INIT('h0001)
	) name10551 (
		\sport0_txctl_Wcnt_reg[0]/NET0131 ,
		\sport0_txctl_Wcnt_reg[1]/NET0131 ,
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		\sport0_txctl_Wcnt_reg[3]/NET0131 ,
		_w14599_
	);
	LUT2 #(
		.INIT('h8)
	) name10552 (
		_w14598_,
		_w14599_,
		_w14600_
	);
	LUT3 #(
		.INIT('hea)
	) name10553 (
		_w14596_,
		_w14597_,
		_w14600_,
		_w14601_
	);
	LUT4 #(
		.INIT('h4c44)
	) name10554 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		\core_c_psq_SSTAT_reg[6]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w14602_
	);
	LUT3 #(
		.INIT('h0e)
	) name10555 (
		_w4971_,
		_w12899_,
		_w14602_,
		_w14603_
	);
	LUT4 #(
		.INIT('h0001)
	) name10556 (
		\core_c_psq_lpstk_ptr_reg[2]/NET0131 ,
		_w4434_,
		_w4971_,
		_w12899_,
		_w14604_
	);
	LUT2 #(
		.INIT('h1)
	) name10557 (
		_w14603_,
		_w14604_,
		_w14605_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10558 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14606_
	);
	LUT4 #(
		.INIT('h8000)
	) name10559 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14607_
	);
	LUT2 #(
		.INIT('he)
	) name10560 (
		_w14606_,
		_w14607_,
		_w14608_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10561 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14609_
	);
	LUT4 #(
		.INIT('h8000)
	) name10562 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14610_
	);
	LUT2 #(
		.INIT('he)
	) name10563 (
		_w14609_,
		_w14610_,
		_w14611_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10564 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14612_
	);
	LUT4 #(
		.INIT('h8000)
	) name10565 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14613_
	);
	LUT2 #(
		.INIT('he)
	) name10566 (
		_w14612_,
		_w14613_,
		_w14614_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10567 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14615_
	);
	LUT4 #(
		.INIT('h8000)
	) name10568 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14616_
	);
	LUT2 #(
		.INIT('he)
	) name10569 (
		_w14615_,
		_w14616_,
		_w14617_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10570 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14618_
	);
	LUT4 #(
		.INIT('h8000)
	) name10571 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14619_
	);
	LUT2 #(
		.INIT('he)
	) name10572 (
		_w14618_,
		_w14619_,
		_w14620_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10573 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14621_
	);
	LUT4 #(
		.INIT('h8000)
	) name10574 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14622_
	);
	LUT2 #(
		.INIT('he)
	) name10575 (
		_w14621_,
		_w14622_,
		_w14623_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10576 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14624_
	);
	LUT4 #(
		.INIT('h8000)
	) name10577 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14625_
	);
	LUT2 #(
		.INIT('he)
	) name10578 (
		_w14624_,
		_w14625_,
		_w14626_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10579 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14627_
	);
	LUT4 #(
		.INIT('h8000)
	) name10580 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14628_
	);
	LUT2 #(
		.INIT('he)
	) name10581 (
		_w14627_,
		_w14628_,
		_w14629_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10582 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14630_
	);
	LUT4 #(
		.INIT('h8000)
	) name10583 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14631_
	);
	LUT2 #(
		.INIT('he)
	) name10584 (
		_w14630_,
		_w14631_,
		_w14632_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10585 (
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14633_
	);
	LUT4 #(
		.INIT('h8000)
	) name10586 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14634_
	);
	LUT2 #(
		.INIT('he)
	) name10587 (
		_w14633_,
		_w14634_,
		_w14635_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10588 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14636_
	);
	LUT4 #(
		.INIT('h8000)
	) name10589 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14637_
	);
	LUT2 #(
		.INIT('he)
	) name10590 (
		_w14636_,
		_w14637_,
		_w14638_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10591 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14639_
	);
	LUT4 #(
		.INIT('h8000)
	) name10592 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14640_
	);
	LUT2 #(
		.INIT('he)
	) name10593 (
		_w14639_,
		_w14640_,
		_w14641_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10594 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14642_
	);
	LUT4 #(
		.INIT('h8000)
	) name10595 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14643_
	);
	LUT2 #(
		.INIT('he)
	) name10596 (
		_w14642_,
		_w14643_,
		_w14644_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10597 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14645_
	);
	LUT4 #(
		.INIT('h8000)
	) name10598 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4073_,
		_w4084_,
		_w13325_,
		_w14646_
	);
	LUT2 #(
		.INIT('he)
	) name10599 (
		_w14645_,
		_w14646_,
		_w14647_
	);
	LUT4 #(
		.INIT('h808c)
	) name10600 (
		\core_c_dec_Post1_E_reg/P0001 ,
		_w4102_,
		_w4104_,
		_w13544_,
		_w14648_
	);
	LUT4 #(
		.INIT('h00bf)
	) name10601 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12390_,
		_w14649_
	);
	LUT3 #(
		.INIT('h3a)
	) name10602 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		_w12978_,
		_w14649_,
		_w14650_
	);
	LUT2 #(
		.INIT('h2)
	) name10603 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		_w14649_,
		_w14651_
	);
	LUT4 #(
		.INIT('h3700)
	) name10604 (
		_w5041_,
		_w6608_,
		_w12984_,
		_w14649_,
		_w14652_
	);
	LUT2 #(
		.INIT('he)
	) name10605 (
		_w14651_,
		_w14652_,
		_w14653_
	);
	LUT3 #(
		.INIT('h23)
	) name10606 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14654_
	);
	LUT3 #(
		.INIT('h1b)
	) name10607 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		_w14655_
	);
	LUT4 #(
		.INIT('h0023)
	) name10608 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14655_,
		_w14656_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name10609 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14657_
	);
	LUT2 #(
		.INIT('he)
	) name10610 (
		_w14656_,
		_w14657_,
		_w14658_
	);
	LUT3 #(
		.INIT('h1b)
	) name10611 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		_w14659_
	);
	LUT4 #(
		.INIT('h0023)
	) name10612 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14659_,
		_w14660_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name10613 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14661_
	);
	LUT2 #(
		.INIT('he)
	) name10614 (
		_w14660_,
		_w14661_,
		_w14662_
	);
	LUT3 #(
		.INIT('h1b)
	) name10615 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		_w14663_
	);
	LUT4 #(
		.INIT('h0023)
	) name10616 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14663_,
		_w14664_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name10617 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14665_
	);
	LUT2 #(
		.INIT('he)
	) name10618 (
		_w14664_,
		_w14665_,
		_w14666_
	);
	LUT3 #(
		.INIT('h1b)
	) name10619 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		_w14667_
	);
	LUT4 #(
		.INIT('h0023)
	) name10620 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14667_,
		_w14668_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name10621 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14669_
	);
	LUT2 #(
		.INIT('he)
	) name10622 (
		_w14668_,
		_w14669_,
		_w14670_
	);
	LUT3 #(
		.INIT('h1b)
	) name10623 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		_w14671_
	);
	LUT4 #(
		.INIT('h0023)
	) name10624 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14671_,
		_w14672_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name10625 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14673_
	);
	LUT2 #(
		.INIT('he)
	) name10626 (
		_w14672_,
		_w14673_,
		_w14674_
	);
	LUT3 #(
		.INIT('h1b)
	) name10627 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		_w14675_
	);
	LUT4 #(
		.INIT('h0023)
	) name10628 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14675_,
		_w14676_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name10629 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14677_
	);
	LUT2 #(
		.INIT('he)
	) name10630 (
		_w14676_,
		_w14677_,
		_w14678_
	);
	LUT3 #(
		.INIT('h1b)
	) name10631 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		_w14679_
	);
	LUT4 #(
		.INIT('h0023)
	) name10632 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14679_,
		_w14680_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name10633 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14681_
	);
	LUT2 #(
		.INIT('he)
	) name10634 (
		_w14680_,
		_w14681_,
		_w14682_
	);
	LUT3 #(
		.INIT('h1b)
	) name10635 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		_w14683_
	);
	LUT4 #(
		.INIT('h0023)
	) name10636 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14683_,
		_w14684_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name10637 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14685_
	);
	LUT2 #(
		.INIT('he)
	) name10638 (
		_w14684_,
		_w14685_,
		_w14686_
	);
	LUT3 #(
		.INIT('h1b)
	) name10639 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w14687_
	);
	LUT4 #(
		.INIT('h0023)
	) name10640 (
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14687_,
		_w14688_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name10641 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4064_,
		_w4084_,
		_w14689_
	);
	LUT2 #(
		.INIT('he)
	) name10642 (
		_w14688_,
		_w14689_,
		_w14690_
	);
	LUT3 #(
		.INIT('ha2)
	) name10643 (
		\emc_IOcst_reg/NET0131 ,
		_w4718_,
		_w9936_,
		_w14691_
	);
	LUT4 #(
		.INIT('he400)
	) name10644 (
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		\memc_IOcmd_E_reg/NET0131 ,
		_w14692_
	);
	LUT3 #(
		.INIT('he4)
	) name10645 (
		_w12057_,
		_w14691_,
		_w14692_,
		_w14693_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name10646 (
		\core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001 ,
		_w12216_,
		_w12219_,
		_w13091_,
		_w14694_
	);
	LUT4 #(
		.INIT('h0040)
	) name10647 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w14695_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name10648 (
		\sice_ICYC_en_reg/NET0131 ,
		\sice_SPC_reg[23]/P0001 ,
		_w14460_,
		_w14695_,
		_w14696_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name10649 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001 ,
		_w12216_,
		_w12219_,
		_w13168_,
		_w14697_
	);
	LUT4 #(
		.INIT('h8000)
	) name10650 (
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[1]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[2]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[3]/NET0131 ,
		_w14698_
	);
	LUT4 #(
		.INIT('h8000)
	) name10651 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		_w14698_,
		_w14699_
	);
	LUT4 #(
		.INIT('h8000)
	) name10652 (
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		_w14699_,
		_w14700_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10653 (
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		_w14699_,
		_w14701_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name10654 (
		\core_c_dec_updMF_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001 ,
		_w9453_,
		_w9894_,
		_w14702_
	);
	LUT4 #(
		.INIT('h4c08)
	) name10655 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w13091_,
		_w14409_,
		_w14561_,
		_w14703_
	);
	LUT2 #(
		.INIT('he)
	) name10656 (
		_w14702_,
		_w14703_,
		_w14704_
	);
	LUT2 #(
		.INIT('h2)
	) name10657 (
		\sport1_rxctl_a_sync1_reg/P0001 ,
		\sport1_rxctl_a_sync2_reg/P0001 ,
		_w14705_
	);
	LUT4 #(
		.INIT('h4044)
	) name10658 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTRX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w14706_
	);
	LUT4 #(
		.INIT('hfc55)
	) name10659 (
		\sport1_rxctl_RX_reg[9]/P0001 ,
		_w7140_,
		_w7240_,
		_w14706_,
		_w14707_
	);
	LUT3 #(
		.INIT('h8b)
	) name10660 (
		\sport1_rxctl_RXSHT_reg[9]/P0001 ,
		_w14705_,
		_w14707_,
		_w14708_
	);
	LUT4 #(
		.INIT('hfc55)
	) name10661 (
		\sport1_rxctl_RX_reg[8]/P0001 ,
		_w7465_,
		_w7565_,
		_w14706_,
		_w14709_
	);
	LUT3 #(
		.INIT('h8b)
	) name10662 (
		\sport1_rxctl_RXSHT_reg[8]/P0001 ,
		_w14705_,
		_w14709_,
		_w14710_
	);
	LUT2 #(
		.INIT('h2)
	) name10663 (
		\sport1_rxctl_RX_reg[7]/P0001 ,
		_w14706_,
		_w14711_
	);
	LUT4 #(
		.INIT('h4500)
	) name10664 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w14706_,
		_w14712_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10665 (
		\sport1_rxctl_RXSHT_reg[7]/P0001 ,
		_w14705_,
		_w14711_,
		_w14712_,
		_w14713_
	);
	LUT2 #(
		.INIT('h2)
	) name10666 (
		\sport1_rxctl_RX_reg[4]/P0001 ,
		_w14706_,
		_w14714_
	);
	LUT4 #(
		.INIT('h4500)
	) name10667 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w14706_,
		_w14715_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10668 (
		\sport1_rxctl_RXSHT_reg[4]/P0001 ,
		_w14705_,
		_w14714_,
		_w14715_,
		_w14716_
	);
	LUT2 #(
		.INIT('h2)
	) name10669 (
		\sport1_rxctl_RX_reg[6]/P0001 ,
		_w14706_,
		_w14717_
	);
	LUT4 #(
		.INIT('h4500)
	) name10670 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w14706_,
		_w14718_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10671 (
		\sport1_rxctl_RXSHT_reg[6]/P0001 ,
		_w14705_,
		_w14717_,
		_w14718_,
		_w14719_
	);
	LUT2 #(
		.INIT('h2)
	) name10672 (
		\sport1_rxctl_RX_reg[3]/P0001 ,
		_w14706_,
		_w14720_
	);
	LUT4 #(
		.INIT('h4500)
	) name10673 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w14706_,
		_w14721_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10674 (
		\sport1_rxctl_RXSHT_reg[3]/P0001 ,
		_w14705_,
		_w14720_,
		_w14721_,
		_w14722_
	);
	LUT2 #(
		.INIT('h2)
	) name10675 (
		\sport1_rxctl_RX_reg[5]/P0001 ,
		_w14706_,
		_w14723_
	);
	LUT4 #(
		.INIT('h4500)
	) name10676 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w14706_,
		_w14724_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10677 (
		\sport1_rxctl_RXSHT_reg[5]/P0001 ,
		_w14705_,
		_w14723_,
		_w14724_,
		_w14725_
	);
	LUT2 #(
		.INIT('h2)
	) name10678 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001 ,
		_w13168_,
		_w14726_
	);
	LUT4 #(
		.INIT('h4c08)
	) name10679 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w13168_,
		_w14409_,
		_w14561_,
		_w14727_
	);
	LUT2 #(
		.INIT('he)
	) name10680 (
		_w14726_,
		_w14727_,
		_w14728_
	);
	LUT2 #(
		.INIT('h2)
	) name10681 (
		\sport1_rxctl_RX_reg[2]/P0001 ,
		_w14706_,
		_w14729_
	);
	LUT4 #(
		.INIT('h4500)
	) name10682 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w14706_,
		_w14730_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10683 (
		\sport1_rxctl_RXSHT_reg[2]/P0001 ,
		_w14705_,
		_w14729_,
		_w14730_,
		_w14731_
	);
	LUT2 #(
		.INIT('h2)
	) name10684 (
		\sport1_rxctl_RX_reg[1]/P0001 ,
		_w14706_,
		_w14732_
	);
	LUT4 #(
		.INIT('h4500)
	) name10685 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w14706_,
		_w14733_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10686 (
		\sport1_rxctl_RXSHT_reg[1]/P0001 ,
		_w14705_,
		_w14732_,
		_w14733_,
		_w14734_
	);
	LUT4 #(
		.INIT('hfc55)
	) name10687 (
		\sport1_rxctl_RX_reg[15]/P0001 ,
		_w8798_,
		_w8801_,
		_w14706_,
		_w14735_
	);
	LUT3 #(
		.INIT('h8b)
	) name10688 (
		\sport1_rxctl_RXSHT_reg[15]/P0001 ,
		_w14705_,
		_w14735_,
		_w14736_
	);
	LUT4 #(
		.INIT('hfc55)
	) name10689 (
		\sport1_rxctl_RX_reg[14]/P0001 ,
		_w8757_,
		_w8760_,
		_w14706_,
		_w14737_
	);
	LUT3 #(
		.INIT('h8b)
	) name10690 (
		\sport1_rxctl_RXSHT_reg[14]/P0001 ,
		_w14705_,
		_w14737_,
		_w14738_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name10691 (
		\sport1_rxctl_RX_reg[13]/P0001 ,
		_w5760_,
		_w14705_,
		_w14706_,
		_w14739_
	);
	LUT3 #(
		.INIT('h08)
	) name10692 (
		\sport1_rxctl_RXSHT_reg[13]/P0001 ,
		\sport1_rxctl_a_sync1_reg/P0001 ,
		\sport1_rxctl_a_sync2_reg/P0001 ,
		_w14740_
	);
	LUT2 #(
		.INIT('he)
	) name10693 (
		_w14739_,
		_w14740_,
		_w14741_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name10694 (
		\sport1_rxctl_RX_reg[12]/P0001 ,
		_w6758_,
		_w14705_,
		_w14706_,
		_w14742_
	);
	LUT3 #(
		.INIT('h08)
	) name10695 (
		\sport1_rxctl_RXSHT_reg[12]/P0001 ,
		\sport1_rxctl_a_sync1_reg/P0001 ,
		\sport1_rxctl_a_sync2_reg/P0001 ,
		_w14743_
	);
	LUT2 #(
		.INIT('he)
	) name10696 (
		_w14742_,
		_w14743_,
		_w14744_
	);
	LUT4 #(
		.INIT('hfc55)
	) name10697 (
		\sport1_rxctl_RX_reg[11]/P0001 ,
		_w6263_,
		_w6362_,
		_w14706_,
		_w14745_
	);
	LUT3 #(
		.INIT('h8b)
	) name10698 (
		\sport1_rxctl_RXSHT_reg[11]/P0001 ,
		_w14705_,
		_w14745_,
		_w14746_
	);
	LUT4 #(
		.INIT('hfc55)
	) name10699 (
		\sport1_rxctl_RX_reg[10]/P0001 ,
		_w5937_,
		_w6038_,
		_w14706_,
		_w14747_
	);
	LUT3 #(
		.INIT('h8b)
	) name10700 (
		\sport1_rxctl_RXSHT_reg[10]/P0001 ,
		_w14705_,
		_w14747_,
		_w14748_
	);
	LUT2 #(
		.INIT('h2)
	) name10701 (
		\sport1_rxctl_RX_reg[0]/P0001 ,
		_w14706_,
		_w14749_
	);
	LUT4 #(
		.INIT('h4500)
	) name10702 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w14706_,
		_w14750_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10703 (
		\sport1_rxctl_RXSHT_reg[0]/P0001 ,
		_w14705_,
		_w14749_,
		_w14750_,
		_w14751_
	);
	LUT4 #(
		.INIT('haa8a)
	) name10704 (
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w14752_
	);
	LUT4 #(
		.INIT('h0051)
	) name10705 (
		\core_c_psq_Iflag_reg[10]/NET0131 ,
		\core_c_psq_T_PWRDN_reg/P0001 ,
		\core_c_psq_T_PWRDN_s1_reg/P0001 ,
		\sport0_regs_AUTO_a_reg[13]/NET0131 ,
		_w14753_
	);
	LUT2 #(
		.INIT('h1)
	) name10706 (
		_w14752_,
		_w14753_,
		_w14754_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10707 (
		\sice_ICYC_reg[7]/NET0131 ,
		\sice_ICYC_reg[8]/NET0131 ,
		\sice_ICYC_reg[9]/NET0131 ,
		_w11932_,
		_w14755_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10708 (
		\sice_IIRC_reg[4]/NET0131 ,
		\sice_IIRC_reg[5]/NET0131 ,
		\sice_IIRC_reg[6]/NET0131 ,
		_w11934_,
		_w14756_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10709 (
		\sice_IIRC_reg[7]/NET0131 ,
		\sice_IIRC_reg[8]/NET0131 ,
		\sice_IIRC_reg[9]/NET0131 ,
		_w11936_,
		_w14757_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10710 (
		\sice_ICYC_reg[4]/NET0131 ,
		\sice_ICYC_reg[5]/NET0131 ,
		\sice_ICYC_reg[6]/NET0131 ,
		_w11931_,
		_w14758_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10711 (
		\T_ED[7]_pad ,
		\emc_DMDreg_reg[7]/P0001 ,
		_w8594_,
		_w9940_,
		_w14759_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10712 (
		\T_ED[6]_pad ,
		\emc_DMDreg_reg[6]/P0001 ,
		_w8594_,
		_w9940_,
		_w14760_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10713 (
		\T_ED[5]_pad ,
		\emc_DMDreg_reg[5]/P0001 ,
		_w8594_,
		_w9940_,
		_w14761_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10714 (
		\T_ED[4]_pad ,
		\emc_DMDreg_reg[4]/P0001 ,
		_w8594_,
		_w9940_,
		_w14762_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10715 (
		\T_ED[3]_pad ,
		\emc_DMDreg_reg[3]/P0001 ,
		_w8594_,
		_w9940_,
		_w14763_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10716 (
		\T_ED[2]_pad ,
		\emc_DMDreg_reg[2]/P0001 ,
		_w8594_,
		_w9940_,
		_w14764_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10717 (
		\T_ED[1]_pad ,
		\emc_DMDreg_reg[1]/P0001 ,
		_w8594_,
		_w9940_,
		_w14765_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10718 (
		\T_ED[15]_pad ,
		\emc_DMDreg_reg[15]/P0001 ,
		_w8594_,
		_w9940_,
		_w14766_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10719 (
		\T_ED[14]_pad ,
		\emc_DMDreg_reg[14]/P0001 ,
		_w8594_,
		_w9940_,
		_w14767_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10720 (
		\T_ED[13]_pad ,
		\emc_DMDreg_reg[13]/P0001 ,
		_w8594_,
		_w9940_,
		_w14768_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10721 (
		\T_ED[12]_pad ,
		\emc_DMDreg_reg[12]/P0001 ,
		_w8594_,
		_w9940_,
		_w14769_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10722 (
		\T_ED[11]_pad ,
		\emc_DMDreg_reg[11]/P0001 ,
		_w8594_,
		_w9940_,
		_w14770_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10723 (
		\T_ED[10]_pad ,
		\emc_DMDreg_reg[10]/P0001 ,
		_w8594_,
		_w9940_,
		_w14771_
	);
	LUT4 #(
		.INIT('hcacc)
	) name10724 (
		\T_ED[0]_pad ,
		\emc_DMDreg_reg[0]/P0001 ,
		_w8594_,
		_w9940_,
		_w14772_
	);
	LUT4 #(
		.INIT('h0002)
	) name10725 (
		_w6884_,
		_w7331_,
		_w7692_,
		_w8008_,
		_w14773_
	);
	LUT3 #(
		.INIT('h80)
	) name10726 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_SHTop_E_reg/P0001 ,
		_w14774_
	);
	LUT2 #(
		.INIT('h8)
	) name10727 (
		_w9498_,
		_w14774_,
		_w14775_
	);
	LUT4 #(
		.INIT('h1000)
	) name10728 (
		_w5744_,
		_w5889_,
		_w6133_,
		_w6469_,
		_w14776_
	);
	LUT4 #(
		.INIT('h4000)
	) name10729 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_SHTop_E_reg/P0001 ,
		_w14777_
	);
	LUT2 #(
		.INIT('h1)
	) name10730 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w14777_,
		_w14778_
	);
	LUT4 #(
		.INIT('h7f00)
	) name10731 (
		_w14775_,
		_w14773_,
		_w14776_,
		_w14778_,
		_w14779_
	);
	LUT4 #(
		.INIT('h0004)
	) name10732 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9452_,
		_w9453_,
		_w14779_,
		_w14780_
	);
	LUT3 #(
		.INIT('h9f)
	) name10733 (
		_w11335_,
		_w11506_,
		_w14774_,
		_w14781_
	);
	LUT3 #(
		.INIT('h9f)
	) name10734 (
		_w11335_,
		_w11510_,
		_w14774_,
		_w14782_
	);
	LUT3 #(
		.INIT('h36)
	) name10735 (
		_w9550_,
		_w11335_,
		_w11486_,
		_w14783_
	);
	LUT3 #(
		.INIT('h98)
	) name10736 (
		_w11335_,
		_w11483_,
		_w14774_,
		_w14784_
	);
	LUT3 #(
		.INIT('h90)
	) name10737 (
		_w11335_,
		_w11483_,
		_w14774_,
		_w14785_
	);
	LUT4 #(
		.INIT('h2a22)
	) name10738 (
		_w14781_,
		_w14782_,
		_w14783_,
		_w14785_,
		_w14786_
	);
	LUT3 #(
		.INIT('h9f)
	) name10739 (
		_w11335_,
		_w11452_,
		_w14774_,
		_w14787_
	);
	LUT3 #(
		.INIT('h60)
	) name10740 (
		_w11335_,
		_w11448_,
		_w14774_,
		_w14788_
	);
	LUT3 #(
		.INIT('h60)
	) name10741 (
		_w11335_,
		_w11468_,
		_w14774_,
		_w14789_
	);
	LUT4 #(
		.INIT('h00f4)
	) name10742 (
		_w14786_,
		_w14787_,
		_w14788_,
		_w14789_,
		_w14790_
	);
	LUT3 #(
		.INIT('h9f)
	) name10743 (
		_w11335_,
		_w11464_,
		_w14774_,
		_w14791_
	);
	LUT3 #(
		.INIT('h9f)
	) name10744 (
		_w11335_,
		_w11514_,
		_w14774_,
		_w14792_
	);
	LUT3 #(
		.INIT('h9f)
	) name10745 (
		_w11335_,
		_w11457_,
		_w14774_,
		_w14793_
	);
	LUT4 #(
		.INIT('h4f00)
	) name10746 (
		_w14790_,
		_w14791_,
		_w14792_,
		_w14793_,
		_w14794_
	);
	LUT3 #(
		.INIT('h9f)
	) name10747 (
		_w11335_,
		_w11498_,
		_w14774_,
		_w14795_
	);
	LUT3 #(
		.INIT('h9f)
	) name10748 (
		_w11335_,
		_w11494_,
		_w14774_,
		_w14796_
	);
	LUT3 #(
		.INIT('h9f)
	) name10749 (
		_w11540_,
		_w11335_,
		_w14774_,
		_w14797_
	);
	LUT4 #(
		.INIT('h4f00)
	) name10750 (
		_w14794_,
		_w14795_,
		_w14796_,
		_w14797_,
		_w14798_
	);
	LUT3 #(
		.INIT('h9f)
	) name10751 (
		_w11536_,
		_w11335_,
		_w14774_,
		_w14799_
	);
	LUT3 #(
		.INIT('h9f)
	) name10752 (
		_w11335_,
		_w11528_,
		_w14774_,
		_w14800_
	);
	LUT3 #(
		.INIT('h20)
	) name10753 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w14801_
	);
	LUT2 #(
		.INIT('h8)
	) name10754 (
		_w14774_,
		_w14801_,
		_w14802_
	);
	LUT4 #(
		.INIT('h8400)
	) name10755 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w9498_,
		_w11335_,
		_w14774_,
		_w14803_
	);
	LUT2 #(
		.INIT('h1)
	) name10756 (
		_w14802_,
		_w14803_,
		_w14804_
	);
	LUT4 #(
		.INIT('h4f00)
	) name10757 (
		_w14798_,
		_w14799_,
		_w14800_,
		_w14804_,
		_w14805_
	);
	LUT4 #(
		.INIT('h7020)
	) name10758 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w12317_,
		_w14780_,
		_w14805_,
		_w14806_
	);
	LUT2 #(
		.INIT('h1)
	) name10759 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001 ,
		_w14780_,
		_w14807_
	);
	LUT2 #(
		.INIT('h1)
	) name10760 (
		_w14806_,
		_w14807_,
		_w14808_
	);
	LUT3 #(
		.INIT('h04)
	) name10761 (
		_w9453_,
		_w9894_,
		_w14779_,
		_w14809_
	);
	LUT4 #(
		.INIT('h7200)
	) name10762 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w12317_,
		_w14805_,
		_w14809_,
		_w14810_
	);
	LUT4 #(
		.INIT('h5545)
	) name10763 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001 ,
		_w9453_,
		_w9894_,
		_w14779_,
		_w14811_
	);
	LUT2 #(
		.INIT('h1)
	) name10764 (
		_w14810_,
		_w14811_,
		_w14812_
	);
	LUT4 #(
		.INIT('h1411)
	) name10765 (
		_w9455_,
		_w14580_,
		_w14581_,
		_w14582_,
		_w14813_
	);
	LUT3 #(
		.INIT('h82)
	) name10766 (
		_w9455_,
		_w9869_,
		_w9872_,
		_w14814_
	);
	LUT4 #(
		.INIT('h222e)
	) name10767 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001 ,
		_w9895_,
		_w14813_,
		_w14814_,
		_w14815_
	);
	LUT4 #(
		.INIT('h222e)
	) name10768 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001 ,
		_w9454_,
		_w14813_,
		_w14814_,
		_w14816_
	);
	LUT2 #(
		.INIT('hd)
	) name10769 (
		_w4140_,
		_w12803_,
		_w14817_
	);
	LUT2 #(
		.INIT('h2)
	) name10770 (
		_w8482_,
		_w14455_,
		_w14818_
	);
	LUT4 #(
		.INIT('h1000)
	) name10771 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14819_
	);
	LUT3 #(
		.INIT('h02)
	) name10772 (
		_w4102_,
		_w9933_,
		_w14819_,
		_w14820_
	);
	LUT4 #(
		.INIT('h0400)
	) name10773 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[9]/NET0131 ,
		_w14821_
	);
	LUT3 #(
		.INIT('h01)
	) name10774 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w14107_,
		_w14113_,
		_w14822_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10775 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w14107_,
		_w14113_,
		_w14823_
	);
	LUT4 #(
		.INIT('h0015)
	) name10776 (
		_w14103_,
		_w14108_,
		_w14114_,
		_w14823_,
		_w14824_
	);
	LUT4 #(
		.INIT('h2333)
	) name10777 (
		\tm_tpr_reg_DO_reg[9]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w14825_
	);
	LUT3 #(
		.INIT('hba)
	) name10778 (
		_w14821_,
		_w14824_,
		_w14825_,
		_w14826_
	);
	LUT4 #(
		.INIT('hb000)
	) name10779 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9437_,
		_w9438_,
		_w14827_
	);
	LUT2 #(
		.INIT('he)
	) name10780 (
		\core_c_psq_SSTAT_reg[3]/NET0131 ,
		_w14827_,
		_w14828_
	);
	LUT4 #(
		.INIT('h2000)
	) name10781 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14829_
	);
	LUT4 #(
		.INIT('h00bf)
	) name10782 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w4818_,
		_w12394_,
		_w14829_,
		_w14830_
	);
	LUT2 #(
		.INIT('h2)
	) name10783 (
		_w4102_,
		_w14830_,
		_w14831_
	);
	LUT4 #(
		.INIT('hb4f0)
	) name10784 (
		\bdma_BSreq_reg/NET0131 ,
		\bdma_BWcnt_reg[0]/NET0131 ,
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w4764_,
		_w14832_
	);
	LUT2 #(
		.INIT('h4)
	) name10785 (
		_w9413_,
		_w14832_,
		_w14833_
	);
	LUT3 #(
		.INIT('h10)
	) name10786 (
		_w4071_,
		_w4072_,
		_w5567_,
		_w14834_
	);
	LUT3 #(
		.INIT('h01)
	) name10787 (
		\clkc_SlowDn_reg/NET0131 ,
		\clkc_SlowDn_s1_reg/P0001 ,
		\clkc_SlowDn_s2_reg/P0001 ,
		_w14835_
	);
	LUT2 #(
		.INIT('h4)
	) name10788 (
		_w14453_,
		_w14835_,
		_w14836_
	);
	LUT4 #(
		.INIT('h4000)
	) name10789 (
		_w4094_,
		_w4097_,
		_w14834_,
		_w14836_,
		_w14837_
	);
	LUT4 #(
		.INIT('h2000)
	) name10790 (
		\core_c_dec_NOP_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14838_
	);
	LUT2 #(
		.INIT('h2)
	) name10791 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w14839_
	);
	LUT3 #(
		.INIT('h80)
	) name10792 (
		_w5028_,
		_w5045_,
		_w14839_,
		_w14840_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name10793 (
		_w4102_,
		_w4834_,
		_w14838_,
		_w14840_,
		_w14841_
	);
	LUT2 #(
		.INIT('h2)
	) name10794 (
		_w14591_,
		_w14594_,
		_w14842_
	);
	LUT2 #(
		.INIT('h8)
	) name10795 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w14843_
	);
	LUT4 #(
		.INIT('hfeaa)
	) name10796 (
		\sport1_rxctl_RSreq_reg/NET0131 ,
		_w14705_,
		_w14706_,
		_w14843_,
		_w14844_
	);
	LUT2 #(
		.INIT('h8)
	) name10797 (
		\emc_eRDY_reg/NET0131 ,
		_w4106_,
		_w14845_
	);
	LUT4 #(
		.INIT('h0400)
	) name10798 (
		\T_TMODE[1]_pad ,
		_w4776_,
		_w4773_,
		_w4780_,
		_w14846_
	);
	LUT3 #(
		.INIT('h40)
	) name10799 (
		_w4747_,
		_w4768_,
		_w14846_,
		_w14847_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name10800 (
		\T_TMODE[1]_pad ,
		_w4776_,
		_w4773_,
		_w4780_,
		_w14848_
	);
	LUT4 #(
		.INIT('hb000)
	) name10801 (
		_w4747_,
		_w4768_,
		_w4796_,
		_w14848_,
		_w14849_
	);
	LUT3 #(
		.INIT('h45)
	) name10802 (
		\emc_eRDY_reg/NET0131 ,
		_w4784_,
		_w4786_,
		_w14850_
	);
	LUT4 #(
		.INIT('hfeaa)
	) name10803 (
		_w14845_,
		_w14847_,
		_w14849_,
		_w14850_,
		_w14851_
	);
	LUT4 #(
		.INIT('h51fb)
	) name10804 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_a_sync1_reg/P0001 ,
		\sport0_rxctl_a_sync2_reg/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w14852_
	);
	LUT2 #(
		.INIT('h2)
	) name10805 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w14852_,
		_w14853_
	);
	LUT2 #(
		.INIT('h8)
	) name10806 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_txctl_b_sync1_reg/P0001 ,
		_w14854_
	);
	LUT2 #(
		.INIT('h2)
	) name10807 (
		_w14597_,
		_w14600_,
		_w14855_
	);
	LUT4 #(
		.INIT('h2000)
	) name10808 (
		\memc_LDaST_Eg_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w14856_
	);
	LUT3 #(
		.INIT('h8a)
	) name10809 (
		_w5056_,
		_w8175_,
		_w8179_,
		_w14857_
	);
	LUT3 #(
		.INIT('h8a)
	) name10810 (
		_w9061_,
		_w9322_,
		_w9324_,
		_w14858_
	);
	LUT2 #(
		.INIT('h1)
	) name10811 (
		_w14857_,
		_w14858_,
		_w14859_
	);
	LUT2 #(
		.INIT('h2)
	) name10812 (
		_w5570_,
		_w14859_,
		_w14860_
	);
	LUT4 #(
		.INIT('h1000)
	) name10813 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4428_,
		_w8172_,
		_w14860_,
		_w14861_
	);
	LUT2 #(
		.INIT('he)
	) name10814 (
		_w14856_,
		_w14861_,
		_w14862_
	);
	LUT3 #(
		.INIT('hac)
	) name10815 (
		\memc_selMIO_E_reg/P0001 ,
		_w8170_,
		_w14573_,
		_w14863_
	);
	LUT2 #(
		.INIT('h8)
	) name10816 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		_w9894_,
		_w14864_
	);
	LUT2 #(
		.INIT('h2)
	) name10817 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8694_,
		_w14865_
	);
	LUT4 #(
		.INIT('h00ab)
	) name10818 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6263_,
		_w6362_,
		_w14865_,
		_w14866_
	);
	LUT3 #(
		.INIT('he2)
	) name10819 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001 ,
		_w14864_,
		_w14866_,
		_w14867_
	);
	LUT3 #(
		.INIT('ha8)
	) name10820 (
		_w5107_,
		_w5937_,
		_w6038_,
		_w14868_
	);
	LUT4 #(
		.INIT('h00ef)
	) name10821 (
		_w5107_,
		_w5920_,
		_w5924_,
		_w14868_,
		_w14869_
	);
	LUT3 #(
		.INIT('hb8)
	) name10822 (
		\core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131 ,
		_w5074_,
		_w14869_,
		_w14870_
	);
	LUT2 #(
		.INIT('h8)
	) name10823 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		_w9894_,
		_w14871_
	);
	LUT3 #(
		.INIT('hca)
	) name10824 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001 ,
		_w13821_,
		_w14871_,
		_w14872_
	);
	LUT3 #(
		.INIT('h3a)
	) name10825 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001 ,
		_w13826_,
		_w14871_,
		_w14873_
	);
	LUT4 #(
		.INIT('h5300)
	) name10826 (
		_w5760_,
		_w8740_,
		_w13819_,
		_w14871_,
		_w14874_
	);
	LUT3 #(
		.INIT('h13)
	) name10827 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001 ,
		_w9894_,
		_w14875_
	);
	LUT2 #(
		.INIT('h1)
	) name10828 (
		_w14874_,
		_w14875_,
		_w14876_
	);
	LUT3 #(
		.INIT('h4c)
	) name10829 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001 ,
		_w9894_,
		_w14877_
	);
	LUT4 #(
		.INIT('hac00)
	) name10830 (
		_w6758_,
		_w8717_,
		_w13819_,
		_w14871_,
		_w14878_
	);
	LUT2 #(
		.INIT('he)
	) name10831 (
		_w14877_,
		_w14878_,
		_w14879_
	);
	LUT3 #(
		.INIT('h3a)
	) name10832 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001 ,
		_w13878_,
		_w14871_,
		_w14880_
	);
	LUT2 #(
		.INIT('h8)
	) name10833 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		_w11300_,
		_w14881_
	);
	LUT3 #(
		.INIT('hca)
	) name10834 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001 ,
		_w13821_,
		_w14881_,
		_w14882_
	);
	LUT4 #(
		.INIT('h5300)
	) name10835 (
		_w5760_,
		_w8740_,
		_w13819_,
		_w14881_,
		_w14883_
	);
	LUT3 #(
		.INIT('h13)
	) name10836 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001 ,
		_w11300_,
		_w14884_
	);
	LUT2 #(
		.INIT('h1)
	) name10837 (
		_w14883_,
		_w14884_,
		_w14885_
	);
	LUT3 #(
		.INIT('h4c)
	) name10838 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001 ,
		_w11300_,
		_w14886_
	);
	LUT4 #(
		.INIT('hac00)
	) name10839 (
		_w6758_,
		_w8717_,
		_w13819_,
		_w14881_,
		_w14887_
	);
	LUT2 #(
		.INIT('he)
	) name10840 (
		_w14886_,
		_w14887_,
		_w14888_
	);
	LUT3 #(
		.INIT('h3a)
	) name10841 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001 ,
		_w13878_,
		_w14881_,
		_w14889_
	);
	LUT3 #(
		.INIT('hca)
	) name10842 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001 ,
		_w13883_,
		_w14881_,
		_w14890_
	);
	LUT2 #(
		.INIT('h8)
	) name10843 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		_w9894_,
		_w14891_
	);
	LUT3 #(
		.INIT('hca)
	) name10844 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001 ,
		_w13821_,
		_w14891_,
		_w14892_
	);
	LUT3 #(
		.INIT('h3a)
	) name10845 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001 ,
		_w13826_,
		_w14891_,
		_w14893_
	);
	LUT3 #(
		.INIT('h4c)
	) name10846 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001 ,
		_w9894_,
		_w14894_
	);
	LUT4 #(
		.INIT('hac00)
	) name10847 (
		_w6758_,
		_w8717_,
		_w13819_,
		_w14891_,
		_w14895_
	);
	LUT2 #(
		.INIT('he)
	) name10848 (
		_w14894_,
		_w14895_,
		_w14896_
	);
	LUT3 #(
		.INIT('h3a)
	) name10849 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001 ,
		_w13878_,
		_w14891_,
		_w14897_
	);
	LUT3 #(
		.INIT('hca)
	) name10850 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001 ,
		_w13883_,
		_w14891_,
		_w14898_
	);
	LUT2 #(
		.INIT('h8)
	) name10851 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		_w11300_,
		_w14899_
	);
	LUT3 #(
		.INIT('hca)
	) name10852 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001 ,
		_w13821_,
		_w14899_,
		_w14900_
	);
	LUT3 #(
		.INIT('h3a)
	) name10853 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001 ,
		_w13826_,
		_w14899_,
		_w14901_
	);
	LUT3 #(
		.INIT('h4c)
	) name10854 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001 ,
		_w11300_,
		_w14902_
	);
	LUT4 #(
		.INIT('hac00)
	) name10855 (
		_w6758_,
		_w8717_,
		_w13819_,
		_w14899_,
		_w14903_
	);
	LUT2 #(
		.INIT('he)
	) name10856 (
		_w14902_,
		_w14903_,
		_w14904_
	);
	LUT3 #(
		.INIT('hca)
	) name10857 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001 ,
		_w13883_,
		_w14899_,
		_w14905_
	);
	LUT3 #(
		.INIT('h80)
	) name10858 (
		_w5658_,
		_w5804_,
		_w9431_,
		_w14906_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10859 (
		\bdma_BOVL_reg[9]/NET0131 ,
		_w7140_,
		_w7240_,
		_w14906_,
		_w14907_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10860 (
		\bdma_BOVL_reg[8]/NET0131 ,
		_w7465_,
		_w7565_,
		_w14906_,
		_w14908_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10861 (
		\bdma_BOVL_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w14906_,
		_w14909_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10862 (
		\bdma_BOVL_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w14906_,
		_w14910_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10863 (
		\bdma_BCTL_reg[9]/NET0131 ,
		_w7140_,
		_w7240_,
		_w13346_,
		_w14911_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10864 (
		\bdma_BCTL_reg[8]/NET0131 ,
		_w7465_,
		_w7565_,
		_w13346_,
		_w14912_
	);
	LUT3 #(
		.INIT('hca)
	) name10865 (
		\bdma_BCTL_reg[13]/NET0131 ,
		_w5760_,
		_w13346_,
		_w14913_
	);
	LUT3 #(
		.INIT('hca)
	) name10866 (
		\bdma_BCTL_reg[12]/NET0131 ,
		_w6758_,
		_w13346_,
		_w14914_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10867 (
		\bdma_BCTL_reg[11]/NET0131 ,
		_w6263_,
		_w6362_,
		_w13346_,
		_w14915_
	);
	LUT4 #(
		.INIT('h03aa)
	) name10868 (
		\bdma_BCTL_reg[10]/NET0131 ,
		_w5937_,
		_w6038_,
		_w13346_,
		_w14916_
	);
	LUT2 #(
		.INIT('h2)
	) name10869 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8998_,
		_w14917_
	);
	LUT4 #(
		.INIT('h00ab)
	) name10870 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w7465_,
		_w7565_,
		_w14917_,
		_w14918_
	);
	LUT3 #(
		.INIT('he2)
	) name10871 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001 ,
		_w14864_,
		_w14918_,
		_w14919_
	);
	LUT4 #(
		.INIT('h4044)
	) name10872 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTTX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w14920_
	);
	LUT2 #(
		.INIT('h1)
	) name10873 (
		\auctl_T1Sack_reg/NET0131 ,
		_w14920_,
		_w14921_
	);
	LUT4 #(
		.INIT('haa03)
	) name10874 (
		\sport1_txctl_TX_reg[9]/P0001 ,
		_w7140_,
		_w7240_,
		_w14921_,
		_w14922_
	);
	LUT4 #(
		.INIT('haa03)
	) name10875 (
		\sport1_txctl_TX_reg[8]/P0001 ,
		_w7465_,
		_w7565_,
		_w14921_,
		_w14923_
	);
	LUT3 #(
		.INIT('hac)
	) name10876 (
		\sport1_txctl_TX_reg[12]/P0001 ,
		_w6758_,
		_w14921_,
		_w14924_
	);
	LUT4 #(
		.INIT('haa03)
	) name10877 (
		\sport1_txctl_TX_reg[11]/P0001 ,
		_w6263_,
		_w6362_,
		_w14921_,
		_w14925_
	);
	LUT4 #(
		.INIT('haa03)
	) name10878 (
		\sport1_txctl_TX_reg[10]/P0001 ,
		_w5937_,
		_w6038_,
		_w14921_,
		_w14926_
	);
	LUT3 #(
		.INIT('h3a)
	) name10879 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001 ,
		_w13826_,
		_w14881_,
		_w14927_
	);
	LUT4 #(
		.INIT('h8a88)
	) name10880 (
		_w5107_,
		_w6054_,
		_w6173_,
		_w6175_,
		_w14928_
	);
	LUT4 #(
		.INIT('h00ef)
	) name10881 (
		_w5107_,
		_w6204_,
		_w6207_,
		_w14928_,
		_w14929_
	);
	LUT3 #(
		.INIT('hb8)
	) name10882 (
		\core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 ,
		_w5074_,
		_w14929_,
		_w14930_
	);
	LUT2 #(
		.INIT('h8)
	) name10883 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		_w9894_,
		_w14931_
	);
	LUT3 #(
		.INIT('hca)
	) name10884 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001 ,
		_w13821_,
		_w14931_,
		_w14932_
	);
	LUT3 #(
		.INIT('h3a)
	) name10885 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001 ,
		_w13826_,
		_w14931_,
		_w14933_
	);
	LUT4 #(
		.INIT('h5300)
	) name10886 (
		_w5760_,
		_w8740_,
		_w13819_,
		_w14931_,
		_w14934_
	);
	LUT3 #(
		.INIT('h13)
	) name10887 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001 ,
		_w9894_,
		_w14935_
	);
	LUT2 #(
		.INIT('h1)
	) name10888 (
		_w14934_,
		_w14935_,
		_w14936_
	);
	LUT3 #(
		.INIT('h4c)
	) name10889 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001 ,
		_w9894_,
		_w14937_
	);
	LUT4 #(
		.INIT('hac00)
	) name10890 (
		_w6758_,
		_w8717_,
		_w13819_,
		_w14931_,
		_w14938_
	);
	LUT2 #(
		.INIT('he)
	) name10891 (
		_w14937_,
		_w14938_,
		_w14939_
	);
	LUT3 #(
		.INIT('h3a)
	) name10892 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001 ,
		_w13878_,
		_w14931_,
		_w14940_
	);
	LUT3 #(
		.INIT('hca)
	) name10893 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001 ,
		_w13883_,
		_w14931_,
		_w14941_
	);
	LUT2 #(
		.INIT('h8)
	) name10894 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		_w9894_,
		_w14942_
	);
	LUT3 #(
		.INIT('hca)
	) name10895 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001 ,
		_w12284_,
		_w14942_,
		_w14943_
	);
	LUT3 #(
		.INIT('hca)
	) name10896 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001 ,
		_w14918_,
		_w14942_,
		_w14944_
	);
	LUT4 #(
		.INIT('h1b00)
	) name10897 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w14942_,
		_w14945_
	);
	LUT3 #(
		.INIT('h13)
	) name10898 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001 ,
		_w9894_,
		_w14946_
	);
	LUT2 #(
		.INIT('h1)
	) name10899 (
		_w14945_,
		_w14946_,
		_w14947_
	);
	LUT2 #(
		.INIT('h2)
	) name10900 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8717_,
		_w14948_
	);
	LUT3 #(
		.INIT('h0e)
	) name10901 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w14948_,
		_w14949_
	);
	LUT4 #(
		.INIT('h1b00)
	) name10902 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w14942_,
		_w14950_
	);
	LUT3 #(
		.INIT('h13)
	) name10903 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001 ,
		_w9894_,
		_w14951_
	);
	LUT2 #(
		.INIT('h1)
	) name10904 (
		_w14950_,
		_w14951_,
		_w14952_
	);
	LUT3 #(
		.INIT('hca)
	) name10905 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001 ,
		_w14866_,
		_w14942_,
		_w14953_
	);
	LUT3 #(
		.INIT('hca)
	) name10906 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001 ,
		_w12486_,
		_w14942_,
		_w14954_
	);
	LUT2 #(
		.INIT('h8)
	) name10907 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		_w9894_,
		_w14955_
	);
	LUT3 #(
		.INIT('hca)
	) name10908 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001 ,
		_w12284_,
		_w14955_,
		_w14956_
	);
	LUT3 #(
		.INIT('hca)
	) name10909 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001 ,
		_w14918_,
		_w14955_,
		_w14957_
	);
	LUT4 #(
		.INIT('h1b00)
	) name10910 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w14955_,
		_w14958_
	);
	LUT3 #(
		.INIT('h13)
	) name10911 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001 ,
		_w9894_,
		_w14959_
	);
	LUT2 #(
		.INIT('h1)
	) name10912 (
		_w14958_,
		_w14959_,
		_w14960_
	);
	LUT4 #(
		.INIT('h1b00)
	) name10913 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w14955_,
		_w14961_
	);
	LUT3 #(
		.INIT('h13)
	) name10914 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001 ,
		_w9894_,
		_w14962_
	);
	LUT2 #(
		.INIT('h1)
	) name10915 (
		_w14961_,
		_w14962_,
		_w14963_
	);
	LUT3 #(
		.INIT('hca)
	) name10916 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001 ,
		_w14866_,
		_w14955_,
		_w14964_
	);
	LUT3 #(
		.INIT('hca)
	) name10917 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001 ,
		_w12486_,
		_w14955_,
		_w14965_
	);
	LUT3 #(
		.INIT('h3a)
	) name10918 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001 ,
		_w13878_,
		_w14899_,
		_w14966_
	);
	LUT4 #(
		.INIT('h5300)
	) name10919 (
		_w5760_,
		_w8740_,
		_w13819_,
		_w14899_,
		_w14967_
	);
	LUT3 #(
		.INIT('h13)
	) name10920 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001 ,
		_w11300_,
		_w14968_
	);
	LUT2 #(
		.INIT('h1)
	) name10921 (
		_w14967_,
		_w14968_,
		_w14969_
	);
	LUT2 #(
		.INIT('h4)
	) name10922 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTIreg_E_reg[7]/P0001 ,
		_w14970_
	);
	LUT4 #(
		.INIT('h00df)
	) name10923 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w5005_,
		_w14970_,
		_w14971_
	);
	LUT2 #(
		.INIT('h4)
	) name10924 (
		_w5002_,
		_w14971_,
		_w14972_
	);
	LUT3 #(
		.INIT('h0e)
	) name10925 (
		_w5004_,
		_w5006_,
		_w14972_,
		_w14973_
	);
	LUT4 #(
		.INIT('haa02)
	) name10926 (
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w14974_
	);
	LUT3 #(
		.INIT('hf4)
	) name10927 (
		_w5007_,
		_w13022_,
		_w14974_,
		_w14975_
	);
	LUT4 #(
		.INIT('haa02)
	) name10928 (
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w14976_
	);
	LUT3 #(
		.INIT('hf4)
	) name10929 (
		_w5007_,
		_w12931_,
		_w14976_,
		_w14977_
	);
	LUT4 #(
		.INIT('haa02)
	) name10930 (
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w14978_
	);
	LUT3 #(
		.INIT('hf4)
	) name10931 (
		_w5007_,
		_w12939_,
		_w14978_,
		_w14979_
	);
	LUT4 #(
		.INIT('haa02)
	) name10932 (
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w14980_
	);
	LUT4 #(
		.INIT('hff54)
	) name10933 (
		_w5007_,
		_w12976_,
		_w12977_,
		_w14980_,
		_w14981_
	);
	LUT4 #(
		.INIT('haa02)
	) name10934 (
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w14982_
	);
	LUT3 #(
		.INIT('hf1)
	) name10935 (
		_w5007_,
		_w12984_,
		_w14982_,
		_w14983_
	);
	LUT3 #(
		.INIT('hb8)
	) name10936 (
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		_w5015_,
		_w13022_,
		_w14984_
	);
	LUT3 #(
		.INIT('hb8)
	) name10937 (
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		_w5015_,
		_w12913_,
		_w14985_
	);
	LUT3 #(
		.INIT('hb8)
	) name10938 (
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		_w5015_,
		_w12923_,
		_w14986_
	);
	LUT3 #(
		.INIT('hb8)
	) name10939 (
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w5015_,
		_w12931_,
		_w14987_
	);
	LUT3 #(
		.INIT('hb8)
	) name10940 (
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w5015_,
		_w12939_,
		_w14988_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10941 (
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		_w5015_,
		_w12976_,
		_w12977_,
		_w14989_
	);
	LUT3 #(
		.INIT('h8b)
	) name10942 (
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		_w5015_,
		_w12984_,
		_w14990_
	);
	LUT3 #(
		.INIT('h8b)
	) name10943 (
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		_w5015_,
		_w12991_,
		_w14991_
	);
	LUT3 #(
		.INIT('hb8)
	) name10944 (
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		_w5015_,
		_w13000_,
		_w14992_
	);
	LUT2 #(
		.INIT('h4)
	) name10945 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTIreg_E_reg[5]/P0001 ,
		_w14993_
	);
	LUT4 #(
		.INIT('h00ef)
	) name10946 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w5005_,
		_w14993_,
		_w14994_
	);
	LUT2 #(
		.INIT('h4)
	) name10947 (
		_w5018_,
		_w14994_,
		_w14995_
	);
	LUT3 #(
		.INIT('h0e)
	) name10948 (
		_w5020_,
		_w5021_,
		_w14995_,
		_w14996_
	);
	LUT4 #(
		.INIT('haa02)
	) name10949 (
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w14997_
	);
	LUT3 #(
		.INIT('hf4)
	) name10950 (
		_w5022_,
		_w13022_,
		_w14997_,
		_w14998_
	);
	LUT4 #(
		.INIT('haa02)
	) name10951 (
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w14999_
	);
	LUT3 #(
		.INIT('hf4)
	) name10952 (
		_w5022_,
		_w12931_,
		_w14999_,
		_w15000_
	);
	LUT4 #(
		.INIT('haa02)
	) name10953 (
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w15001_
	);
	LUT3 #(
		.INIT('hf4)
	) name10954 (
		_w5022_,
		_w12939_,
		_w15001_,
		_w15002_
	);
	LUT4 #(
		.INIT('haa02)
	) name10955 (
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w15003_
	);
	LUT4 #(
		.INIT('hff54)
	) name10956 (
		_w5022_,
		_w12976_,
		_w12977_,
		_w15003_,
		_w15004_
	);
	LUT4 #(
		.INIT('haa02)
	) name10957 (
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w15005_
	);
	LUT3 #(
		.INIT('hf1)
	) name10958 (
		_w5022_,
		_w12984_,
		_w15005_,
		_w15006_
	);
	LUT2 #(
		.INIT('h4)
	) name10959 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTIreg_E_reg[4]/P0001 ,
		_w15007_
	);
	LUT4 #(
		.INIT('h00ef)
	) name10960 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4973_,
		_w4977_,
		_w15007_,
		_w15008_
	);
	LUT2 #(
		.INIT('h4)
	) name10961 (
		_w4974_,
		_w15008_,
		_w15009_
	);
	LUT3 #(
		.INIT('h0e)
	) name10962 (
		_w4976_,
		_w4978_,
		_w15009_,
		_w15010_
	);
	LUT4 #(
		.INIT('haa02)
	) name10963 (
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15011_
	);
	LUT3 #(
		.INIT('hf4)
	) name10964 (
		_w4979_,
		_w13022_,
		_w15011_,
		_w15012_
	);
	LUT3 #(
		.INIT('hca)
	) name10965 (
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		_w12913_,
		_w15010_,
		_w15013_
	);
	LUT3 #(
		.INIT('hca)
	) name10966 (
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		_w12923_,
		_w15010_,
		_w15014_
	);
	LUT4 #(
		.INIT('haa02)
	) name10967 (
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15015_
	);
	LUT3 #(
		.INIT('hf4)
	) name10968 (
		_w4979_,
		_w12931_,
		_w15015_,
		_w15016_
	);
	LUT4 #(
		.INIT('haa02)
	) name10969 (
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15017_
	);
	LUT3 #(
		.INIT('hf4)
	) name10970 (
		_w4979_,
		_w12939_,
		_w15017_,
		_w15018_
	);
	LUT4 #(
		.INIT('haa02)
	) name10971 (
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15019_
	);
	LUT4 #(
		.INIT('hff54)
	) name10972 (
		_w4979_,
		_w12976_,
		_w12977_,
		_w15019_,
		_w15020_
	);
	LUT4 #(
		.INIT('haa02)
	) name10973 (
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15021_
	);
	LUT3 #(
		.INIT('hf1)
	) name10974 (
		_w4979_,
		_w12984_,
		_w15021_,
		_w15022_
	);
	LUT3 #(
		.INIT('h3a)
	) name10975 (
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		_w12991_,
		_w15010_,
		_w15023_
	);
	LUT3 #(
		.INIT('hca)
	) name10976 (
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		_w13000_,
		_w15010_,
		_w15024_
	);
	LUT3 #(
		.INIT('hca)
	) name10977 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001 ,
		_w12284_,
		_w14864_,
		_w15025_
	);
	LUT4 #(
		.INIT('h1b00)
	) name10978 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w14864_,
		_w15026_
	);
	LUT3 #(
		.INIT('h13)
	) name10979 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001 ,
		_w9894_,
		_w15027_
	);
	LUT2 #(
		.INIT('h1)
	) name10980 (
		_w15026_,
		_w15027_,
		_w15028_
	);
	LUT4 #(
		.INIT('h5300)
	) name10981 (
		_w5760_,
		_w8740_,
		_w13819_,
		_w14891_,
		_w15029_
	);
	LUT3 #(
		.INIT('h13)
	) name10982 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001 ,
		_w9894_,
		_w15030_
	);
	LUT2 #(
		.INIT('h1)
	) name10983 (
		_w15029_,
		_w15030_,
		_w15031_
	);
	LUT4 #(
		.INIT('h4501)
	) name10984 (
		_w5091_,
		_w5107_,
		_w7400_,
		_w7566_,
		_w15032_
	);
	LUT3 #(
		.INIT('h02)
	) name10985 (
		\core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 ,
		_w5087_,
		_w5090_,
		_w15033_
	);
	LUT2 #(
		.INIT('he)
	) name10986 (
		_w15032_,
		_w15033_,
		_w15034_
	);
	LUT4 #(
		.INIT('h1054)
	) name10987 (
		_w5091_,
		_w5107_,
		_w7579_,
		_w7710_,
		_w15035_
	);
	LUT3 #(
		.INIT('h01)
	) name10988 (
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w5087_,
		_w5090_,
		_w15036_
	);
	LUT2 #(
		.INIT('h1)
	) name10989 (
		_w15035_,
		_w15036_,
		_w15037_
	);
	LUT4 #(
		.INIT('h1054)
	) name10990 (
		_w5091_,
		_w5107_,
		_w6591_,
		_w6897_,
		_w15038_
	);
	LUT3 #(
		.INIT('h01)
	) name10991 (
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w5087_,
		_w5090_,
		_w15039_
	);
	LUT2 #(
		.INIT('h1)
	) name10992 (
		_w15038_,
		_w15039_,
		_w15040_
	);
	LUT2 #(
		.INIT('h2)
	) name10993 (
		_w5107_,
		_w5760_,
		_w15041_
	);
	LUT4 #(
		.INIT('h00ef)
	) name10994 (
		_w5107_,
		_w5312_,
		_w5315_,
		_w15041_,
		_w15042_
	);
	LUT3 #(
		.INIT('hb8)
	) name10995 (
		\core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 ,
		_w5091_,
		_w15042_,
		_w15043_
	);
	LUT2 #(
		.INIT('h8)
	) name10996 (
		_w5107_,
		_w6758_,
		_w15044_
	);
	LUT4 #(
		.INIT('h00ba)
	) name10997 (
		_w5107_,
		_w6643_,
		_w6646_,
		_w15044_,
		_w15045_
	);
	LUT3 #(
		.INIT('h8b)
	) name10998 (
		\core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 ,
		_w5091_,
		_w15045_,
		_w15046_
	);
	LUT3 #(
		.INIT('h02)
	) name10999 (
		_w5107_,
		_w6263_,
		_w6362_,
		_w15047_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11000 (
		_w5107_,
		_w6245_,
		_w6250_,
		_w15047_,
		_w15048_
	);
	LUT3 #(
		.INIT('h8b)
	) name11001 (
		\core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 ,
		_w5091_,
		_w15048_,
		_w15049_
	);
	LUT3 #(
		.INIT('hb8)
	) name11002 (
		\core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 ,
		_w5091_,
		_w14869_,
		_w15050_
	);
	LUT3 #(
		.INIT('h02)
	) name11003 (
		_w5107_,
		_w7140_,
		_w7240_,
		_w15051_
	);
	LUT4 #(
		.INIT('h00ab)
	) name11004 (
		_w5107_,
		_w7062_,
		_w7067_,
		_w15051_,
		_w15052_
	);
	LUT4 #(
		.INIT('hff54)
	) name11005 (
		_w5107_,
		_w7062_,
		_w7067_,
		_w15051_,
		_w15053_
	);
	LUT3 #(
		.INIT('h8b)
	) name11006 (
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		_w5074_,
		_w15052_,
		_w15054_
	);
	LUT4 #(
		.INIT('h4501)
	) name11007 (
		_w5074_,
		_w5107_,
		_w7400_,
		_w7566_,
		_w15055_
	);
	LUT2 #(
		.INIT('he)
	) name11008 (
		_w7437_,
		_w15055_,
		_w15056_
	);
	LUT4 #(
		.INIT('h2022)
	) name11009 (
		_w5107_,
		_w7793_,
		_w7903_,
		_w7905_,
		_w15057_
	);
	LUT3 #(
		.INIT('hf1)
	) name11010 (
		_w5107_,
		_w7731_,
		_w15057_,
		_w15058_
	);
	LUT4 #(
		.INIT('h4501)
	) name11011 (
		_w5074_,
		_w5107_,
		_w7731_,
		_w7906_,
		_w15059_
	);
	LUT2 #(
		.INIT('he)
	) name11012 (
		_w7766_,
		_w15059_,
		_w15060_
	);
	LUT4 #(
		.INIT('h2022)
	) name11013 (
		_w5107_,
		_w7927_,
		_w8040_,
		_w8042_,
		_w15061_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11014 (
		_w5107_,
		_w7911_,
		_w7914_,
		_w15061_,
		_w15062_
	);
	LUT4 #(
		.INIT('hff45)
	) name11015 (
		_w5107_,
		_w7911_,
		_w7914_,
		_w15061_,
		_w15063_
	);
	LUT3 #(
		.INIT('h8b)
	) name11016 (
		\core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 ,
		_w5074_,
		_w15062_,
		_w15064_
	);
	LUT4 #(
		.INIT('h4501)
	) name11017 (
		_w5074_,
		_w5107_,
		_w7579_,
		_w7710_,
		_w15065_
	);
	LUT2 #(
		.INIT('he)
	) name11018 (
		_w7406_,
		_w15065_,
		_w15066_
	);
	LUT4 #(
		.INIT('h2022)
	) name11019 (
		_w5107_,
		_w7257_,
		_w7375_,
		_w7377_,
		_w15067_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11020 (
		_w5107_,
		_w7122_,
		_w7126_,
		_w15067_,
		_w15068_
	);
	LUT4 #(
		.INIT('hff45)
	) name11021 (
		_w5107_,
		_w7122_,
		_w7126_,
		_w15067_,
		_w15069_
	);
	LUT3 #(
		.INIT('h8b)
	) name11022 (
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w5074_,
		_w15068_,
		_w15070_
	);
	LUT4 #(
		.INIT('h2022)
	) name11023 (
		_w5107_,
		_w6378_,
		_w6498_,
		_w6500_,
		_w15071_
	);
	LUT3 #(
		.INIT('hf1)
	) name11024 (
		_w5107_,
		_w6555_,
		_w15071_,
		_w15072_
	);
	LUT4 #(
		.INIT('h4051)
	) name11025 (
		_w5074_,
		_w5107_,
		_w6501_,
		_w6555_,
		_w15073_
	);
	LUT2 #(
		.INIT('he)
	) name11026 (
		_w6561_,
		_w15073_,
		_w15074_
	);
	LUT4 #(
		.INIT('h1054)
	) name11027 (
		_w5074_,
		_w5107_,
		_w6591_,
		_w6897_,
		_w15075_
	);
	LUT3 #(
		.INIT('h01)
	) name11028 (
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w5070_,
		_w5073_,
		_w15076_
	);
	LUT2 #(
		.INIT('h1)
	) name11029 (
		_w15075_,
		_w15076_,
		_w15077_
	);
	LUT3 #(
		.INIT('hb8)
	) name11030 (
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		_w5074_,
		_w15042_,
		_w15078_
	);
	LUT3 #(
		.INIT('h8b)
	) name11031 (
		\core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 ,
		_w5074_,
		_w15045_,
		_w15079_
	);
	LUT3 #(
		.INIT('h8b)
	) name11032 (
		\core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131 ,
		_w5074_,
		_w15048_,
		_w15080_
	);
	LUT3 #(
		.INIT('hac)
	) name11033 (
		\sport1_txctl_TX_reg[13]/P0001 ,
		_w5760_,
		_w14921_,
		_w15081_
	);
	LUT4 #(
		.INIT('h2022)
	) name11034 (
		_w5107_,
		_w5784_,
		_w5911_,
		_w5913_,
		_w15082_
	);
	LUT3 #(
		.INIT('hf1)
	) name11035 (
		_w5107_,
		_w5771_,
		_w15082_,
		_w15083_
	);
	LUT4 #(
		.INIT('h4051)
	) name11036 (
		_w5074_,
		_w5107_,
		_w5914_,
		_w5771_,
		_w15084_
	);
	LUT3 #(
		.INIT('h02)
	) name11037 (
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w5070_,
		_w5073_,
		_w15085_
	);
	LUT2 #(
		.INIT('he)
	) name11038 (
		_w15084_,
		_w15085_,
		_w15086_
	);
	LUT4 #(
		.INIT('h4501)
	) name11039 (
		_w5083_,
		_w5107_,
		_w7400_,
		_w7566_,
		_w15087_
	);
	LUT2 #(
		.INIT('he)
	) name11040 (
		_w7439_,
		_w15087_,
		_w15088_
	);
	LUT3 #(
		.INIT('h02)
	) name11041 (
		\core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 ,
		_w5079_,
		_w5082_,
		_w15089_
	);
	LUT4 #(
		.INIT('h4501)
	) name11042 (
		_w5083_,
		_w5107_,
		_w7579_,
		_w7710_,
		_w15090_
	);
	LUT2 #(
		.INIT('he)
	) name11043 (
		_w15089_,
		_w15090_,
		_w15091_
	);
	LUT4 #(
		.INIT('h4501)
	) name11044 (
		_w5083_,
		_w5107_,
		_w6591_,
		_w6897_,
		_w15092_
	);
	LUT2 #(
		.INIT('he)
	) name11045 (
		_w6627_,
		_w15092_,
		_w15093_
	);
	LUT3 #(
		.INIT('hb8)
	) name11046 (
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		_w5083_,
		_w15042_,
		_w15094_
	);
	LUT3 #(
		.INIT('h8b)
	) name11047 (
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		_w5083_,
		_w15045_,
		_w15095_
	);
	LUT3 #(
		.INIT('h8b)
	) name11048 (
		\core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 ,
		_w5083_,
		_w15048_,
		_w15096_
	);
	LUT3 #(
		.INIT('hb8)
	) name11049 (
		\core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 ,
		_w5083_,
		_w14869_,
		_w15097_
	);
	LUT3 #(
		.INIT('h8b)
	) name11050 (
		\core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 ,
		_w5066_,
		_w15052_,
		_w15098_
	);
	LUT3 #(
		.INIT('h02)
	) name11051 (
		\core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 ,
		_w5061_,
		_w5065_,
		_w15099_
	);
	LUT4 #(
		.INIT('h4501)
	) name11052 (
		_w5066_,
		_w5107_,
		_w7400_,
		_w7566_,
		_w15100_
	);
	LUT2 #(
		.INIT('he)
	) name11053 (
		_w15099_,
		_w15100_,
		_w15101_
	);
	LUT4 #(
		.INIT('h4501)
	) name11054 (
		_w5066_,
		_w5107_,
		_w7731_,
		_w7906_,
		_w15102_
	);
	LUT3 #(
		.INIT('h02)
	) name11055 (
		\core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 ,
		_w5061_,
		_w5065_,
		_w15103_
	);
	LUT2 #(
		.INIT('he)
	) name11056 (
		_w15102_,
		_w15103_,
		_w15104_
	);
	LUT3 #(
		.INIT('h8b)
	) name11057 (
		\core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 ,
		_w5066_,
		_w15062_,
		_w15105_
	);
	LUT4 #(
		.INIT('h4501)
	) name11058 (
		_w5066_,
		_w5107_,
		_w7579_,
		_w7710_,
		_w15106_
	);
	LUT2 #(
		.INIT('he)
	) name11059 (
		_w7404_,
		_w15106_,
		_w15107_
	);
	LUT3 #(
		.INIT('h8b)
	) name11060 (
		\core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 ,
		_w5066_,
		_w15068_,
		_w15108_
	);
	LUT3 #(
		.INIT('hb8)
	) name11061 (
		\core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 ,
		_w5066_,
		_w14929_,
		_w15109_
	);
	LUT4 #(
		.INIT('h4051)
	) name11062 (
		_w5066_,
		_w5107_,
		_w6501_,
		_w6555_,
		_w15110_
	);
	LUT3 #(
		.INIT('h02)
	) name11063 (
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		_w5061_,
		_w5065_,
		_w15111_
	);
	LUT2 #(
		.INIT('he)
	) name11064 (
		_w15110_,
		_w15111_,
		_w15112_
	);
	LUT4 #(
		.INIT('h4501)
	) name11065 (
		_w5066_,
		_w5107_,
		_w6591_,
		_w6897_,
		_w15113_
	);
	LUT2 #(
		.INIT('he)
	) name11066 (
		_w6629_,
		_w15113_,
		_w15114_
	);
	LUT3 #(
		.INIT('hb8)
	) name11067 (
		\core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 ,
		_w5066_,
		_w15042_,
		_w15115_
	);
	LUT3 #(
		.INIT('h8b)
	) name11068 (
		\core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 ,
		_w5066_,
		_w15045_,
		_w15116_
	);
	LUT3 #(
		.INIT('h8b)
	) name11069 (
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		_w5066_,
		_w15048_,
		_w15117_
	);
	LUT3 #(
		.INIT('hb8)
	) name11070 (
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		_w5066_,
		_w14869_,
		_w15118_
	);
	LUT4 #(
		.INIT('h4051)
	) name11071 (
		_w5066_,
		_w5107_,
		_w5914_,
		_w5771_,
		_w15119_
	);
	LUT2 #(
		.INIT('he)
	) name11072 (
		_w5552_,
		_w15119_,
		_w15120_
	);
	LUT3 #(
		.INIT('hca)
	) name11073 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001 ,
		_w13883_,
		_w14871_,
		_w15121_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11074 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w14864_,
		_w15122_
	);
	LUT3 #(
		.INIT('h13)
	) name11075 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001 ,
		_w9894_,
		_w15123_
	);
	LUT2 #(
		.INIT('h1)
	) name11076 (
		_w15122_,
		_w15123_,
		_w15124_
	);
	LUT3 #(
		.INIT('hca)
	) name11077 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001 ,
		_w12486_,
		_w14864_,
		_w15125_
	);
	LUT4 #(
		.INIT('haa02)
	) name11078 (
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w15126_
	);
	LUT3 #(
		.INIT('hf4)
	) name11079 (
		_w5007_,
		_w12947_,
		_w15126_,
		_w15127_
	);
	LUT4 #(
		.INIT('haa02)
	) name11080 (
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w15128_
	);
	LUT3 #(
		.INIT('hf4)
	) name11081 (
		_w5007_,
		_w9156_,
		_w15128_,
		_w15129_
	);
	LUT4 #(
		.INIT('haa02)
	) name11082 (
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w15130_
	);
	LUT3 #(
		.INIT('hf1)
	) name11083 (
		_w5007_,
		_w12961_,
		_w15130_,
		_w15131_
	);
	LUT4 #(
		.INIT('haa02)
	) name11084 (
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w15132_
	);
	LUT3 #(
		.INIT('hf1)
	) name11085 (
		_w5007_,
		_w12969_,
		_w15132_,
		_w15133_
	);
	LUT4 #(
		.INIT('haa02)
	) name11086 (
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w5004_,
		_w5006_,
		_w14972_,
		_w15134_
	);
	LUT3 #(
		.INIT('hf1)
	) name11087 (
		_w5007_,
		_w13008_,
		_w15134_,
		_w15135_
	);
	LUT3 #(
		.INIT('hb8)
	) name11088 (
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w5015_,
		_w12947_,
		_w15136_
	);
	LUT3 #(
		.INIT('hb8)
	) name11089 (
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w5015_,
		_w9156_,
		_w15137_
	);
	LUT3 #(
		.INIT('h8b)
	) name11090 (
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w5015_,
		_w12961_,
		_w15138_
	);
	LUT3 #(
		.INIT('h8b)
	) name11091 (
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w5015_,
		_w12969_,
		_w15139_
	);
	LUT3 #(
		.INIT('h8b)
	) name11092 (
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w5015_,
		_w13008_,
		_w15140_
	);
	LUT4 #(
		.INIT('haa02)
	) name11093 (
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w15141_
	);
	LUT3 #(
		.INIT('hf4)
	) name11094 (
		_w5022_,
		_w12947_,
		_w15141_,
		_w15142_
	);
	LUT4 #(
		.INIT('haa02)
	) name11095 (
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w15143_
	);
	LUT3 #(
		.INIT('hf4)
	) name11096 (
		_w5022_,
		_w9156_,
		_w15143_,
		_w15144_
	);
	LUT4 #(
		.INIT('haa02)
	) name11097 (
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w15145_
	);
	LUT3 #(
		.INIT('hf1)
	) name11098 (
		_w5022_,
		_w12961_,
		_w15145_,
		_w15146_
	);
	LUT4 #(
		.INIT('haa02)
	) name11099 (
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w15147_
	);
	LUT3 #(
		.INIT('hf1)
	) name11100 (
		_w5022_,
		_w12969_,
		_w15147_,
		_w15148_
	);
	LUT4 #(
		.INIT('haa02)
	) name11101 (
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		_w5020_,
		_w5021_,
		_w14995_,
		_w15149_
	);
	LUT3 #(
		.INIT('hf1)
	) name11102 (
		_w5022_,
		_w13008_,
		_w15149_,
		_w15150_
	);
	LUT4 #(
		.INIT('haa02)
	) name11103 (
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15151_
	);
	LUT3 #(
		.INIT('hf4)
	) name11104 (
		_w4979_,
		_w12947_,
		_w15151_,
		_w15152_
	);
	LUT4 #(
		.INIT('haa02)
	) name11105 (
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15153_
	);
	LUT3 #(
		.INIT('hf4)
	) name11106 (
		_w4979_,
		_w9156_,
		_w15153_,
		_w15154_
	);
	LUT4 #(
		.INIT('haa02)
	) name11107 (
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15155_
	);
	LUT3 #(
		.INIT('hf1)
	) name11108 (
		_w4979_,
		_w12961_,
		_w15155_,
		_w15156_
	);
	LUT4 #(
		.INIT('haa02)
	) name11109 (
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15157_
	);
	LUT3 #(
		.INIT('hf1)
	) name11110 (
		_w4979_,
		_w12969_,
		_w15157_,
		_w15158_
	);
	LUT4 #(
		.INIT('haa02)
	) name11111 (
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		_w4976_,
		_w4978_,
		_w15009_,
		_w15159_
	);
	LUT3 #(
		.INIT('hf1)
	) name11112 (
		_w4979_,
		_w13008_,
		_w15159_,
		_w15160_
	);
	LUT4 #(
		.INIT('h0080)
	) name11113 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w15161_
	);
	LUT2 #(
		.INIT('h4)
	) name11114 (
		\sice_ICYC_clr_reg/NET0131 ,
		\sice_SPC_reg[23]/P0001 ,
		_w15162_
	);
	LUT3 #(
		.INIT('h80)
	) name11115 (
		_w14460_,
		_w15161_,
		_w15162_,
		_w15163_
	);
	LUT4 #(
		.INIT('hc444)
	) name11116 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[9]/NET0131 ,
		_w4073_,
		_w4084_,
		_w15164_
	);
	LUT4 #(
		.INIT('h0020)
	) name11117 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_Iflag_reg[10]/NET0131 ,
		\core_c_psq_Iflag_reg[8]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w15165_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11118 (
		\core_c_psq_INT_en_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15165_,
		_w15166_
	);
	LUT2 #(
		.INIT('he)
	) name11119 (
		_w15164_,
		_w15166_,
		_w15167_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11120 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001 ,
		_w13835_,
		_w13836_,
		_w14881_,
		_w15168_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11121 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15169_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11122 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15170_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11123 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15171_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11124 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15172_
	);
	LUT4 #(
		.INIT('hccac)
	) name11125 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15173_
	);
	LUT4 #(
		.INIT('hccac)
	) name11126 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15174_
	);
	LUT4 #(
		.INIT('hccca)
	) name11127 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15175_
	);
	LUT4 #(
		.INIT('hccca)
	) name11128 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15176_
	);
	LUT4 #(
		.INIT('haccc)
	) name11129 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15177_
	);
	LUT4 #(
		.INIT('haccc)
	) name11130 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15178_
	);
	LUT4 #(
		.INIT('haccc)
	) name11131 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15179_
	);
	LUT4 #(
		.INIT('hccac)
	) name11132 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15180_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11133 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15181_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11134 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15182_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11135 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15183_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11136 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15184_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11137 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15185_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11138 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15186_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11139 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15187_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11140 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15188_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11141 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15189_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11142 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15190_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11143 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15191_
	);
	LUT4 #(
		.INIT('hccac)
	) name11144 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15192_
	);
	LUT4 #(
		.INIT('hccac)
	) name11145 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15193_
	);
	LUT4 #(
		.INIT('hccac)
	) name11146 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15194_
	);
	LUT4 #(
		.INIT('hccac)
	) name11147 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15195_
	);
	LUT4 #(
		.INIT('hccac)
	) name11148 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15196_
	);
	LUT4 #(
		.INIT('hccac)
	) name11149 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15197_
	);
	LUT4 #(
		.INIT('hccca)
	) name11150 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15198_
	);
	LUT4 #(
		.INIT('hccca)
	) name11151 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15199_
	);
	LUT4 #(
		.INIT('hccca)
	) name11152 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15200_
	);
	LUT4 #(
		.INIT('hccca)
	) name11153 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15201_
	);
	LUT4 #(
		.INIT('hccca)
	) name11154 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15202_
	);
	LUT4 #(
		.INIT('hccca)
	) name11155 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15203_
	);
	LUT4 #(
		.INIT('hccca)
	) name11156 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15204_
	);
	LUT4 #(
		.INIT('hccca)
	) name11157 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15205_
	);
	LUT4 #(
		.INIT('hccca)
	) name11158 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15206_
	);
	LUT4 #(
		.INIT('haccc)
	) name11159 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15207_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11160 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w14864_,
		_w15208_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11161 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001 ,
		_w13850_,
		_w13851_,
		_w14899_,
		_w15209_
	);
	LUT4 #(
		.INIT('h4044)
	) name11162 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTPMOVL_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15210_
	);
	LUT4 #(
		.INIT('h8000)
	) name11163 (
		_w5914_,
		_w6176_,
		_w6501_,
		_w6897_,
		_w15211_
	);
	LUT4 #(
		.INIT('hba00)
	) name11164 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w15210_,
		_w15212_
	);
	LUT4 #(
		.INIT('h00ae)
	) name11165 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w15210_,
		_w15211_,
		_w15212_,
		_w15213_
	);
	LUT4 #(
		.INIT('hba00)
	) name11166 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w15210_,
		_w15214_
	);
	LUT4 #(
		.INIT('h00ae)
	) name11167 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w15210_,
		_w15211_,
		_w15214_,
		_w15215_
	);
	LUT4 #(
		.INIT('haaca)
	) name11168 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w6897_,
		_w15210_,
		_w15211_,
		_w15216_
	);
	LUT4 #(
		.INIT('haaca)
	) name11169 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w5914_,
		_w15210_,
		_w15211_,
		_w15217_
	);
	LUT4 #(
		.INIT('h8000)
	) name11170 (
		_w7378_,
		_w7710_,
		_w7906_,
		_w8043_,
		_w15218_
	);
	LUT4 #(
		.INIT('hba00)
	) name11171 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w15210_,
		_w15219_
	);
	LUT4 #(
		.INIT('h00ae)
	) name11172 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w15210_,
		_w15218_,
		_w15219_,
		_w15220_
	);
	LUT4 #(
		.INIT('haaca)
	) name11173 (
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		_w8043_,
		_w15210_,
		_w15218_,
		_w15221_
	);
	LUT4 #(
		.INIT('hba00)
	) name11174 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w15210_,
		_w15222_
	);
	LUT4 #(
		.INIT('h00ae)
	) name11175 (
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		_w15210_,
		_w15218_,
		_w15222_,
		_w15223_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11176 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w14864_,
		_w15224_
	);
	LUT4 #(
		.INIT('hccca)
	) name11177 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15225_
	);
	LUT4 #(
		.INIT('haccc)
	) name11178 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15226_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name11179 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w15227_
	);
	LUT4 #(
		.INIT('hbf00)
	) name11180 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15227_,
		_w15228_
	);
	LUT4 #(
		.INIT('h1000)
	) name11181 (
		\core_c_dec_imm16_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15229_
	);
	LUT2 #(
		.INIT('h1)
	) name11182 (
		_w15228_,
		_w15229_,
		_w15230_
	);
	LUT4 #(
		.INIT('haaca)
	) name11183 (
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		_w7378_,
		_w15210_,
		_w15218_,
		_w15231_
	);
	LUT4 #(
		.INIT('hccac)
	) name11184 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15232_
	);
	LUT4 #(
		.INIT('haccc)
	) name11185 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15233_
	);
	LUT4 #(
		.INIT('haccc)
	) name11186 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15234_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11187 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001 ,
		_w13830_,
		_w13831_,
		_w14871_,
		_w15235_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11188 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001 ,
		_w13835_,
		_w13836_,
		_w14871_,
		_w15236_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11189 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001 ,
		_w13840_,
		_w13841_,
		_w14871_,
		_w15237_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11190 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001 ,
		_w13845_,
		_w13846_,
		_w14871_,
		_w15238_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11191 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001 ,
		_w13850_,
		_w13851_,
		_w14871_,
		_w15239_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11192 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001 ,
		_w13855_,
		_w13856_,
		_w14871_,
		_w15240_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11193 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001 ,
		_w13897_,
		_w13898_,
		_w14871_,
		_w15241_
	);
	LUT3 #(
		.INIT('hca)
	) name11194 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001 ,
		_w13861_,
		_w14871_,
		_w15242_
	);
	LUT3 #(
		.INIT('hca)
	) name11195 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001 ,
		_w13866_,
		_w14871_,
		_w15243_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11196 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001 ,
		_w13830_,
		_w13831_,
		_w14881_,
		_w15244_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11197 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001 ,
		_w13845_,
		_w13846_,
		_w14881_,
		_w15245_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11198 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001 ,
		_w13850_,
		_w13851_,
		_w14881_,
		_w15246_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11199 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001 ,
		_w13897_,
		_w13898_,
		_w14881_,
		_w15247_
	);
	LUT3 #(
		.INIT('hca)
	) name11200 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001 ,
		_w13861_,
		_w14881_,
		_w15248_
	);
	LUT3 #(
		.INIT('hca)
	) name11201 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001 ,
		_w13866_,
		_w14881_,
		_w15249_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11202 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001 ,
		_w13845_,
		_w13846_,
		_w14891_,
		_w15250_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11203 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001 ,
		_w13835_,
		_w13836_,
		_w14891_,
		_w15251_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11204 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001 ,
		_w13850_,
		_w13851_,
		_w14891_,
		_w15252_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11205 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001 ,
		_w13897_,
		_w13898_,
		_w14891_,
		_w15253_
	);
	LUT4 #(
		.INIT('hba00)
	) name11206 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13819_,
		_w15254_
	);
	LUT2 #(
		.INIT('h1)
	) name11207 (
		_w8647_,
		_w13819_,
		_w15255_
	);
	LUT4 #(
		.INIT('h222e)
	) name11208 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001 ,
		_w14891_,
		_w15254_,
		_w15255_,
		_w15256_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11209 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001 ,
		_w13830_,
		_w13831_,
		_w14899_,
		_w15257_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11210 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001 ,
		_w13840_,
		_w13841_,
		_w14899_,
		_w15258_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11211 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001 ,
		_w13845_,
		_w13846_,
		_w14899_,
		_w15259_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11212 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001 ,
		_w13855_,
		_w13856_,
		_w14899_,
		_w15260_
	);
	LUT4 #(
		.INIT('hccca)
	) name11213 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15261_
	);
	LUT3 #(
		.INIT('hca)
	) name11214 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001 ,
		_w13866_,
		_w14899_,
		_w15262_
	);
	LUT4 #(
		.INIT('h222e)
	) name11215 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001 ,
		_w14899_,
		_w15254_,
		_w15255_,
		_w15263_
	);
	LUT4 #(
		.INIT('hccca)
	) name11216 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15264_
	);
	LUT4 #(
		.INIT('hba00)
	) name11217 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w14906_,
		_w15265_
	);
	LUT4 #(
		.INIT('h1555)
	) name11218 (
		\bdma_BOVL_reg[7]/NET0131 ,
		_w5658_,
		_w5804_,
		_w9431_,
		_w15266_
	);
	LUT2 #(
		.INIT('h1)
	) name11219 (
		_w15265_,
		_w15266_,
		_w15267_
	);
	LUT4 #(
		.INIT('hba00)
	) name11220 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w14906_,
		_w15268_
	);
	LUT4 #(
		.INIT('h1555)
	) name11221 (
		\bdma_BOVL_reg[6]/NET0131 ,
		_w5658_,
		_w5804_,
		_w9431_,
		_w15269_
	);
	LUT2 #(
		.INIT('h1)
	) name11222 (
		_w15268_,
		_w15269_,
		_w15270_
	);
	LUT4 #(
		.INIT('hba00)
	) name11223 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w14906_,
		_w15271_
	);
	LUT4 #(
		.INIT('h1555)
	) name11224 (
		\bdma_BOVL_reg[5]/NET0131 ,
		_w5658_,
		_w5804_,
		_w9431_,
		_w15272_
	);
	LUT2 #(
		.INIT('h1)
	) name11225 (
		_w15271_,
		_w15272_,
		_w15273_
	);
	LUT4 #(
		.INIT('hba00)
	) name11226 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w14906_,
		_w15274_
	);
	LUT4 #(
		.INIT('h1555)
	) name11227 (
		\bdma_BOVL_reg[4]/NET0131 ,
		_w5658_,
		_w5804_,
		_w9431_,
		_w15275_
	);
	LUT2 #(
		.INIT('h1)
	) name11228 (
		_w15274_,
		_w15275_,
		_w15276_
	);
	LUT4 #(
		.INIT('hba00)
	) name11229 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w14906_,
		_w15277_
	);
	LUT4 #(
		.INIT('h1555)
	) name11230 (
		\bdma_BOVL_reg[3]/NET0131 ,
		_w5658_,
		_w5804_,
		_w9431_,
		_w15278_
	);
	LUT2 #(
		.INIT('h1)
	) name11231 (
		_w15277_,
		_w15278_,
		_w15279_
	);
	LUT4 #(
		.INIT('hba00)
	) name11232 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w14906_,
		_w15280_
	);
	LUT4 #(
		.INIT('h1555)
	) name11233 (
		\bdma_BOVL_reg[2]/NET0131 ,
		_w5658_,
		_w5804_,
		_w9431_,
		_w15281_
	);
	LUT2 #(
		.INIT('h1)
	) name11234 (
		_w15280_,
		_w15281_,
		_w15282_
	);
	LUT4 #(
		.INIT('hba00)
	) name11235 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w14906_,
		_w15283_
	);
	LUT4 #(
		.INIT('h1555)
	) name11236 (
		\bdma_BOVL_reg[1]/NET0131 ,
		_w5658_,
		_w5804_,
		_w9431_,
		_w15284_
	);
	LUT2 #(
		.INIT('h1)
	) name11237 (
		_w15283_,
		_w15284_,
		_w15285_
	);
	LUT4 #(
		.INIT('hba00)
	) name11238 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w14906_,
		_w15286_
	);
	LUT4 #(
		.INIT('h1555)
	) name11239 (
		\bdma_BOVL_reg[0]/NET0131 ,
		_w5658_,
		_w5804_,
		_w9431_,
		_w15287_
	);
	LUT2 #(
		.INIT('h1)
	) name11240 (
		_w15286_,
		_w15287_,
		_w15288_
	);
	LUT4 #(
		.INIT('hba00)
	) name11241 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13346_,
		_w15289_
	);
	LUT4 #(
		.INIT('h1555)
	) name11242 (
		\bdma_BCTL_reg[3]/NET0131 ,
		_w5658_,
		_w9431_,
		_w12824_,
		_w15290_
	);
	LUT2 #(
		.INIT('h1)
	) name11243 (
		_w15289_,
		_w15290_,
		_w15291_
	);
	LUT4 #(
		.INIT('hba00)
	) name11244 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13346_,
		_w15292_
	);
	LUT4 #(
		.INIT('h1555)
	) name11245 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w5658_,
		_w9431_,
		_w12824_,
		_w15293_
	);
	LUT2 #(
		.INIT('h1)
	) name11246 (
		_w15292_,
		_w15293_,
		_w15294_
	);
	LUT4 #(
		.INIT('hba00)
	) name11247 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w13346_,
		_w15295_
	);
	LUT4 #(
		.INIT('h1555)
	) name11248 (
		\bdma_BCTL_reg[1]/NET0131 ,
		_w5658_,
		_w9431_,
		_w12824_,
		_w15296_
	);
	LUT2 #(
		.INIT('h1)
	) name11249 (
		_w15295_,
		_w15296_,
		_w15297_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11250 (
		\bdma_BCTL_reg[15]/NET0131 ,
		_w8798_,
		_w8801_,
		_w13346_,
		_w15298_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11251 (
		\bdma_BCTL_reg[14]/NET0131 ,
		_w8757_,
		_w8760_,
		_w13346_,
		_w15299_
	);
	LUT4 #(
		.INIT('hba00)
	) name11252 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13346_,
		_w15300_
	);
	LUT4 #(
		.INIT('h1555)
	) name11253 (
		\bdma_BCTL_reg[0]/NET0131 ,
		_w5658_,
		_w9431_,
		_w12824_,
		_w15301_
	);
	LUT2 #(
		.INIT('h1)
	) name11254 (
		_w15300_,
		_w15301_,
		_w15302_
	);
	LUT4 #(
		.INIT('hccac)
	) name11255 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15303_
	);
	LUT4 #(
		.INIT('hccac)
	) name11256 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15304_
	);
	LUT4 #(
		.INIT('haccc)
	) name11257 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15305_
	);
	LUT3 #(
		.INIT('h6c)
	) name11258 (
		\sice_ICYC_reg[4]/NET0131 ,
		\sice_ICYC_reg[5]/NET0131 ,
		_w11931_,
		_w15306_
	);
	LUT4 #(
		.INIT('hccca)
	) name11259 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001 ,
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w15307_
	);
	LUT4 #(
		.INIT('hccac)
	) name11260 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15308_
	);
	LUT4 #(
		.INIT('hccac)
	) name11261 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15309_
	);
	LUT4 #(
		.INIT('h222e)
	) name11262 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001 ,
		_w14871_,
		_w15254_,
		_w15255_,
		_w15310_
	);
	LUT4 #(
		.INIT('haccc)
	) name11263 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15311_
	);
	LUT4 #(
		.INIT('haccc)
	) name11264 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15312_
	);
	LUT4 #(
		.INIT('hccac)
	) name11265 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15313_
	);
	LUT4 #(
		.INIT('hccac)
	) name11266 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15314_
	);
	LUT4 #(
		.INIT('haccc)
	) name11267 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15315_
	);
	LUT4 #(
		.INIT('hccac)
	) name11268 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15316_
	);
	LUT3 #(
		.INIT('hca)
	) name11269 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001 ,
		_w12673_,
		_w14864_,
		_w15317_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11270 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w14864_,
		_w15318_
	);
	LUT4 #(
		.INIT('haccc)
	) name11271 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15319_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11272 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w14864_,
		_w15320_
	);
	LUT4 #(
		.INIT('haccc)
	) name11273 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15321_
	);
	LUT4 #(
		.INIT('h2000)
	) name11274 (
		\memc_Dwrite_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15322_
	);
	LUT4 #(
		.INIT('h8000)
	) name11275 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w5044_,
		_w5045_,
		_w5046_,
		_w15323_
	);
	LUT3 #(
		.INIT('h08)
	) name11276 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w4090_,
		_w4091_,
		_w15324_
	);
	LUT4 #(
		.INIT('h0080)
	) name11277 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w15325_
	);
	LUT4 #(
		.INIT('h0f7f)
	) name11278 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w15326_
	);
	LUT4 #(
		.INIT('hf700)
	) name11279 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w4090_,
		_w4091_,
		_w15326_,
		_w15327_
	);
	LUT2 #(
		.INIT('h4)
	) name11280 (
		_w15323_,
		_w15327_,
		_w15328_
	);
	LUT3 #(
		.INIT('hce)
	) name11281 (
		_w8174_,
		_w15322_,
		_w15328_,
		_w15329_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11282 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15330_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11283 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w14864_,
		_w15331_
	);
	LUT4 #(
		.INIT('hccca)
	) name11284 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15332_
	);
	LUT4 #(
		.INIT('h0045)
	) name11285 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w14921_,
		_w15333_
	);
	LUT3 #(
		.INIT('h04)
	) name11286 (
		\auctl_T1Sack_reg/NET0131 ,
		\sport1_txctl_TX_reg[7]/P0001 ,
		_w14920_,
		_w15334_
	);
	LUT2 #(
		.INIT('he)
	) name11287 (
		_w15333_,
		_w15334_,
		_w15335_
	);
	LUT4 #(
		.INIT('hccca)
	) name11288 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15336_
	);
	LUT4 #(
		.INIT('h0045)
	) name11289 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w14921_,
		_w15337_
	);
	LUT3 #(
		.INIT('h04)
	) name11290 (
		\auctl_T1Sack_reg/NET0131 ,
		\sport1_txctl_TX_reg[6]/P0001 ,
		_w14920_,
		_w15338_
	);
	LUT2 #(
		.INIT('he)
	) name11291 (
		_w15337_,
		_w15338_,
		_w15339_
	);
	LUT4 #(
		.INIT('h0045)
	) name11292 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w14921_,
		_w15340_
	);
	LUT3 #(
		.INIT('h04)
	) name11293 (
		\auctl_T1Sack_reg/NET0131 ,
		\sport1_txctl_TX_reg[5]/P0001 ,
		_w14920_,
		_w15341_
	);
	LUT2 #(
		.INIT('he)
	) name11294 (
		_w15340_,
		_w15341_,
		_w15342_
	);
	LUT4 #(
		.INIT('h0045)
	) name11295 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w14921_,
		_w15343_
	);
	LUT3 #(
		.INIT('h04)
	) name11296 (
		\auctl_T1Sack_reg/NET0131 ,
		\sport1_txctl_TX_reg[4]/P0001 ,
		_w14920_,
		_w15344_
	);
	LUT2 #(
		.INIT('he)
	) name11297 (
		_w15343_,
		_w15344_,
		_w15345_
	);
	LUT4 #(
		.INIT('h0045)
	) name11298 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w14921_,
		_w15346_
	);
	LUT3 #(
		.INIT('h04)
	) name11299 (
		\auctl_T1Sack_reg/NET0131 ,
		\sport1_txctl_TX_reg[3]/P0001 ,
		_w14920_,
		_w15347_
	);
	LUT2 #(
		.INIT('he)
	) name11300 (
		_w15346_,
		_w15347_,
		_w15348_
	);
	LUT4 #(
		.INIT('h0045)
	) name11301 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w14921_,
		_w15349_
	);
	LUT3 #(
		.INIT('h04)
	) name11302 (
		\auctl_T1Sack_reg/NET0131 ,
		\sport1_txctl_TX_reg[2]/P0001 ,
		_w14920_,
		_w15350_
	);
	LUT2 #(
		.INIT('he)
	) name11303 (
		_w15349_,
		_w15350_,
		_w15351_
	);
	LUT4 #(
		.INIT('h0045)
	) name11304 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w14921_,
		_w15352_
	);
	LUT3 #(
		.INIT('h04)
	) name11305 (
		\auctl_T1Sack_reg/NET0131 ,
		\sport1_txctl_TX_reg[1]/P0001 ,
		_w14920_,
		_w15353_
	);
	LUT2 #(
		.INIT('he)
	) name11306 (
		_w15352_,
		_w15353_,
		_w15354_
	);
	LUT4 #(
		.INIT('haa03)
	) name11307 (
		\sport1_txctl_TX_reg[15]/P0001 ,
		_w8798_,
		_w8801_,
		_w14921_,
		_w15355_
	);
	LUT4 #(
		.INIT('haa03)
	) name11308 (
		\sport1_txctl_TX_reg[14]/P0001 ,
		_w8757_,
		_w8760_,
		_w14921_,
		_w15356_
	);
	LUT4 #(
		.INIT('h0045)
	) name11309 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w14921_,
		_w15357_
	);
	LUT3 #(
		.INIT('h04)
	) name11310 (
		\auctl_T1Sack_reg/NET0131 ,
		\sport1_txctl_TX_reg[0]/P0001 ,
		_w14920_,
		_w15358_
	);
	LUT2 #(
		.INIT('he)
	) name11311 (
		_w15357_,
		_w15358_,
		_w15359_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11312 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w14864_,
		_w15360_
	);
	LUT4 #(
		.INIT('haccc)
	) name11313 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15361_
	);
	LUT4 #(
		.INIT('haccc)
	) name11314 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15362_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11315 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001 ,
		_w13835_,
		_w13836_,
		_w14899_,
		_w15363_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11316 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001 ,
		_w13840_,
		_w13841_,
		_w14891_,
		_w15364_
	);
	LUT3 #(
		.INIT('h20)
	) name11317 (
		\core_eu_ec_cun_updateMV_C_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15365_
	);
	LUT2 #(
		.INIT('he)
	) name11318 (
		_w13380_,
		_w15365_,
		_w15366_
	);
	LUT3 #(
		.INIT('h28)
	) name11319 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14324_,
		_w14390_,
		_w15367_
	);
	LUT2 #(
		.INIT('h9)
	) name11320 (
		_w14314_,
		_w14319_,
		_w15368_
	);
	LUT2 #(
		.INIT('h1)
	) name11321 (
		_w14317_,
		_w14321_,
		_w15369_
	);
	LUT2 #(
		.INIT('h8)
	) name11322 (
		_w14317_,
		_w14321_,
		_w15370_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name11323 (
		_w14289_,
		_w14292_,
		_w15369_,
		_w15370_,
		_w15371_
	);
	LUT3 #(
		.INIT('h41)
	) name11324 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15368_,
		_w15371_,
		_w15372_
	);
	LUT2 #(
		.INIT('h1)
	) name11325 (
		_w15367_,
		_w15372_,
		_w15373_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11326 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001 ,
		_w13830_,
		_w13831_,
		_w14931_,
		_w15374_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11327 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001 ,
		_w13835_,
		_w13836_,
		_w14931_,
		_w15375_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11328 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001 ,
		_w13840_,
		_w13841_,
		_w14931_,
		_w15376_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11329 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001 ,
		_w13845_,
		_w13846_,
		_w14931_,
		_w15377_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11330 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001 ,
		_w13850_,
		_w13851_,
		_w14931_,
		_w15378_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11331 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001 ,
		_w13855_,
		_w13856_,
		_w14931_,
		_w15379_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11332 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001 ,
		_w13897_,
		_w13898_,
		_w14931_,
		_w15380_
	);
	LUT3 #(
		.INIT('hca)
	) name11333 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001 ,
		_w13861_,
		_w14931_,
		_w15381_
	);
	LUT3 #(
		.INIT('hca)
	) name11334 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001 ,
		_w13866_,
		_w14931_,
		_w15382_
	);
	LUT4 #(
		.INIT('h222e)
	) name11335 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001 ,
		_w14931_,
		_w15254_,
		_w15255_,
		_w15383_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11336 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w14942_,
		_w15384_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11337 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w14942_,
		_w15385_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11338 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w14942_,
		_w15386_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11339 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w14942_,
		_w15387_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11340 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w14942_,
		_w15388_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11341 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w14942_,
		_w15389_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11342 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w14942_,
		_w15390_
	);
	LUT3 #(
		.INIT('hca)
	) name11343 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001 ,
		_w11318_,
		_w14942_,
		_w15391_
	);
	LUT3 #(
		.INIT('hca)
	) name11344 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001 ,
		_w12673_,
		_w14942_,
		_w15392_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11345 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w14942_,
		_w15393_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11346 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w14955_,
		_w15394_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11347 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w14955_,
		_w15395_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11348 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w14955_,
		_w15396_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11349 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w14955_,
		_w15397_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11350 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w14955_,
		_w15398_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11351 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w14955_,
		_w15399_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11352 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w14955_,
		_w15400_
	);
	LUT3 #(
		.INIT('hca)
	) name11353 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001 ,
		_w11318_,
		_w14955_,
		_w15401_
	);
	LUT3 #(
		.INIT('hca)
	) name11354 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001 ,
		_w12673_,
		_w14955_,
		_w15402_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11355 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w14955_,
		_w15403_
	);
	LUT3 #(
		.INIT('hca)
	) name11356 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001 ,
		_w13861_,
		_w14891_,
		_w15404_
	);
	LUT3 #(
		.INIT('h80)
	) name11357 (
		_w5028_,
		_w12393_,
		_w13333_,
		_w15405_
	);
	LUT2 #(
		.INIT('h8)
	) name11358 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w4106_,
		_w15406_
	);
	LUT3 #(
		.INIT('hf8)
	) name11359 (
		_w14570_,
		_w15405_,
		_w15406_,
		_w15407_
	);
	LUT3 #(
		.INIT('hca)
	) name11360 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001 ,
		_w13861_,
		_w14899_,
		_w15408_
	);
	LUT4 #(
		.INIT('haccc)
	) name11361 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15409_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11362 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001 ,
		_w13897_,
		_w13898_,
		_w14899_,
		_w15410_
	);
	LUT4 #(
		.INIT('hcacc)
	) name11363 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15411_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11364 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w14864_,
		_w15412_
	);
	LUT4 #(
		.INIT('haccc)
	) name11365 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w15413_
	);
	LUT3 #(
		.INIT('hca)
	) name11366 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001 ,
		_w13866_,
		_w14891_,
		_w15414_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11367 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001 ,
		_w13855_,
		_w13856_,
		_w14891_,
		_w15415_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11368 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001 ,
		_w13830_,
		_w13831_,
		_w14891_,
		_w15416_
	);
	LUT4 #(
		.INIT('h222e)
	) name11369 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001 ,
		_w14881_,
		_w15254_,
		_w15255_,
		_w15417_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11370 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001 ,
		_w13855_,
		_w13856_,
		_w14881_,
		_w15418_
	);
	LUT3 #(
		.INIT('hca)
	) name11371 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001 ,
		_w11318_,
		_w14864_,
		_w15419_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11372 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w14864_,
		_w15420_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11373 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001 ,
		_w13840_,
		_w13841_,
		_w14881_,
		_w15421_
	);
	LUT3 #(
		.INIT('h40)
	) name11374 (
		\sice_GO_NX_reg/NET0131 ,
		\sice_IDONE_reg/NET0131 ,
		_w4084_,
		_w15422_
	);
	LUT4 #(
		.INIT('h0001)
	) name11375 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_NOP_E_reg/P0001 ,
		_w4971_,
		_w9453_,
		_w15423_
	);
	LUT2 #(
		.INIT('he)
	) name11376 (
		_w15422_,
		_w15423_,
		_w15424_
	);
	LUT3 #(
		.INIT('h78)
	) name11377 (
		\sice_IIRC_reg[0]/NET0131 ,
		\sice_IIRC_reg[1]/NET0131 ,
		\sice_IIRC_reg[2]/NET0131 ,
		_w15425_
	);
	LUT3 #(
		.INIT('h78)
	) name11378 (
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[1]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[2]/NET0131 ,
		_w15426_
	);
	LUT3 #(
		.INIT('h78)
	) name11379 (
		\sice_ICYC_reg[0]/NET0131 ,
		\sice_ICYC_reg[1]/NET0131 ,
		\sice_ICYC_reg[2]/NET0131 ,
		_w15427_
	);
	LUT2 #(
		.INIT('h8)
	) name11380 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		_w11300_,
		_w15428_
	);
	LUT3 #(
		.INIT('hca)
	) name11381 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001 ,
		_w13821_,
		_w15428_,
		_w15429_
	);
	LUT3 #(
		.INIT('h3a)
	) name11382 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001 ,
		_w13826_,
		_w15428_,
		_w15430_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11383 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001 ,
		_w13830_,
		_w13831_,
		_w15428_,
		_w15431_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11384 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001 ,
		_w13835_,
		_w13836_,
		_w15428_,
		_w15432_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11385 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001 ,
		_w13840_,
		_w13841_,
		_w15428_,
		_w15433_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11386 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001 ,
		_w13845_,
		_w13846_,
		_w15428_,
		_w15434_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11387 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001 ,
		_w13850_,
		_w13851_,
		_w15428_,
		_w15435_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11388 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001 ,
		_w13855_,
		_w13856_,
		_w15428_,
		_w15436_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11389 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001 ,
		_w13897_,
		_w13898_,
		_w15428_,
		_w15437_
	);
	LUT3 #(
		.INIT('hca)
	) name11390 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001 ,
		_w13861_,
		_w15428_,
		_w15438_
	);
	LUT3 #(
		.INIT('hca)
	) name11391 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001 ,
		_w13866_,
		_w15428_,
		_w15439_
	);
	LUT4 #(
		.INIT('h5300)
	) name11392 (
		_w5760_,
		_w8740_,
		_w13819_,
		_w15428_,
		_w15440_
	);
	LUT3 #(
		.INIT('h13)
	) name11393 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001 ,
		_w11300_,
		_w15441_
	);
	LUT2 #(
		.INIT('h1)
	) name11394 (
		_w15440_,
		_w15441_,
		_w15442_
	);
	LUT3 #(
		.INIT('h4c)
	) name11395 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001 ,
		_w11300_,
		_w15443_
	);
	LUT4 #(
		.INIT('hac00)
	) name11396 (
		_w6758_,
		_w8717_,
		_w13819_,
		_w15428_,
		_w15444_
	);
	LUT2 #(
		.INIT('he)
	) name11397 (
		_w15443_,
		_w15444_,
		_w15445_
	);
	LUT3 #(
		.INIT('h3a)
	) name11398 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001 ,
		_w13878_,
		_w15428_,
		_w15446_
	);
	LUT3 #(
		.INIT('hca)
	) name11399 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001 ,
		_w13883_,
		_w15428_,
		_w15447_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11400 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001 ,
		_w15254_,
		_w15255_,
		_w15428_,
		_w15448_
	);
	LUT3 #(
		.INIT('h13)
	) name11401 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 ,
		_w9894_,
		_w15449_
	);
	LUT4 #(
		.INIT('h0002)
	) name11402 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w15449_,
		_w15450_
	);
	LUT4 #(
		.INIT('h313b)
	) name11403 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 ,
		_w11308_,
		_w11635_,
		_w15451_
	);
	LUT4 #(
		.INIT('h2f00)
	) name11404 (
		_w12282_,
		_w14918_,
		_w15450_,
		_w15451_,
		_w15452_
	);
	LUT2 #(
		.INIT('h1)
	) name11405 (
		_w11624_,
		_w15452_,
		_w15453_
	);
	LUT3 #(
		.INIT('h41)
	) name11406 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12246_,
		_w14404_,
		_w15454_
	);
	LUT3 #(
		.INIT('hf8)
	) name11407 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12293_,
		_w15454_,
		_w15455_
	);
	LUT4 #(
		.INIT('hc480)
	) name11408 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w12293_,
		_w14405_,
		_w15456_
	);
	LUT2 #(
		.INIT('he)
	) name11409 (
		_w15453_,
		_w15456_,
		_w15457_
	);
	LUT4 #(
		.INIT('h1011)
	) name11410 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w6378_,
		_w6498_,
		_w6500_,
		_w15458_
	);
	LUT4 #(
		.INIT('h5455)
	) name11411 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w13129_,
		_w13130_,
		_w13138_,
		_w15459_
	);
	LUT3 #(
		.INIT('h40)
	) name11412 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w15460_
	);
	LUT2 #(
		.INIT('h1)
	) name11413 (
		_w13158_,
		_w15460_,
		_w15461_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11414 (
		_w13155_,
		_w13137_,
		_w15459_,
		_w15461_,
		_w15462_
	);
	LUT4 #(
		.INIT('hafac)
	) name11415 (
		\sport0_rxctl_RXSHT_reg[2]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w15463_
	);
	LUT4 #(
		.INIT('h0002)
	) name11416 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w15464_
	);
	LUT4 #(
		.INIT('hffb0)
	) name11417 (
		_w15458_,
		_w15462_,
		_w15463_,
		_w15464_,
		_w15465_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11418 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w12282_,
		_w15466_
	);
	LUT3 #(
		.INIT('h13)
	) name11419 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 ,
		_w9894_,
		_w15467_
	);
	LUT4 #(
		.INIT('h0002)
	) name11420 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w15467_,
		_w15468_
	);
	LUT4 #(
		.INIT('h313b)
	) name11421 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 ,
		_w11308_,
		_w11635_,
		_w15469_
	);
	LUT4 #(
		.INIT('h1055)
	) name11422 (
		_w11624_,
		_w15466_,
		_w15468_,
		_w15469_,
		_w15470_
	);
	LUT2 #(
		.INIT('h9)
	) name11423 (
		_w11264_,
		_w11270_,
		_w15471_
	);
	LUT4 #(
		.INIT('h718e)
	) name11424 (
		_w11250_,
		_w11268_,
		_w11272_,
		_w15471_,
		_w15472_
	);
	LUT3 #(
		.INIT('h8d)
	) name11425 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14432_,
		_w15472_,
		_w15473_
	);
	LUT4 #(
		.INIT('h80c4)
	) name11426 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w14432_,
		_w15472_,
		_w15474_
	);
	LUT2 #(
		.INIT('he)
	) name11427 (
		_w15470_,
		_w15474_,
		_w15475_
	);
	LUT3 #(
		.INIT('h6c)
	) name11428 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		_w14698_,
		_w15476_
	);
	LUT2 #(
		.INIT('hd)
	) name11429 (
		\clkc_CTR_cnt_reg[0]/NET0131 ,
		\clkc_CTR_cnt_reg[1]/NET0131 ,
		_w15477_
	);
	LUT3 #(
		.INIT('h13)
	) name11430 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001 ,
		_w9894_,
		_w15478_
	);
	LUT4 #(
		.INIT('h0002)
	) name11431 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w15478_,
		_w15479_
	);
	LUT4 #(
		.INIT('h5700)
	) name11432 (
		_w11625_,
		_w13610_,
		_w13611_,
		_w15479_,
		_w15480_
	);
	LUT4 #(
		.INIT('h313b)
	) name11433 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001 ,
		_w11631_,
		_w11635_,
		_w15481_
	);
	LUT2 #(
		.INIT('h2)
	) name11434 (
		_w11624_,
		_w12362_,
		_w15482_
	);
	LUT4 #(
		.INIT('hff45)
	) name11435 (
		_w11624_,
		_w15480_,
		_w15481_,
		_w15482_,
		_w15483_
	);
	LUT2 #(
		.INIT('h8)
	) name11436 (
		_w9946_,
		_w12362_,
		_w15484_
	);
	LUT2 #(
		.INIT('h2)
	) name11437 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001 ,
		_w11656_,
		_w15485_
	);
	LUT3 #(
		.INIT('h01)
	) name11438 (
		_w9946_,
		_w11659_,
		_w15485_,
		_w15486_
	);
	LUT4 #(
		.INIT('hfd00)
	) name11439 (
		_w11655_,
		_w13610_,
		_w13611_,
		_w15486_,
		_w15487_
	);
	LUT2 #(
		.INIT('h1)
	) name11440 (
		_w15484_,
		_w15487_,
		_w15488_
	);
	LUT4 #(
		.INIT('h2700)
	) name11441 (
		_w9455_,
		_w9860_,
		_w9878_,
		_w9895_,
		_w15489_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11442 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001 ,
		_w9451_,
		_w9453_,
		_w9894_,
		_w15490_
	);
	LUT2 #(
		.INIT('he)
	) name11443 (
		_w15489_,
		_w15490_,
		_w15491_
	);
	LUT4 #(
		.INIT('h082a)
	) name11444 (
		_w9454_,
		_w9455_,
		_w9860_,
		_w9878_,
		_w15492_
	);
	LUT2 #(
		.INIT('h2)
	) name11445 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001 ,
		_w9454_,
		_w15493_
	);
	LUT2 #(
		.INIT('he)
	) name11446 (
		_w15492_,
		_w15493_,
		_w15494_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11447 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w12282_,
		_w15495_
	);
	LUT3 #(
		.INIT('h13)
	) name11448 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 ,
		_w9894_,
		_w15496_
	);
	LUT4 #(
		.INIT('h0002)
	) name11449 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w15496_,
		_w15497_
	);
	LUT4 #(
		.INIT('h313b)
	) name11450 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 ,
		_w11308_,
		_w11635_,
		_w15498_
	);
	LUT4 #(
		.INIT('h1055)
	) name11451 (
		_w11624_,
		_w15495_,
		_w15497_,
		_w15498_,
		_w15499_
	);
	LUT4 #(
		.INIT('h1441)
	) name11452 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11250_,
		_w11268_,
		_w11272_,
		_w15500_
	);
	LUT3 #(
		.INIT('h07)
	) name11453 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15472_,
		_w15500_,
		_w15501_
	);
	LUT4 #(
		.INIT('h048c)
	) name11454 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w12243_,
		_w15472_,
		_w15502_
	);
	LUT2 #(
		.INIT('he)
	) name11455 (
		_w15499_,
		_w15502_,
		_w15503_
	);
	LUT3 #(
		.INIT('h37)
	) name11456 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w15504_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11457 (
		_w5044_,
		_w5045_,
		_w5046_,
		_w15504_,
		_w15505_
	);
	LUT2 #(
		.INIT('h8)
	) name11458 (
		_w11917_,
		_w15505_,
		_w15506_
	);
	LUT2 #(
		.INIT('h7)
	) name11459 (
		_w11917_,
		_w15505_,
		_w15507_
	);
	LUT4 #(
		.INIT('h2000)
	) name11460 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w15508_
	);
	LUT2 #(
		.INIT('h8)
	) name11461 (
		_w14460_,
		_w15508_,
		_w15509_
	);
	LUT4 #(
		.INIT('h084c)
	) name11462 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w12293_,
		_w14405_,
		_w15510_
	);
	LUT2 #(
		.INIT('h2)
	) name11463 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001 ,
		_w11310_,
		_w15511_
	);
	LUT3 #(
		.INIT('h01)
	) name11464 (
		_w9946_,
		_w12442_,
		_w15511_,
		_w15512_
	);
	LUT3 #(
		.INIT('h70)
	) name11465 (
		_w12440_,
		_w14918_,
		_w15512_,
		_w15513_
	);
	LUT2 #(
		.INIT('h1)
	) name11466 (
		_w15510_,
		_w15513_,
		_w15514_
	);
	LUT4 #(
		.INIT('h8000)
	) name11467 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w5028_,
		_w5044_,
		_w12393_,
		_w15515_
	);
	LUT4 #(
		.INIT('h8c80)
	) name11468 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		_w4102_,
		_w4104_,
		_w15515_,
		_w15516_
	);
	LUT3 #(
		.INIT('h80)
	) name11469 (
		_w4761_,
		_w9080_,
		_w12533_,
		_w15517_
	);
	LUT3 #(
		.INIT('h7f)
	) name11470 (
		_w4761_,
		_w9080_,
		_w12533_,
		_w15518_
	);
	LUT4 #(
		.INIT('h8000)
	) name11471 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w15519_
	);
	LUT2 #(
		.INIT('h8)
	) name11472 (
		_w14460_,
		_w15519_,
		_w15520_
	);
	LUT4 #(
		.INIT('h4c08)
	) name11473 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w14432_,
		_w15472_,
		_w15521_
	);
	LUT4 #(
		.INIT('he400)
	) name11474 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w12440_,
		_w15522_
	);
	LUT2 #(
		.INIT('h2)
	) name11475 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001 ,
		_w11310_,
		_w15523_
	);
	LUT3 #(
		.INIT('h01)
	) name11476 (
		_w9946_,
		_w12442_,
		_w15523_,
		_w15524_
	);
	LUT2 #(
		.INIT('h4)
	) name11477 (
		_w15522_,
		_w15524_,
		_w15525_
	);
	LUT2 #(
		.INIT('h1)
	) name11478 (
		_w15521_,
		_w15525_,
		_w15526_
	);
	LUT4 #(
		.INIT('h0800)
	) name11479 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w15527_
	);
	LUT2 #(
		.INIT('h8)
	) name11480 (
		_w14460_,
		_w15527_,
		_w15528_
	);
	LUT4 #(
		.INIT('hc840)
	) name11481 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w12243_,
		_w15472_,
		_w15529_
	);
	LUT4 #(
		.INIT('he400)
	) name11482 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w12440_,
		_w15530_
	);
	LUT2 #(
		.INIT('h2)
	) name11483 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001 ,
		_w11310_,
		_w15531_
	);
	LUT3 #(
		.INIT('h01)
	) name11484 (
		_w9946_,
		_w12442_,
		_w15531_,
		_w15532_
	);
	LUT2 #(
		.INIT('h4)
	) name11485 (
		_w15530_,
		_w15532_,
		_w15533_
	);
	LUT2 #(
		.INIT('h1)
	) name11486 (
		_w15529_,
		_w15533_,
		_w15534_
	);
	LUT3 #(
		.INIT('h08)
	) name11487 (
		T_ICE_RSTn_pad,
		T_RSTn_pad,
		\clkc_RSTtext_reg/P0001 ,
		_w15535_
	);
	LUT2 #(
		.INIT('h7)
	) name11488 (
		_w14449_,
		_w15535_,
		_w15536_
	);
	LUT4 #(
		.INIT('h8a00)
	) name11489 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w12895_,
		_w15537_
	);
	LUT2 #(
		.INIT('he)
	) name11490 (
		\core_c_psq_SSTAT_reg[7]/NET0131 ,
		_w15537_,
		_w15538_
	);
	LUT4 #(
		.INIT('hbf00)
	) name11491 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12389_,
		_w15539_
	);
	LUT4 #(
		.INIT('h1000)
	) name11492 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15540_
	);
	LUT3 #(
		.INIT('h02)
	) name11493 (
		_w4102_,
		_w15540_,
		_w15539_,
		_w15541_
	);
	LUT4 #(
		.INIT('h2000)
	) name11494 (
		\core_c_dec_RET_Ed_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15542_
	);
	LUT4 #(
		.INIT('haa80)
	) name11495 (
		_w4102_,
		_w8174_,
		_w13450_,
		_w15542_,
		_w15543_
	);
	LUT4 #(
		.INIT('h1000)
	) name11496 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w15544_
	);
	LUT2 #(
		.INIT('h8)
	) name11497 (
		_w14460_,
		_w15544_,
		_w15545_
	);
	LUT2 #(
		.INIT('h2)
	) name11498 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_txctl_TCS_reg[1]/NET0131 ,
		_w15546_
	);
	LUT2 #(
		.INIT('h4)
	) name11499 (
		_w12552_,
		_w15546_,
		_w15547_
	);
	LUT4 #(
		.INIT('hcecc)
	) name11500 (
		\sport0_regs_AUTOreg_DO_reg[1]/NET0131 ,
		\sport0_txctl_TSreqi_reg/NET0131 ,
		_w12552_,
		_w15546_,
		_w15548_
	);
	LUT3 #(
		.INIT('h9c)
	) name11501 (
		\bdma_BSreq_reg/NET0131 ,
		\bdma_BWcnt_reg[0]/NET0131 ,
		_w4764_,
		_w15549_
	);
	LUT2 #(
		.INIT('h4)
	) name11502 (
		_w9413_,
		_w15549_,
		_w15550_
	);
	LUT2 #(
		.INIT('h6)
	) name11503 (
		_w14317_,
		_w14321_,
		_w15551_
	);
	LUT3 #(
		.INIT('h4b)
	) name11504 (
		_w14289_,
		_w14292_,
		_w15551_,
		_w15552_
	);
	LUT4 #(
		.INIT('h1045)
	) name11505 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14289_,
		_w14292_,
		_w15551_,
		_w15553_
	);
	LUT4 #(
		.INIT('h00d7)
	) name11506 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15368_,
		_w15371_,
		_w15553_,
		_w15554_
	);
	LUT4 #(
		.INIT('hff28)
	) name11507 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15368_,
		_w15371_,
		_w15553_,
		_w15555_
	);
	LUT2 #(
		.INIT('h2)
	) name11508 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_txctl_TCS_reg[1]/NET0131 ,
		_w15556_
	);
	LUT2 #(
		.INIT('h4)
	) name11509 (
		_w14269_,
		_w15556_,
		_w15557_
	);
	LUT4 #(
		.INIT('hcecc)
	) name11510 (
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		\sport1_txctl_TSreqi_reg/NET0131 ,
		_w14269_,
		_w15556_,
		_w15558_
	);
	LUT4 #(
		.INIT('h0200)
	) name11511 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w15559_
	);
	LUT2 #(
		.INIT('h8)
	) name11512 (
		_w14460_,
		_w15559_,
		_w15560_
	);
	LUT3 #(
		.INIT('h01)
	) name11513 (
		\bdma_BWcnt_reg[2]/NET0131 ,
		\bdma_BWcnt_reg[3]/NET0131 ,
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w15561_
	);
	LUT4 #(
		.INIT('h8000)
	) name11514 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWcnt_reg[0]/NET0131 ,
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w15562_
	);
	LUT2 #(
		.INIT('h8)
	) name11515 (
		_w15561_,
		_w15562_,
		_w15563_
	);
	LUT3 #(
		.INIT('h10)
	) name11516 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w15564_
	);
	LUT3 #(
		.INIT('h80)
	) name11517 (
		_w5028_,
		_w5045_,
		_w15564_,
		_w15565_
	);
	LUT4 #(
		.INIT('h1000)
	) name11518 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4428_,
		_w8172_,
		_w15565_,
		_w15566_
	);
	LUT3 #(
		.INIT('h01)
	) name11519 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w15567_
	);
	LUT4 #(
		.INIT('h0010)
	) name11520 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w15568_
	);
	LUT2 #(
		.INIT('h8)
	) name11521 (
		_w14460_,
		_w15568_,
		_w15569_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11522 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10132_,
		_w11290_,
		_w12237_,
		_w15570_
	);
	LUT3 #(
		.INIT('h14)
	) name11523 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10132_,
		_w12215_,
		_w15571_
	);
	LUT2 #(
		.INIT('h1)
	) name11524 (
		_w15570_,
		_w15571_,
		_w15572_
	);
	LUT3 #(
		.INIT('he8)
	) name11525 (
		\core_c_psq_T_IRQ1p_reg/P0001 ,
		\core_c_psq_irq1_de_IN_syn_reg/P0001 ,
		\core_c_psq_irq1_de_OUT_reg/P0001 ,
		_w15573_
	);
	LUT3 #(
		.INIT('he8)
	) name11526 (
		\core_c_psq_T_IRQ0p_reg/P0001 ,
		\core_c_psq_irq0_de_IN_syn_reg/P0001 ,
		\core_c_psq_irq0_de_OUT_reg/P0001 ,
		_w15574_
	);
	LUT3 #(
		.INIT('h8a)
	) name11527 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15575_
	);
	LUT2 #(
		.INIT('h2)
	) name11528 (
		\core_c_psq_IFC_reg[10]/NET0131 ,
		\core_c_psq_IFC_reg[11]/NET0131 ,
		_w15576_
	);
	LUT4 #(
		.INIT('h7500)
	) name11529 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15576_,
		_w15577_
	);
	LUT4 #(
		.INIT('hff10)
	) name11530 (
		_w6263_,
		_w6362_,
		_w15575_,
		_w15577_,
		_w15578_
	);
	LUT3 #(
		.INIT('he8)
	) name11531 (
		\core_c_psq_T_IRQ2p_reg/P0001 ,
		\core_c_psq_irq2_de_IN_syn_reg/P0001 ,
		\core_c_psq_irq2_de_OUT_reg/P0001 ,
		_w15579_
	);
	LUT2 #(
		.INIT('h2)
	) name11532 (
		\core_c_psq_IFC_reg[8]/NET0131 ,
		\core_c_psq_IFC_reg[9]/NET0131 ,
		_w15580_
	);
	LUT4 #(
		.INIT('h7500)
	) name11533 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15580_,
		_w15581_
	);
	LUT4 #(
		.INIT('hff10)
	) name11534 (
		_w7140_,
		_w7240_,
		_w15575_,
		_w15581_,
		_w15582_
	);
	LUT3 #(
		.INIT('he8)
	) name11535 (
		\core_c_psq_T_IRQL1p_reg/P0001 ,
		\core_c_psq_irql1_de_IN_syn_reg/P0001 ,
		\core_c_psq_irql1_de_OUT_reg/P0001 ,
		_w15583_
	);
	LUT2 #(
		.INIT('h8)
	) name11536 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		_w11300_,
		_w15584_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11537 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w15584_,
		_w15585_
	);
	LUT3 #(
		.INIT('h13)
	) name11538 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001 ,
		_w11300_,
		_w15586_
	);
	LUT2 #(
		.INIT('h1)
	) name11539 (
		_w15585_,
		_w15586_,
		_w15587_
	);
	LUT2 #(
		.INIT('h8)
	) name11540 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		_w11300_,
		_w15588_
	);
	LUT3 #(
		.INIT('hca)
	) name11541 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001 ,
		_w12486_,
		_w15588_,
		_w15589_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11542 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w15588_,
		_w15590_
	);
	LUT3 #(
		.INIT('h13)
	) name11543 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001 ,
		_w11300_,
		_w15591_
	);
	LUT2 #(
		.INIT('h1)
	) name11544 (
		_w15590_,
		_w15591_,
		_w15592_
	);
	LUT2 #(
		.INIT('h8)
	) name11545 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		_w9894_,
		_w15593_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11546 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w15593_,
		_w15594_
	);
	LUT3 #(
		.INIT('h13)
	) name11547 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001 ,
		_w9894_,
		_w15595_
	);
	LUT2 #(
		.INIT('h1)
	) name11548 (
		_w15594_,
		_w15595_,
		_w15596_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11549 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w15584_,
		_w15597_
	);
	LUT3 #(
		.INIT('h13)
	) name11550 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001 ,
		_w11300_,
		_w15598_
	);
	LUT2 #(
		.INIT('h1)
	) name11551 (
		_w15597_,
		_w15598_,
		_w15599_
	);
	LUT2 #(
		.INIT('h8)
	) name11552 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		_w9894_,
		_w15600_
	);
	LUT3 #(
		.INIT('hca)
	) name11553 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001 ,
		_w12284_,
		_w15600_,
		_w15601_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11554 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w15600_,
		_w15602_
	);
	LUT3 #(
		.INIT('h13)
	) name11555 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001 ,
		_w9894_,
		_w15603_
	);
	LUT2 #(
		.INIT('h1)
	) name11556 (
		_w15602_,
		_w15603_,
		_w15604_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11557 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w15600_,
		_w15605_
	);
	LUT3 #(
		.INIT('h13)
	) name11558 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001 ,
		_w9894_,
		_w15606_
	);
	LUT2 #(
		.INIT('h1)
	) name11559 (
		_w15605_,
		_w15606_,
		_w15607_
	);
	LUT3 #(
		.INIT('hca)
	) name11560 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001 ,
		_w12486_,
		_w15600_,
		_w15608_
	);
	LUT3 #(
		.INIT('hca)
	) name11561 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001 ,
		_w14918_,
		_w15584_,
		_w15609_
	);
	LUT3 #(
		.INIT('hca)
	) name11562 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001 ,
		_w14918_,
		_w15593_,
		_w15610_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11563 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w15593_,
		_w15611_
	);
	LUT3 #(
		.INIT('h13)
	) name11564 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001 ,
		_w9894_,
		_w15612_
	);
	LUT2 #(
		.INIT('h1)
	) name11565 (
		_w15611_,
		_w15612_,
		_w15613_
	);
	LUT3 #(
		.INIT('hca)
	) name11566 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001 ,
		_w14866_,
		_w15593_,
		_w15614_
	);
	LUT3 #(
		.INIT('hca)
	) name11567 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001 ,
		_w14918_,
		_w15588_,
		_w15615_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11568 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w15588_,
		_w15616_
	);
	LUT3 #(
		.INIT('h13)
	) name11569 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001 ,
		_w11300_,
		_w15617_
	);
	LUT2 #(
		.INIT('h1)
	) name11570 (
		_w15616_,
		_w15617_,
		_w15618_
	);
	LUT3 #(
		.INIT('hca)
	) name11571 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001 ,
		_w12284_,
		_w15588_,
		_w15619_
	);
	LUT3 #(
		.INIT('hca)
	) name11572 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001 ,
		_w14866_,
		_w15588_,
		_w15620_
	);
	LUT3 #(
		.INIT('hca)
	) name11573 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001 ,
		_w14866_,
		_w15600_,
		_w15621_
	);
	LUT3 #(
		.INIT('hca)
	) name11574 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001 ,
		_w12486_,
		_w15593_,
		_w15622_
	);
	LUT3 #(
		.INIT('hca)
	) name11575 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001 ,
		_w12284_,
		_w15593_,
		_w15623_
	);
	LUT3 #(
		.INIT('hca)
	) name11576 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001 ,
		_w14918_,
		_w15600_,
		_w15624_
	);
	LUT3 #(
		.INIT('hca)
	) name11577 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001 ,
		_w14866_,
		_w15584_,
		_w15625_
	);
	LUT3 #(
		.INIT('hca)
	) name11578 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001 ,
		_w12486_,
		_w15584_,
		_w15626_
	);
	LUT3 #(
		.INIT('hca)
	) name11579 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001 ,
		_w12284_,
		_w15584_,
		_w15627_
	);
	LUT4 #(
		.INIT('h0015)
	) name11580 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4971_,
		_w15628_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11581 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8914_,
		_w8915_,
		_w8913_,
		_w15629_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11582 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w7634_,
		_w7705_,
		_w15629_,
		_w15630_
	);
	LUT3 #(
		.INIT('h2e)
	) name11583 (
		\regout_STD_C_reg[5]/P0001 ,
		_w15628_,
		_w15630_,
		_w15631_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11584 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w15600_,
		_w15632_
	);
	LUT4 #(
		.INIT('h4555)
	) name11585 (
		T_BRn_pad,
		\core_c_psq_PCS_reg[10]/NET0131 ,
		_w4073_,
		_w4084_,
		_w15633_
	);
	LUT2 #(
		.INIT('h8)
	) name11586 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w4873_,
		_w15634_
	);
	LUT4 #(
		.INIT('h2000)
	) name11587 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w4094_,
		_w4097_,
		_w4873_,
		_w15635_
	);
	LUT4 #(
		.INIT('h4000)
	) name11588 (
		\core_c_psq_PCS_reg[10]/NET0131 ,
		_w4073_,
		_w4084_,
		_w15635_,
		_w15636_
	);
	LUT2 #(
		.INIT('he)
	) name11589 (
		_w15633_,
		_w15636_,
		_w15637_
	);
	LUT2 #(
		.INIT('h8)
	) name11590 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w15638_
	);
	LUT4 #(
		.INIT('h20aa)
	) name11591 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15638_,
		_w15639_
	);
	LUT4 #(
		.INIT('h8a00)
	) name11592 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15638_,
		_w15640_
	);
	LUT2 #(
		.INIT('he)
	) name11593 (
		_w15639_,
		_w15640_,
		_w15641_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11594 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8387_,
		_w8807_,
		_w15628_,
		_w15642_
	);
	LUT2 #(
		.INIT('h2)
	) name11595 (
		\regout_STD_C_reg[15]/P0001 ,
		_w15628_,
		_w15643_
	);
	LUT2 #(
		.INIT('he)
	) name11596 (
		_w15642_,
		_w15643_,
		_w15644_
	);
	LUT2 #(
		.INIT('h4)
	) name11597 (
		\core_c_psq_IFC_reg[8]/NET0131 ,
		\core_c_psq_IFC_reg[9]/NET0131 ,
		_w15645_
	);
	LUT4 #(
		.INIT('h7500)
	) name11598 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15645_,
		_w15646_
	);
	LUT4 #(
		.INIT('hff10)
	) name11599 (
		_w7465_,
		_w7565_,
		_w15575_,
		_w15646_,
		_w15647_
	);
	LUT4 #(
		.INIT('h4500)
	) name11600 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w15575_,
		_w15648_
	);
	LUT2 #(
		.INIT('h2)
	) name11601 (
		\core_c_psq_IFC_reg[6]/NET0131 ,
		\core_c_psq_IFC_reg[7]/NET0131 ,
		_w15649_
	);
	LUT4 #(
		.INIT('h7500)
	) name11602 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15649_,
		_w15650_
	);
	LUT2 #(
		.INIT('he)
	) name11603 (
		_w15648_,
		_w15650_,
		_w15651_
	);
	LUT4 #(
		.INIT('h4044)
	) name11604 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTDMOVL_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15652_
	);
	LUT4 #(
		.INIT('hba00)
	) name11605 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w15652_,
		_w15653_
	);
	LUT2 #(
		.INIT('h1)
	) name11606 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		_w15652_,
		_w15654_
	);
	LUT2 #(
		.INIT('h1)
	) name11607 (
		_w15653_,
		_w15654_,
		_w15655_
	);
	LUT4 #(
		.INIT('hba00)
	) name11608 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w15652_,
		_w15656_
	);
	LUT2 #(
		.INIT('h1)
	) name11609 (
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		_w15652_,
		_w15657_
	);
	LUT2 #(
		.INIT('h1)
	) name11610 (
		_w15656_,
		_w15657_,
		_w15658_
	);
	LUT4 #(
		.INIT('hba00)
	) name11611 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w15652_,
		_w15659_
	);
	LUT2 #(
		.INIT('h1)
	) name11612 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		_w15652_,
		_w15660_
	);
	LUT2 #(
		.INIT('h1)
	) name11613 (
		_w15659_,
		_w15660_,
		_w15661_
	);
	LUT4 #(
		.INIT('hba00)
	) name11614 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w15652_,
		_w15662_
	);
	LUT2 #(
		.INIT('h1)
	) name11615 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		_w15652_,
		_w15663_
	);
	LUT2 #(
		.INIT('h1)
	) name11616 (
		_w15662_,
		_w15663_,
		_w15664_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11617 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8725_,
		_w8726_,
		_w8724_,
		_w15665_
	);
	LUT4 #(
		.INIT('h5455)
	) name11618 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w5686_,
		_w5680_,
		_w5756_,
		_w15666_
	);
	LUT4 #(
		.INIT('heee2)
	) name11619 (
		\regout_STD_C_reg[13]/P0001 ,
		_w15628_,
		_w15665_,
		_w15666_,
		_w15667_
	);
	LUT2 #(
		.INIT('h8)
	) name11620 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w9931_,
		_w15668_
	);
	LUT4 #(
		.INIT('hbf00)
	) name11621 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15668_,
		_w15669_
	);
	LUT4 #(
		.INIT('h2000)
	) name11622 (
		\core_c_dec_imm14_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15670_
	);
	LUT2 #(
		.INIT('he)
	) name11623 (
		_w15669_,
		_w15670_,
		_w15671_
	);
	LUT2 #(
		.INIT('h8)
	) name11624 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		_w4106_,
		_w15672_
	);
	LUT2 #(
		.INIT('h8)
	) name11625 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w5046_,
		_w15673_
	);
	LUT3 #(
		.INIT('hec)
	) name11626 (
		_w14570_,
		_w15672_,
		_w15673_,
		_w15674_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11627 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w15584_,
		_w15675_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11628 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w15588_,
		_w15676_
	);
	LUT3 #(
		.INIT('hca)
	) name11629 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001 ,
		_w12673_,
		_w15593_,
		_w15677_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11630 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w15600_,
		_w15678_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11631 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w15600_,
		_w15679_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11632 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w15600_,
		_w15680_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11633 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w15600_,
		_w15681_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11634 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w15584_,
		_w15682_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11635 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w15584_,
		_w15683_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11636 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w15584_,
		_w15684_
	);
	LUT3 #(
		.INIT('hca)
	) name11637 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001 ,
		_w11318_,
		_w15584_,
		_w15685_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11638 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w15584_,
		_w15686_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11639 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w15593_,
		_w15687_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11640 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w15593_,
		_w15688_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11641 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w15593_,
		_w15689_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11642 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w15593_,
		_w15690_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11643 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w15588_,
		_w15691_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11644 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w15588_,
		_w15692_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11645 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w15588_,
		_w15693_
	);
	LUT3 #(
		.INIT('hca)
	) name11646 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001 ,
		_w12673_,
		_w15588_,
		_w15694_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11647 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w15588_,
		_w15695_
	);
	LUT2 #(
		.INIT('h8)
	) name11648 (
		\core_c_dec_RTI_Ed_reg/P0001 ,
		_w4106_,
		_w15696_
	);
	LUT4 #(
		.INIT('h0020)
	) name11649 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w15697_
	);
	LUT4 #(
		.INIT('hf8f0)
	) name11650 (
		_w8174_,
		_w13450_,
		_w15696_,
		_w15697_,
		_w15698_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11651 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w7237_,
		_w9007_,
		_w15628_,
		_w15699_
	);
	LUT2 #(
		.INIT('h2)
	) name11652 (
		\regout_STD_C_reg[9]/P0001 ,
		_w15628_,
		_w15700_
	);
	LUT2 #(
		.INIT('he)
	) name11653 (
		_w15699_,
		_w15700_,
		_w15701_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11654 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8870_,
		_w8871_,
		_w8869_,
		_w15702_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11655 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w6095_,
		_w6171_,
		_w15702_,
		_w15703_
	);
	LUT3 #(
		.INIT('h2e)
	) name11656 (
		\regout_STD_C_reg[3]/P0001 ,
		_w15628_,
		_w15703_,
		_w15704_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11657 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w6359_,
		_w8680_,
		_w15628_,
		_w15705_
	);
	LUT2 #(
		.INIT('h2)
	) name11658 (
		\regout_STD_C_reg[11]/P0001 ,
		_w15628_,
		_w15706_
	);
	LUT2 #(
		.INIT('he)
	) name11659 (
		_w15705_,
		_w15706_,
		_w15707_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11660 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w15593_,
		_w15708_
	);
	LUT2 #(
		.INIT('h4)
	) name11661 (
		\core_c_psq_IFC_reg[10]/NET0131 ,
		\core_c_psq_IFC_reg[11]/NET0131 ,
		_w15709_
	);
	LUT4 #(
		.INIT('h7500)
	) name11662 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15709_,
		_w15710_
	);
	LUT4 #(
		.INIT('hff10)
	) name11663 (
		_w5937_,
		_w6038_,
		_w15575_,
		_w15710_,
		_w15711_
	);
	LUT3 #(
		.INIT('hca)
	) name11664 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001 ,
		_w12673_,
		_w15584_,
		_w15712_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11665 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w15600_,
		_w15713_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11666 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w15593_,
		_w15714_
	);
	LUT4 #(
		.INIT('h4500)
	) name11667 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w15575_,
		_w15715_
	);
	LUT2 #(
		.INIT('h2)
	) name11668 (
		\core_c_psq_IFC_reg[2]/NET0131 ,
		\core_c_psq_IFC_reg[3]/NET0131 ,
		_w15716_
	);
	LUT4 #(
		.INIT('h7500)
	) name11669 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15716_,
		_w15717_
	);
	LUT2 #(
		.INIT('he)
	) name11670 (
		_w15715_,
		_w15717_,
		_w15718_
	);
	LUT4 #(
		.INIT('h4500)
	) name11671 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w15575_,
		_w15719_
	);
	LUT2 #(
		.INIT('h2)
	) name11672 (
		\core_c_psq_IFC_reg[4]/NET0131 ,
		\core_c_psq_IFC_reg[5]/NET0131 ,
		_w15720_
	);
	LUT4 #(
		.INIT('h7500)
	) name11673 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15720_,
		_w15721_
	);
	LUT2 #(
		.INIT('he)
	) name11674 (
		_w15719_,
		_w15721_,
		_w15722_
	);
	LUT3 #(
		.INIT('hca)
	) name11675 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001 ,
		_w11318_,
		_w15593_,
		_w15723_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11676 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8308_,
		_w8767_,
		_w15628_,
		_w15724_
	);
	LUT2 #(
		.INIT('h2)
	) name11677 (
		\regout_STD_C_reg[14]/P0001 ,
		_w15628_,
		_w15725_
	);
	LUT2 #(
		.INIT('he)
	) name11678 (
		_w15724_,
		_w15725_,
		_w15726_
	);
	LUT3 #(
		.INIT('hca)
	) name11679 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001 ,
		_w11318_,
		_w15588_,
		_w15727_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11680 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8826_,
		_w8827_,
		_w8825_,
		_w15728_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11681 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w6815_,
		_w6892_,
		_w15728_,
		_w15729_
	);
	LUT3 #(
		.INIT('h2e)
	) name11682 (
		\regout_STD_C_reg[1]/P0001 ,
		_w15628_,
		_w15729_,
		_w15730_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11683 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w15588_,
		_w15731_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11684 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w15593_,
		_w15732_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11685 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w15584_,
		_w15733_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11686 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w7562_,
		_w8984_,
		_w15628_,
		_w15734_
	);
	LUT2 #(
		.INIT('h2)
	) name11687 (
		\regout_STD_C_reg[8]/P0001 ,
		_w15628_,
		_w15735_
	);
	LUT2 #(
		.INIT('he)
	) name11688 (
		_w15734_,
		_w15735_,
		_w15736_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11689 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8892_,
		_w8893_,
		_w8891_,
		_w15737_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11690 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w7298_,
		_w7373_,
		_w15737_,
		_w15738_
	);
	LUT3 #(
		.INIT('h2e)
	) name11691 (
		\regout_STD_C_reg[4]/P0001 ,
		_w15628_,
		_w15738_,
		_w15739_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11692 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w15600_,
		_w15740_
	);
	LUT3 #(
		.INIT('hca)
	) name11693 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001 ,
		_w12673_,
		_w15600_,
		_w15741_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11694 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8608_,
		_w8610_,
		_w8606_,
		_w15742_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11695 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w5832_,
		_w5909_,
		_w15742_,
		_w15743_
	);
	LUT3 #(
		.INIT('h2e)
	) name11696 (
		\regout_STD_C_reg[0]/P0001 ,
		_w15628_,
		_w15743_,
		_w15744_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11697 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8959_,
		_w8960_,
		_w8958_,
		_w15745_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11698 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w7834_,
		_w7901_,
		_w15745_,
		_w15746_
	);
	LUT3 #(
		.INIT('h2e)
	) name11699 (
		\regout_STD_C_reg[7]/P0001 ,
		_w15628_,
		_w15746_,
		_w15747_
	);
	LUT4 #(
		.INIT('h4500)
	) name11700 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w15575_,
		_w15748_
	);
	LUT2 #(
		.INIT('h2)
	) name11701 (
		\core_c_psq_IFC_reg[0]/NET0131 ,
		\core_c_psq_IFC_reg[1]/NET0131 ,
		_w15749_
	);
	LUT4 #(
		.INIT('h7500)
	) name11702 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15749_,
		_w15750_
	);
	LUT2 #(
		.INIT('he)
	) name11703 (
		_w15748_,
		_w15750_,
		_w15751_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11704 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8702_,
		_w8703_,
		_w8701_,
		_w15752_
	);
	LUT4 #(
		.INIT('h5455)
	) name11705 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w6696_,
		_w6665_,
		_w6754_,
		_w15753_
	);
	LUT4 #(
		.INIT('heee2)
	) name11706 (
		\regout_STD_C_reg[12]/P0001 ,
		_w15628_,
		_w15752_,
		_w15753_,
		_w15754_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11707 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8848_,
		_w8849_,
		_w8847_,
		_w15755_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11708 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w6419_,
		_w6496_,
		_w15755_,
		_w15756_
	);
	LUT3 #(
		.INIT('h2e)
	) name11709 (
		\regout_STD_C_reg[2]/P0001 ,
		_w15628_,
		_w15756_,
		_w15757_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11710 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w15600_,
		_w15758_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11711 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w6035_,
		_w8657_,
		_w15628_,
		_w15759_
	);
	LUT2 #(
		.INIT('h2)
	) name11712 (
		\regout_STD_C_reg[10]/P0001 ,
		_w15628_,
		_w15760_
	);
	LUT2 #(
		.INIT('he)
	) name11713 (
		_w15759_,
		_w15760_,
		_w15761_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11714 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w15588_,
		_w15762_
	);
	LUT2 #(
		.INIT('h2)
	) name11715 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8949_,
		_w15763_
	);
	LUT4 #(
		.INIT('h00ba)
	) name11716 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w7941_,
		_w8038_,
		_w15763_,
		_w15764_
	);
	LUT3 #(
		.INIT('h2e)
	) name11717 (
		\regout_STD_C_reg[6]/P0001 ,
		_w15628_,
		_w15764_,
		_w15765_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11718 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w15584_,
		_w15766_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11719 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w15584_,
		_w15767_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11720 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w15593_,
		_w15768_
	);
	LUT3 #(
		.INIT('hca)
	) name11721 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001 ,
		_w11318_,
		_w15600_,
		_w15769_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11722 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w15588_,
		_w15770_
	);
	LUT4 #(
		.INIT('h2000)
	) name11723 (
		\memc_Pwrite_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15771_
	);
	LUT4 #(
		.INIT('h8000)
	) name11724 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w5045_,
		_w5046_,
		_w15772_
	);
	LUT2 #(
		.INIT('h8)
	) name11725 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w9323_,
		_w15773_
	);
	LUT2 #(
		.INIT('h1)
	) name11726 (
		_w15772_,
		_w15773_,
		_w15774_
	);
	LUT3 #(
		.INIT('hce)
	) name11727 (
		_w8174_,
		_w15771_,
		_w15774_,
		_w15775_
	);
	LUT4 #(
		.INIT('h4500)
	) name11728 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w15575_,
		_w15776_
	);
	LUT2 #(
		.INIT('h4)
	) name11729 (
		\core_c_psq_IFC_reg[6]/NET0131 ,
		\core_c_psq_IFC_reg[7]/NET0131 ,
		_w15777_
	);
	LUT4 #(
		.INIT('h7500)
	) name11730 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15777_,
		_w15778_
	);
	LUT2 #(
		.INIT('he)
	) name11731 (
		_w15776_,
		_w15778_,
		_w15779_
	);
	LUT4 #(
		.INIT('h4500)
	) name11732 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w15575_,
		_w15780_
	);
	LUT2 #(
		.INIT('h4)
	) name11733 (
		\core_c_psq_IFC_reg[4]/NET0131 ,
		\core_c_psq_IFC_reg[5]/NET0131 ,
		_w15781_
	);
	LUT4 #(
		.INIT('h7500)
	) name11734 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15781_,
		_w15782_
	);
	LUT2 #(
		.INIT('he)
	) name11735 (
		_w15780_,
		_w15782_,
		_w15783_
	);
	LUT4 #(
		.INIT('h4500)
	) name11736 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w15575_,
		_w15784_
	);
	LUT2 #(
		.INIT('h4)
	) name11737 (
		\core_c_psq_IFC_reg[2]/NET0131 ,
		\core_c_psq_IFC_reg[3]/NET0131 ,
		_w15785_
	);
	LUT4 #(
		.INIT('h7500)
	) name11738 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15785_,
		_w15786_
	);
	LUT2 #(
		.INIT('he)
	) name11739 (
		_w15784_,
		_w15786_,
		_w15787_
	);
	LUT4 #(
		.INIT('h4500)
	) name11740 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w15575_,
		_w15788_
	);
	LUT2 #(
		.INIT('h4)
	) name11741 (
		\core_c_psq_IFC_reg[0]/NET0131 ,
		\core_c_psq_IFC_reg[1]/NET0131 ,
		_w15789_
	);
	LUT4 #(
		.INIT('h7500)
	) name11742 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15789_,
		_w15790_
	);
	LUT2 #(
		.INIT('he)
	) name11743 (
		_w15788_,
		_w15790_,
		_w15791_
	);
	LUT4 #(
		.INIT('h5111)
	) name11744 (
		\T_TMODE[0]_pad ,
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w14105_,
		_w14106_,
		_w15792_
	);
	LUT2 #(
		.INIT('h1)
	) name11745 (
		_w12802_,
		_w15792_,
		_w15793_
	);
	LUT4 #(
		.INIT('h0302)
	) name11746 (
		\T_TMODE[0]_pad ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TSR_TMP_reg[4]/NET0131 ,
		_w14105_,
		_w15794_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name11747 (
		\tm_TSR_TMP_reg[5]/NET0131 ,
		\tm_TSR_TMP_reg[6]/NET0131 ,
		\tm_TSR_TMP_reg[7]/NET0131 ,
		_w15794_,
		_w15795_
	);
	LUT3 #(
		.INIT('h2e)
	) name11748 (
		\tm_tsr_reg_DO_reg[7]/NET0131 ,
		_w15793_,
		_w15795_,
		_w15796_
	);
	LUT2 #(
		.INIT('h8)
	) name11749 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		_w11300_,
		_w15797_
	);
	LUT3 #(
		.INIT('hca)
	) name11750 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001 ,
		_w12284_,
		_w15797_,
		_w15798_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11751 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w15797_,
		_w15799_
	);
	LUT3 #(
		.INIT('h13)
	) name11752 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001 ,
		_w11300_,
		_w15800_
	);
	LUT2 #(
		.INIT('h1)
	) name11753 (
		_w15799_,
		_w15800_,
		_w15801_
	);
	LUT3 #(
		.INIT('hca)
	) name11754 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001 ,
		_w14918_,
		_w15797_,
		_w15802_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11755 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w15797_,
		_w15803_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11756 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w15797_,
		_w15804_
	);
	LUT3 #(
		.INIT('hca)
	) name11757 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001 ,
		_w14866_,
		_w15797_,
		_w15805_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11758 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w15797_,
		_w15806_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11759 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w15797_,
		_w15807_
	);
	LUT2 #(
		.INIT('h8)
	) name11760 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		_w11300_,
		_w15808_
	);
	LUT3 #(
		.INIT('hca)
	) name11761 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001 ,
		_w14918_,
		_w15808_,
		_w15809_
	);
	LUT3 #(
		.INIT('hca)
	) name11762 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001 ,
		_w11318_,
		_w15797_,
		_w15810_
	);
	LUT2 #(
		.INIT('h8)
	) name11763 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		_w11300_,
		_w15811_
	);
	LUT3 #(
		.INIT('hca)
	) name11764 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001 ,
		_w12284_,
		_w15811_,
		_w15812_
	);
	LUT3 #(
		.INIT('hca)
	) name11765 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001 ,
		_w14918_,
		_w15811_,
		_w15813_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11766 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w15811_,
		_w15814_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11767 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w15811_,
		_w15815_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11768 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w15811_,
		_w15816_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11769 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w15811_,
		_w15817_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11770 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w15811_,
		_w15818_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11771 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w15811_,
		_w15819_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11772 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w15811_,
		_w15820_
	);
	LUT3 #(
		.INIT('hca)
	) name11773 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001 ,
		_w11318_,
		_w15811_,
		_w15821_
	);
	LUT3 #(
		.INIT('hca)
	) name11774 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001 ,
		_w12673_,
		_w15811_,
		_w15822_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11775 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w15811_,
		_w15823_
	);
	LUT3 #(
		.INIT('h13)
	) name11776 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001 ,
		_w11300_,
		_w15824_
	);
	LUT2 #(
		.INIT('h1)
	) name11777 (
		_w15823_,
		_w15824_,
		_w15825_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11778 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w15811_,
		_w15826_
	);
	LUT3 #(
		.INIT('h13)
	) name11779 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001 ,
		_w11300_,
		_w15827_
	);
	LUT2 #(
		.INIT('h1)
	) name11780 (
		_w15826_,
		_w15827_,
		_w15828_
	);
	LUT3 #(
		.INIT('hca)
	) name11781 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001 ,
		_w14866_,
		_w15811_,
		_w15829_
	);
	LUT3 #(
		.INIT('hca)
	) name11782 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001 ,
		_w12486_,
		_w15811_,
		_w15830_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11783 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w15811_,
		_w15831_
	);
	LUT3 #(
		.INIT('hca)
	) name11784 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001 ,
		_w12284_,
		_w15808_,
		_w15832_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11785 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w15808_,
		_w15833_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11786 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001 ,
		_w11626_,
		_w11627_,
		_w15808_,
		_w15834_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11787 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001 ,
		_w12736_,
		_w12737_,
		_w15808_,
		_w15835_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11788 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w15808_,
		_w15836_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11789 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w15808_,
		_w15837_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11790 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001 ,
		_w11313_,
		_w11314_,
		_w15808_,
		_w15838_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11791 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w15808_,
		_w15839_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11792 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w15808_,
		_w15840_
	);
	LUT3 #(
		.INIT('h13)
	) name11793 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001 ,
		_w11300_,
		_w15841_
	);
	LUT2 #(
		.INIT('h1)
	) name11794 (
		_w15840_,
		_w15841_,
		_w15842_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11795 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w15808_,
		_w15843_
	);
	LUT3 #(
		.INIT('h13)
	) name11796 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001 ,
		_w11300_,
		_w15844_
	);
	LUT2 #(
		.INIT('h1)
	) name11797 (
		_w15843_,
		_w15844_,
		_w15845_
	);
	LUT3 #(
		.INIT('hca)
	) name11798 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001 ,
		_w14866_,
		_w15808_,
		_w15846_
	);
	LUT3 #(
		.INIT('hca)
	) name11799 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001 ,
		_w12486_,
		_w15808_,
		_w15847_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11800 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001 ,
		_w12315_,
		_w12316_,
		_w15808_,
		_w15848_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11801 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001 ,
		_w12560_,
		_w12561_,
		_w15797_,
		_w15849_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11802 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001 ,
		_w12626_,
		_w12627_,
		_w15797_,
		_w15850_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11803 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001 ,
		_w13610_,
		_w13611_,
		_w15797_,
		_w15851_
	);
	LUT4 #(
		.INIT('h03aa)
	) name11804 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001 ,
		_w12006_,
		_w12007_,
		_w15797_,
		_w15852_
	);
	LUT3 #(
		.INIT('hca)
	) name11805 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001 ,
		_w12673_,
		_w15797_,
		_w15853_
	);
	LUT4 #(
		.INIT('h1b00)
	) name11806 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w15797_,
		_w15854_
	);
	LUT3 #(
		.INIT('h13)
	) name11807 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001 ,
		_w11300_,
		_w15855_
	);
	LUT2 #(
		.INIT('h1)
	) name11808 (
		_w15854_,
		_w15855_,
		_w15856_
	);
	LUT3 #(
		.INIT('hca)
	) name11809 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001 ,
		_w12486_,
		_w15797_,
		_w15857_
	);
	LUT3 #(
		.INIT('hca)
	) name11810 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001 ,
		_w12673_,
		_w15808_,
		_w15858_
	);
	LUT3 #(
		.INIT('hca)
	) name11811 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001 ,
		_w11318_,
		_w15808_,
		_w15859_
	);
	LUT3 #(
		.INIT('h80)
	) name11812 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15860_
	);
	LUT3 #(
		.INIT('h7f)
	) name11813 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15861_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11814 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[9]/NET0131 ,
		_w15862_
	);
	LUT4 #(
		.INIT('h8000)
	) name11815 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[9]/P0001 ,
		_w15863_
	);
	LUT2 #(
		.INIT('he)
	) name11816 (
		_w15862_,
		_w15863_,
		_w15864_
	);
	LUT3 #(
		.INIT('h80)
	) name11817 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15865_
	);
	LUT3 #(
		.INIT('h7f)
	) name11818 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15866_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11819 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[1]/NET0131 ,
		_w15867_
	);
	LUT4 #(
		.INIT('h8000)
	) name11820 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[1]/P0001 ,
		_w15868_
	);
	LUT2 #(
		.INIT('he)
	) name11821 (
		_w15867_,
		_w15868_,
		_w15869_
	);
	LUT3 #(
		.INIT('h80)
	) name11822 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15870_
	);
	LUT3 #(
		.INIT('h7f)
	) name11823 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15871_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11824 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[11]/NET0131 ,
		_w15872_
	);
	LUT4 #(
		.INIT('h8000)
	) name11825 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[11]/P0001 ,
		_w15873_
	);
	LUT2 #(
		.INIT('he)
	) name11826 (
		_w15872_,
		_w15873_,
		_w15874_
	);
	LUT3 #(
		.INIT('h80)
	) name11827 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15875_
	);
	LUT3 #(
		.INIT('h7f)
	) name11828 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15876_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11829 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[3]/NET0131 ,
		_w15877_
	);
	LUT4 #(
		.INIT('h8000)
	) name11830 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[3]/P0001 ,
		_w15878_
	);
	LUT2 #(
		.INIT('he)
	) name11831 (
		_w15877_,
		_w15878_,
		_w15879_
	);
	LUT3 #(
		.INIT('h80)
	) name11832 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15880_
	);
	LUT3 #(
		.INIT('h7f)
	) name11833 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15881_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11834 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[7]/NET0131 ,
		_w15882_
	);
	LUT4 #(
		.INIT('h8000)
	) name11835 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[7]/P0001 ,
		_w15883_
	);
	LUT2 #(
		.INIT('he)
	) name11836 (
		_w15882_,
		_w15883_,
		_w15884_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11837 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[8]/NET0131 ,
		_w15885_
	);
	LUT4 #(
		.INIT('h8000)
	) name11838 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[8]/P0001 ,
		_w15886_
	);
	LUT2 #(
		.INIT('he)
	) name11839 (
		_w15885_,
		_w15886_,
		_w15887_
	);
	LUT3 #(
		.INIT('h80)
	) name11840 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15888_
	);
	LUT3 #(
		.INIT('h7f)
	) name11841 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w15889_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11842 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[5]/NET0131 ,
		_w15890_
	);
	LUT4 #(
		.INIT('h8000)
	) name11843 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[5]/P0001 ,
		_w15891_
	);
	LUT2 #(
		.INIT('he)
	) name11844 (
		_w15890_,
		_w15891_,
		_w15892_
	);
	LUT3 #(
		.INIT('h20)
	) name11845 (
		PWDACK_pad,
		\clkc_SLEEP_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w15893_
	);
	LUT4 #(
		.INIT('hd2f0)
	) name11846 (
		PWDACK_pad,
		\clkc_SLEEP_reg/NET0131 ,
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w15894_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name11847 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w15895_
	);
	LUT4 #(
		.INIT('h2000)
	) name11848 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w15896_
	);
	LUT2 #(
		.INIT('h1)
	) name11849 (
		_w15895_,
		_w15896_,
		_w15897_
	);
	LUT4 #(
		.INIT('h00bf)
	) name11850 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15897_,
		_w15898_
	);
	LUT4 #(
		.INIT('h2000)
	) name11851 (
		\core_dag_ilm2reg_M_E_reg[1]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15899_
	);
	LUT2 #(
		.INIT('he)
	) name11852 (
		_w15898_,
		_w15899_,
		_w15900_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name11853 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w15901_
	);
	LUT4 #(
		.INIT('h2000)
	) name11854 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w15902_
	);
	LUT2 #(
		.INIT('h1)
	) name11855 (
		_w15901_,
		_w15902_,
		_w15903_
	);
	LUT4 #(
		.INIT('h00bf)
	) name11856 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15903_,
		_w15904_
	);
	LUT4 #(
		.INIT('h2000)
	) name11857 (
		\core_dag_ilm2reg_M_E_reg[0]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15905_
	);
	LUT2 #(
		.INIT('he)
	) name11858 (
		_w15904_,
		_w15905_,
		_w15906_
	);
	LUT2 #(
		.INIT('h4)
	) name11859 (
		_w9332_,
		_w9341_,
		_w15907_
	);
	LUT2 #(
		.INIT('h2)
	) name11860 (
		_w9321_,
		_w9332_,
		_w15908_
	);
	LUT2 #(
		.INIT('h4)
	) name11861 (
		_w9332_,
		_w9339_,
		_w15909_
	);
	LUT4 #(
		.INIT('h0800)
	) name11862 (
		_w9313_,
		_w9319_,
		_w9332_,
		_w9345_,
		_w15910_
	);
	LUT4 #(
		.INIT('h0400)
	) name11863 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[8]/NET0131 ,
		_w15911_
	);
	LUT3 #(
		.INIT('hc8)
	) name11864 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TCR_TMP_reg[8]/NET0131 ,
		_w14107_,
		_w15912_
	);
	LUT4 #(
		.INIT('h2333)
	) name11865 (
		\tm_tpr_reg_DO_reg[8]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w15913_
	);
	LUT4 #(
		.INIT('hfe00)
	) name11866 (
		_w14103_,
		_w14822_,
		_w15912_,
		_w15913_,
		_w15914_
	);
	LUT2 #(
		.INIT('he)
	) name11867 (
		_w15911_,
		_w15914_,
		_w15915_
	);
	LUT4 #(
		.INIT('h0200)
	) name11868 (
		_w6944_,
		_w8187_,
		_w8470_,
		_w8478_,
		_w15916_
	);
	LUT4 #(
		.INIT('h0200)
	) name11869 (
		_w6944_,
		_w8187_,
		_w8470_,
		_w8476_,
		_w15917_
	);
	LUT4 #(
		.INIT('h2000)
	) name11870 (
		_w6944_,
		_w8187_,
		_w8470_,
		_w8478_,
		_w15918_
	);
	LUT4 #(
		.INIT('h2000)
	) name11871 (
		_w6944_,
		_w8187_,
		_w8470_,
		_w8476_,
		_w15919_
	);
	LUT4 #(
		.INIT('h0200)
	) name11872 (
		_w6944_,
		_w8187_,
		_w8470_,
		_w8472_,
		_w15920_
	);
	LUT4 #(
		.INIT('h0020)
	) name11873 (
		_w6944_,
		_w8187_,
		_w8468_,
		_w8470_,
		_w15921_
	);
	LUT4 #(
		.INIT('h2000)
	) name11874 (
		_w6944_,
		_w8187_,
		_w8470_,
		_w8472_,
		_w15922_
	);
	LUT4 #(
		.INIT('h2000)
	) name11875 (
		_w6944_,
		_w8187_,
		_w8468_,
		_w8470_,
		_w15923_
	);
	LUT3 #(
		.INIT('h01)
	) name11876 (
		_w6944_,
		_w8170_,
		_w8187_,
		_w15924_
	);
	LUT4 #(
		.INIT('h0100)
	) name11877 (
		_w9313_,
		_w9319_,
		_w9332_,
		_w9345_,
		_w15925_
	);
	LUT2 #(
		.INIT('h4)
	) name11878 (
		_w9332_,
		_w9343_,
		_w15926_
	);
	LUT4 #(
		.INIT('h0200)
	) name11879 (
		_w9313_,
		_w9319_,
		_w9332_,
		_w9345_,
		_w15927_
	);
	LUT4 #(
		.INIT('h0400)
	) name11880 (
		_w9313_,
		_w9319_,
		_w9332_,
		_w9345_,
		_w15928_
	);
	LUT4 #(
		.INIT('hbf00)
	) name11881 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4967_,
		_w15929_
	);
	LUT4 #(
		.INIT('h2000)
	) name11882 (
		\core_c_dec_Double_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15930_
	);
	LUT3 #(
		.INIT('ha8)
	) name11883 (
		_w4102_,
		_w15929_,
		_w15930_,
		_w15931_
	);
	LUT4 #(
		.INIT('h1000)
	) name11884 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15932_
	);
	LUT4 #(
		.INIT('h4555)
	) name11885 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15933_
	);
	LUT3 #(
		.INIT('h02)
	) name11886 (
		_w4142_,
		_w15933_,
		_w15932_,
		_w15934_
	);
	LUT4 #(
		.INIT('h2000)
	) name11887 (
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15935_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name11888 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15936_
	);
	LUT3 #(
		.INIT('ha8)
	) name11889 (
		_w4142_,
		_w15935_,
		_w15936_,
		_w15937_
	);
	LUT4 #(
		.INIT('h0008)
	) name11890 (
		T_ICE_RSTn_pad,
		T_RSTn_pad,
		\clkc_Awake_reg/NET0131 ,
		\clkc_RSTtext_reg/P0001 ,
		_w15938_
	);
	LUT3 #(
		.INIT('h08)
	) name11891 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_rxctl_a_sync1_reg/P0001 ,
		\sport1_rxctl_a_sync2_reg/P0001 ,
		_w15939_
	);
	LUT3 #(
		.INIT('hae)
	) name11892 (
		_w8171_,
		_w8174_,
		_w8180_,
		_w15940_
	);
	LUT3 #(
		.INIT('hf2)
	) name11893 (
		_w8174_,
		_w9325_,
		_w9330_,
		_w15941_
	);
	LUT4 #(
		.INIT('h7000)
	) name11894 (
		_w14420_,
		_w14421_,
		_w14514_,
		_w14515_,
		_w15942_
	);
	LUT4 #(
		.INIT('h8000)
	) name11895 (
		_w14414_,
		_w14415_,
		_w14520_,
		_w14521_,
		_w15943_
	);
	LUT2 #(
		.INIT('h8)
	) name11896 (
		_w15942_,
		_w15943_,
		_w15944_
	);
	LUT4 #(
		.INIT('h4b00)
	) name11897 (
		_w12121_,
		_w12134_,
		_w12149_,
		_w15944_,
		_w15945_
	);
	LUT4 #(
		.INIT('h0888)
	) name11898 (
		_w14414_,
		_w14415_,
		_w14520_,
		_w14521_,
		_w15946_
	);
	LUT2 #(
		.INIT('h8)
	) name11899 (
		_w15942_,
		_w15946_,
		_w15947_
	);
	LUT4 #(
		.INIT('hb400)
	) name11900 (
		_w12121_,
		_w12134_,
		_w12149_,
		_w15947_,
		_w15948_
	);
	LUT4 #(
		.INIT('h0777)
	) name11901 (
		_w14420_,
		_w14421_,
		_w14514_,
		_w14515_,
		_w15949_
	);
	LUT2 #(
		.INIT('h8)
	) name11902 (
		_w15946_,
		_w15949_,
		_w15950_
	);
	LUT2 #(
		.INIT('h8)
	) name11903 (
		_w15943_,
		_w15949_,
		_w15951_
	);
	LUT4 #(
		.INIT('h8000)
	) name11904 (
		_w14420_,
		_w14421_,
		_w14514_,
		_w14515_,
		_w15952_
	);
	LUT4 #(
		.INIT('h7000)
	) name11905 (
		_w14414_,
		_w14415_,
		_w14520_,
		_w14521_,
		_w15953_
	);
	LUT2 #(
		.INIT('h8)
	) name11906 (
		_w15952_,
		_w15953_,
		_w15954_
	);
	LUT4 #(
		.INIT('h0777)
	) name11907 (
		_w14414_,
		_w14415_,
		_w14520_,
		_w14521_,
		_w15955_
	);
	LUT2 #(
		.INIT('h8)
	) name11908 (
		_w15952_,
		_w15955_,
		_w15956_
	);
	LUT4 #(
		.INIT('h04bf)
	) name11909 (
		_w12164_,
		_w12177_,
		_w15954_,
		_w15956_,
		_w15957_
	);
	LUT4 #(
		.INIT('h2700)
	) name11910 (
		_w12149_,
		_w15951_,
		_w15950_,
		_w15957_,
		_w15958_
	);
	LUT4 #(
		.INIT('h5455)
	) name11911 (
		_w12114_,
		_w15948_,
		_w15945_,
		_w15958_,
		_w15959_
	);
	LUT4 #(
		.INIT('h5554)
	) name11912 (
		_w12185_,
		_w12199_,
		_w12200_,
		_w12198_,
		_w15960_
	);
	LUT3 #(
		.INIT('h08)
	) name11913 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w12112_,
		_w12184_,
		_w15961_
	);
	LUT4 #(
		.INIT('h7000)
	) name11914 (
		_w14414_,
		_w14415_,
		_w14420_,
		_w14421_,
		_w15962_
	);
	LUT2 #(
		.INIT('h4)
	) name11915 (
		_w14516_,
		_w15962_,
		_w15963_
	);
	LUT4 #(
		.INIT('h5600)
	) name11916 (
		_w14522_,
		_w15960_,
		_w15961_,
		_w15963_,
		_w15964_
	);
	LUT4 #(
		.INIT('h4800)
	) name11917 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w14416_,
		_w14522_,
		_w15949_,
		_w15965_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name11918 (
		_w4161_,
		_w14416_,
		_w14522_,
		_w15942_,
		_w15966_
	);
	LUT4 #(
		.INIT('hedff)
	) name11919 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w14416_,
		_w14522_,
		_w15952_,
		_w15967_
	);
	LUT3 #(
		.INIT('h40)
	) name11920 (
		_w15965_,
		_w15966_,
		_w15967_,
		_w15968_
	);
	LUT3 #(
		.INIT('h51)
	) name11921 (
		_w4104_,
		_w12114_,
		_w15968_,
		_w15969_
	);
	LUT2 #(
		.INIT('h4)
	) name11922 (
		_w15964_,
		_w15969_,
		_w15970_
	);
	LUT4 #(
		.INIT('h1000)
	) name11923 (
		\core_eu_ec_cun_termOK_CE_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15971_
	);
	LUT2 #(
		.INIT('h2)
	) name11924 (
		_w4140_,
		_w15971_,
		_w15972_
	);
	LUT3 #(
		.INIT('hb0)
	) name11925 (
		_w15959_,
		_w15970_,
		_w15972_,
		_w15973_
	);
	LUT3 #(
		.INIT('he8)
	) name11926 (
		\T_PIOin[3]_pad ,
		\pio_PIO_IN_P_reg[3]/P0001 ,
		\pio_PIO_RES_reg[3]/NET0131 ,
		_w15974_
	);
	LUT3 #(
		.INIT('he8)
	) name11927 (
		\T_PIOin[1]_pad ,
		\pio_PIO_IN_P_reg[1]/P0001 ,
		\pio_PIO_RES_reg[1]/NET0131 ,
		_w15975_
	);
	LUT3 #(
		.INIT('he8)
	) name11928 (
		\T_PIOin[10]_pad ,
		\pio_PIO_IN_P_reg[10]/P0001 ,
		\pio_PIO_RES_reg[10]/NET0131 ,
		_w15976_
	);
	LUT3 #(
		.INIT('h10)
	) name11929 (
		\core_c_dec_Long_Cg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w15977_
	);
	LUT4 #(
		.INIT('hba00)
	) name11930 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w4102_,
		_w15978_
	);
	LUT2 #(
		.INIT('h4)
	) name11931 (
		_w15977_,
		_w15978_,
		_w15979_
	);
	LUT3 #(
		.INIT('h10)
	) name11932 (
		\auctl_T0Sack_reg/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w15980_
	);
	LUT2 #(
		.INIT('h4)
	) name11933 (
		_w4088_,
		_w15980_,
		_w15981_
	);
	LUT3 #(
		.INIT('h10)
	) name11934 (
		\auctl_R1Sack_reg/NET0131 ,
		_w4088_,
		_w4980_,
		_w15982_
	);
	LUT3 #(
		.INIT('he8)
	) name11935 (
		\T_PIOin[8]_pad ,
		\pio_PIO_IN_P_reg[8]/P0001 ,
		\pio_PIO_RES_reg[8]/NET0131 ,
		_w15983_
	);
	LUT3 #(
		.INIT('he8)
	) name11936 (
		\T_PIOin[5]_pad ,
		\pio_PIO_IN_P_reg[5]/P0001 ,
		\pio_PIO_RES_reg[5]/NET0131 ,
		_w15984_
	);
	LUT3 #(
		.INIT('he8)
	) name11937 (
		\T_PIOin[6]_pad ,
		\pio_PIO_IN_P_reg[6]/P0001 ,
		\pio_PIO_RES_reg[6]/NET0131 ,
		_w15985_
	);
	LUT3 #(
		.INIT('he8)
	) name11938 (
		\T_PIOin[11]_pad ,
		\pio_PIO_IN_P_reg[11]/P0001 ,
		\pio_PIO_RES_reg[11]/NET0131 ,
		_w15986_
	);
	LUT3 #(
		.INIT('h10)
	) name11939 (
		\auctl_R0Sack_reg/NET0131 ,
		_w4088_,
		_w4984_,
		_w15987_
	);
	LUT2 #(
		.INIT('h4)
	) name11940 (
		\auctl_T1Sack_reg/NET0131 ,
		_w4982_,
		_w15988_
	);
	LUT2 #(
		.INIT('h4)
	) name11941 (
		_w4088_,
		_w15988_,
		_w15989_
	);
	LUT4 #(
		.INIT('h0400)
	) name11942 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[15]/NET0131 ,
		_w15990_
	);
	LUT4 #(
		.INIT('h1333)
	) name11943 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		\tm_TCR_TMP_reg[11]/NET0131 ,
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w14110_,
		_w15991_
	);
	LUT2 #(
		.INIT('h8)
	) name11944 (
		_w14115_,
		_w15991_,
		_w15992_
	);
	LUT4 #(
		.INIT('h8000)
	) name11945 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		\tm_TCR_TMP_reg[11]/NET0131 ,
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w14110_,
		_w15993_
	);
	LUT3 #(
		.INIT('h45)
	) name11946 (
		\T_TMODE[0]_pad ,
		_w14114_,
		_w15993_,
		_w15994_
	);
	LUT3 #(
		.INIT('h8a)
	) name11947 (
		_w14108_,
		_w15992_,
		_w15994_,
		_w15995_
	);
	LUT4 #(
		.INIT('h4044)
	) name11948 (
		\tm_TCR_TMP_reg[12]/NET0131 ,
		_w14108_,
		_w15992_,
		_w15994_,
		_w15996_
	);
	LUT4 #(
		.INIT('he1f0)
	) name11949 (
		\tm_TCR_TMP_reg[13]/NET0131 ,
		\tm_TCR_TMP_reg[14]/NET0131 ,
		\tm_TCR_TMP_reg[15]/NET0131 ,
		_w15996_,
		_w15997_
	);
	LUT4 #(
		.INIT('h2333)
	) name11950 (
		\tm_tpr_reg_DO_reg[15]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w15998_
	);
	LUT4 #(
		.INIT('hfecc)
	) name11951 (
		_w14103_,
		_w15990_,
		_w15997_,
		_w15998_,
		_w15999_
	);
	LUT2 #(
		.INIT('hb)
	) name11952 (
		\T_TMODE[1]_pad ,
		\core_c_dec_PPclr_reg/P0001 ,
		_w16000_
	);
	LUT4 #(
		.INIT('h2000)
	) name11953 (
		\core_eu_ec_cun_COND_E_reg[2]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16001_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name11954 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16002_
	);
	LUT3 #(
		.INIT('ha8)
	) name11955 (
		_w4142_,
		_w16001_,
		_w16002_,
		_w16003_
	);
	LUT3 #(
		.INIT('he8)
	) name11956 (
		\T_PIOin[4]_pad ,
		\pio_PIO_IN_P_reg[4]/P0001 ,
		\pio_PIO_RES_reg[4]/NET0131 ,
		_w16004_
	);
	LUT3 #(
		.INIT('he8)
	) name11957 (
		\T_PIOin[7]_pad ,
		\pio_PIO_IN_P_reg[7]/P0001 ,
		\pio_PIO_RES_reg[7]/NET0131 ,
		_w16005_
	);
	LUT4 #(
		.INIT('h2000)
	) name11958 (
		\core_eu_ec_cun_COND_E_reg[3]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16006_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name11959 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16007_
	);
	LUT3 #(
		.INIT('ha8)
	) name11960 (
		_w4142_,
		_w16006_,
		_w16007_,
		_w16008_
	);
	LUT3 #(
		.INIT('he8)
	) name11961 (
		\T_PIOin[9]_pad ,
		\pio_PIO_IN_P_reg[9]/P0001 ,
		\pio_PIO_RES_reg[9]/NET0131 ,
		_w16009_
	);
	LUT3 #(
		.INIT('h2a)
	) name11962 (
		_w11713_,
		_w11736_,
		_w14468_,
		_w16010_
	);
	LUT3 #(
		.INIT('h08)
	) name11963 (
		_w11726_,
		_w14472_,
		_w14477_,
		_w16011_
	);
	LUT4 #(
		.INIT('hcf80)
	) name11964 (
		_w11721_,
		_w11725_,
		_w14472_,
		_w14531_,
		_w16012_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name11965 (
		_w11725_,
		_w14489_,
		_w14484_,
		_w14472_,
		_w16013_
	);
	LUT3 #(
		.INIT('h23)
	) name11966 (
		_w11721_,
		_w14483_,
		_w14484_,
		_w16014_
	);
	LUT4 #(
		.INIT('h4f00)
	) name11967 (
		_w16011_,
		_w16012_,
		_w16013_,
		_w16014_,
		_w16015_
	);
	LUT3 #(
		.INIT('hb3)
	) name11968 (
		_w11710_,
		_w11713_,
		_w11718_,
		_w16016_
	);
	LUT3 #(
		.INIT('hb0)
	) name11969 (
		_w11725_,
		_w14483_,
		_w16016_,
		_w16017_
	);
	LUT4 #(
		.INIT('h0400)
	) name11970 (
		_w11698_,
		_w11705_,
		_w11709_,
		_w11733_,
		_w16018_
	);
	LUT4 #(
		.INIT('h0800)
	) name11971 (
		_w11710_,
		_w11713_,
		_w11718_,
		_w11729_,
		_w16019_
	);
	LUT2 #(
		.INIT('h1)
	) name11972 (
		_w16018_,
		_w16019_,
		_w16020_
	);
	LUT4 #(
		.INIT('h20aa)
	) name11973 (
		_w16010_,
		_w16015_,
		_w16017_,
		_w16020_,
		_w16021_
	);
	LUT2 #(
		.INIT('h4)
	) name11974 (
		_w11713_,
		_w11718_,
		_w16022_
	);
	LUT4 #(
		.INIT('h00f7)
	) name11975 (
		_w11736_,
		_w14468_,
		_w14477_,
		_w16022_,
		_w16023_
	);
	LUT4 #(
		.INIT('h0004)
	) name11976 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[2]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w16024_
	);
	LUT4 #(
		.INIT('h4500)
	) name11977 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13382_,
		_w16025_
	);
	LUT2 #(
		.INIT('h1)
	) name11978 (
		_w16024_,
		_w16025_,
		_w16026_
	);
	LUT4 #(
		.INIT('h8aff)
	) name11979 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w16021_,
		_w16023_,
		_w16026_,
		_w16027_
	);
	LUT3 #(
		.INIT('he8)
	) name11980 (
		\T_PIOin[2]_pad ,
		\pio_PIO_IN_P_reg[2]/P0001 ,
		\pio_PIO_RES_reg[2]/NET0131 ,
		_w16028_
	);
	LUT3 #(
		.INIT('h80)
	) name11981 (
		\T_TMODE[1]_pad ,
		_w4787_,
		_w12703_,
		_w16029_
	);
	LUT3 #(
		.INIT('h7f)
	) name11982 (
		\T_TMODE[1]_pad ,
		_w4787_,
		_w12703_,
		_w16030_
	);
	LUT3 #(
		.INIT('h80)
	) name11983 (
		\T_TMODE[1]_pad ,
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w16031_
	);
	LUT3 #(
		.INIT('h2a)
	) name11984 (
		\emc_ECMcs_reg/NET0131 ,
		_w4793_,
		_w16031_,
		_w16032_
	);
	LUT4 #(
		.INIT('hff80)
	) name11985 (
		\T_TMODE[1]_pad ,
		_w4787_,
		_w12703_,
		_w16032_,
		_w16033_
	);
	LUT3 #(
		.INIT('he8)
	) name11986 (
		\T_PIOin[0]_pad ,
		\pio_PIO_IN_P_reg[0]/P0001 ,
		\pio_PIO_RES_reg[0]/NET0131 ,
		_w16034_
	);
	LUT3 #(
		.INIT('h80)
	) name11987 (
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		_w4073_,
		_w4084_,
		_w16035_
	);
	LUT3 #(
		.INIT('h2a)
	) name11988 (
		\core_c_psq_Eqend_D_reg/P0001 ,
		_w4073_,
		_w4084_,
		_w16036_
	);
	LUT4 #(
		.INIT('h1000)
	) name11989 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4428_,
		_w8172_,
		_w16036_,
		_w16037_
	);
	LUT3 #(
		.INIT('ha8)
	) name11990 (
		_w4102_,
		_w16035_,
		_w16037_,
		_w16038_
	);
	LUT4 #(
		.INIT('hd98c)
	) name11991 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w16039_
	);
	LUT3 #(
		.INIT('h70)
	) name11992 (
		_w11726_,
		_w14472_,
		_w16039_,
		_w16040_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name11993 (
		_w11721_,
		_w11725_,
		_w14472_,
		_w14527_,
		_w16041_
	);
	LUT4 #(
		.INIT('h2333)
	) name11994 (
		_w11725_,
		_w14484_,
		_w14472_,
		_w14530_,
		_w16042_
	);
	LUT3 #(
		.INIT('h51)
	) name11995 (
		_w14483_,
		_w14484_,
		_w14476_,
		_w16043_
	);
	LUT4 #(
		.INIT('h4f00)
	) name11996 (
		_w16040_,
		_w16041_,
		_w16042_,
		_w16043_,
		_w16044_
	);
	LUT3 #(
		.INIT('h2a)
	) name11997 (
		_w11706_,
		_w14479_,
		_w14483_,
		_w16045_
	);
	LUT4 #(
		.INIT('h0400)
	) name11998 (
		_w11698_,
		_w11705_,
		_w11709_,
		_w11724_,
		_w16046_
	);
	LUT4 #(
		.INIT('h0008)
	) name11999 (
		_w11710_,
		_w11713_,
		_w11718_,
		_w11721_,
		_w16047_
	);
	LUT2 #(
		.INIT('h1)
	) name12000 (
		_w16046_,
		_w16047_,
		_w16048_
	);
	LUT4 #(
		.INIT('h7500)
	) name12001 (
		_w16016_,
		_w16044_,
		_w16045_,
		_w16048_,
		_w16049_
	);
	LUT2 #(
		.INIT('h4)
	) name12002 (
		_w11713_,
		_w11729_,
		_w16050_
	);
	LUT4 #(
		.INIT('h00f7)
	) name12003 (
		_w11736_,
		_w14468_,
		_w14528_,
		_w16050_,
		_w16051_
	);
	LUT4 #(
		.INIT('h08aa)
	) name12004 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w16010_,
		_w16049_,
		_w16051_,
		_w16052_
	);
	LUT4 #(
		.INIT('h0004)
	) name12005 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w16053_
	);
	LUT4 #(
		.INIT('h4500)
	) name12006 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13382_,
		_w16054_
	);
	LUT2 #(
		.INIT('h1)
	) name12007 (
		_w16053_,
		_w16054_,
		_w16055_
	);
	LUT2 #(
		.INIT('hb)
	) name12008 (
		_w16052_,
		_w16055_,
		_w16056_
	);
	LUT2 #(
		.INIT('h2)
	) name12009 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w16057_
	);
	LUT3 #(
		.INIT('h20)
	) name12010 (
		PWDACK_pad,
		\clkc_Awake_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w16058_
	);
	LUT4 #(
		.INIT('hff40)
	) name12011 (
		_w4099_,
		_w4100_,
		_w16057_,
		_w16058_,
		_w16059_
	);
	LUT4 #(
		.INIT('h4044)
	) name12012 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTLreg_E_reg[4]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16060_
	);
	LUT4 #(
		.INIT('h4044)
	) name12013 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTLreg_E_reg[5]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16061_
	);
	LUT4 #(
		.INIT('h2000)
	) name12014 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16062_
	);
	LUT3 #(
		.INIT('hf4)
	) name12015 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w4942_,
		_w16062_,
		_w16063_
	);
	LUT4 #(
		.INIT('h4044)
	) name12016 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTLreg_E_reg[7]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16064_
	);
	LUT4 #(
		.INIT('h0400)
	) name12017 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_Dwrite_C_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16065_
	);
	LUT2 #(
		.INIT('he)
	) name12018 (
		_w9430_,
		_w16065_,
		_w16066_
	);
	LUT4 #(
		.INIT('hff08)
	) name12019 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_txctl_SP_EN_D1_reg/P0001 ,
		\sport1_txctl_TSreqi_reg/NET0131 ,
		_w16067_
	);
	LUT4 #(
		.INIT('h4044)
	) name12020 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTLreg_E_reg[6]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16068_
	);
	LUT4 #(
		.INIT('hff08)
	) name12021 (
		\memc_usysr_DO_reg[12]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_txctl_SP_EN_D1_reg/P0001 ,
		\sport0_txctl_TSreqi_reg/NET0131 ,
		_w16069_
	);
	LUT3 #(
		.INIT('h34)
	) name12022 (
		IACKn_pad,
		\sice_RCS_reg[0]/NET0131 ,
		\sice_RCS_reg[1]/NET0131 ,
		_w16070_
	);
	LUT4 #(
		.INIT('h4044)
	) name12023 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTLreg_E_reg[2]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16071_
	);
	LUT4 #(
		.INIT('h4044)
	) name12024 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTLreg_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16072_
	);
	LUT4 #(
		.INIT('h4044)
	) name12025 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTLreg_E_reg[0]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16073_
	);
	LUT4 #(
		.INIT('h4044)
	) name12026 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTLreg_E_reg[3]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16074_
	);
	LUT4 #(
		.INIT('hc444)
	) name12027 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		_w4073_,
		_w4084_,
		_w16075_
	);
	LUT2 #(
		.INIT('h2)
	) name12028 (
		\core_c_psq_Iflag_reg[10]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w16076_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12029 (
		\core_c_psq_INT_en_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16076_,
		_w16077_
	);
	LUT2 #(
		.INIT('he)
	) name12030 (
		_w16075_,
		_w16077_,
		_w16078_
	);
	LUT2 #(
		.INIT('h8)
	) name12031 (
		\clkc_SLEEP_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w16079_
	);
	LUT4 #(
		.INIT('hff40)
	) name12032 (
		_w4099_,
		_w4100_,
		_w16057_,
		_w16079_,
		_w16080_
	);
	LUT4 #(
		.INIT('ha802)
	) name12033 (
		_w9455_,
		_w9456_,
		_w9570_,
		_w9852_,
		_w16081_
	);
	LUT4 #(
		.INIT('h00eb)
	) name12034 (
		_w9455_,
		_w9862_,
		_w9865_,
		_w16081_,
		_w16082_
	);
	LUT3 #(
		.INIT('h2e)
	) name12035 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001 ,
		_w9895_,
		_w16082_,
		_w16083_
	);
	LUT3 #(
		.INIT('h8a)
	) name12036 (
		\core_c_dec_MTICNTL_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16084_
	);
	LUT4 #(
		.INIT('hba00)
	) name12037 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w16084_,
		_w16085_
	);
	LUT4 #(
		.INIT('h1311)
	) name12038 (
		\core_c_dec_MTICNTL_Eg_reg/P0001 ,
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16086_
	);
	LUT2 #(
		.INIT('h1)
	) name12039 (
		_w16085_,
		_w16086_,
		_w16087_
	);
	LUT4 #(
		.INIT('hba00)
	) name12040 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w16084_,
		_w16088_
	);
	LUT4 #(
		.INIT('h1311)
	) name12041 (
		\core_c_dec_MTICNTL_Eg_reg/P0001 ,
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16089_
	);
	LUT2 #(
		.INIT('h1)
	) name12042 (
		_w16088_,
		_w16089_,
		_w16090_
	);
	LUT3 #(
		.INIT('h2e)
	) name12043 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001 ,
		_w9454_,
		_w16082_,
		_w16091_
	);
	LUT3 #(
		.INIT('h20)
	) name12044 (
		\memc_STI_Cg_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16092_
	);
	LUT2 #(
		.INIT('h1)
	) name12045 (
		_w5056_,
		_w9061_,
		_w16093_
	);
	LUT4 #(
		.INIT('h0045)
	) name12046 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16093_,
		_w16094_
	);
	LUT2 #(
		.INIT('he)
	) name12047 (
		_w16092_,
		_w16094_,
		_w16095_
	);
	LUT3 #(
		.INIT('h13)
	) name12048 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 ,
		_w9894_,
		_w16096_
	);
	LUT4 #(
		.INIT('h0002)
	) name12049 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w16096_,
		_w16097_
	);
	LUT4 #(
		.INIT('h5700)
	) name12050 (
		_w12282_,
		_w12736_,
		_w12737_,
		_w16097_,
		_w16098_
	);
	LUT4 #(
		.INIT('h313b)
	) name12051 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 ,
		_w11308_,
		_w11635_,
		_w16099_
	);
	LUT3 #(
		.INIT('h45)
	) name12052 (
		_w11624_,
		_w16098_,
		_w16099_,
		_w16100_
	);
	LUT4 #(
		.INIT('h0a0e)
	) name12053 (
		_w11174_,
		_w11243_,
		_w11233_,
		_w12245_,
		_w16101_
	);
	LUT2 #(
		.INIT('h6)
	) name12054 (
		_w11080_,
		_w11145_,
		_w16102_
	);
	LUT3 #(
		.INIT('h41)
	) name12055 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16101_,
		_w16102_,
		_w16103_
	);
	LUT3 #(
		.INIT('h82)
	) name12056 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14407_,
		_w14560_,
		_w16104_
	);
	LUT4 #(
		.INIT('heeec)
	) name12057 (
		_w11624_,
		_w16100_,
		_w16103_,
		_w16104_,
		_w16105_
	);
	LUT3 #(
		.INIT('h63)
	) name12058 (
		\tm_TSR_TMP_reg[5]/NET0131 ,
		\tm_TSR_TMP_reg[6]/NET0131 ,
		_w15794_,
		_w16106_
	);
	LUT3 #(
		.INIT('h2e)
	) name12059 (
		\tm_tsr_reg_DO_reg[6]/NET0131 ,
		_w15793_,
		_w16106_,
		_w16107_
	);
	LUT3 #(
		.INIT('h8a)
	) name12060 (
		\memc_Pwrite_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16108_
	);
	LUT4 #(
		.INIT('h0400)
	) name12061 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\memc_Pwrite_C_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16109_
	);
	LUT2 #(
		.INIT('he)
	) name12062 (
		_w16108_,
		_w16109_,
		_w16110_
	);
	LUT3 #(
		.INIT('h08)
	) name12063 (
		\clkc_STBY_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_c_psq_TRAP_R_L_reg/NET0131 ,
		_w16111_
	);
	LUT2 #(
		.INIT('h1)
	) name12064 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w16112_
	);
	LUT4 #(
		.INIT('hf4f0)
	) name12065 (
		_w4099_,
		_w4100_,
		_w16111_,
		_w16112_,
		_w16113_
	);
	LUT2 #(
		.INIT('h2)
	) name12066 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001 ,
		_w11310_,
		_w16114_
	);
	LUT3 #(
		.INIT('h01)
	) name12067 (
		_w9946_,
		_w12442_,
		_w16114_,
		_w16115_
	);
	LUT4 #(
		.INIT('hfd00)
	) name12068 (
		_w12440_,
		_w12736_,
		_w12737_,
		_w16115_,
		_w16116_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12069 (
		_w9946_,
		_w16103_,
		_w16104_,
		_w16116_,
		_w16117_
	);
	LUT2 #(
		.INIT('h6)
	) name12070 (
		\sice_IIRC_reg[0]/NET0131 ,
		\sice_IIRC_reg[1]/NET0131 ,
		_w16118_
	);
	LUT2 #(
		.INIT('h6)
	) name12071 (
		\sice_ICYC_reg[0]/NET0131 ,
		\sice_ICYC_reg[1]/NET0131 ,
		_w16119_
	);
	LUT2 #(
		.INIT('h6)
	) name12072 (
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[1]/NET0131 ,
		_w16120_
	);
	LUT4 #(
		.INIT('heee2)
	) name12073 (
		\core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001 ,
		_w13091_,
		_w16103_,
		_w16104_,
		_w16121_
	);
	LUT3 #(
		.INIT('h10)
	) name12074 (
		_w8798_,
		_w8801_,
		_w15575_,
		_w16122_
	);
	LUT2 #(
		.INIT('h8)
	) name12075 (
		_w12054_,
		_w15634_,
		_w16123_
	);
	LUT2 #(
		.INIT('h8)
	) name12076 (
		_w4749_,
		_w4778_,
		_w16124_
	);
	LUT3 #(
		.INIT('h10)
	) name12077 (
		_w8757_,
		_w8760_,
		_w15575_,
		_w16125_
	);
	LUT2 #(
		.INIT('h1)
	) name12078 (
		\clkc_SIDLE_s2_reg/NET0131 ,
		\clkc_STBY_reg/NET0131 ,
		_w16126_
	);
	LUT3 #(
		.INIT('h04)
	) name12079 (
		_w8486_,
		_w8488_,
		_w16126_,
		_w16127_
	);
	LUT4 #(
		.INIT('heee2)
	) name12080 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001 ,
		_w13168_,
		_w16103_,
		_w16104_,
		_w16128_
	);
	LUT4 #(
		.INIT('h4044)
	) name12081 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMreg_E_reg[6]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16129_
	);
	LUT4 #(
		.INIT('h4044)
	) name12082 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMreg_E_reg[5]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16130_
	);
	LUT4 #(
		.INIT('h0400)
	) name12083 (
		\auctl_DSack_reg/NET0131 ,
		\idma_DSreq_reg/NET0131 ,
		_w4061_,
		_w4062_,
		_w16131_
	);
	LUT4 #(
		.INIT('hbf00)
	) name12084 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4067_,
		_w4088_,
		_w16131_,
		_w16132_
	);
	LUT3 #(
		.INIT('h04)
	) name12085 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w16133_
	);
	LUT2 #(
		.INIT('h8)
	) name12086 (
		_w5760_,
		_w15575_,
		_w16134_
	);
	LUT4 #(
		.INIT('h1500)
	) name12087 (
		\auctl_BSack_reg/NET0131 ,
		_w4067_,
		_w4088_,
		_w4519_,
		_w16135_
	);
	LUT2 #(
		.INIT('he)
	) name12088 (
		\auctl_DSack_reg/NET0131 ,
		\auctl_RST_reg/P0001 ,
		_w16136_
	);
	LUT3 #(
		.INIT('h80)
	) name12089 (
		\clkc_DSPoff_reg/NET0131 ,
		\clkc_SLEEP_reg/NET0131 ,
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w16137_
	);
	LUT2 #(
		.INIT('h8)
	) name12090 (
		_w6758_,
		_w15575_,
		_w16138_
	);
	LUT4 #(
		.INIT('h3b33)
	) name12091 (
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4140_,
		_w8484_,
		_w8490_,
		_w16139_
	);
	LUT4 #(
		.INIT('h4044)
	) name12092 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMreg_E_reg[7]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16140_
	);
	LUT4 #(
		.INIT('h4044)
	) name12093 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMreg_E_reg[4]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16141_
	);
	LUT4 #(
		.INIT('h4044)
	) name12094 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMreg_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16142_
	);
	LUT4 #(
		.INIT('h4044)
	) name12095 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMreg_E_reg[3]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16143_
	);
	LUT2 #(
		.INIT('h1)
	) name12096 (
		\auctl_BSack_reg/NET0131 ,
		\auctl_RST_reg/P0001 ,
		_w16144_
	);
	LUT4 #(
		.INIT('h4044)
	) name12097 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMreg_E_reg[2]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16145_
	);
	LUT4 #(
		.INIT('h4044)
	) name12098 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMreg_E_reg[0]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16146_
	);
	LUT3 #(
		.INIT('ha8)
	) name12099 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[4]/NET0131 ,
		_w16147_
	);
	LUT3 #(
		.INIT('hb0)
	) name12100 (
		\clkc_SIDLE_s1_reg/NET0131 ,
		\clkc_SIDLE_s2_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w16148_
	);
	LUT3 #(
		.INIT('h1f)
	) name12101 (
		T_BMODE_pad,
		T_MMAP_pad,
		\bdma_RST_pin_reg/P0001 ,
		_w16149_
	);
	LUT4 #(
		.INIT('h2000)
	) name12102 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16150_
	);
	LUT2 #(
		.INIT('he)
	) name12103 (
		_w16007_,
		_w16150_,
		_w16151_
	);
	LUT3 #(
		.INIT('hd0)
	) name12104 (
		T_BMODE_pad,
		T_MMAP_pad,
		\bdma_RST_pin_reg/P0001 ,
		_w16152_
	);
	LUT3 #(
		.INIT('h20)
	) name12105 (
		T_BMODE_pad,
		T_MMAP_pad,
		\bdma_RST_pin_reg/P0001 ,
		_w16153_
	);
	LUT4 #(
		.INIT('h2000)
	) name12106 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16154_
	);
	LUT2 #(
		.INIT('he)
	) name12107 (
		_w16002_,
		_w16154_,
		_w16155_
	);
	LUT4 #(
		.INIT('h5545)
	) name12108 (
		\bdma_BDMAmode_reg/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w16156_
	);
	LUT2 #(
		.INIT('hd)
	) name12109 (
		_w4140_,
		_w16156_,
		_w16157_
	);
	LUT4 #(
		.INIT('h1000)
	) name12110 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16158_
	);
	LUT2 #(
		.INIT('h1)
	) name12111 (
		_w8174_,
		_w16158_,
		_w16159_
	);
	LUT3 #(
		.INIT('he4)
	) name12112 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		_w16160_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12113 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16161_
	);
	LUT4 #(
		.INIT('h2000)
	) name12114 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16162_
	);
	LUT2 #(
		.INIT('he)
	) name12115 (
		_w16161_,
		_w16162_,
		_w16163_
	);
	LUT4 #(
		.INIT('h2000)
	) name12116 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16164_
	);
	LUT2 #(
		.INIT('he)
	) name12117 (
		_w15936_,
		_w16164_,
		_w16165_
	);
	LUT3 #(
		.INIT('he4)
	) name12118 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		_w16166_
	);
	LUT3 #(
		.INIT('he4)
	) name12119 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		_w16167_
	);
	LUT3 #(
		.INIT('he4)
	) name12120 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		_w16168_
	);
	LUT3 #(
		.INIT('he4)
	) name12121 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		_w16169_
	);
	LUT3 #(
		.INIT('h8a)
	) name12122 (
		\tm_tsr_reg_DO_reg[8]/NET0131 ,
		_w8486_,
		_w8488_,
		_w16170_
	);
	LUT4 #(
		.INIT('h00ba)
	) name12123 (
		\tm_tsr_reg_DO_reg[8]/NET0131 ,
		_w8484_,
		_w8490_,
		_w16170_,
		_w16171_
	);
	LUT3 #(
		.INIT('h74)
	) name12124 (
		\clkc_Cnt4096_reg/NET0131 ,
		\clkc_DSPoff_reg/NET0131 ,
		\clkc_SLEEP_reg/NET0131 ,
		_w16172_
	);
	LUT3 #(
		.INIT('hca)
	) name12125 (
		\sport1_txctl_TXSHT_reg[13]/P0001 ,
		\sport1_txctl_TX_reg[14]/P0001 ,
		_w14269_,
		_w16173_
	);
	LUT3 #(
		.INIT('h80)
	) name12126 (
		_w4073_,
		_w4084_,
		_w4102_,
		_w16174_
	);
	LUT4 #(
		.INIT('haacf)
	) name12127 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w4809_,
		_w4817_,
		_w16174_,
		_w16175_
	);
	LUT4 #(
		.INIT('haacf)
	) name12128 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w4703_,
		_w4709_,
		_w16174_,
		_w16176_
	);
	LUT4 #(
		.INIT('haacf)
	) name12129 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w4658_,
		_w4664_,
		_w16174_,
		_w16177_
	);
	LUT4 #(
		.INIT('haacf)
	) name12130 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w4640_,
		_w4649_,
		_w16174_,
		_w16178_
	);
	LUT4 #(
		.INIT('haacf)
	) name12131 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w4577_,
		_w4591_,
		_w16174_,
		_w16179_
	);
	LUT4 #(
		.INIT('haacf)
	) name12132 (
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w4562_,
		_w4568_,
		_w16174_,
		_w16180_
	);
	LUT4 #(
		.INIT('haacf)
	) name12133 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w4547_,
		_w4553_,
		_w16174_,
		_w16181_
	);
	LUT4 #(
		.INIT('haacf)
	) name12134 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w4503_,
		_w4515_,
		_w16174_,
		_w16182_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12135 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		\core_c_psq_EXA_reg[7]/P0001 ,
		_w4073_,
		_w4084_,
		_w16183_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12136 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		\core_c_psq_EXA_reg[6]/P0001 ,
		_w4073_,
		_w4084_,
		_w16184_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12137 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		\core_c_psq_EXA_reg[3]/P0001 ,
		_w4073_,
		_w4084_,
		_w16185_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12138 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		\core_c_psq_EXA_reg[2]/P0001 ,
		_w4073_,
		_w4084_,
		_w16186_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12139 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		\core_c_psq_EXA_reg[13]/P0001 ,
		_w4073_,
		_w4084_,
		_w16187_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12140 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		\core_c_psq_EXA_reg[12]/P0001 ,
		_w4073_,
		_w4084_,
		_w16188_
	);
	LUT4 #(
		.INIT('h2000)
	) name12141 (
		\core_c_dec_accCM_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16189_
	);
	LUT2 #(
		.INIT('he)
	) name12142 (
		_w4942_,
		_w16189_,
		_w16190_
	);
	LUT4 #(
		.INIT('haacf)
	) name12143 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w4600_,
		_w4612_,
		_w16174_,
		_w16191_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12144 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		\core_c_psq_EXA_reg[0]/P0001 ,
		_w4073_,
		_w4084_,
		_w16192_
	);
	LUT3 #(
		.INIT('hac)
	) name12145 (
		\core_c_dec_Prderr_Cg_reg/NET0131 ,
		_w4428_,
		_w4971_,
		_w16193_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12146 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		\core_c_psq_EXA_reg[9]/P0001 ,
		_w4073_,
		_w4084_,
		_w16194_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12147 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16195_
	);
	LUT4 #(
		.INIT('h2000)
	) name12148 (
		\core_c_dec_IRE_reg[18]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16196_
	);
	LUT2 #(
		.INIT('he)
	) name12149 (
		_w16195_,
		_w16196_,
		_w16197_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12150 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16198_
	);
	LUT4 #(
		.INIT('h2000)
	) name12151 (
		\core_c_dec_IRE_reg[19]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16199_
	);
	LUT2 #(
		.INIT('he)
	) name12152 (
		_w16198_,
		_w16199_,
		_w16200_
	);
	LUT4 #(
		.INIT('haacf)
	) name12153 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w4673_,
		_w4679_,
		_w16174_,
		_w16201_
	);
	LUT3 #(
		.INIT('hca)
	) name12154 (
		\sport1_txctl_TXSHT_reg[14]/P0001 ,
		\sport1_txctl_TX_reg[15]/P0001 ,
		_w14269_,
		_w16202_
	);
	LUT4 #(
		.INIT('h00bf)
	) name12155 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w5031_,
		_w16203_
	);
	LUT4 #(
		.INIT('h2000)
	) name12156 (
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16204_
	);
	LUT2 #(
		.INIT('he)
	) name12157 (
		_w16203_,
		_w16204_,
		_w16205_
	);
	LUT4 #(
		.INIT('h00bf)
	) name12158 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w5032_,
		_w16206_
	);
	LUT4 #(
		.INIT('h2000)
	) name12159 (
		\core_dag_ilm2reg_IL_E_reg[0]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w16207_
	);
	LUT2 #(
		.INIT('he)
	) name12160 (
		_w16206_,
		_w16207_,
		_w16208_
	);
	LUT4 #(
		.INIT('h0015)
	) name12161 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4992_,
		_w16209_
	);
	LUT4 #(
		.INIT('ha888)
	) name12162 (
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w4064_,
		_w4067_,
		_w4088_,
		_w16210_
	);
	LUT2 #(
		.INIT('he)
	) name12163 (
		_w16209_,
		_w16210_,
		_w16211_
	);
	LUT4 #(
		.INIT('h0015)
	) name12164 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4987_,
		_w16212_
	);
	LUT4 #(
		.INIT('ha888)
	) name12165 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4064_,
		_w4067_,
		_w4088_,
		_w16213_
	);
	LUT2 #(
		.INIT('he)
	) name12166 (
		_w16212_,
		_w16213_,
		_w16214_
	);
	LUT4 #(
		.INIT('h0015)
	) name12167 (
		_w4064_,
		_w4067_,
		_w4088_,
		_w4998_,
		_w16215_
	);
	LUT4 #(
		.INIT('ha888)
	) name12168 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		_w4064_,
		_w4067_,
		_w4088_,
		_w16216_
	);
	LUT2 #(
		.INIT('he)
	) name12169 (
		_w16215_,
		_w16216_,
		_w16217_
	);
	LUT3 #(
		.INIT('hca)
	) name12170 (
		\sport1_txctl_TXSHT_reg[12]/P0001 ,
		\sport1_txctl_TX_reg[13]/P0001 ,
		_w14269_,
		_w16218_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12171 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		\core_c_psq_EXA_reg[1]/P0001 ,
		_w4073_,
		_w4084_,
		_w16219_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12172 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		\core_c_psq_EXA_reg[10]/P0001 ,
		_w4073_,
		_w4084_,
		_w16220_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12173 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		\core_c_psq_EXA_reg[11]/P0001 ,
		_w4073_,
		_w4084_,
		_w16221_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12174 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		\core_c_psq_EXA_reg[5]/P0001 ,
		_w4073_,
		_w4084_,
		_w16222_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12175 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		\core_c_psq_EXA_reg[4]/P0001 ,
		_w4073_,
		_w4084_,
		_w16223_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name12176 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		\core_c_psq_EXA_reg[8]/P0001 ,
		_w4073_,
		_w4084_,
		_w16224_
	);
	LUT4 #(
		.INIT('haacf)
	) name12177 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w4526_,
		_w4538_,
		_w16174_,
		_w16225_
	);
	LUT4 #(
		.INIT('haacf)
	) name12178 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w4827_,
		_w4833_,
		_w16174_,
		_w16226_
	);
	LUT4 #(
		.INIT('haacf)
	) name12179 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w4621_,
		_w4631_,
		_w16174_,
		_w16227_
	);
	LUT4 #(
		.INIT('haacf)
	) name12180 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w4688_,
		_w4694_,
		_w16174_,
		_w16228_
	);
	LUT4 #(
		.INIT('h1011)
	) name12181 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w6774_,
		_w6894_,
		_w6896_,
		_w16229_
	);
	LUT4 #(
		.INIT('h4445)
	) name12182 (
		_w13096_,
		_w13132_,
		_w13129_,
		_w13130_,
		_w16230_
	);
	LUT2 #(
		.INIT('h1)
	) name12183 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w13138_,
		_w16231_
	);
	LUT3 #(
		.INIT('h40)
	) name12184 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w16232_
	);
	LUT2 #(
		.INIT('h1)
	) name12185 (
		_w13158_,
		_w16232_,
		_w16233_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12186 (
		_w13155_,
		_w16230_,
		_w16231_,
		_w16233_,
		_w16234_
	);
	LUT4 #(
		.INIT('hafac)
	) name12187 (
		\sport0_rxctl_RXSHT_reg[1]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w16235_
	);
	LUT4 #(
		.INIT('h0002)
	) name12188 (
		\sport0_rxctl_RX_reg[1]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w16236_
	);
	LUT4 #(
		.INIT('hffb0)
	) name12189 (
		_w16229_,
		_w16234_,
		_w16235_,
		_w16236_,
		_w16237_
	);
	LUT4 #(
		.INIT('h81ff)
	) name12190 (
		_w11335_,
		_w11464_,
		_w11468_,
		_w14774_,
		_w16238_
	);
	LUT4 #(
		.INIT('h81ff)
	) name12191 (
		_w11335_,
		_w11448_,
		_w11452_,
		_w14774_,
		_w16239_
	);
	LUT4 #(
		.INIT('h81ff)
	) name12192 (
		_w11335_,
		_w11506_,
		_w11510_,
		_w14774_,
		_w16240_
	);
	LUT4 #(
		.INIT('h8100)
	) name12193 (
		_w11335_,
		_w11506_,
		_w11510_,
		_w14774_,
		_w16241_
	);
	LUT4 #(
		.INIT('h80f0)
	) name12194 (
		_w14784_,
		_w14783_,
		_w16239_,
		_w16241_,
		_w16242_
	);
	LUT4 #(
		.INIT('h81ff)
	) name12195 (
		_w11335_,
		_w11514_,
		_w11457_,
		_w14774_,
		_w16243_
	);
	LUT4 #(
		.INIT('h81ff)
	) name12196 (
		_w11335_,
		_w11494_,
		_w11498_,
		_w14774_,
		_w16244_
	);
	LUT4 #(
		.INIT('h2f00)
	) name12197 (
		_w16238_,
		_w16242_,
		_w16243_,
		_w16244_,
		_w16245_
	);
	LUT4 #(
		.INIT('h81ff)
	) name12198 (
		_w11536_,
		_w11540_,
		_w11335_,
		_w14774_,
		_w16246_
	);
	LUT3 #(
		.INIT('h02)
	) name12199 (
		_w14800_,
		_w14802_,
		_w14803_,
		_w16247_
	);
	LUT4 #(
		.INIT('h1055)
	) name12200 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w16245_,
		_w16246_,
		_w16247_,
		_w16248_
	);
	LUT4 #(
		.INIT('h0057)
	) name12201 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w12006_,
		_w12007_,
		_w16248_,
		_w16249_
	);
	LUT3 #(
		.INIT('he2)
	) name12202 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001 ,
		_w14809_,
		_w16249_,
		_w16250_
	);
	LUT3 #(
		.INIT('he2)
	) name12203 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001 ,
		_w14780_,
		_w16249_,
		_w16251_
	);
	LUT2 #(
		.INIT('h6)
	) name12204 (
		\clkc_CTR_cnt_reg[0]/NET0131 ,
		\clkc_CTR_cnt_reg[1]/NET0131 ,
		_w16252_
	);
	LUT2 #(
		.INIT('h1)
	) name12205 (
		\auctl_R0Sack_reg/NET0131 ,
		\auctl_RST_reg/P0001 ,
		_w16253_
	);
	LUT2 #(
		.INIT('h1)
	) name12206 (
		\auctl_RST_reg/P0001 ,
		\auctl_T0Sack_reg/NET0131 ,
		_w16254_
	);
	LUT2 #(
		.INIT('h1)
	) name12207 (
		\auctl_R1Sack_reg/NET0131 ,
		\auctl_RST_reg/P0001 ,
		_w16255_
	);
	LUT3 #(
		.INIT('h20)
	) name12208 (
		\sice_ICYC_en_syn_reg/P0001 ,
		_w8484_,
		_w8490_,
		_w16256_
	);
	LUT2 #(
		.INIT('h1)
	) name12209 (
		\auctl_RST_reg/P0001 ,
		\auctl_T1Sack_reg/NET0131 ,
		_w16257_
	);
	LUT4 #(
		.INIT('hfbff)
	) name12210 (
		_w4094_,
		_w4097_,
		_w4101_,
		_w4140_,
		_w16258_
	);
	LUT4 #(
		.INIT('hd700)
	) name12211 (
		T_IMS_pad,
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w16259_
	);
	LUT4 #(
		.INIT('h287b)
	) name12212 (
		T_IMS_pad,
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w16260_
	);
	LUT2 #(
		.INIT('h2)
	) name12213 (
		_w8482_,
		_w16260_,
		_w16261_
	);
	LUT3 #(
		.INIT('h13)
	) name12214 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 ,
		_w9894_,
		_w16262_
	);
	LUT4 #(
		.INIT('h0002)
	) name12215 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w16262_,
		_w16263_
	);
	LUT4 #(
		.INIT('h5700)
	) name12216 (
		_w12282_,
		_w12626_,
		_w12627_,
		_w16263_,
		_w16264_
	);
	LUT4 #(
		.INIT('h313b)
	) name12217 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 ,
		_w11308_,
		_w11635_,
		_w16265_
	);
	LUT3 #(
		.INIT('h45)
	) name12218 (
		_w11624_,
		_w16264_,
		_w16265_,
		_w16266_
	);
	LUT2 #(
		.INIT('h6)
	) name12219 (
		_w11146_,
		_w11173_,
		_w16267_
	);
	LUT4 #(
		.INIT('h0451)
	) name12220 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11243_,
		_w12245_,
		_w16267_,
		_w16268_
	);
	LUT4 #(
		.INIT('h007d)
	) name12221 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16101_,
		_w16102_,
		_w16268_,
		_w16269_
	);
	LUT4 #(
		.INIT('hff82)
	) name12222 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16101_,
		_w16102_,
		_w16268_,
		_w16270_
	);
	LUT3 #(
		.INIT('hce)
	) name12223 (
		_w11624_,
		_w16266_,
		_w16269_,
		_w16271_
	);
	LUT3 #(
		.INIT('hef)
	) name12224 (
		\clkc_ckr_reg_DO_reg[15]/NET0131 ,
		_w8484_,
		_w8490_,
		_w16272_
	);
	LUT2 #(
		.INIT('h2)
	) name12225 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001 ,
		_w11310_,
		_w16273_
	);
	LUT3 #(
		.INIT('h01)
	) name12226 (
		_w9946_,
		_w12442_,
		_w16273_,
		_w16274_
	);
	LUT4 #(
		.INIT('hfd00)
	) name12227 (
		_w12440_,
		_w12626_,
		_w12627_,
		_w16274_,
		_w16275_
	);
	LUT3 #(
		.INIT('h07)
	) name12228 (
		_w9946_,
		_w16269_,
		_w16275_,
		_w16276_
	);
	LUT2 #(
		.INIT('h1)
	) name12229 (
		T_ISn_pad,
		T_IWRn_pad,
		_w16277_
	);
	LUT4 #(
		.INIT('hd258)
	) name12230 (
		T_IMS_pad,
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w16278_
	);
	LUT2 #(
		.INIT('h8)
	) name12231 (
		_w8482_,
		_w16278_,
		_w16279_
	);
	LUT4 #(
		.INIT('h5551)
	) name12232 (
		T_IMS_pad,
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w16280_
	);
	LUT2 #(
		.INIT('h8)
	) name12233 (
		_w8482_,
		_w16280_,
		_w16281_
	);
	LUT3 #(
		.INIT('hfe)
	) name12234 (
		\bdma_RST_pin_reg/P0001 ,
		\sice_ICYC_clr_reg/NET0131 ,
		\sice_RCS_reg[1]/NET0131 ,
		_w16282_
	);
	LUT4 #(
		.INIT('hbbab)
	) name12235 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTSR1_E_reg/P0001 ,
		\core_c_dec_updSR_E_reg/P0001 ,
		_w9453_,
		_w16283_
	);
	LUT2 #(
		.INIT('h8)
	) name12236 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w16284_
	);
	LUT3 #(
		.INIT('h80)
	) name12237 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w16285_
	);
	LUT2 #(
		.INIT('h4)
	) name12238 (
		_w16283_,
		_w16285_,
		_w16286_
	);
	LUT4 #(
		.INIT('hd500)
	) name12239 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w11924_,
		_w13505_,
		_w16284_,
		_w16287_
	);
	LUT4 #(
		.INIT('h0400)
	) name12240 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_updSR_E_reg/P0001 ,
		_w9453_,
		_w16287_,
		_w16288_
	);
	LUT3 #(
		.INIT('h10)
	) name12241 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w16289_
	);
	LUT4 #(
		.INIT('h0100)
	) name12242 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w16290_
	);
	LUT4 #(
		.INIT('hae00)
	) name12243 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_dec_updAR_E_reg/P0001 ,
		_w9453_,
		_w16290_,
		_w16291_
	);
	LUT2 #(
		.INIT('h4)
	) name12244 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w16292_
	);
	LUT4 #(
		.INIT('h5400)
	) name12245 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR0_E_reg/P0001 ,
		_w11305_,
		_w16292_,
		_w16293_
	);
	LUT4 #(
		.INIT('h0400)
	) name12246 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w16294_
	);
	LUT3 #(
		.INIT('ha8)
	) name12247 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w16293_,
		_w16294_,
		_w16295_
	);
	LUT2 #(
		.INIT('h2)
	) name12248 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w16296_
	);
	LUT3 #(
		.INIT('h40)
	) name12249 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTMR2_E_reg/P0001 ,
		_w16297_
	);
	LUT4 #(
		.INIT('h00ab)
	) name12250 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w11305_,
		_w16297_,
		_w16298_
	);
	LUT2 #(
		.INIT('h2)
	) name12251 (
		_w16296_,
		_w16298_,
		_w16299_
	);
	LUT4 #(
		.INIT('h0001)
	) name12252 (
		_w16295_,
		_w16299_,
		_w16291_,
		_w16288_,
		_w16300_
	);
	LUT3 #(
		.INIT('h40)
	) name12253 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w16301_
	);
	LUT2 #(
		.INIT('h1)
	) name12254 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w16302_
	);
	LUT3 #(
		.INIT('h40)
	) name12255 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w16303_
	);
	LUT4 #(
		.INIT('h0777)
	) name12256 (
		_w11630_,
		_w16301_,
		_w16302_,
		_w16303_,
		_w16304_
	);
	LUT4 #(
		.INIT('h008a)
	) name12257 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w16304_,
		_w16305_
	);
	LUT2 #(
		.INIT('h4)
	) name12258 (
		_w4856_,
		_w16305_,
		_w16306_
	);
	LUT4 #(
		.INIT('ha200)
	) name12259 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w16296_,
		_w16307_
	);
	LUT2 #(
		.INIT('h8)
	) name12260 (
		_w11304_,
		_w16307_,
		_w16308_
	);
	LUT4 #(
		.INIT('h8a00)
	) name12261 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w16308_,
		_w16309_
	);
	LUT3 #(
		.INIT('h0b)
	) name12262 (
		_w4856_,
		_w16305_,
		_w16309_,
		_w16310_
	);
	LUT2 #(
		.INIT('h8)
	) name12263 (
		_w16296_,
		_w16297_,
		_w16311_
	);
	LUT4 #(
		.INIT('h7000)
	) name12264 (
		_w11917_,
		_w11920_,
		_w11924_,
		_w16311_,
		_w16312_
	);
	LUT3 #(
		.INIT('h20)
	) name12265 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w4856_,
		_w16312_,
		_w16313_
	);
	LUT4 #(
		.INIT('h000b)
	) name12266 (
		_w4856_,
		_w16305_,
		_w16309_,
		_w16313_,
		_w16314_
	);
	LUT4 #(
		.INIT('h0b00)
	) name12267 (
		_w4856_,
		_w16305_,
		_w16309_,
		_w16313_,
		_w16315_
	);
	LUT3 #(
		.INIT('h31)
	) name12268 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		\core_c_dec_accPM_E_reg/P0001 ,
		_w4855_,
		_w16316_
	);
	LUT2 #(
		.INIT('h8)
	) name12269 (
		_w16312_,
		_w16316_,
		_w16317_
	);
	LUT3 #(
		.INIT('h4f)
	) name12270 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w4856_,
		_w16312_,
		_w16318_
	);
	LUT2 #(
		.INIT('h8)
	) name12271 (
		_w16309_,
		_w16318_,
		_w16319_
	);
	LUT2 #(
		.INIT('h1)
	) name12272 (
		_w16315_,
		_w16319_,
		_w16320_
	);
	LUT2 #(
		.INIT('he)
	) name12273 (
		_w16315_,
		_w16319_,
		_w16321_
	);
	LUT4 #(
		.INIT('h0001)
	) name12274 (
		_w16306_,
		_w16314_,
		_w16315_,
		_w16319_,
		_w16322_
	);
	LUT3 #(
		.INIT('hca)
	) name12275 (
		\sport0_txctl_TXSHT_reg[12]/P0001 ,
		\sport0_txctl_TX_reg[13]/P0001 ,
		_w12552_,
		_w16323_
	);
	LUT3 #(
		.INIT('h02)
	) name12276 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		\sice_DBR1_reg[10]/P0001 ,
		\sice_DMR1_reg[10]/NET0131 ,
		_w16324_
	);
	LUT2 #(
		.INIT('h6)
	) name12277 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[17]/P0001 ,
		_w16325_
	);
	LUT3 #(
		.INIT('h04)
	) name12278 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		\sice_DBR1_reg[10]/P0001 ,
		\sice_DMR1_reg[10]/NET0131 ,
		_w16326_
	);
	LUT3 #(
		.INIT('h04)
	) name12279 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR1_reg[11]/P0001 ,
		\sice_DMR1_reg[11]/NET0131 ,
		_w16327_
	);
	LUT4 #(
		.INIT('h0001)
	) name12280 (
		_w16324_,
		_w16325_,
		_w16326_,
		_w16327_,
		_w16328_
	);
	LUT3 #(
		.INIT('h06)
	) name12281 (
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[16]/P0001 ,
		\sice_DMR1_reg[16]/NET0131 ,
		_w16329_
	);
	LUT3 #(
		.INIT('h02)
	) name12282 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR1_reg[11]/P0001 ,
		\sice_DMR1_reg[11]/NET0131 ,
		_w16330_
	);
	LUT2 #(
		.INIT('h4)
	) name12283 (
		\sice_DBR1_reg[18]/P0001 ,
		\sice_DMR1_reg[17]/NET0131 ,
		_w16331_
	);
	LUT3 #(
		.INIT('h10)
	) name12284 (
		_w16330_,
		_w16329_,
		_w16331_,
		_w16332_
	);
	LUT3 #(
		.INIT('h06)
	) name12285 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[1]/P0001 ,
		\sice_DMR1_reg[1]/NET0131 ,
		_w16333_
	);
	LUT3 #(
		.INIT('h06)
	) name12286 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[3]/P0001 ,
		\sice_DMR1_reg[3]/NET0131 ,
		_w16334_
	);
	LUT2 #(
		.INIT('h1)
	) name12287 (
		_w16333_,
		_w16334_,
		_w16335_
	);
	LUT3 #(
		.INIT('h80)
	) name12288 (
		_w16328_,
		_w16332_,
		_w16335_,
		_w16336_
	);
	LUT3 #(
		.INIT('h06)
	) name12289 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[0]/P0001 ,
		\sice_DMR1_reg[0]/NET0131 ,
		_w16337_
	);
	LUT3 #(
		.INIT('h06)
	) name12290 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR1_reg[6]/P0001 ,
		\sice_DMR1_reg[6]/NET0131 ,
		_w16338_
	);
	LUT3 #(
		.INIT('h06)
	) name12291 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR1_reg[9]/P0001 ,
		\sice_DMR1_reg[9]/NET0131 ,
		_w16339_
	);
	LUT3 #(
		.INIT('h06)
	) name12292 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR1_reg[7]/P0001 ,
		\sice_DMR1_reg[7]/NET0131 ,
		_w16340_
	);
	LUT4 #(
		.INIT('h0001)
	) name12293 (
		_w16337_,
		_w16338_,
		_w16339_,
		_w16340_,
		_w16341_
	);
	LUT3 #(
		.INIT('h06)
	) name12294 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR1_reg[13]/P0001 ,
		\sice_DMR1_reg[13]/NET0131 ,
		_w16342_
	);
	LUT3 #(
		.INIT('h06)
	) name12295 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR1_reg[5]/P0001 ,
		\sice_DMR1_reg[5]/NET0131 ,
		_w16343_
	);
	LUT3 #(
		.INIT('h06)
	) name12296 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR1_reg[12]/P0001 ,
		\sice_DMR1_reg[12]/NET0131 ,
		_w16344_
	);
	LUT3 #(
		.INIT('h06)
	) name12297 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR1_reg[8]/P0001 ,
		\sice_DMR1_reg[8]/NET0131 ,
		_w16345_
	);
	LUT4 #(
		.INIT('h0001)
	) name12298 (
		_w16342_,
		_w16343_,
		_w16344_,
		_w16345_,
		_w16346_
	);
	LUT3 #(
		.INIT('h06)
	) name12299 (
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[15]/P0001 ,
		\sice_DMR1_reg[15]/NET0131 ,
		_w16347_
	);
	LUT3 #(
		.INIT('h06)
	) name12300 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[2]/P0001 ,
		\sice_DMR1_reg[2]/NET0131 ,
		_w16348_
	);
	LUT3 #(
		.INIT('h06)
	) name12301 (
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[14]/P0001 ,
		\sice_DMR1_reg[14]/NET0131 ,
		_w16349_
	);
	LUT3 #(
		.INIT('h06)
	) name12302 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR1_reg[4]/P0001 ,
		\sice_DMR1_reg[4]/NET0131 ,
		_w16350_
	);
	LUT4 #(
		.INIT('h0001)
	) name12303 (
		_w16347_,
		_w16348_,
		_w16349_,
		_w16350_,
		_w16351_
	);
	LUT3 #(
		.INIT('h80)
	) name12304 (
		_w16341_,
		_w16346_,
		_w16351_,
		_w16352_
	);
	LUT3 #(
		.INIT('h02)
	) name12305 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR2_reg[5]/P0001 ,
		\sice_DMR2_reg[5]/NET0131 ,
		_w16353_
	);
	LUT3 #(
		.INIT('h02)
	) name12306 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		\sice_DBR2_reg[10]/P0001 ,
		\sice_DMR2_reg[10]/NET0131 ,
		_w16354_
	);
	LUT3 #(
		.INIT('h04)
	) name12307 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		\sice_DBR2_reg[10]/P0001 ,
		\sice_DMR2_reg[10]/NET0131 ,
		_w16355_
	);
	LUT3 #(
		.INIT('h04)
	) name12308 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR2_reg[5]/P0001 ,
		\sice_DMR2_reg[5]/NET0131 ,
		_w16356_
	);
	LUT4 #(
		.INIT('h0001)
	) name12309 (
		_w16353_,
		_w16354_,
		_w16355_,
		_w16356_,
		_w16357_
	);
	LUT3 #(
		.INIT('h06)
	) name12310 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR2_reg[9]/P0001 ,
		\sice_DMR2_reg[9]/NET0131 ,
		_w16358_
	);
	LUT4 #(
		.INIT('h0900)
	) name12311 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[17]/P0001 ,
		\sice_DBR2_reg[18]/P0001 ,
		\sice_DMR2_reg[17]/NET0131 ,
		_w16359_
	);
	LUT3 #(
		.INIT('h06)
	) name12312 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR2_reg[11]/P0001 ,
		\sice_DMR2_reg[11]/NET0131 ,
		_w16360_
	);
	LUT3 #(
		.INIT('h06)
	) name12313 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR2_reg[4]/P0001 ,
		\sice_DMR2_reg[4]/NET0131 ,
		_w16361_
	);
	LUT4 #(
		.INIT('h0100)
	) name12314 (
		_w16358_,
		_w16360_,
		_w16361_,
		_w16359_,
		_w16362_
	);
	LUT2 #(
		.INIT('h8)
	) name12315 (
		_w16357_,
		_w16362_,
		_w16363_
	);
	LUT3 #(
		.INIT('h06)
	) name12316 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR2_reg[7]/P0001 ,
		\sice_DMR2_reg[7]/NET0131 ,
		_w16364_
	);
	LUT3 #(
		.INIT('h06)
	) name12317 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[2]/P0001 ,
		\sice_DMR2_reg[2]/NET0131 ,
		_w16365_
	);
	LUT3 #(
		.INIT('h06)
	) name12318 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[0]/P0001 ,
		\sice_DMR2_reg[0]/NET0131 ,
		_w16366_
	);
	LUT3 #(
		.INIT('h06)
	) name12319 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR2_reg[13]/P0001 ,
		\sice_DMR2_reg[13]/NET0131 ,
		_w16367_
	);
	LUT4 #(
		.INIT('h0001)
	) name12320 (
		_w16364_,
		_w16365_,
		_w16366_,
		_w16367_,
		_w16368_
	);
	LUT3 #(
		.INIT('h06)
	) name12321 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[3]/P0001 ,
		\sice_DMR2_reg[3]/NET0131 ,
		_w16369_
	);
	LUT3 #(
		.INIT('h06)
	) name12322 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR2_reg[12]/P0001 ,
		\sice_DMR2_reg[12]/NET0131 ,
		_w16370_
	);
	LUT3 #(
		.INIT('h06)
	) name12323 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[1]/P0001 ,
		\sice_DMR2_reg[1]/NET0131 ,
		_w16371_
	);
	LUT3 #(
		.INIT('h06)
	) name12324 (
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[16]/P0001 ,
		\sice_DMR2_reg[16]/NET0131 ,
		_w16372_
	);
	LUT4 #(
		.INIT('h0001)
	) name12325 (
		_w16369_,
		_w16370_,
		_w16371_,
		_w16372_,
		_w16373_
	);
	LUT3 #(
		.INIT('h06)
	) name12326 (
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[14]/P0001 ,
		\sice_DMR2_reg[14]/NET0131 ,
		_w16374_
	);
	LUT3 #(
		.INIT('h06)
	) name12327 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR2_reg[8]/P0001 ,
		\sice_DMR2_reg[8]/NET0131 ,
		_w16375_
	);
	LUT3 #(
		.INIT('h06)
	) name12328 (
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[15]/P0001 ,
		\sice_DMR2_reg[15]/NET0131 ,
		_w16376_
	);
	LUT3 #(
		.INIT('h06)
	) name12329 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR2_reg[6]/P0001 ,
		\sice_DMR2_reg[6]/NET0131 ,
		_w16377_
	);
	LUT4 #(
		.INIT('h0001)
	) name12330 (
		_w16374_,
		_w16375_,
		_w16376_,
		_w16377_,
		_w16378_
	);
	LUT3 #(
		.INIT('h80)
	) name12331 (
		_w16368_,
		_w16373_,
		_w16378_,
		_w16379_
	);
	LUT4 #(
		.INIT('h0777)
	) name12332 (
		_w16336_,
		_w16352_,
		_w16363_,
		_w16379_,
		_w16380_
	);
	LUT2 #(
		.INIT('h4)
	) name12333 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\memc_accPM_E_reg/NET0131 ,
		_w16381_
	);
	LUT3 #(
		.INIT('h04)
	) name12334 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		\sice_DBR2_reg[10]/P0001 ,
		\sice_DMR2_reg[10]/NET0131 ,
		_w16382_
	);
	LUT3 #(
		.INIT('h04)
	) name12335 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR2_reg[5]/P0001 ,
		\sice_DMR2_reg[5]/NET0131 ,
		_w16383_
	);
	LUT3 #(
		.INIT('h02)
	) name12336 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		\sice_DBR2_reg[10]/P0001 ,
		\sice_DMR2_reg[10]/NET0131 ,
		_w16384_
	);
	LUT3 #(
		.INIT('h02)
	) name12337 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR2_reg[5]/P0001 ,
		\sice_DMR2_reg[5]/NET0131 ,
		_w16385_
	);
	LUT4 #(
		.INIT('h0001)
	) name12338 (
		_w16382_,
		_w16383_,
		_w16384_,
		_w16385_,
		_w16386_
	);
	LUT3 #(
		.INIT('h06)
	) name12339 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[3]/P0001 ,
		\sice_DMR2_reg[3]/NET0131 ,
		_w16387_
	);
	LUT4 #(
		.INIT('hb000)
	) name12340 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[17]/P0001 ,
		\sice_DBR2_reg[18]/P0001 ,
		\sice_DMR2_reg[17]/NET0131 ,
		_w16388_
	);
	LUT4 #(
		.INIT('h5010)
	) name12341 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\memc_accDM_E_reg/NET0131 ,
		\sice_DBR2_reg[17]/P0001 ,
		_w16389_
	);
	LUT3 #(
		.INIT('h40)
	) name12342 (
		_w16387_,
		_w16388_,
		_w16389_,
		_w16390_
	);
	LUT3 #(
		.INIT('h06)
	) name12343 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[1]/P0001 ,
		\sice_DMR2_reg[1]/NET0131 ,
		_w16391_
	);
	LUT3 #(
		.INIT('h06)
	) name12344 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR2_reg[11]/P0001 ,
		\sice_DMR2_reg[11]/NET0131 ,
		_w16392_
	);
	LUT2 #(
		.INIT('h1)
	) name12345 (
		_w16391_,
		_w16392_,
		_w16393_
	);
	LUT3 #(
		.INIT('h80)
	) name12346 (
		_w16386_,
		_w16390_,
		_w16393_,
		_w16394_
	);
	LUT3 #(
		.INIT('h06)
	) name12347 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR2_reg[13]/P0001 ,
		\sice_DMR2_reg[13]/NET0131 ,
		_w16395_
	);
	LUT3 #(
		.INIT('h06)
	) name12348 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR2_reg[7]/P0001 ,
		\sice_DMR2_reg[7]/NET0131 ,
		_w16396_
	);
	LUT3 #(
		.INIT('h06)
	) name12349 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[2]/P0001 ,
		\sice_DMR2_reg[2]/NET0131 ,
		_w16397_
	);
	LUT3 #(
		.INIT('h06)
	) name12350 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR2_reg[4]/P0001 ,
		\sice_DMR2_reg[4]/NET0131 ,
		_w16398_
	);
	LUT4 #(
		.INIT('h0001)
	) name12351 (
		_w16395_,
		_w16396_,
		_w16397_,
		_w16398_,
		_w16399_
	);
	LUT3 #(
		.INIT('h06)
	) name12352 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR2_reg[9]/P0001 ,
		\sice_DMR2_reg[9]/NET0131 ,
		_w16400_
	);
	LUT3 #(
		.INIT('h06)
	) name12353 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[0]/P0001 ,
		\sice_DMR2_reg[0]/NET0131 ,
		_w16401_
	);
	LUT3 #(
		.INIT('h06)
	) name12354 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[15]/P0001 ,
		\sice_DMR2_reg[15]/NET0131 ,
		_w16402_
	);
	LUT3 #(
		.INIT('h06)
	) name12355 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[14]/P0001 ,
		\sice_DMR2_reg[14]/NET0131 ,
		_w16403_
	);
	LUT4 #(
		.INIT('h0001)
	) name12356 (
		_w16400_,
		_w16401_,
		_w16402_,
		_w16403_,
		_w16404_
	);
	LUT3 #(
		.INIT('h06)
	) name12357 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR2_reg[12]/P0001 ,
		\sice_DMR2_reg[12]/NET0131 ,
		_w16405_
	);
	LUT3 #(
		.INIT('h06)
	) name12358 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR2_reg[6]/P0001 ,
		\sice_DMR2_reg[6]/NET0131 ,
		_w16406_
	);
	LUT3 #(
		.INIT('h06)
	) name12359 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR2_reg[8]/P0001 ,
		\sice_DMR2_reg[8]/NET0131 ,
		_w16407_
	);
	LUT3 #(
		.INIT('h06)
	) name12360 (
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[16]/P0001 ,
		\sice_DMR2_reg[16]/NET0131 ,
		_w16408_
	);
	LUT4 #(
		.INIT('h0001)
	) name12361 (
		_w16405_,
		_w16406_,
		_w16407_,
		_w16408_,
		_w16409_
	);
	LUT3 #(
		.INIT('h80)
	) name12362 (
		_w16399_,
		_w16404_,
		_w16409_,
		_w16410_
	);
	LUT3 #(
		.INIT('h04)
	) name12363 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		\sice_DBR1_reg[10]/P0001 ,
		\sice_DMR1_reg[10]/NET0131 ,
		_w16411_
	);
	LUT3 #(
		.INIT('h04)
	) name12364 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR1_reg[11]/P0001 ,
		\sice_DMR1_reg[11]/NET0131 ,
		_w16412_
	);
	LUT2 #(
		.INIT('h6)
	) name12365 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[17]/P0001 ,
		_w16413_
	);
	LUT3 #(
		.INIT('h02)
	) name12366 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR1_reg[11]/P0001 ,
		\sice_DMR1_reg[11]/NET0131 ,
		_w16414_
	);
	LUT4 #(
		.INIT('h0001)
	) name12367 (
		_w16411_,
		_w16412_,
		_w16413_,
		_w16414_,
		_w16415_
	);
	LUT3 #(
		.INIT('h06)
	) name12368 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[2]/P0001 ,
		\sice_DMR1_reg[2]/NET0131 ,
		_w16416_
	);
	LUT3 #(
		.INIT('h02)
	) name12369 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		\sice_DBR1_reg[10]/P0001 ,
		\sice_DMR1_reg[10]/NET0131 ,
		_w16417_
	);
	LUT4 #(
		.INIT('h4000)
	) name12370 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\memc_accDM_E_reg/NET0131 ,
		\sice_DBR1_reg[18]/P0001 ,
		\sice_DMR1_reg[17]/NET0131 ,
		_w16418_
	);
	LUT3 #(
		.INIT('h10)
	) name12371 (
		_w16417_,
		_w16416_,
		_w16418_,
		_w16419_
	);
	LUT3 #(
		.INIT('h06)
	) name12372 (
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[16]/P0001 ,
		\sice_DMR1_reg[16]/NET0131 ,
		_w16420_
	);
	LUT3 #(
		.INIT('h06)
	) name12373 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR1_reg[5]/P0001 ,
		\sice_DMR1_reg[5]/NET0131 ,
		_w16421_
	);
	LUT2 #(
		.INIT('h1)
	) name12374 (
		_w16420_,
		_w16421_,
		_w16422_
	);
	LUT3 #(
		.INIT('h80)
	) name12375 (
		_w16415_,
		_w16419_,
		_w16422_,
		_w16423_
	);
	LUT3 #(
		.INIT('h06)
	) name12376 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR1_reg[8]/P0001 ,
		\sice_DMR1_reg[8]/NET0131 ,
		_w16424_
	);
	LUT3 #(
		.INIT('h06)
	) name12377 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR1_reg[4]/P0001 ,
		\sice_DMR1_reg[4]/NET0131 ,
		_w16425_
	);
	LUT3 #(
		.INIT('h06)
	) name12378 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR1_reg[6]/P0001 ,
		\sice_DMR1_reg[6]/NET0131 ,
		_w16426_
	);
	LUT3 #(
		.INIT('h06)
	) name12379 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[0]/P0001 ,
		\sice_DMR1_reg[0]/NET0131 ,
		_w16427_
	);
	LUT4 #(
		.INIT('h0001)
	) name12380 (
		_w16424_,
		_w16425_,
		_w16426_,
		_w16427_,
		_w16428_
	);
	LUT3 #(
		.INIT('h06)
	) name12381 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR1_reg[13]/P0001 ,
		\sice_DMR1_reg[13]/NET0131 ,
		_w16429_
	);
	LUT3 #(
		.INIT('h06)
	) name12382 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[15]/P0001 ,
		\sice_DMR1_reg[15]/NET0131 ,
		_w16430_
	);
	LUT3 #(
		.INIT('h06)
	) name12383 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[14]/P0001 ,
		\sice_DMR1_reg[14]/NET0131 ,
		_w16431_
	);
	LUT3 #(
		.INIT('h06)
	) name12384 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[3]/P0001 ,
		\sice_DMR1_reg[3]/NET0131 ,
		_w16432_
	);
	LUT4 #(
		.INIT('h0001)
	) name12385 (
		_w16429_,
		_w16430_,
		_w16431_,
		_w16432_,
		_w16433_
	);
	LUT3 #(
		.INIT('h06)
	) name12386 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR1_reg[7]/P0001 ,
		\sice_DMR1_reg[7]/NET0131 ,
		_w16434_
	);
	LUT3 #(
		.INIT('h06)
	) name12387 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR1_reg[12]/P0001 ,
		\sice_DMR1_reg[12]/NET0131 ,
		_w16435_
	);
	LUT3 #(
		.INIT('h06)
	) name12388 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[1]/P0001 ,
		\sice_DMR1_reg[1]/NET0131 ,
		_w16436_
	);
	LUT3 #(
		.INIT('h06)
	) name12389 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR1_reg[9]/P0001 ,
		\sice_DMR1_reg[9]/NET0131 ,
		_w16437_
	);
	LUT4 #(
		.INIT('h0001)
	) name12390 (
		_w16434_,
		_w16435_,
		_w16436_,
		_w16437_,
		_w16438_
	);
	LUT3 #(
		.INIT('h80)
	) name12391 (
		_w16428_,
		_w16433_,
		_w16438_,
		_w16439_
	);
	LUT4 #(
		.INIT('h0777)
	) name12392 (
		_w16394_,
		_w16410_,
		_w16423_,
		_w16439_,
		_w16440_
	);
	LUT4 #(
		.INIT('h20aa)
	) name12393 (
		\sice_ITR_reg[2]/NET0131 ,
		_w16380_,
		_w16381_,
		_w16440_,
		_w16441_
	);
	LUT3 #(
		.INIT('h06)
	) name12394 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		\sice_IBR2_reg[6]/P0001 ,
		\sice_IMR2_reg[6]/NET0131 ,
		_w16442_
	);
	LUT4 #(
		.INIT('h9000)
	) name12395 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\sice_IBR2_reg[17]/P0001 ,
		\sice_IMR2_reg[17]/NET0131 ,
		\sice_ITR_reg[1]/NET0131 ,
		_w16443_
	);
	LUT2 #(
		.INIT('h4)
	) name12396 (
		_w16442_,
		_w16443_,
		_w16444_
	);
	LUT3 #(
		.INIT('h06)
	) name12397 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		\sice_IBR2_reg[12]/P0001 ,
		\sice_IMR2_reg[12]/NET0131 ,
		_w16445_
	);
	LUT3 #(
		.INIT('h06)
	) name12398 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		\sice_IBR2_reg[9]/P0001 ,
		\sice_IMR2_reg[9]/NET0131 ,
		_w16446_
	);
	LUT3 #(
		.INIT('h06)
	) name12399 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		\sice_IBR2_reg[4]/P0001 ,
		\sice_IMR2_reg[4]/NET0131 ,
		_w16447_
	);
	LUT3 #(
		.INIT('h06)
	) name12400 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\sice_IBR2_reg[16]/P0001 ,
		\sice_IMR2_reg[16]/NET0131 ,
		_w16448_
	);
	LUT4 #(
		.INIT('h0001)
	) name12401 (
		_w16445_,
		_w16446_,
		_w16447_,
		_w16448_,
		_w16449_
	);
	LUT2 #(
		.INIT('h8)
	) name12402 (
		_w16444_,
		_w16449_,
		_w16450_
	);
	LUT3 #(
		.INIT('h06)
	) name12403 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		\sice_IBR2_reg[11]/P0001 ,
		\sice_IMR2_reg[11]/NET0131 ,
		_w16451_
	);
	LUT3 #(
		.INIT('h06)
	) name12404 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		\sice_IBR2_reg[3]/P0001 ,
		\sice_IMR2_reg[3]/NET0131 ,
		_w16452_
	);
	LUT3 #(
		.INIT('h06)
	) name12405 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\sice_IBR2_reg[15]/P0001 ,
		\sice_IMR2_reg[15]/NET0131 ,
		_w16453_
	);
	LUT3 #(
		.INIT('h06)
	) name12406 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		\sice_IBR2_reg[10]/P0001 ,
		\sice_IMR2_reg[10]/NET0131 ,
		_w16454_
	);
	LUT4 #(
		.INIT('h0001)
	) name12407 (
		_w16451_,
		_w16452_,
		_w16453_,
		_w16454_,
		_w16455_
	);
	LUT3 #(
		.INIT('h06)
	) name12408 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		\sice_IBR2_reg[13]/P0001 ,
		\sice_IMR2_reg[13]/NET0131 ,
		_w16456_
	);
	LUT3 #(
		.INIT('h06)
	) name12409 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		\sice_IBR2_reg[5]/P0001 ,
		\sice_IMR2_reg[5]/NET0131 ,
		_w16457_
	);
	LUT3 #(
		.INIT('h06)
	) name12410 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\sice_IBR2_reg[14]/P0001 ,
		\sice_IMR2_reg[14]/NET0131 ,
		_w16458_
	);
	LUT3 #(
		.INIT('h06)
	) name12411 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		\sice_IBR2_reg[7]/P0001 ,
		\sice_IMR2_reg[7]/NET0131 ,
		_w16459_
	);
	LUT4 #(
		.INIT('h0001)
	) name12412 (
		_w16456_,
		_w16457_,
		_w16458_,
		_w16459_,
		_w16460_
	);
	LUT3 #(
		.INIT('h06)
	) name12413 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		\sice_IBR2_reg[1]/P0001 ,
		\sice_IMR2_reg[1]/NET0131 ,
		_w16461_
	);
	LUT3 #(
		.INIT('h06)
	) name12414 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		\sice_IBR2_reg[2]/P0001 ,
		\sice_IMR2_reg[2]/NET0131 ,
		_w16462_
	);
	LUT3 #(
		.INIT('h06)
	) name12415 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		\sice_IBR2_reg[0]/P0001 ,
		\sice_IMR2_reg[0]/NET0131 ,
		_w16463_
	);
	LUT3 #(
		.INIT('h06)
	) name12416 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		\sice_IBR2_reg[8]/P0001 ,
		\sice_IMR2_reg[8]/NET0131 ,
		_w16464_
	);
	LUT4 #(
		.INIT('h0001)
	) name12417 (
		_w16461_,
		_w16462_,
		_w16463_,
		_w16464_,
		_w16465_
	);
	LUT3 #(
		.INIT('h80)
	) name12418 (
		_w16455_,
		_w16460_,
		_w16465_,
		_w16466_
	);
	LUT2 #(
		.INIT('h8)
	) name12419 (
		_w16450_,
		_w16466_,
		_w16467_
	);
	LUT3 #(
		.INIT('h06)
	) name12420 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\sice_IBR1_reg[16]/P0001 ,
		\sice_IMR1_reg[16]/NET0131 ,
		_w16468_
	);
	LUT4 #(
		.INIT('h9000)
	) name12421 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\sice_IBR1_reg[17]/P0001 ,
		\sice_IMR1_reg[17]/NET0131 ,
		\sice_ITR_reg[1]/NET0131 ,
		_w16469_
	);
	LUT2 #(
		.INIT('h4)
	) name12422 (
		_w16468_,
		_w16469_,
		_w16470_
	);
	LUT3 #(
		.INIT('h06)
	) name12423 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		\sice_IBR1_reg[13]/P0001 ,
		\sice_IMR1_reg[13]/NET0131 ,
		_w16471_
	);
	LUT3 #(
		.INIT('h06)
	) name12424 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		\sice_IBR1_reg[6]/P0001 ,
		\sice_IMR1_reg[6]/NET0131 ,
		_w16472_
	);
	LUT3 #(
		.INIT('h06)
	) name12425 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		\sice_IBR1_reg[12]/P0001 ,
		\sice_IMR1_reg[12]/NET0131 ,
		_w16473_
	);
	LUT3 #(
		.INIT('h06)
	) name12426 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		\sice_IBR1_reg[8]/P0001 ,
		\sice_IMR1_reg[8]/NET0131 ,
		_w16474_
	);
	LUT4 #(
		.INIT('h0001)
	) name12427 (
		_w16471_,
		_w16472_,
		_w16473_,
		_w16474_,
		_w16475_
	);
	LUT2 #(
		.INIT('h8)
	) name12428 (
		_w16470_,
		_w16475_,
		_w16476_
	);
	LUT3 #(
		.INIT('h06)
	) name12429 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		\sice_IBR1_reg[3]/P0001 ,
		\sice_IMR1_reg[3]/NET0131 ,
		_w16477_
	);
	LUT3 #(
		.INIT('h06)
	) name12430 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		\sice_IBR1_reg[0]/P0001 ,
		\sice_IMR1_reg[0]/NET0131 ,
		_w16478_
	);
	LUT3 #(
		.INIT('h06)
	) name12431 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		\sice_IBR1_reg[9]/P0001 ,
		\sice_IMR1_reg[9]/NET0131 ,
		_w16479_
	);
	LUT3 #(
		.INIT('h06)
	) name12432 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		\sice_IBR1_reg[2]/P0001 ,
		\sice_IMR1_reg[2]/NET0131 ,
		_w16480_
	);
	LUT4 #(
		.INIT('h0001)
	) name12433 (
		_w16477_,
		_w16478_,
		_w16479_,
		_w16480_,
		_w16481_
	);
	LUT3 #(
		.INIT('h06)
	) name12434 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		\sice_IBR1_reg[1]/P0001 ,
		\sice_IMR1_reg[1]/NET0131 ,
		_w16482_
	);
	LUT3 #(
		.INIT('h06)
	) name12435 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		\sice_IBR1_reg[4]/P0001 ,
		\sice_IMR1_reg[4]/NET0131 ,
		_w16483_
	);
	LUT3 #(
		.INIT('h06)
	) name12436 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		\sice_IBR1_reg[11]/P0001 ,
		\sice_IMR1_reg[11]/NET0131 ,
		_w16484_
	);
	LUT3 #(
		.INIT('h06)
	) name12437 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\sice_IBR1_reg[14]/P0001 ,
		\sice_IMR1_reg[14]/NET0131 ,
		_w16485_
	);
	LUT4 #(
		.INIT('h0001)
	) name12438 (
		_w16482_,
		_w16483_,
		_w16484_,
		_w16485_,
		_w16486_
	);
	LUT3 #(
		.INIT('h06)
	) name12439 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		\sice_IBR1_reg[5]/P0001 ,
		\sice_IMR1_reg[5]/NET0131 ,
		_w16487_
	);
	LUT3 #(
		.INIT('h06)
	) name12440 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		\sice_IBR1_reg[10]/P0001 ,
		\sice_IMR1_reg[10]/NET0131 ,
		_w16488_
	);
	LUT3 #(
		.INIT('h06)
	) name12441 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\sice_IBR1_reg[15]/P0001 ,
		\sice_IMR1_reg[15]/NET0131 ,
		_w16489_
	);
	LUT3 #(
		.INIT('h06)
	) name12442 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		\sice_IBR1_reg[7]/P0001 ,
		\sice_IMR1_reg[7]/NET0131 ,
		_w16490_
	);
	LUT4 #(
		.INIT('h0001)
	) name12443 (
		_w16487_,
		_w16488_,
		_w16489_,
		_w16490_,
		_w16491_
	);
	LUT3 #(
		.INIT('h80)
	) name12444 (
		_w16481_,
		_w16486_,
		_w16491_,
		_w16492_
	);
	LUT4 #(
		.INIT('h0100)
	) name12445 (
		\core_c_psq_PCS_reg[0]/NET0131 ,
		\core_c_psq_PCS_reg[15]/NET0131 ,
		\core_c_psq_PCS_reg[1]/NET0131 ,
		\sice_GOICE_syn_reg/P0001 ,
		_w16493_
	);
	LUT2 #(
		.INIT('h8)
	) name12446 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\sice_ITR_reg[0]/NET0131 ,
		_w16494_
	);
	LUT4 #(
		.INIT('h8000)
	) name12447 (
		_w5026_,
		_w5028_,
		_w5045_,
		_w16494_,
		_w16495_
	);
	LUT2 #(
		.INIT('h1)
	) name12448 (
		_w16493_,
		_w16495_,
		_w16496_
	);
	LUT3 #(
		.INIT('h70)
	) name12449 (
		_w16476_,
		_w16492_,
		_w16496_,
		_w16497_
	);
	LUT2 #(
		.INIT('h4)
	) name12450 (
		_w16467_,
		_w16497_,
		_w16498_
	);
	LUT3 #(
		.INIT('h45)
	) name12451 (
		_w4084_,
		_w16441_,
		_w16498_,
		_w16499_
	);
	LUT4 #(
		.INIT('h1000)
	) name12452 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4428_,
		_w8172_,
		_w16499_,
		_w16500_
	);
	LUT4 #(
		.INIT('h4000)
	) name12453 (
		_w4094_,
		_w4097_,
		_w8482_,
		_w14834_,
		_w16501_
	);
	LUT3 #(
		.INIT('he0)
	) name12454 (
		\sice_HALT_E_reg/P0001 ,
		_w16500_,
		_w16501_,
		_w16502_
	);
	LUT2 #(
		.INIT('h8)
	) name12455 (
		_w16305_,
		_w16316_,
		_w16503_
	);
	LUT4 #(
		.INIT('h0075)
	) name12456 (
		_w16310_,
		_w16313_,
		_w16317_,
		_w16503_,
		_w16504_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12457 (
		_w16310_,
		_w16313_,
		_w16317_,
		_w16503_,
		_w16505_
	);
	LUT2 #(
		.INIT('h2)
	) name12458 (
		\sice_UpdDR_sd1_reg/P0001 ,
		\sice_UpdDR_sd2_reg/P0001 ,
		_w16506_
	);
	LUT4 #(
		.INIT('h0004)
	) name12459 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w16507_
	);
	LUT2 #(
		.INIT('h8)
	) name12460 (
		_w16506_,
		_w16507_,
		_w16508_
	);
	LUT2 #(
		.INIT('h4)
	) name12461 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTIDR_E_reg/P0001 ,
		_w16509_
	);
	LUT3 #(
		.INIT('h0b)
	) name12462 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTIDR_E_reg/P0001 ,
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16510_
	);
	LUT4 #(
		.INIT('h0f04)
	) name12463 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16508_,
		_w16510_,
		_w16511_
	);
	LUT4 #(
		.INIT('hf0fb)
	) name12464 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w16508_,
		_w16510_,
		_w16512_
	);
	LUT2 #(
		.INIT('h8)
	) name12465 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[15]/P0001 ,
		_w16513_
	);
	LUT4 #(
		.INIT('h0001)
	) name12466 (
		\idma_CMo_oe3_reg/P0001 ,
		\idma_CMo_oe4_reg/P0001 ,
		\idma_CMo_oe5_reg/P0001 ,
		\idma_CMo_oe6_reg/P0001 ,
		_w16514_
	);
	LUT2 #(
		.INIT('h1)
	) name12467 (
		\idma_CMo_oe1_reg/P0001 ,
		\idma_CMo_oe2_reg/P0001 ,
		_w16515_
	);
	LUT3 #(
		.INIT('h04)
	) name12468 (
		\idma_CM_oe_reg/P0001 ,
		\idma_CMo_oe0_reg/P0001 ,
		\idma_CMo_oe7_reg/P0001 ,
		_w16516_
	);
	LUT3 #(
		.INIT('h10)
	) name12469 (
		\idma_CM_oe_reg/P0001 ,
		\idma_CMo_oe0_reg/P0001 ,
		\idma_CMo_oe7_reg/P0001 ,
		_w16517_
	);
	LUT4 #(
		.INIT('h777f)
	) name12470 (
		_w16514_,
		_w16515_,
		_w16516_,
		_w16517_,
		_w16518_
	);
	LUT3 #(
		.INIT('h01)
	) name12471 (
		\idma_CM_oe_reg/P0001 ,
		\idma_CMo_oe0_reg/P0001 ,
		\idma_CMo_oe7_reg/P0001 ,
		_w16519_
	);
	LUT2 #(
		.INIT('h4)
	) name12472 (
		\idma_CMo_oe1_reg/P0001 ,
		\idma_CMo_oe2_reg/P0001 ,
		_w16520_
	);
	LUT3 #(
		.INIT('h80)
	) name12473 (
		_w16514_,
		_w16519_,
		_w16520_,
		_w16521_
	);
	LUT3 #(
		.INIT('h10)
	) name12474 (
		\idma_CMo_oe3_reg/P0001 ,
		\idma_CMo_oe4_reg/P0001 ,
		\idma_CMo_oe5_reg/P0001 ,
		_w16522_
	);
	LUT4 #(
		.INIT('h4000)
	) name12475 (
		\idma_CMo_oe6_reg/P0001 ,
		_w16519_,
		_w16515_,
		_w16522_,
		_w16523_
	);
	LUT3 #(
		.INIT('h10)
	) name12476 (
		_w16521_,
		_w16523_,
		_w16518_,
		_w16524_
	);
	LUT4 #(
		.INIT('h1000)
	) name12477 (
		\idma_CMo_oe5_reg/P0001 ,
		\idma_CMo_oe6_reg/P0001 ,
		_w16519_,
		_w16515_,
		_w16525_
	);
	LUT2 #(
		.INIT('h2)
	) name12478 (
		\idma_CMo_oe3_reg/P0001 ,
		\idma_CMo_oe4_reg/P0001 ,
		_w16526_
	);
	LUT2 #(
		.INIT('h8)
	) name12479 (
		_w16525_,
		_w16526_,
		_w16527_
	);
	LUT2 #(
		.INIT('h4)
	) name12480 (
		\idma_CMo_oe3_reg/P0001 ,
		\idma_CMo_oe4_reg/P0001 ,
		_w16528_
	);
	LUT2 #(
		.INIT('h2)
	) name12481 (
		\idma_CMo_oe1_reg/P0001 ,
		\idma_CMo_oe2_reg/P0001 ,
		_w16529_
	);
	LUT3 #(
		.INIT('h80)
	) name12482 (
		_w16514_,
		_w16519_,
		_w16529_,
		_w16530_
	);
	LUT4 #(
		.INIT('h0100)
	) name12483 (
		\idma_CMo_oe3_reg/P0001 ,
		\idma_CMo_oe4_reg/P0001 ,
		\idma_CMo_oe5_reg/P0001 ,
		\idma_CMo_oe6_reg/P0001 ,
		_w16531_
	);
	LUT3 #(
		.INIT('h80)
	) name12484 (
		_w16519_,
		_w16515_,
		_w16531_,
		_w16532_
	);
	LUT4 #(
		.INIT('h0111)
	) name12485 (
		_w16530_,
		_w16532_,
		_w16525_,
		_w16528_,
		_w16533_
	);
	LUT4 #(
		.INIT('h2000)
	) name12486 (
		\CM_rdm[15]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16534_
	);
	LUT4 #(
		.INIT('h8000)
	) name12487 (
		\CM_rd0[15]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16535_
	);
	LUT4 #(
		.INIT('h8000)
	) name12488 (
		\CM_rd7[15]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16536_
	);
	LUT2 #(
		.INIT('h1)
	) name12489 (
		_w16535_,
		_w16536_,
		_w16537_
	);
	LUT4 #(
		.INIT('h8000)
	) name12490 (
		\CM_rd2[15]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16538_
	);
	LUT3 #(
		.INIT('h13)
	) name12491 (
		\CM_rd5[15]_pad ,
		_w16538_,
		_w16523_,
		_w16539_
	);
	LUT2 #(
		.INIT('h8)
	) name12492 (
		_w16537_,
		_w16539_,
		_w16540_
	);
	LUT3 #(
		.INIT('h80)
	) name12493 (
		\CM_rd3[15]_pad ,
		_w16525_,
		_w16526_,
		_w16541_
	);
	LUT3 #(
		.INIT('h80)
	) name12494 (
		\CM_rd4[15]_pad ,
		_w16525_,
		_w16528_,
		_w16542_
	);
	LUT4 #(
		.INIT('h8000)
	) name12495 (
		\CM_rd1[15]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16543_
	);
	LUT4 #(
		.INIT('h8000)
	) name12496 (
		\CM_rd6[15]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16544_
	);
	LUT2 #(
		.INIT('h1)
	) name12497 (
		_w16543_,
		_w16544_,
		_w16545_
	);
	LUT3 #(
		.INIT('h10)
	) name12498 (
		_w16542_,
		_w16541_,
		_w16545_,
		_w16546_
	);
	LUT4 #(
		.INIT('h4555)
	) name12499 (
		\T_TMODE[1]_pad ,
		_w16534_,
		_w16540_,
		_w16546_,
		_w16547_
	);
	LUT3 #(
		.INIT('ha8)
	) name12500 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16513_,
		_w16547_,
		_w16548_
	);
	LUT4 #(
		.INIT('h00ef)
	) name12501 (
		_w8798_,
		_w8801_,
		_w16509_,
		_w16548_,
		_w16549_
	);
	LUT3 #(
		.INIT('h80)
	) name12502 (
		\sice_SPC_reg[15]/P0001 ,
		_w16506_,
		_w16507_,
		_w16550_
	);
	LUT3 #(
		.INIT('h07)
	) name12503 (
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w16511_,
		_w16550_,
		_w16551_
	);
	LUT3 #(
		.INIT('h1f)
	) name12504 (
		_w16511_,
		_w16549_,
		_w16551_,
		_w16552_
	);
	LUT3 #(
		.INIT('h13)
	) name12505 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 ,
		_w9894_,
		_w16553_
	);
	LUT4 #(
		.INIT('h0002)
	) name12506 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w16553_,
		_w16554_
	);
	LUT4 #(
		.INIT('h1f00)
	) name12507 (
		_w12006_,
		_w12007_,
		_w12282_,
		_w16554_,
		_w16555_
	);
	LUT4 #(
		.INIT('h313b)
	) name12508 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 ,
		_w11308_,
		_w11635_,
		_w16556_
	);
	LUT3 #(
		.INIT('h45)
	) name12509 (
		_w11624_,
		_w16555_,
		_w16556_,
		_w16557_
	);
	LUT4 #(
		.INIT('h0514)
	) name12510 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11239_,
		_w12383_,
		_w12384_,
		_w16558_
	);
	LUT2 #(
		.INIT('h6)
	) name12511 (
		_w11207_,
		_w11216_,
		_w16559_
	);
	LUT4 #(
		.INIT('h4f00)
	) name12512 (
		_w10433_,
		_w10640_,
		_w10645_,
		_w11230_,
		_w16560_
	);
	LUT4 #(
		.INIT('h0a28)
	) name12513 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11240_,
		_w16559_,
		_w16560_,
		_w16561_
	);
	LUT2 #(
		.INIT('he)
	) name12514 (
		_w16558_,
		_w16561_,
		_w16562_
	);
	LUT4 #(
		.INIT('heeec)
	) name12515 (
		_w11624_,
		_w16557_,
		_w16558_,
		_w16561_,
		_w16563_
	);
	LUT2 #(
		.INIT('h8)
	) name12516 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[14]/P0001 ,
		_w16564_
	);
	LUT4 #(
		.INIT('h2000)
	) name12517 (
		\CM_rdm[14]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16565_
	);
	LUT4 #(
		.INIT('h8000)
	) name12518 (
		\CM_rd0[14]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16566_
	);
	LUT4 #(
		.INIT('h8000)
	) name12519 (
		\CM_rd7[14]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16567_
	);
	LUT2 #(
		.INIT('h1)
	) name12520 (
		_w16566_,
		_w16567_,
		_w16568_
	);
	LUT4 #(
		.INIT('h8000)
	) name12521 (
		\CM_rd2[14]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16569_
	);
	LUT3 #(
		.INIT('h07)
	) name12522 (
		\CM_rd5[14]_pad ,
		_w16523_,
		_w16569_,
		_w16570_
	);
	LUT2 #(
		.INIT('h8)
	) name12523 (
		_w16568_,
		_w16570_,
		_w16571_
	);
	LUT3 #(
		.INIT('h80)
	) name12524 (
		\CM_rd3[14]_pad ,
		_w16525_,
		_w16526_,
		_w16572_
	);
	LUT3 #(
		.INIT('h80)
	) name12525 (
		\CM_rd4[14]_pad ,
		_w16525_,
		_w16528_,
		_w16573_
	);
	LUT4 #(
		.INIT('h8000)
	) name12526 (
		\CM_rd1[14]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16574_
	);
	LUT4 #(
		.INIT('h8000)
	) name12527 (
		\CM_rd6[14]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16575_
	);
	LUT2 #(
		.INIT('h1)
	) name12528 (
		_w16574_,
		_w16575_,
		_w16576_
	);
	LUT3 #(
		.INIT('h10)
	) name12529 (
		_w16573_,
		_w16572_,
		_w16576_,
		_w16577_
	);
	LUT4 #(
		.INIT('h4555)
	) name12530 (
		\T_TMODE[1]_pad ,
		_w16565_,
		_w16571_,
		_w16577_,
		_w16578_
	);
	LUT3 #(
		.INIT('ha8)
	) name12531 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16564_,
		_w16578_,
		_w16579_
	);
	LUT4 #(
		.INIT('h00ef)
	) name12532 (
		_w8757_,
		_w8760_,
		_w16509_,
		_w16579_,
		_w16580_
	);
	LUT3 #(
		.INIT('h80)
	) name12533 (
		\sice_SPC_reg[14]/P0001 ,
		_w16506_,
		_w16507_,
		_w16581_
	);
	LUT3 #(
		.INIT('h07)
	) name12534 (
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w16511_,
		_w16581_,
		_w16582_
	);
	LUT3 #(
		.INIT('h1f)
	) name12535 (
		_w16511_,
		_w16580_,
		_w16582_,
		_w16583_
	);
	LUT4 #(
		.INIT('h4500)
	) name12536 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w16509_,
		_w16584_
	);
	LUT2 #(
		.INIT('h8)
	) name12537 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[7]/P0001 ,
		_w16585_
	);
	LUT4 #(
		.INIT('h2000)
	) name12538 (
		\CM_rdm[7]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16586_
	);
	LUT4 #(
		.INIT('h8000)
	) name12539 (
		\CM_rd0[7]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16587_
	);
	LUT4 #(
		.INIT('h8000)
	) name12540 (
		\CM_rd7[7]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16588_
	);
	LUT2 #(
		.INIT('h1)
	) name12541 (
		_w16587_,
		_w16588_,
		_w16589_
	);
	LUT4 #(
		.INIT('h8000)
	) name12542 (
		\CM_rd2[7]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16590_
	);
	LUT3 #(
		.INIT('h07)
	) name12543 (
		\CM_rd5[7]_pad ,
		_w16523_,
		_w16590_,
		_w16591_
	);
	LUT2 #(
		.INIT('h8)
	) name12544 (
		_w16589_,
		_w16591_,
		_w16592_
	);
	LUT3 #(
		.INIT('h80)
	) name12545 (
		\CM_rd3[7]_pad ,
		_w16525_,
		_w16526_,
		_w16593_
	);
	LUT3 #(
		.INIT('h80)
	) name12546 (
		\CM_rd4[7]_pad ,
		_w16525_,
		_w16528_,
		_w16594_
	);
	LUT4 #(
		.INIT('h8000)
	) name12547 (
		\CM_rd1[7]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16595_
	);
	LUT4 #(
		.INIT('h8000)
	) name12548 (
		\CM_rd6[7]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16596_
	);
	LUT2 #(
		.INIT('h1)
	) name12549 (
		_w16595_,
		_w16596_,
		_w16597_
	);
	LUT3 #(
		.INIT('h10)
	) name12550 (
		_w16594_,
		_w16593_,
		_w16597_,
		_w16598_
	);
	LUT4 #(
		.INIT('h4555)
	) name12551 (
		\T_TMODE[1]_pad ,
		_w16586_,
		_w16592_,
		_w16598_,
		_w16599_
	);
	LUT3 #(
		.INIT('ha8)
	) name12552 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16585_,
		_w16599_,
		_w16600_
	);
	LUT3 #(
		.INIT('h80)
	) name12553 (
		\sice_SPC_reg[7]/P0001 ,
		_w16506_,
		_w16507_,
		_w16601_
	);
	LUT3 #(
		.INIT('h07)
	) name12554 (
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w16511_,
		_w16601_,
		_w16602_
	);
	LUT4 #(
		.INIT('h54ff)
	) name12555 (
		_w16511_,
		_w16584_,
		_w16600_,
		_w16602_,
		_w16603_
	);
	LUT4 #(
		.INIT('h4500)
	) name12556 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w16509_,
		_w16604_
	);
	LUT2 #(
		.INIT('h8)
	) name12557 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[6]/P0001 ,
		_w16605_
	);
	LUT4 #(
		.INIT('h2000)
	) name12558 (
		\CM_rdm[6]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16606_
	);
	LUT4 #(
		.INIT('h8000)
	) name12559 (
		\CM_rd0[6]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16607_
	);
	LUT4 #(
		.INIT('h8000)
	) name12560 (
		\CM_rd7[6]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16608_
	);
	LUT2 #(
		.INIT('h1)
	) name12561 (
		_w16607_,
		_w16608_,
		_w16609_
	);
	LUT4 #(
		.INIT('h8000)
	) name12562 (
		\CM_rd2[6]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16610_
	);
	LUT3 #(
		.INIT('h07)
	) name12563 (
		\CM_rd5[6]_pad ,
		_w16523_,
		_w16610_,
		_w16611_
	);
	LUT2 #(
		.INIT('h8)
	) name12564 (
		_w16609_,
		_w16611_,
		_w16612_
	);
	LUT3 #(
		.INIT('h80)
	) name12565 (
		\CM_rd3[6]_pad ,
		_w16525_,
		_w16526_,
		_w16613_
	);
	LUT3 #(
		.INIT('h80)
	) name12566 (
		\CM_rd4[6]_pad ,
		_w16525_,
		_w16528_,
		_w16614_
	);
	LUT4 #(
		.INIT('h8000)
	) name12567 (
		\CM_rd1[6]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16615_
	);
	LUT4 #(
		.INIT('h8000)
	) name12568 (
		\CM_rd6[6]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16616_
	);
	LUT2 #(
		.INIT('h1)
	) name12569 (
		_w16615_,
		_w16616_,
		_w16617_
	);
	LUT3 #(
		.INIT('h10)
	) name12570 (
		_w16614_,
		_w16613_,
		_w16617_,
		_w16618_
	);
	LUT4 #(
		.INIT('h4555)
	) name12571 (
		\T_TMODE[1]_pad ,
		_w16606_,
		_w16612_,
		_w16618_,
		_w16619_
	);
	LUT3 #(
		.INIT('ha8)
	) name12572 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16605_,
		_w16619_,
		_w16620_
	);
	LUT3 #(
		.INIT('h80)
	) name12573 (
		\sice_SPC_reg[6]/P0001 ,
		_w16506_,
		_w16507_,
		_w16621_
	);
	LUT3 #(
		.INIT('h07)
	) name12574 (
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w16511_,
		_w16621_,
		_w16622_
	);
	LUT4 #(
		.INIT('h54ff)
	) name12575 (
		_w16511_,
		_w16604_,
		_w16620_,
		_w16622_,
		_w16623_
	);
	LUT4 #(
		.INIT('h4500)
	) name12576 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w16509_,
		_w16624_
	);
	LUT2 #(
		.INIT('h8)
	) name12577 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[5]/P0001 ,
		_w16625_
	);
	LUT4 #(
		.INIT('h2000)
	) name12578 (
		\CM_rdm[5]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16626_
	);
	LUT4 #(
		.INIT('h8000)
	) name12579 (
		\CM_rd0[5]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16627_
	);
	LUT4 #(
		.INIT('h8000)
	) name12580 (
		\CM_rd7[5]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16628_
	);
	LUT2 #(
		.INIT('h1)
	) name12581 (
		_w16627_,
		_w16628_,
		_w16629_
	);
	LUT4 #(
		.INIT('h8000)
	) name12582 (
		\CM_rd2[5]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16630_
	);
	LUT3 #(
		.INIT('h07)
	) name12583 (
		\CM_rd5[5]_pad ,
		_w16523_,
		_w16630_,
		_w16631_
	);
	LUT2 #(
		.INIT('h8)
	) name12584 (
		_w16629_,
		_w16631_,
		_w16632_
	);
	LUT3 #(
		.INIT('h80)
	) name12585 (
		\CM_rd3[5]_pad ,
		_w16525_,
		_w16526_,
		_w16633_
	);
	LUT3 #(
		.INIT('h80)
	) name12586 (
		\CM_rd4[5]_pad ,
		_w16525_,
		_w16528_,
		_w16634_
	);
	LUT4 #(
		.INIT('h8000)
	) name12587 (
		\CM_rd1[5]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16635_
	);
	LUT4 #(
		.INIT('h8000)
	) name12588 (
		\CM_rd6[5]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16636_
	);
	LUT2 #(
		.INIT('h1)
	) name12589 (
		_w16635_,
		_w16636_,
		_w16637_
	);
	LUT3 #(
		.INIT('h10)
	) name12590 (
		_w16634_,
		_w16633_,
		_w16637_,
		_w16638_
	);
	LUT4 #(
		.INIT('h4555)
	) name12591 (
		\T_TMODE[1]_pad ,
		_w16626_,
		_w16632_,
		_w16638_,
		_w16639_
	);
	LUT3 #(
		.INIT('ha8)
	) name12592 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16625_,
		_w16639_,
		_w16640_
	);
	LUT3 #(
		.INIT('h80)
	) name12593 (
		\sice_SPC_reg[5]/P0001 ,
		_w16506_,
		_w16507_,
		_w16641_
	);
	LUT3 #(
		.INIT('h07)
	) name12594 (
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w16511_,
		_w16641_,
		_w16642_
	);
	LUT4 #(
		.INIT('h54ff)
	) name12595 (
		_w16511_,
		_w16624_,
		_w16640_,
		_w16642_,
		_w16643_
	);
	LUT4 #(
		.INIT('h4500)
	) name12596 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w16509_,
		_w16644_
	);
	LUT2 #(
		.INIT('h8)
	) name12597 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[4]/P0001 ,
		_w16645_
	);
	LUT4 #(
		.INIT('h2000)
	) name12598 (
		\CM_rdm[4]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16646_
	);
	LUT4 #(
		.INIT('h8000)
	) name12599 (
		\CM_rd0[4]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16647_
	);
	LUT4 #(
		.INIT('h8000)
	) name12600 (
		\CM_rd7[4]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16648_
	);
	LUT2 #(
		.INIT('h1)
	) name12601 (
		_w16647_,
		_w16648_,
		_w16649_
	);
	LUT4 #(
		.INIT('h8000)
	) name12602 (
		\CM_rd2[4]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16650_
	);
	LUT3 #(
		.INIT('h07)
	) name12603 (
		\CM_rd5[4]_pad ,
		_w16523_,
		_w16650_,
		_w16651_
	);
	LUT2 #(
		.INIT('h8)
	) name12604 (
		_w16649_,
		_w16651_,
		_w16652_
	);
	LUT3 #(
		.INIT('h80)
	) name12605 (
		\CM_rd3[4]_pad ,
		_w16525_,
		_w16526_,
		_w16653_
	);
	LUT3 #(
		.INIT('h80)
	) name12606 (
		\CM_rd4[4]_pad ,
		_w16525_,
		_w16528_,
		_w16654_
	);
	LUT4 #(
		.INIT('h8000)
	) name12607 (
		\CM_rd1[4]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16655_
	);
	LUT4 #(
		.INIT('h8000)
	) name12608 (
		\CM_rd6[4]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16656_
	);
	LUT2 #(
		.INIT('h1)
	) name12609 (
		_w16655_,
		_w16656_,
		_w16657_
	);
	LUT3 #(
		.INIT('h10)
	) name12610 (
		_w16654_,
		_w16653_,
		_w16657_,
		_w16658_
	);
	LUT4 #(
		.INIT('h4555)
	) name12611 (
		\T_TMODE[1]_pad ,
		_w16646_,
		_w16652_,
		_w16658_,
		_w16659_
	);
	LUT3 #(
		.INIT('ha8)
	) name12612 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16645_,
		_w16659_,
		_w16660_
	);
	LUT3 #(
		.INIT('h80)
	) name12613 (
		\sice_SPC_reg[4]/P0001 ,
		_w16506_,
		_w16507_,
		_w16661_
	);
	LUT3 #(
		.INIT('h07)
	) name12614 (
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w16511_,
		_w16661_,
		_w16662_
	);
	LUT4 #(
		.INIT('h54ff)
	) name12615 (
		_w16511_,
		_w16644_,
		_w16660_,
		_w16662_,
		_w16663_
	);
	LUT4 #(
		.INIT('h4500)
	) name12616 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w16509_,
		_w16664_
	);
	LUT2 #(
		.INIT('h8)
	) name12617 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[3]/P0001 ,
		_w16665_
	);
	LUT4 #(
		.INIT('h2000)
	) name12618 (
		\CM_rdm[3]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16666_
	);
	LUT4 #(
		.INIT('h8000)
	) name12619 (
		\CM_rd0[3]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16667_
	);
	LUT4 #(
		.INIT('h8000)
	) name12620 (
		\CM_rd7[3]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16668_
	);
	LUT2 #(
		.INIT('h1)
	) name12621 (
		_w16667_,
		_w16668_,
		_w16669_
	);
	LUT4 #(
		.INIT('h8000)
	) name12622 (
		\CM_rd2[3]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16670_
	);
	LUT3 #(
		.INIT('h07)
	) name12623 (
		\CM_rd5[3]_pad ,
		_w16523_,
		_w16670_,
		_w16671_
	);
	LUT2 #(
		.INIT('h8)
	) name12624 (
		_w16669_,
		_w16671_,
		_w16672_
	);
	LUT3 #(
		.INIT('h80)
	) name12625 (
		\CM_rd3[3]_pad ,
		_w16525_,
		_w16526_,
		_w16673_
	);
	LUT3 #(
		.INIT('h80)
	) name12626 (
		\CM_rd4[3]_pad ,
		_w16525_,
		_w16528_,
		_w16674_
	);
	LUT4 #(
		.INIT('h8000)
	) name12627 (
		\CM_rd1[3]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16675_
	);
	LUT4 #(
		.INIT('h8000)
	) name12628 (
		\CM_rd6[3]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16676_
	);
	LUT2 #(
		.INIT('h1)
	) name12629 (
		_w16675_,
		_w16676_,
		_w16677_
	);
	LUT3 #(
		.INIT('h10)
	) name12630 (
		_w16674_,
		_w16673_,
		_w16677_,
		_w16678_
	);
	LUT4 #(
		.INIT('h4555)
	) name12631 (
		\T_TMODE[1]_pad ,
		_w16666_,
		_w16672_,
		_w16678_,
		_w16679_
	);
	LUT3 #(
		.INIT('ha8)
	) name12632 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16665_,
		_w16679_,
		_w16680_
	);
	LUT3 #(
		.INIT('h80)
	) name12633 (
		\sice_SPC_reg[3]/P0001 ,
		_w16506_,
		_w16507_,
		_w16681_
	);
	LUT3 #(
		.INIT('h07)
	) name12634 (
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w16511_,
		_w16681_,
		_w16682_
	);
	LUT4 #(
		.INIT('h54ff)
	) name12635 (
		_w16511_,
		_w16664_,
		_w16680_,
		_w16682_,
		_w16683_
	);
	LUT4 #(
		.INIT('h4500)
	) name12636 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w16509_,
		_w16684_
	);
	LUT2 #(
		.INIT('h8)
	) name12637 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[2]/P0001 ,
		_w16685_
	);
	LUT4 #(
		.INIT('h2000)
	) name12638 (
		\CM_rdm[2]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16686_
	);
	LUT4 #(
		.INIT('h8000)
	) name12639 (
		\CM_rd0[2]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16687_
	);
	LUT4 #(
		.INIT('h8000)
	) name12640 (
		\CM_rd7[2]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16688_
	);
	LUT2 #(
		.INIT('h1)
	) name12641 (
		_w16687_,
		_w16688_,
		_w16689_
	);
	LUT4 #(
		.INIT('h8000)
	) name12642 (
		\CM_rd2[2]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16690_
	);
	LUT3 #(
		.INIT('h07)
	) name12643 (
		\CM_rd5[2]_pad ,
		_w16523_,
		_w16690_,
		_w16691_
	);
	LUT2 #(
		.INIT('h8)
	) name12644 (
		_w16689_,
		_w16691_,
		_w16692_
	);
	LUT3 #(
		.INIT('h80)
	) name12645 (
		\CM_rd3[2]_pad ,
		_w16525_,
		_w16526_,
		_w16693_
	);
	LUT3 #(
		.INIT('h80)
	) name12646 (
		\CM_rd4[2]_pad ,
		_w16525_,
		_w16528_,
		_w16694_
	);
	LUT4 #(
		.INIT('h8000)
	) name12647 (
		\CM_rd1[2]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16695_
	);
	LUT4 #(
		.INIT('h8000)
	) name12648 (
		\CM_rd6[2]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16696_
	);
	LUT2 #(
		.INIT('h1)
	) name12649 (
		_w16695_,
		_w16696_,
		_w16697_
	);
	LUT3 #(
		.INIT('h10)
	) name12650 (
		_w16694_,
		_w16693_,
		_w16697_,
		_w16698_
	);
	LUT4 #(
		.INIT('h4555)
	) name12651 (
		\T_TMODE[1]_pad ,
		_w16686_,
		_w16692_,
		_w16698_,
		_w16699_
	);
	LUT3 #(
		.INIT('ha8)
	) name12652 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16685_,
		_w16699_,
		_w16700_
	);
	LUT3 #(
		.INIT('h80)
	) name12653 (
		\sice_SPC_reg[2]/P0001 ,
		_w16506_,
		_w16507_,
		_w16701_
	);
	LUT3 #(
		.INIT('h07)
	) name12654 (
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w16511_,
		_w16701_,
		_w16702_
	);
	LUT4 #(
		.INIT('h54ff)
	) name12655 (
		_w16511_,
		_w16684_,
		_w16700_,
		_w16702_,
		_w16703_
	);
	LUT4 #(
		.INIT('h4500)
	) name12656 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w16509_,
		_w16704_
	);
	LUT2 #(
		.INIT('h8)
	) name12657 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[1]/P0001 ,
		_w16705_
	);
	LUT4 #(
		.INIT('h2000)
	) name12658 (
		\CM_rdm[1]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16706_
	);
	LUT4 #(
		.INIT('h8000)
	) name12659 (
		\CM_rd0[1]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16707_
	);
	LUT4 #(
		.INIT('h8000)
	) name12660 (
		\CM_rd7[1]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16708_
	);
	LUT2 #(
		.INIT('h1)
	) name12661 (
		_w16707_,
		_w16708_,
		_w16709_
	);
	LUT4 #(
		.INIT('h8000)
	) name12662 (
		\CM_rd2[1]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16710_
	);
	LUT3 #(
		.INIT('h07)
	) name12663 (
		\CM_rd5[1]_pad ,
		_w16523_,
		_w16710_,
		_w16711_
	);
	LUT2 #(
		.INIT('h8)
	) name12664 (
		_w16709_,
		_w16711_,
		_w16712_
	);
	LUT3 #(
		.INIT('h80)
	) name12665 (
		\CM_rd3[1]_pad ,
		_w16525_,
		_w16526_,
		_w16713_
	);
	LUT3 #(
		.INIT('h80)
	) name12666 (
		\CM_rd4[1]_pad ,
		_w16525_,
		_w16528_,
		_w16714_
	);
	LUT4 #(
		.INIT('h8000)
	) name12667 (
		\CM_rd1[1]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16715_
	);
	LUT4 #(
		.INIT('h8000)
	) name12668 (
		\CM_rd6[1]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16716_
	);
	LUT2 #(
		.INIT('h1)
	) name12669 (
		_w16715_,
		_w16716_,
		_w16717_
	);
	LUT3 #(
		.INIT('h10)
	) name12670 (
		_w16714_,
		_w16713_,
		_w16717_,
		_w16718_
	);
	LUT4 #(
		.INIT('h4555)
	) name12671 (
		\T_TMODE[1]_pad ,
		_w16706_,
		_w16712_,
		_w16718_,
		_w16719_
	);
	LUT3 #(
		.INIT('ha8)
	) name12672 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16705_,
		_w16719_,
		_w16720_
	);
	LUT3 #(
		.INIT('h80)
	) name12673 (
		\sice_SPC_reg[1]/P0001 ,
		_w16506_,
		_w16507_,
		_w16721_
	);
	LUT3 #(
		.INIT('h07)
	) name12674 (
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w16511_,
		_w16721_,
		_w16722_
	);
	LUT4 #(
		.INIT('h54ff)
	) name12675 (
		_w16511_,
		_w16704_,
		_w16720_,
		_w16722_,
		_w16723_
	);
	LUT4 #(
		.INIT('h4500)
	) name12676 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w16509_,
		_w16724_
	);
	LUT2 #(
		.INIT('h8)
	) name12677 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[0]/P0001 ,
		_w16725_
	);
	LUT4 #(
		.INIT('h2000)
	) name12678 (
		\CM_rdm[0]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16726_
	);
	LUT4 #(
		.INIT('h8000)
	) name12679 (
		\CM_rd0[0]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16727_
	);
	LUT4 #(
		.INIT('h8000)
	) name12680 (
		\CM_rd7[0]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16728_
	);
	LUT2 #(
		.INIT('h1)
	) name12681 (
		_w16727_,
		_w16728_,
		_w16729_
	);
	LUT4 #(
		.INIT('h8000)
	) name12682 (
		\CM_rd2[0]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16730_
	);
	LUT3 #(
		.INIT('h07)
	) name12683 (
		\CM_rd5[0]_pad ,
		_w16523_,
		_w16730_,
		_w16731_
	);
	LUT2 #(
		.INIT('h8)
	) name12684 (
		_w16729_,
		_w16731_,
		_w16732_
	);
	LUT3 #(
		.INIT('h80)
	) name12685 (
		\CM_rd3[0]_pad ,
		_w16525_,
		_w16526_,
		_w16733_
	);
	LUT3 #(
		.INIT('h80)
	) name12686 (
		\CM_rd4[0]_pad ,
		_w16525_,
		_w16528_,
		_w16734_
	);
	LUT4 #(
		.INIT('h8000)
	) name12687 (
		\CM_rd1[0]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16735_
	);
	LUT4 #(
		.INIT('h8000)
	) name12688 (
		\CM_rd6[0]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16736_
	);
	LUT2 #(
		.INIT('h1)
	) name12689 (
		_w16735_,
		_w16736_,
		_w16737_
	);
	LUT3 #(
		.INIT('h10)
	) name12690 (
		_w16734_,
		_w16733_,
		_w16737_,
		_w16738_
	);
	LUT4 #(
		.INIT('h4555)
	) name12691 (
		\T_TMODE[1]_pad ,
		_w16726_,
		_w16732_,
		_w16738_,
		_w16739_
	);
	LUT3 #(
		.INIT('ha8)
	) name12692 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16725_,
		_w16739_,
		_w16740_
	);
	LUT3 #(
		.INIT('h80)
	) name12693 (
		\sice_SPC_reg[0]/P0001 ,
		_w16506_,
		_w16507_,
		_w16741_
	);
	LUT3 #(
		.INIT('h07)
	) name12694 (
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w16511_,
		_w16741_,
		_w16742_
	);
	LUT4 #(
		.INIT('h54ff)
	) name12695 (
		_w16511_,
		_w16724_,
		_w16740_,
		_w16742_,
		_w16743_
	);
	LUT2 #(
		.INIT('h2)
	) name12696 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001 ,
		_w11310_,
		_w16744_
	);
	LUT3 #(
		.INIT('h01)
	) name12697 (
		_w9946_,
		_w12442_,
		_w16744_,
		_w16745_
	);
	LUT4 #(
		.INIT('hef00)
	) name12698 (
		_w12006_,
		_w12007_,
		_w12440_,
		_w16745_,
		_w16746_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12699 (
		_w9946_,
		_w16558_,
		_w16561_,
		_w16746_,
		_w16747_
	);
	LUT2 #(
		.INIT('h8)
	) name12700 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[13]/P0001 ,
		_w16748_
	);
	LUT4 #(
		.INIT('h2000)
	) name12701 (
		\CM_rdm[13]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16749_
	);
	LUT4 #(
		.INIT('h8000)
	) name12702 (
		\CM_rd0[13]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16750_
	);
	LUT4 #(
		.INIT('h8000)
	) name12703 (
		\CM_rd7[13]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16751_
	);
	LUT2 #(
		.INIT('h1)
	) name12704 (
		_w16750_,
		_w16751_,
		_w16752_
	);
	LUT4 #(
		.INIT('h8000)
	) name12705 (
		\CM_rd2[13]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16753_
	);
	LUT3 #(
		.INIT('h07)
	) name12706 (
		\CM_rd5[13]_pad ,
		_w16523_,
		_w16753_,
		_w16754_
	);
	LUT2 #(
		.INIT('h8)
	) name12707 (
		_w16752_,
		_w16754_,
		_w16755_
	);
	LUT3 #(
		.INIT('h80)
	) name12708 (
		\CM_rd3[13]_pad ,
		_w16525_,
		_w16526_,
		_w16756_
	);
	LUT3 #(
		.INIT('h80)
	) name12709 (
		\CM_rd4[13]_pad ,
		_w16525_,
		_w16528_,
		_w16757_
	);
	LUT4 #(
		.INIT('h8000)
	) name12710 (
		\CM_rd1[13]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16758_
	);
	LUT4 #(
		.INIT('h8000)
	) name12711 (
		\CM_rd6[13]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16759_
	);
	LUT2 #(
		.INIT('h1)
	) name12712 (
		_w16758_,
		_w16759_,
		_w16760_
	);
	LUT3 #(
		.INIT('h10)
	) name12713 (
		_w16757_,
		_w16756_,
		_w16760_,
		_w16761_
	);
	LUT4 #(
		.INIT('h4555)
	) name12714 (
		\T_TMODE[1]_pad ,
		_w16749_,
		_w16755_,
		_w16761_,
		_w16762_
	);
	LUT3 #(
		.INIT('ha8)
	) name12715 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16748_,
		_w16762_,
		_w16763_
	);
	LUT4 #(
		.INIT('h0f08)
	) name12716 (
		_w5760_,
		_w16509_,
		_w16511_,
		_w16763_,
		_w16764_
	);
	LUT3 #(
		.INIT('h80)
	) name12717 (
		\sice_SPC_reg[13]/P0001 ,
		_w16506_,
		_w16507_,
		_w16765_
	);
	LUT3 #(
		.INIT('h07)
	) name12718 (
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w16511_,
		_w16765_,
		_w16766_
	);
	LUT2 #(
		.INIT('hb)
	) name12719 (
		_w16764_,
		_w16766_,
		_w16767_
	);
	LUT2 #(
		.INIT('h8)
	) name12720 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[12]/P0001 ,
		_w16768_
	);
	LUT4 #(
		.INIT('h2000)
	) name12721 (
		\CM_rdm[12]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16769_
	);
	LUT4 #(
		.INIT('h8000)
	) name12722 (
		\CM_rd0[12]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16770_
	);
	LUT4 #(
		.INIT('h8000)
	) name12723 (
		\CM_rd7[12]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16771_
	);
	LUT2 #(
		.INIT('h1)
	) name12724 (
		_w16770_,
		_w16771_,
		_w16772_
	);
	LUT4 #(
		.INIT('h8000)
	) name12725 (
		\CM_rd2[12]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16773_
	);
	LUT3 #(
		.INIT('h07)
	) name12726 (
		\CM_rd5[12]_pad ,
		_w16523_,
		_w16773_,
		_w16774_
	);
	LUT2 #(
		.INIT('h8)
	) name12727 (
		_w16772_,
		_w16774_,
		_w16775_
	);
	LUT3 #(
		.INIT('h80)
	) name12728 (
		\CM_rd3[12]_pad ,
		_w16525_,
		_w16526_,
		_w16776_
	);
	LUT3 #(
		.INIT('h80)
	) name12729 (
		\CM_rd4[12]_pad ,
		_w16525_,
		_w16528_,
		_w16777_
	);
	LUT4 #(
		.INIT('h8000)
	) name12730 (
		\CM_rd1[12]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16778_
	);
	LUT4 #(
		.INIT('h8000)
	) name12731 (
		\CM_rd6[12]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16779_
	);
	LUT2 #(
		.INIT('h1)
	) name12732 (
		_w16778_,
		_w16779_,
		_w16780_
	);
	LUT3 #(
		.INIT('h10)
	) name12733 (
		_w16777_,
		_w16776_,
		_w16780_,
		_w16781_
	);
	LUT4 #(
		.INIT('h4555)
	) name12734 (
		\T_TMODE[1]_pad ,
		_w16769_,
		_w16775_,
		_w16781_,
		_w16782_
	);
	LUT3 #(
		.INIT('ha8)
	) name12735 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16768_,
		_w16782_,
		_w16783_
	);
	LUT4 #(
		.INIT('h0f08)
	) name12736 (
		_w6758_,
		_w16509_,
		_w16511_,
		_w16783_,
		_w16784_
	);
	LUT3 #(
		.INIT('h80)
	) name12737 (
		\sice_SPC_reg[12]/P0001 ,
		_w16506_,
		_w16507_,
		_w16785_
	);
	LUT3 #(
		.INIT('h07)
	) name12738 (
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w16511_,
		_w16785_,
		_w16786_
	);
	LUT2 #(
		.INIT('hb)
	) name12739 (
		_w16784_,
		_w16786_,
		_w16787_
	);
	LUT2 #(
		.INIT('h8)
	) name12740 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[8]/P0001 ,
		_w16788_
	);
	LUT4 #(
		.INIT('h2000)
	) name12741 (
		\CM_rdm[8]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16789_
	);
	LUT4 #(
		.INIT('h8000)
	) name12742 (
		\CM_rd0[8]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16790_
	);
	LUT4 #(
		.INIT('h8000)
	) name12743 (
		\CM_rd7[8]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16791_
	);
	LUT2 #(
		.INIT('h1)
	) name12744 (
		_w16790_,
		_w16791_,
		_w16792_
	);
	LUT4 #(
		.INIT('h8000)
	) name12745 (
		\CM_rd2[8]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16793_
	);
	LUT3 #(
		.INIT('h07)
	) name12746 (
		\CM_rd5[8]_pad ,
		_w16523_,
		_w16793_,
		_w16794_
	);
	LUT2 #(
		.INIT('h8)
	) name12747 (
		_w16792_,
		_w16794_,
		_w16795_
	);
	LUT3 #(
		.INIT('h80)
	) name12748 (
		\CM_rd3[8]_pad ,
		_w16525_,
		_w16526_,
		_w16796_
	);
	LUT3 #(
		.INIT('h80)
	) name12749 (
		\CM_rd4[8]_pad ,
		_w16525_,
		_w16528_,
		_w16797_
	);
	LUT4 #(
		.INIT('h8000)
	) name12750 (
		\CM_rd1[8]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16798_
	);
	LUT4 #(
		.INIT('h8000)
	) name12751 (
		\CM_rd6[8]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16799_
	);
	LUT2 #(
		.INIT('h1)
	) name12752 (
		_w16798_,
		_w16799_,
		_w16800_
	);
	LUT3 #(
		.INIT('h10)
	) name12753 (
		_w16797_,
		_w16796_,
		_w16800_,
		_w16801_
	);
	LUT4 #(
		.INIT('h4555)
	) name12754 (
		\T_TMODE[1]_pad ,
		_w16789_,
		_w16795_,
		_w16801_,
		_w16802_
	);
	LUT3 #(
		.INIT('ha8)
	) name12755 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16788_,
		_w16802_,
		_w16803_
	);
	LUT4 #(
		.INIT('h00ef)
	) name12756 (
		_w7465_,
		_w7565_,
		_w16509_,
		_w16803_,
		_w16804_
	);
	LUT3 #(
		.INIT('h80)
	) name12757 (
		\sice_SPC_reg[8]/P0001 ,
		_w16506_,
		_w16507_,
		_w16805_
	);
	LUT3 #(
		.INIT('h07)
	) name12758 (
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w16511_,
		_w16805_,
		_w16806_
	);
	LUT3 #(
		.INIT('h1f)
	) name12759 (
		_w16511_,
		_w16804_,
		_w16806_,
		_w16807_
	);
	LUT2 #(
		.INIT('h8)
	) name12760 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[9]/P0001 ,
		_w16808_
	);
	LUT4 #(
		.INIT('h2000)
	) name12761 (
		\CM_rdm[9]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16809_
	);
	LUT4 #(
		.INIT('h8000)
	) name12762 (
		\CM_rd0[9]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16810_
	);
	LUT4 #(
		.INIT('h8000)
	) name12763 (
		\CM_rd7[9]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16811_
	);
	LUT2 #(
		.INIT('h1)
	) name12764 (
		_w16810_,
		_w16811_,
		_w16812_
	);
	LUT4 #(
		.INIT('h8000)
	) name12765 (
		\CM_rd2[9]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16813_
	);
	LUT3 #(
		.INIT('h07)
	) name12766 (
		\CM_rd5[9]_pad ,
		_w16523_,
		_w16813_,
		_w16814_
	);
	LUT2 #(
		.INIT('h8)
	) name12767 (
		_w16812_,
		_w16814_,
		_w16815_
	);
	LUT3 #(
		.INIT('h80)
	) name12768 (
		\CM_rd3[9]_pad ,
		_w16525_,
		_w16526_,
		_w16816_
	);
	LUT3 #(
		.INIT('h80)
	) name12769 (
		\CM_rd4[9]_pad ,
		_w16525_,
		_w16528_,
		_w16817_
	);
	LUT4 #(
		.INIT('h8000)
	) name12770 (
		\CM_rd1[9]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16818_
	);
	LUT4 #(
		.INIT('h8000)
	) name12771 (
		\CM_rd6[9]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16819_
	);
	LUT2 #(
		.INIT('h1)
	) name12772 (
		_w16818_,
		_w16819_,
		_w16820_
	);
	LUT3 #(
		.INIT('h10)
	) name12773 (
		_w16817_,
		_w16816_,
		_w16820_,
		_w16821_
	);
	LUT4 #(
		.INIT('h4555)
	) name12774 (
		\T_TMODE[1]_pad ,
		_w16809_,
		_w16815_,
		_w16821_,
		_w16822_
	);
	LUT3 #(
		.INIT('ha8)
	) name12775 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16808_,
		_w16822_,
		_w16823_
	);
	LUT4 #(
		.INIT('h00ef)
	) name12776 (
		_w7140_,
		_w7240_,
		_w16509_,
		_w16823_,
		_w16824_
	);
	LUT3 #(
		.INIT('h80)
	) name12777 (
		\sice_SPC_reg[9]/P0001 ,
		_w16506_,
		_w16507_,
		_w16825_
	);
	LUT3 #(
		.INIT('h07)
	) name12778 (
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w16511_,
		_w16825_,
		_w16826_
	);
	LUT3 #(
		.INIT('h1f)
	) name12779 (
		_w16511_,
		_w16824_,
		_w16826_,
		_w16827_
	);
	LUT2 #(
		.INIT('h8)
	) name12780 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[11]/P0001 ,
		_w16828_
	);
	LUT4 #(
		.INIT('h2000)
	) name12781 (
		\CM_rdm[11]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16829_
	);
	LUT4 #(
		.INIT('h8000)
	) name12782 (
		\CM_rd0[11]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16830_
	);
	LUT4 #(
		.INIT('h8000)
	) name12783 (
		\CM_rd7[11]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16831_
	);
	LUT2 #(
		.INIT('h1)
	) name12784 (
		_w16830_,
		_w16831_,
		_w16832_
	);
	LUT4 #(
		.INIT('h8000)
	) name12785 (
		\CM_rd2[11]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16833_
	);
	LUT3 #(
		.INIT('h07)
	) name12786 (
		\CM_rd5[11]_pad ,
		_w16523_,
		_w16833_,
		_w16834_
	);
	LUT2 #(
		.INIT('h8)
	) name12787 (
		_w16832_,
		_w16834_,
		_w16835_
	);
	LUT3 #(
		.INIT('h80)
	) name12788 (
		\CM_rd3[11]_pad ,
		_w16525_,
		_w16526_,
		_w16836_
	);
	LUT3 #(
		.INIT('h80)
	) name12789 (
		\CM_rd4[11]_pad ,
		_w16525_,
		_w16528_,
		_w16837_
	);
	LUT4 #(
		.INIT('h8000)
	) name12790 (
		\CM_rd1[11]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16838_
	);
	LUT4 #(
		.INIT('h8000)
	) name12791 (
		\CM_rd6[11]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16839_
	);
	LUT2 #(
		.INIT('h1)
	) name12792 (
		_w16838_,
		_w16839_,
		_w16840_
	);
	LUT3 #(
		.INIT('h10)
	) name12793 (
		_w16837_,
		_w16836_,
		_w16840_,
		_w16841_
	);
	LUT4 #(
		.INIT('h4555)
	) name12794 (
		\T_TMODE[1]_pad ,
		_w16829_,
		_w16835_,
		_w16841_,
		_w16842_
	);
	LUT3 #(
		.INIT('ha8)
	) name12795 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16828_,
		_w16842_,
		_w16843_
	);
	LUT4 #(
		.INIT('h00ef)
	) name12796 (
		_w6263_,
		_w6362_,
		_w16509_,
		_w16843_,
		_w16844_
	);
	LUT3 #(
		.INIT('h80)
	) name12797 (
		\sice_SPC_reg[11]/P0001 ,
		_w16506_,
		_w16507_,
		_w16845_
	);
	LUT3 #(
		.INIT('h07)
	) name12798 (
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w16511_,
		_w16845_,
		_w16846_
	);
	LUT3 #(
		.INIT('h1f)
	) name12799 (
		_w16511_,
		_w16844_,
		_w16846_,
		_w16847_
	);
	LUT2 #(
		.INIT('h8)
	) name12800 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[10]/P0001 ,
		_w16848_
	);
	LUT4 #(
		.INIT('h2000)
	) name12801 (
		\CM_rdm[10]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16849_
	);
	LUT4 #(
		.INIT('h8000)
	) name12802 (
		\CM_rd0[10]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16850_
	);
	LUT4 #(
		.INIT('h8000)
	) name12803 (
		\CM_rd7[10]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16851_
	);
	LUT2 #(
		.INIT('h1)
	) name12804 (
		_w16850_,
		_w16851_,
		_w16852_
	);
	LUT4 #(
		.INIT('h8000)
	) name12805 (
		\CM_rd2[10]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16853_
	);
	LUT3 #(
		.INIT('h07)
	) name12806 (
		\CM_rd5[10]_pad ,
		_w16523_,
		_w16853_,
		_w16854_
	);
	LUT2 #(
		.INIT('h8)
	) name12807 (
		_w16852_,
		_w16854_,
		_w16855_
	);
	LUT3 #(
		.INIT('h80)
	) name12808 (
		\CM_rd3[10]_pad ,
		_w16525_,
		_w16526_,
		_w16856_
	);
	LUT3 #(
		.INIT('h80)
	) name12809 (
		\CM_rd4[10]_pad ,
		_w16525_,
		_w16528_,
		_w16857_
	);
	LUT4 #(
		.INIT('h8000)
	) name12810 (
		\CM_rd1[10]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16858_
	);
	LUT4 #(
		.INIT('h8000)
	) name12811 (
		\CM_rd6[10]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16859_
	);
	LUT2 #(
		.INIT('h1)
	) name12812 (
		_w16858_,
		_w16859_,
		_w16860_
	);
	LUT3 #(
		.INIT('h10)
	) name12813 (
		_w16857_,
		_w16856_,
		_w16860_,
		_w16861_
	);
	LUT4 #(
		.INIT('h4555)
	) name12814 (
		\T_TMODE[1]_pad ,
		_w16849_,
		_w16855_,
		_w16861_,
		_w16862_
	);
	LUT3 #(
		.INIT('ha8)
	) name12815 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w16848_,
		_w16862_,
		_w16863_
	);
	LUT4 #(
		.INIT('h00ef)
	) name12816 (
		_w5937_,
		_w6038_,
		_w16509_,
		_w16863_,
		_w16864_
	);
	LUT3 #(
		.INIT('h80)
	) name12817 (
		\sice_SPC_reg[10]/P0001 ,
		_w16506_,
		_w16507_,
		_w16865_
	);
	LUT3 #(
		.INIT('h07)
	) name12818 (
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w16511_,
		_w16865_,
		_w16866_
	);
	LUT3 #(
		.INIT('h1f)
	) name12819 (
		_w16511_,
		_w16864_,
		_w16866_,
		_w16867_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12820 (
		_w16238_,
		_w16239_,
		_w16240_,
		_w16243_,
		_w16868_
	);
	LUT2 #(
		.INIT('h8)
	) name12821 (
		_w16244_,
		_w16246_,
		_w16869_
	);
	LUT4 #(
		.INIT('h1511)
	) name12822 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w16247_,
		_w16868_,
		_w16869_,
		_w16870_
	);
	LUT4 #(
		.INIT('h0057)
	) name12823 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w11313_,
		_w11314_,
		_w16870_,
		_w16871_
	);
	LUT3 #(
		.INIT('he2)
	) name12824 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001 ,
		_w14809_,
		_w16871_,
		_w16872_
	);
	LUT3 #(
		.INIT('he2)
	) name12825 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001 ,
		_w14780_,
		_w16871_,
		_w16873_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12826 (
		_w9326_,
		_w16534_,
		_w16540_,
		_w16546_,
		_w16874_
	);
	LUT2 #(
		.INIT('h4)
	) name12827 (
		_w4937_,
		_w9326_,
		_w16875_
	);
	LUT3 #(
		.INIT('h8a)
	) name12828 (
		\idma_IADi_reg[7]/P0001 ,
		_w4937_,
		_w9326_,
		_w16876_
	);
	LUT3 #(
		.INIT('h35)
	) name12829 (
		\idma_IADi_reg[7]/P0001 ,
		_w4937_,
		_w9326_,
		_w16877_
	);
	LUT2 #(
		.INIT('h4)
	) name12830 (
		_w16874_,
		_w16877_,
		_w16878_
	);
	LUT3 #(
		.INIT('h45)
	) name12831 (
		_w8182_,
		_w8974_,
		_w9327_,
		_w16879_
	);
	LUT2 #(
		.INIT('h4)
	) name12832 (
		_w16878_,
		_w16879_,
		_w16880_
	);
	LUT4 #(
		.INIT('h4500)
	) name12833 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w8182_,
		_w16881_
	);
	LUT2 #(
		.INIT('he)
	) name12834 (
		_w16880_,
		_w16881_,
		_w16882_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12835 (
		_w9326_,
		_w16565_,
		_w16571_,
		_w16577_,
		_w16883_
	);
	LUT3 #(
		.INIT('h8a)
	) name12836 (
		\idma_IADi_reg[6]/P0001 ,
		_w4937_,
		_w9326_,
		_w16884_
	);
	LUT3 #(
		.INIT('h35)
	) name12837 (
		\idma_IADi_reg[6]/P0001 ,
		_w4937_,
		_w9326_,
		_w16885_
	);
	LUT3 #(
		.INIT('h45)
	) name12838 (
		_w8182_,
		_w16883_,
		_w16885_,
		_w16886_
	);
	LUT3 #(
		.INIT('hb0)
	) name12839 (
		_w8952_,
		_w9327_,
		_w16886_,
		_w16887_
	);
	LUT4 #(
		.INIT('h4500)
	) name12840 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w8182_,
		_w16888_
	);
	LUT2 #(
		.INIT('he)
	) name12841 (
		_w16887_,
		_w16888_,
		_w16889_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12842 (
		_w9326_,
		_w16749_,
		_w16755_,
		_w16761_,
		_w16890_
	);
	LUT3 #(
		.INIT('h8a)
	) name12843 (
		\idma_IADi_reg[5]/P0001 ,
		_w4937_,
		_w9326_,
		_w16891_
	);
	LUT3 #(
		.INIT('h35)
	) name12844 (
		\idma_IADi_reg[5]/P0001 ,
		_w4937_,
		_w9326_,
		_w16892_
	);
	LUT2 #(
		.INIT('h4)
	) name12845 (
		_w16890_,
		_w16892_,
		_w16893_
	);
	LUT3 #(
		.INIT('h45)
	) name12846 (
		_w8182_,
		_w8929_,
		_w9327_,
		_w16894_
	);
	LUT2 #(
		.INIT('h4)
	) name12847 (
		_w16893_,
		_w16894_,
		_w16895_
	);
	LUT4 #(
		.INIT('h4500)
	) name12848 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w8182_,
		_w16896_
	);
	LUT2 #(
		.INIT('he)
	) name12849 (
		_w16895_,
		_w16896_,
		_w16897_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12850 (
		_w9326_,
		_w16769_,
		_w16775_,
		_w16781_,
		_w16898_
	);
	LUT3 #(
		.INIT('h8a)
	) name12851 (
		\idma_IADi_reg[4]/P0001 ,
		_w4937_,
		_w9326_,
		_w16899_
	);
	LUT3 #(
		.INIT('h35)
	) name12852 (
		\idma_IADi_reg[4]/P0001 ,
		_w4937_,
		_w9326_,
		_w16900_
	);
	LUT2 #(
		.INIT('h4)
	) name12853 (
		_w16898_,
		_w16900_,
		_w16901_
	);
	LUT3 #(
		.INIT('h45)
	) name12854 (
		_w8182_,
		_w8907_,
		_w9327_,
		_w16902_
	);
	LUT2 #(
		.INIT('h4)
	) name12855 (
		_w16901_,
		_w16902_,
		_w16903_
	);
	LUT4 #(
		.INIT('h4500)
	) name12856 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w8182_,
		_w16904_
	);
	LUT2 #(
		.INIT('he)
	) name12857 (
		_w16903_,
		_w16904_,
		_w16905_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12858 (
		_w9326_,
		_w16829_,
		_w16835_,
		_w16841_,
		_w16906_
	);
	LUT3 #(
		.INIT('h8a)
	) name12859 (
		\idma_IADi_reg[3]/P0001 ,
		_w4937_,
		_w9326_,
		_w16907_
	);
	LUT3 #(
		.INIT('h35)
	) name12860 (
		\idma_IADi_reg[3]/P0001 ,
		_w4937_,
		_w9326_,
		_w16908_
	);
	LUT2 #(
		.INIT('h4)
	) name12861 (
		_w16906_,
		_w16908_,
		_w16909_
	);
	LUT3 #(
		.INIT('h45)
	) name12862 (
		_w8182_,
		_w8885_,
		_w9327_,
		_w16910_
	);
	LUT2 #(
		.INIT('h4)
	) name12863 (
		_w16909_,
		_w16910_,
		_w16911_
	);
	LUT4 #(
		.INIT('h4500)
	) name12864 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w8182_,
		_w16912_
	);
	LUT2 #(
		.INIT('he)
	) name12865 (
		_w16911_,
		_w16912_,
		_w16913_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12866 (
		_w9326_,
		_w16849_,
		_w16855_,
		_w16861_,
		_w16914_
	);
	LUT3 #(
		.INIT('h8a)
	) name12867 (
		\idma_IADi_reg[2]/P0001 ,
		_w4937_,
		_w9326_,
		_w16915_
	);
	LUT3 #(
		.INIT('h35)
	) name12868 (
		\idma_IADi_reg[2]/P0001 ,
		_w4937_,
		_w9326_,
		_w16916_
	);
	LUT2 #(
		.INIT('h4)
	) name12869 (
		_w16914_,
		_w16916_,
		_w16917_
	);
	LUT3 #(
		.INIT('h45)
	) name12870 (
		_w8182_,
		_w8863_,
		_w9327_,
		_w16918_
	);
	LUT2 #(
		.INIT('h4)
	) name12871 (
		_w16917_,
		_w16918_,
		_w16919_
	);
	LUT4 #(
		.INIT('h4500)
	) name12872 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w8182_,
		_w16920_
	);
	LUT2 #(
		.INIT('he)
	) name12873 (
		_w16919_,
		_w16920_,
		_w16921_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12874 (
		_w9326_,
		_w16809_,
		_w16815_,
		_w16821_,
		_w16922_
	);
	LUT3 #(
		.INIT('h8a)
	) name12875 (
		\idma_IADi_reg[1]/P0001 ,
		_w4937_,
		_w9326_,
		_w16923_
	);
	LUT3 #(
		.INIT('h35)
	) name12876 (
		\idma_IADi_reg[1]/P0001 ,
		_w4937_,
		_w9326_,
		_w16924_
	);
	LUT2 #(
		.INIT('h4)
	) name12877 (
		_w16922_,
		_w16924_,
		_w16925_
	);
	LUT3 #(
		.INIT('h45)
	) name12878 (
		_w8182_,
		_w8841_,
		_w9327_,
		_w16926_
	);
	LUT2 #(
		.INIT('h4)
	) name12879 (
		_w16925_,
		_w16926_,
		_w16927_
	);
	LUT4 #(
		.INIT('h4500)
	) name12880 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w8182_,
		_w16928_
	);
	LUT2 #(
		.INIT('he)
	) name12881 (
		_w16927_,
		_w16928_,
		_w16929_
	);
	LUT4 #(
		.INIT('h2000)
	) name12882 (
		\CM_rdm[23]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16930_
	);
	LUT4 #(
		.INIT('h8000)
	) name12883 (
		\CM_rd0[23]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16931_
	);
	LUT4 #(
		.INIT('h8000)
	) name12884 (
		\CM_rd7[23]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16932_
	);
	LUT2 #(
		.INIT('h1)
	) name12885 (
		_w16931_,
		_w16932_,
		_w16933_
	);
	LUT4 #(
		.INIT('h8000)
	) name12886 (
		\CM_rd2[23]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16934_
	);
	LUT3 #(
		.INIT('h07)
	) name12887 (
		\CM_rd5[23]_pad ,
		_w16523_,
		_w16934_,
		_w16935_
	);
	LUT2 #(
		.INIT('h8)
	) name12888 (
		_w16933_,
		_w16935_,
		_w16936_
	);
	LUT3 #(
		.INIT('h80)
	) name12889 (
		\CM_rd3[23]_pad ,
		_w16525_,
		_w16526_,
		_w16937_
	);
	LUT3 #(
		.INIT('h80)
	) name12890 (
		\CM_rd4[23]_pad ,
		_w16525_,
		_w16528_,
		_w16938_
	);
	LUT4 #(
		.INIT('h8000)
	) name12891 (
		\CM_rd1[23]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16939_
	);
	LUT4 #(
		.INIT('h8000)
	) name12892 (
		\CM_rd6[23]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16940_
	);
	LUT2 #(
		.INIT('h1)
	) name12893 (
		_w16939_,
		_w16940_,
		_w16941_
	);
	LUT3 #(
		.INIT('h10)
	) name12894 (
		_w16938_,
		_w16937_,
		_w16941_,
		_w16942_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12895 (
		_w16875_,
		_w16930_,
		_w16936_,
		_w16942_,
		_w16943_
	);
	LUT3 #(
		.INIT('h8a)
	) name12896 (
		\idma_IADi_reg[15]/P0001 ,
		_w4937_,
		_w9326_,
		_w16944_
	);
	LUT4 #(
		.INIT('h4447)
	) name12897 (
		_w8821_,
		_w9327_,
		_w16943_,
		_w16944_,
		_w16945_
	);
	LUT4 #(
		.INIT('h0257)
	) name12898 (
		_w8182_,
		_w8798_,
		_w8801_,
		_w16945_,
		_w16946_
	);
	LUT4 #(
		.INIT('h2000)
	) name12899 (
		\CM_rdm[22]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16947_
	);
	LUT4 #(
		.INIT('h8000)
	) name12900 (
		\CM_rd0[22]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16948_
	);
	LUT4 #(
		.INIT('h8000)
	) name12901 (
		\CM_rd7[22]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16949_
	);
	LUT2 #(
		.INIT('h1)
	) name12902 (
		_w16948_,
		_w16949_,
		_w16950_
	);
	LUT4 #(
		.INIT('h8000)
	) name12903 (
		\CM_rd2[22]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16951_
	);
	LUT3 #(
		.INIT('h07)
	) name12904 (
		\CM_rd5[22]_pad ,
		_w16523_,
		_w16951_,
		_w16952_
	);
	LUT2 #(
		.INIT('h8)
	) name12905 (
		_w16950_,
		_w16952_,
		_w16953_
	);
	LUT3 #(
		.INIT('h80)
	) name12906 (
		\CM_rd3[22]_pad ,
		_w16525_,
		_w16526_,
		_w16954_
	);
	LUT3 #(
		.INIT('h80)
	) name12907 (
		\CM_rd4[22]_pad ,
		_w16525_,
		_w16528_,
		_w16955_
	);
	LUT4 #(
		.INIT('h8000)
	) name12908 (
		\CM_rd1[22]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16956_
	);
	LUT4 #(
		.INIT('h8000)
	) name12909 (
		\CM_rd6[22]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16957_
	);
	LUT2 #(
		.INIT('h1)
	) name12910 (
		_w16956_,
		_w16957_,
		_w16958_
	);
	LUT3 #(
		.INIT('h10)
	) name12911 (
		_w16955_,
		_w16954_,
		_w16958_,
		_w16959_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12912 (
		_w16875_,
		_w16947_,
		_w16953_,
		_w16959_,
		_w16960_
	);
	LUT3 #(
		.INIT('h8a)
	) name12913 (
		\idma_IADi_reg[14]/P0001 ,
		_w4937_,
		_w9326_,
		_w16961_
	);
	LUT4 #(
		.INIT('h4447)
	) name12914 (
		_w8781_,
		_w9327_,
		_w16960_,
		_w16961_,
		_w16962_
	);
	LUT4 #(
		.INIT('h0257)
	) name12915 (
		_w8182_,
		_w8757_,
		_w8760_,
		_w16962_,
		_w16963_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12916 (
		_w9326_,
		_w16789_,
		_w16795_,
		_w16801_,
		_w16964_
	);
	LUT3 #(
		.INIT('h8a)
	) name12917 (
		\idma_IADi_reg[0]/P0001 ,
		_w4937_,
		_w9326_,
		_w16965_
	);
	LUT3 #(
		.INIT('h35)
	) name12918 (
		\idma_IADi_reg[0]/P0001 ,
		_w4937_,
		_w9326_,
		_w16966_
	);
	LUT2 #(
		.INIT('h4)
	) name12919 (
		_w16964_,
		_w16966_,
		_w16967_
	);
	LUT3 #(
		.INIT('h45)
	) name12920 (
		_w8182_,
		_w8647_,
		_w9327_,
		_w16968_
	);
	LUT2 #(
		.INIT('h4)
	) name12921 (
		_w16967_,
		_w16968_,
		_w16969_
	);
	LUT4 #(
		.INIT('h4500)
	) name12922 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w8182_,
		_w16970_
	);
	LUT2 #(
		.INIT('he)
	) name12923 (
		_w16969_,
		_w16970_,
		_w16971_
	);
	LUT4 #(
		.INIT('h0102)
	) name12924 (
		\tm_TSR_TMP_reg[5]/NET0131 ,
		_w12802_,
		_w15792_,
		_w15794_,
		_w16972_
	);
	LUT3 #(
		.INIT('ha8)
	) name12925 (
		\tm_tsr_reg_DO_reg[5]/NET0131 ,
		_w12802_,
		_w15792_,
		_w16973_
	);
	LUT2 #(
		.INIT('he)
	) name12926 (
		_w16972_,
		_w16973_,
		_w16974_
	);
	LUT4 #(
		.INIT('h2000)
	) name12927 (
		\CM_rdm[17]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16975_
	);
	LUT4 #(
		.INIT('h8000)
	) name12928 (
		\CM_rd0[17]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16976_
	);
	LUT4 #(
		.INIT('h8000)
	) name12929 (
		\CM_rd7[17]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16977_
	);
	LUT2 #(
		.INIT('h1)
	) name12930 (
		_w16976_,
		_w16977_,
		_w16978_
	);
	LUT4 #(
		.INIT('h8000)
	) name12931 (
		\CM_rd2[17]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16979_
	);
	LUT3 #(
		.INIT('h07)
	) name12932 (
		\CM_rd5[17]_pad ,
		_w16523_,
		_w16979_,
		_w16980_
	);
	LUT2 #(
		.INIT('h8)
	) name12933 (
		_w16978_,
		_w16980_,
		_w16981_
	);
	LUT3 #(
		.INIT('h80)
	) name12934 (
		\CM_rd3[17]_pad ,
		_w16525_,
		_w16526_,
		_w16982_
	);
	LUT3 #(
		.INIT('h80)
	) name12935 (
		\CM_rd4[17]_pad ,
		_w16525_,
		_w16528_,
		_w16983_
	);
	LUT4 #(
		.INIT('h8000)
	) name12936 (
		\CM_rd1[17]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w16984_
	);
	LUT4 #(
		.INIT('h8000)
	) name12937 (
		\CM_rd6[17]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w16985_
	);
	LUT2 #(
		.INIT('h1)
	) name12938 (
		_w16984_,
		_w16985_,
		_w16986_
	);
	LUT3 #(
		.INIT('h10)
	) name12939 (
		_w16983_,
		_w16982_,
		_w16986_,
		_w16987_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12940 (
		_w16875_,
		_w16975_,
		_w16981_,
		_w16987_,
		_w16988_
	);
	LUT3 #(
		.INIT('h8a)
	) name12941 (
		\idma_IADi_reg[9]/P0001 ,
		_w4937_,
		_w9326_,
		_w16989_
	);
	LUT4 #(
		.INIT('h4447)
	) name12942 (
		_w9021_,
		_w9327_,
		_w16988_,
		_w16989_,
		_w16990_
	);
	LUT2 #(
		.INIT('h1)
	) name12943 (
		_w8182_,
		_w16990_,
		_w16991_
	);
	LUT4 #(
		.INIT('hff10)
	) name12944 (
		_w7140_,
		_w7240_,
		_w8182_,
		_w16991_,
		_w16992_
	);
	LUT4 #(
		.INIT('h2000)
	) name12945 (
		\CM_rdm[16]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w16993_
	);
	LUT4 #(
		.INIT('h8000)
	) name12946 (
		\CM_rd0[16]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w16994_
	);
	LUT4 #(
		.INIT('h8000)
	) name12947 (
		\CM_rd7[16]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w16995_
	);
	LUT2 #(
		.INIT('h1)
	) name12948 (
		_w16994_,
		_w16995_,
		_w16996_
	);
	LUT4 #(
		.INIT('h8000)
	) name12949 (
		\CM_rd2[16]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w16997_
	);
	LUT3 #(
		.INIT('h07)
	) name12950 (
		\CM_rd5[16]_pad ,
		_w16523_,
		_w16997_,
		_w16998_
	);
	LUT2 #(
		.INIT('h8)
	) name12951 (
		_w16996_,
		_w16998_,
		_w16999_
	);
	LUT3 #(
		.INIT('h80)
	) name12952 (
		\CM_rd3[16]_pad ,
		_w16525_,
		_w16526_,
		_w17000_
	);
	LUT3 #(
		.INIT('h80)
	) name12953 (
		\CM_rd4[16]_pad ,
		_w16525_,
		_w16528_,
		_w17001_
	);
	LUT4 #(
		.INIT('h8000)
	) name12954 (
		\CM_rd1[16]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w17002_
	);
	LUT4 #(
		.INIT('h8000)
	) name12955 (
		\CM_rd6[16]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w17003_
	);
	LUT2 #(
		.INIT('h1)
	) name12956 (
		_w17002_,
		_w17003_,
		_w17004_
	);
	LUT3 #(
		.INIT('h10)
	) name12957 (
		_w17001_,
		_w17000_,
		_w17004_,
		_w17005_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12958 (
		_w16875_,
		_w16993_,
		_w16999_,
		_w17005_,
		_w17006_
	);
	LUT3 #(
		.INIT('h8a)
	) name12959 (
		\idma_IADi_reg[8]/P0001 ,
		_w4937_,
		_w9326_,
		_w17007_
	);
	LUT4 #(
		.INIT('h4447)
	) name12960 (
		_w8998_,
		_w9327_,
		_w17006_,
		_w17007_,
		_w17008_
	);
	LUT2 #(
		.INIT('h1)
	) name12961 (
		_w8182_,
		_w17008_,
		_w17009_
	);
	LUT4 #(
		.INIT('hff10)
	) name12962 (
		_w7465_,
		_w7565_,
		_w8182_,
		_w17009_,
		_w17010_
	);
	LUT4 #(
		.INIT('h2000)
	) name12963 (
		\CM_rdm[21]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w17011_
	);
	LUT4 #(
		.INIT('h8000)
	) name12964 (
		\CM_rd0[21]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w17012_
	);
	LUT4 #(
		.INIT('h8000)
	) name12965 (
		\CM_rd7[21]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w17013_
	);
	LUT2 #(
		.INIT('h1)
	) name12966 (
		_w17012_,
		_w17013_,
		_w17014_
	);
	LUT4 #(
		.INIT('h8000)
	) name12967 (
		\CM_rd2[21]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w17015_
	);
	LUT3 #(
		.INIT('h07)
	) name12968 (
		\CM_rd5[21]_pad ,
		_w16523_,
		_w17015_,
		_w17016_
	);
	LUT2 #(
		.INIT('h8)
	) name12969 (
		_w17014_,
		_w17016_,
		_w17017_
	);
	LUT3 #(
		.INIT('h80)
	) name12970 (
		\CM_rd3[21]_pad ,
		_w16525_,
		_w16526_,
		_w17018_
	);
	LUT3 #(
		.INIT('h80)
	) name12971 (
		\CM_rd4[21]_pad ,
		_w16525_,
		_w16528_,
		_w17019_
	);
	LUT4 #(
		.INIT('h8000)
	) name12972 (
		\CM_rd1[21]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w17020_
	);
	LUT4 #(
		.INIT('h8000)
	) name12973 (
		\CM_rd6[21]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w17021_
	);
	LUT2 #(
		.INIT('h1)
	) name12974 (
		_w17020_,
		_w17021_,
		_w17022_
	);
	LUT3 #(
		.INIT('h10)
	) name12975 (
		_w17019_,
		_w17018_,
		_w17022_,
		_w17023_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12976 (
		_w16875_,
		_w17011_,
		_w17017_,
		_w17023_,
		_w17024_
	);
	LUT3 #(
		.INIT('h8a)
	) name12977 (
		\idma_IADi_reg[13]/P0001 ,
		_w4937_,
		_w9326_,
		_w17025_
	);
	LUT4 #(
		.INIT('h4447)
	) name12978 (
		_w8740_,
		_w9327_,
		_w17024_,
		_w17025_,
		_w17026_
	);
	LUT2 #(
		.INIT('h1)
	) name12979 (
		_w8182_,
		_w17026_,
		_w17027_
	);
	LUT3 #(
		.INIT('hf8)
	) name12980 (
		_w5760_,
		_w8182_,
		_w17027_,
		_w17028_
	);
	LUT4 #(
		.INIT('h2000)
	) name12981 (
		\CM_rdm[20]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w17029_
	);
	LUT4 #(
		.INIT('h8000)
	) name12982 (
		\CM_rd0[20]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w17030_
	);
	LUT4 #(
		.INIT('h8000)
	) name12983 (
		\CM_rd7[20]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w17031_
	);
	LUT2 #(
		.INIT('h1)
	) name12984 (
		_w17030_,
		_w17031_,
		_w17032_
	);
	LUT4 #(
		.INIT('h8000)
	) name12985 (
		\CM_rd2[20]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w17033_
	);
	LUT3 #(
		.INIT('h07)
	) name12986 (
		\CM_rd5[20]_pad ,
		_w16523_,
		_w17033_,
		_w17034_
	);
	LUT2 #(
		.INIT('h8)
	) name12987 (
		_w17032_,
		_w17034_,
		_w17035_
	);
	LUT3 #(
		.INIT('h80)
	) name12988 (
		\CM_rd3[20]_pad ,
		_w16525_,
		_w16526_,
		_w17036_
	);
	LUT3 #(
		.INIT('h80)
	) name12989 (
		\CM_rd4[20]_pad ,
		_w16525_,
		_w16528_,
		_w17037_
	);
	LUT4 #(
		.INIT('h8000)
	) name12990 (
		\CM_rd1[20]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w17038_
	);
	LUT4 #(
		.INIT('h8000)
	) name12991 (
		\CM_rd6[20]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w17039_
	);
	LUT2 #(
		.INIT('h1)
	) name12992 (
		_w17038_,
		_w17039_,
		_w17040_
	);
	LUT3 #(
		.INIT('h10)
	) name12993 (
		_w17037_,
		_w17036_,
		_w17040_,
		_w17041_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12994 (
		_w16875_,
		_w17029_,
		_w17035_,
		_w17041_,
		_w17042_
	);
	LUT3 #(
		.INIT('h8a)
	) name12995 (
		\idma_IADi_reg[12]/P0001 ,
		_w4937_,
		_w9326_,
		_w17043_
	);
	LUT4 #(
		.INIT('h4447)
	) name12996 (
		_w8717_,
		_w9327_,
		_w17042_,
		_w17043_,
		_w17044_
	);
	LUT2 #(
		.INIT('h1)
	) name12997 (
		_w8182_,
		_w17044_,
		_w17045_
	);
	LUT3 #(
		.INIT('hf8)
	) name12998 (
		_w6758_,
		_w8182_,
		_w17045_,
		_w17046_
	);
	LUT4 #(
		.INIT('h2000)
	) name12999 (
		\CM_rdm[19]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w17047_
	);
	LUT4 #(
		.INIT('h8000)
	) name13000 (
		\CM_rd0[19]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w17048_
	);
	LUT4 #(
		.INIT('h8000)
	) name13001 (
		\CM_rd7[19]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w17049_
	);
	LUT2 #(
		.INIT('h1)
	) name13002 (
		_w17048_,
		_w17049_,
		_w17050_
	);
	LUT4 #(
		.INIT('h8000)
	) name13003 (
		\CM_rd2[19]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w17051_
	);
	LUT3 #(
		.INIT('h07)
	) name13004 (
		\CM_rd5[19]_pad ,
		_w16523_,
		_w17051_,
		_w17052_
	);
	LUT2 #(
		.INIT('h8)
	) name13005 (
		_w17050_,
		_w17052_,
		_w17053_
	);
	LUT3 #(
		.INIT('h80)
	) name13006 (
		\CM_rd3[19]_pad ,
		_w16525_,
		_w16526_,
		_w17054_
	);
	LUT3 #(
		.INIT('h80)
	) name13007 (
		\CM_rd4[19]_pad ,
		_w16525_,
		_w16528_,
		_w17055_
	);
	LUT4 #(
		.INIT('h8000)
	) name13008 (
		\CM_rd1[19]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w17056_
	);
	LUT4 #(
		.INIT('h8000)
	) name13009 (
		\CM_rd6[19]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w17057_
	);
	LUT2 #(
		.INIT('h1)
	) name13010 (
		_w17056_,
		_w17057_,
		_w17058_
	);
	LUT3 #(
		.INIT('h10)
	) name13011 (
		_w17055_,
		_w17054_,
		_w17058_,
		_w17059_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name13012 (
		_w16875_,
		_w17047_,
		_w17053_,
		_w17059_,
		_w17060_
	);
	LUT3 #(
		.INIT('h8a)
	) name13013 (
		\idma_IADi_reg[11]/P0001 ,
		_w4937_,
		_w9326_,
		_w17061_
	);
	LUT4 #(
		.INIT('h4447)
	) name13014 (
		_w8694_,
		_w9327_,
		_w17060_,
		_w17061_,
		_w17062_
	);
	LUT2 #(
		.INIT('h1)
	) name13015 (
		_w8182_,
		_w17062_,
		_w17063_
	);
	LUT4 #(
		.INIT('hff10)
	) name13016 (
		_w6263_,
		_w6362_,
		_w8182_,
		_w17063_,
		_w17064_
	);
	LUT4 #(
		.INIT('h2000)
	) name13017 (
		\CM_rdm[18]_pad ,
		_w16527_,
		_w16524_,
		_w16533_,
		_w17065_
	);
	LUT4 #(
		.INIT('h8000)
	) name13018 (
		\CM_rd0[18]_pad ,
		_w16514_,
		_w16515_,
		_w16516_,
		_w17066_
	);
	LUT4 #(
		.INIT('h8000)
	) name13019 (
		\CM_rd7[18]_pad ,
		_w16514_,
		_w16515_,
		_w16517_,
		_w17067_
	);
	LUT2 #(
		.INIT('h1)
	) name13020 (
		_w17066_,
		_w17067_,
		_w17068_
	);
	LUT4 #(
		.INIT('h8000)
	) name13021 (
		\CM_rd2[18]_pad ,
		_w16514_,
		_w16519_,
		_w16520_,
		_w17069_
	);
	LUT3 #(
		.INIT('h07)
	) name13022 (
		\CM_rd5[18]_pad ,
		_w16523_,
		_w17069_,
		_w17070_
	);
	LUT2 #(
		.INIT('h8)
	) name13023 (
		_w17068_,
		_w17070_,
		_w17071_
	);
	LUT3 #(
		.INIT('h80)
	) name13024 (
		\CM_rd3[18]_pad ,
		_w16525_,
		_w16526_,
		_w17072_
	);
	LUT3 #(
		.INIT('h80)
	) name13025 (
		\CM_rd4[18]_pad ,
		_w16525_,
		_w16528_,
		_w17073_
	);
	LUT4 #(
		.INIT('h8000)
	) name13026 (
		\CM_rd1[18]_pad ,
		_w16514_,
		_w16519_,
		_w16529_,
		_w17074_
	);
	LUT4 #(
		.INIT('h8000)
	) name13027 (
		\CM_rd6[18]_pad ,
		_w16519_,
		_w16515_,
		_w16531_,
		_w17075_
	);
	LUT2 #(
		.INIT('h1)
	) name13028 (
		_w17074_,
		_w17075_,
		_w17076_
	);
	LUT3 #(
		.INIT('h10)
	) name13029 (
		_w17073_,
		_w17072_,
		_w17076_,
		_w17077_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name13030 (
		_w16875_,
		_w17065_,
		_w17071_,
		_w17077_,
		_w17078_
	);
	LUT3 #(
		.INIT('h8a)
	) name13031 (
		\idma_IADi_reg[10]/P0001 ,
		_w4937_,
		_w9326_,
		_w17079_
	);
	LUT4 #(
		.INIT('h4447)
	) name13032 (
		_w8671_,
		_w9327_,
		_w17078_,
		_w17079_,
		_w17080_
	);
	LUT2 #(
		.INIT('h1)
	) name13033 (
		_w8182_,
		_w17080_,
		_w17081_
	);
	LUT4 #(
		.INIT('hff10)
	) name13034 (
		_w5937_,
		_w6038_,
		_w8182_,
		_w17081_,
		_w17082_
	);
	LUT2 #(
		.INIT('h1)
	) name13035 (
		_w5570_,
		_w5575_,
		_w17083_
	);
	LUT4 #(
		.INIT('h00b8)
	) name13036 (
		\memc_Pwrite_C_reg/NET0131 ,
		_w4971_,
		_w9085_,
		_w17083_,
		_w17084_
	);
	LUT2 #(
		.INIT('h2)
	) name13037 (
		_w9333_,
		_w17084_,
		_w17085_
	);
	LUT4 #(
		.INIT('hffef)
	) name13038 (
		_w9297_,
		_w9310_,
		_w9315_,
		_w17085_,
		_w17086_
	);
	LUT3 #(
		.INIT('h13)
	) name13039 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 ,
		_w9894_,
		_w17087_
	);
	LUT4 #(
		.INIT('h0002)
	) name13040 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w17087_,
		_w17088_
	);
	LUT4 #(
		.INIT('h1f00)
	) name13041 (
		_w11313_,
		_w11314_,
		_w12282_,
		_w17088_,
		_w17089_
	);
	LUT4 #(
		.INIT('h313b)
	) name13042 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 ,
		_w11308_,
		_w11635_,
		_w17090_
	);
	LUT3 #(
		.INIT('h45)
	) name13043 (
		_w11624_,
		_w17089_,
		_w17090_,
		_w17091_
	);
	LUT4 #(
		.INIT('h5041)
	) name13044 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11240_,
		_w16559_,
		_w16560_,
		_w17092_
	);
	LUT2 #(
		.INIT('h9)
	) name13045 (
		_w11188_,
		_w11206_,
		_w17093_
	);
	LUT4 #(
		.INIT('h2223)
	) name13046 (
		_w11217_,
		_w11241_,
		_w11240_,
		_w16560_,
		_w17094_
	);
	LUT4 #(
		.INIT('h3113)
	) name13047 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17092_,
		_w17093_,
		_w17094_,
		_w17095_
	);
	LUT3 #(
		.INIT('hec)
	) name13048 (
		_w11624_,
		_w17091_,
		_w17095_,
		_w17096_
	);
	LUT3 #(
		.INIT('h13)
	) name13049 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 ,
		_w9894_,
		_w17097_
	);
	LUT4 #(
		.INIT('h0002)
	) name13050 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w17097_,
		_w17098_
	);
	LUT4 #(
		.INIT('h5700)
	) name13051 (
		_w12282_,
		_w13610_,
		_w13611_,
		_w17098_,
		_w17099_
	);
	LUT4 #(
		.INIT('h313b)
	) name13052 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 ,
		_w11308_,
		_w11635_,
		_w17100_
	);
	LUT3 #(
		.INIT('h45)
	) name13053 (
		_w11624_,
		_w17099_,
		_w17100_,
		_w17101_
	);
	LUT4 #(
		.INIT('h08a2)
	) name13054 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11243_,
		_w12245_,
		_w16267_,
		_w17102_
	);
	LUT4 #(
		.INIT('h00be)
	) name13055 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17093_,
		_w17094_,
		_w17102_,
		_w17103_
	);
	LUT4 #(
		.INIT('hff41)
	) name13056 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17093_,
		_w17094_,
		_w17102_,
		_w17104_
	);
	LUT3 #(
		.INIT('hce)
	) name13057 (
		_w11624_,
		_w17101_,
		_w17103_,
		_w17105_
	);
	LUT2 #(
		.INIT('h2)
	) name13058 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001 ,
		_w11310_,
		_w17106_
	);
	LUT3 #(
		.INIT('h01)
	) name13059 (
		_w9946_,
		_w12442_,
		_w17106_,
		_w17107_
	);
	LUT4 #(
		.INIT('hfd00)
	) name13060 (
		_w12440_,
		_w13610_,
		_w13611_,
		_w17107_,
		_w17108_
	);
	LUT3 #(
		.INIT('h07)
	) name13061 (
		_w9946_,
		_w17103_,
		_w17108_,
		_w17109_
	);
	LUT2 #(
		.INIT('h2)
	) name13062 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001 ,
		_w11310_,
		_w17110_
	);
	LUT3 #(
		.INIT('h01)
	) name13063 (
		_w9946_,
		_w12442_,
		_w17110_,
		_w17111_
	);
	LUT4 #(
		.INIT('hef00)
	) name13064 (
		_w11313_,
		_w11314_,
		_w12440_,
		_w17111_,
		_w17112_
	);
	LUT3 #(
		.INIT('h0d)
	) name13065 (
		_w9946_,
		_w17095_,
		_w17112_,
		_w17113_
	);
	LUT3 #(
		.INIT('h13)
	) name13066 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001 ,
		_w9894_,
		_w17114_
	);
	LUT4 #(
		.INIT('h0002)
	) name13067 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w17114_,
		_w17115_
	);
	LUT4 #(
		.INIT('h313b)
	) name13068 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001 ,
		_w11631_,
		_w11635_,
		_w17116_
	);
	LUT4 #(
		.INIT('h2f00)
	) name13069 (
		_w11625_,
		_w12673_,
		_w17115_,
		_w17116_,
		_w17117_
	);
	LUT2 #(
		.INIT('h1)
	) name13070 (
		_w11624_,
		_w17117_,
		_w17118_
	);
	LUT3 #(
		.INIT('hf2)
	) name13071 (
		_w11624_,
		_w12331_,
		_w17118_,
		_w17119_
	);
	LUT2 #(
		.INIT('h2)
	) name13072 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001 ,
		_w11656_,
		_w17120_
	);
	LUT3 #(
		.INIT('h01)
	) name13073 (
		_w9946_,
		_w11659_,
		_w17120_,
		_w17121_
	);
	LUT3 #(
		.INIT('h70)
	) name13074 (
		_w11655_,
		_w12673_,
		_w17121_,
		_w17122_
	);
	LUT3 #(
		.INIT('h07)
	) name13075 (
		_w9946_,
		_w12331_,
		_w17122_,
		_w17123_
	);
	LUT3 #(
		.INIT('h13)
	) name13076 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001 ,
		_w9894_,
		_w17124_
	);
	LUT4 #(
		.INIT('h0002)
	) name13077 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w17124_,
		_w17125_
	);
	LUT4 #(
		.INIT('h1f00)
	) name13078 (
		_w11313_,
		_w11314_,
		_w11625_,
		_w17125_,
		_w17126_
	);
	LUT4 #(
		.INIT('h313b)
	) name13079 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001 ,
		_w11631_,
		_w11635_,
		_w17127_
	);
	LUT4 #(
		.INIT('h0020)
	) name13080 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w9453_,
		_w9894_,
		_w12364_,
		_w17128_
	);
	LUT4 #(
		.INIT('hff45)
	) name13081 (
		_w11624_,
		_w17126_,
		_w17127_,
		_w17128_,
		_w17129_
	);
	LUT2 #(
		.INIT('h8)
	) name13082 (
		_w9946_,
		_w12364_,
		_w17130_
	);
	LUT2 #(
		.INIT('h2)
	) name13083 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001 ,
		_w11656_,
		_w17131_
	);
	LUT3 #(
		.INIT('h01)
	) name13084 (
		_w9946_,
		_w11659_,
		_w17131_,
		_w17132_
	);
	LUT4 #(
		.INIT('hef00)
	) name13085 (
		_w11313_,
		_w11314_,
		_w11655_,
		_w17132_,
		_w17133_
	);
	LUT2 #(
		.INIT('h1)
	) name13086 (
		_w17130_,
		_w17133_,
		_w17134_
	);
	LUT3 #(
		.INIT('h13)
	) name13087 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001 ,
		_w9894_,
		_w17135_
	);
	LUT4 #(
		.INIT('h0002)
	) name13088 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w17135_,
		_w17136_
	);
	LUT4 #(
		.INIT('h313b)
	) name13089 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001 ,
		_w11631_,
		_w11635_,
		_w17137_
	);
	LUT4 #(
		.INIT('h4f00)
	) name13090 (
		_w11318_,
		_w11625_,
		_w17136_,
		_w17137_,
		_w17138_
	);
	LUT2 #(
		.INIT('h1)
	) name13091 (
		_w11624_,
		_w17138_,
		_w17139_
	);
	LUT3 #(
		.INIT('hf2)
	) name13092 (
		_w11624_,
		_w12328_,
		_w17139_,
		_w17140_
	);
	LUT4 #(
		.INIT('h1411)
	) name13093 (
		_w9455_,
		_w9838_,
		_w9839_,
		_w9840_,
		_w17141_
	);
	LUT2 #(
		.INIT('h8)
	) name13094 (
		_w8351_,
		_w9455_,
		_w17142_
	);
	LUT4 #(
		.INIT('h222e)
	) name13095 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001 ,
		_w9895_,
		_w17141_,
		_w17142_,
		_w17143_
	);
	LUT4 #(
		.INIT('h222e)
	) name13096 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001 ,
		_w9454_,
		_w17141_,
		_w17142_,
		_w17144_
	);
	LUT2 #(
		.INIT('h2)
	) name13097 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001 ,
		_w11656_,
		_w17145_
	);
	LUT3 #(
		.INIT('h01)
	) name13098 (
		_w9946_,
		_w11659_,
		_w17145_,
		_w17146_
	);
	LUT3 #(
		.INIT('h70)
	) name13099 (
		_w11318_,
		_w11655_,
		_w17146_,
		_w17147_
	);
	LUT3 #(
		.INIT('h07)
	) name13100 (
		_w9946_,
		_w12328_,
		_w17147_,
		_w17148_
	);
	LUT4 #(
		.INIT('h0400)
	) name13101 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[7]/NET0131 ,
		_w17149_
	);
	LUT4 #(
		.INIT('h0302)
	) name13102 (
		\T_TMODE[0]_pad ,
		\tm_TCR_TMP_reg[4]/NET0131 ,
		\tm_TCR_TMP_reg[5]/NET0131 ,
		_w12797_,
		_w17150_
	);
	LUT3 #(
		.INIT('h10)
	) name13103 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w14107_,
		_w17150_,
		_w17151_
	);
	LUT4 #(
		.INIT('h0100)
	) name13104 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TCR_TMP_reg[6]/NET0131 ,
		_w14107_,
		_w17150_,
		_w17152_
	);
	LUT3 #(
		.INIT('he0)
	) name13105 (
		\T_TMODE[0]_pad ,
		_w12797_,
		_w12798_,
		_w17153_
	);
	LUT3 #(
		.INIT('h10)
	) name13106 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w14107_,
		_w17153_,
		_w17154_
	);
	LUT4 #(
		.INIT('h0301)
	) name13107 (
		\tm_TCR_TMP_reg[7]/NET0131 ,
		_w14103_,
		_w17154_,
		_w17152_,
		_w17155_
	);
	LUT4 #(
		.INIT('h2333)
	) name13108 (
		\tm_tpr_reg_DO_reg[7]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w17156_
	);
	LUT3 #(
		.INIT('hba)
	) name13109 (
		_w17149_,
		_w17155_,
		_w17156_,
		_w17157_
	);
	LUT4 #(
		.INIT('h4000)
	) name13110 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w17158_
	);
	LUT2 #(
		.INIT('h8)
	) name13111 (
		_w14460_,
		_w17158_,
		_w17159_
	);
	LUT2 #(
		.INIT('h8)
	) name13112 (
		_w15953_,
		_w15949_,
		_w17160_
	);
	LUT3 #(
		.INIT('h20)
	) name13113 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_dec_IRE_reg[0]/NET0131 ,
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w17161_
	);
	LUT2 #(
		.INIT('h8)
	) name13114 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w17162_
	);
	LUT2 #(
		.INIT('h1)
	) name13115 (
		\core_c_dec_MTCNTR_Eg_reg/P0001 ,
		\core_c_dec_MTOWRCNTR_Eg_reg/P0001 ,
		_w17163_
	);
	LUT4 #(
		.INIT('h0103)
	) name13116 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_MTCNTR_Eg_reg/P0001 ,
		\core_c_dec_MTOWRCNTR_Eg_reg/P0001 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w17164_
	);
	LUT3 #(
		.INIT('h70)
	) name13117 (
		_w5088_,
		_w17161_,
		_w17164_,
		_w17165_
	);
	LUT4 #(
		.INIT('hdf00)
	) name13118 (
		_w4169_,
		_w4430_,
		_w17160_,
		_w17165_,
		_w17166_
	);
	LUT2 #(
		.INIT('h1)
	) name13119 (
		_w4971_,
		_w17166_,
		_w17167_
	);
	LUT3 #(
		.INIT('ha8)
	) name13120 (
		\core_c_psq_CE_reg/NET0131 ,
		_w4971_,
		_w17166_,
		_w17168_
	);
	LUT4 #(
		.INIT('h0200)
	) name13121 (
		_w4169_,
		_w4430_,
		_w4178_,
		_w17160_,
		_w17169_
	);
	LUT4 #(
		.INIT('h070f)
	) name13122 (
		\core_c_psq_CE_reg/NET0131 ,
		_w5088_,
		_w17162_,
		_w17161_,
		_w17170_
	);
	LUT4 #(
		.INIT('h0001)
	) name13123 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w17171_
	);
	LUT4 #(
		.INIT('h0100)
	) name13124 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w17171_,
		_w17172_
	);
	LUT4 #(
		.INIT('h0100)
	) name13125 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w17172_,
		_w17173_
	);
	LUT4 #(
		.INIT('h0100)
	) name13126 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w17173_,
		_w17174_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name13127 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w17173_,
		_w17175_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13128 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17175_,
		_w17176_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name13129 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17177_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name13130 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17178_
	);
	LUT2 #(
		.INIT('h8)
	) name13131 (
		_w17177_,
		_w17178_,
		_w17179_
	);
	LUT4 #(
		.INIT('h0045)
	) name13132 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17179_,
		_w17180_
	);
	LUT4 #(
		.INIT('h111d)
	) name13133 (
		_w6758_,
		_w17163_,
		_w17176_,
		_w17180_,
		_w17181_
	);
	LUT2 #(
		.INIT('h9)
	) name13134 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w17173_,
		_w17182_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13135 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17182_,
		_w17183_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13136 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17184_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13137 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17185_
	);
	LUT2 #(
		.INIT('h8)
	) name13138 (
		_w17184_,
		_w17185_,
		_w17186_
	);
	LUT4 #(
		.INIT('h0045)
	) name13139 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17186_,
		_w17187_
	);
	LUT3 #(
		.INIT('ha8)
	) name13140 (
		_w17163_,
		_w17183_,
		_w17187_,
		_w17188_
	);
	LUT3 #(
		.INIT('h01)
	) name13141 (
		_w5937_,
		_w6038_,
		_w17163_,
		_w17189_
	);
	LUT3 #(
		.INIT('h02)
	) name13142 (
		_w17181_,
		_w17188_,
		_w17189_,
		_w17190_
	);
	LUT3 #(
		.INIT('h63)
	) name13143 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w17172_,
		_w17191_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13144 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17191_,
		_w17192_
	);
	LUT4 #(
		.INIT('h35ff)
	) name13145 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17193_
	);
	LUT4 #(
		.INIT('hff35)
	) name13146 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17194_
	);
	LUT2 #(
		.INIT('h8)
	) name13147 (
		_w17193_,
		_w17194_,
		_w17195_
	);
	LUT4 #(
		.INIT('h0045)
	) name13148 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17195_,
		_w17196_
	);
	LUT3 #(
		.INIT('ha8)
	) name13149 (
		_w17163_,
		_w17192_,
		_w17196_,
		_w17197_
	);
	LUT3 #(
		.INIT('h01)
	) name13150 (
		_w7465_,
		_w7565_,
		_w17163_,
		_w17198_
	);
	LUT2 #(
		.INIT('h9)
	) name13151 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w17171_,
		_w17199_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13152 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17199_,
		_w17200_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13153 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17201_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13154 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17202_
	);
	LUT2 #(
		.INIT('h8)
	) name13155 (
		_w17201_,
		_w17202_,
		_w17203_
	);
	LUT4 #(
		.INIT('h0045)
	) name13156 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17203_,
		_w17204_
	);
	LUT3 #(
		.INIT('ha8)
	) name13157 (
		_w17163_,
		_w17200_,
		_w17204_,
		_w17205_
	);
	LUT4 #(
		.INIT('h0045)
	) name13158 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w17163_,
		_w17206_
	);
	LUT4 #(
		.INIT('h0001)
	) name13159 (
		_w17197_,
		_w17198_,
		_w17205_,
		_w17206_,
		_w17207_
	);
	LUT4 #(
		.INIT('h0045)
	) name13160 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w17163_,
		_w17208_
	);
	LUT2 #(
		.INIT('h6)
	) name13161 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w17209_
	);
	LUT4 #(
		.INIT('hba00)
	) name13162 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17209_,
		_w17210_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13163 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17211_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13164 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17212_
	);
	LUT2 #(
		.INIT('h8)
	) name13165 (
		_w17211_,
		_w17212_,
		_w17213_
	);
	LUT4 #(
		.INIT('h4500)
	) name13166 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17213_,
		_w17214_
	);
	LUT3 #(
		.INIT('h02)
	) name13167 (
		_w17163_,
		_w17214_,
		_w17210_,
		_w17215_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name13168 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w17172_,
		_w17216_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13169 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17216_,
		_w17217_
	);
	LUT4 #(
		.INIT('h35ff)
	) name13170 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17218_
	);
	LUT4 #(
		.INIT('hff35)
	) name13171 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17219_
	);
	LUT2 #(
		.INIT('h8)
	) name13172 (
		_w17218_,
		_w17219_,
		_w17220_
	);
	LUT4 #(
		.INIT('h0045)
	) name13173 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17220_,
		_w17221_
	);
	LUT3 #(
		.INIT('ha8)
	) name13174 (
		_w17163_,
		_w17217_,
		_w17221_,
		_w17222_
	);
	LUT3 #(
		.INIT('h01)
	) name13175 (
		_w7140_,
		_w7240_,
		_w17163_,
		_w17223_
	);
	LUT4 #(
		.INIT('h0001)
	) name13176 (
		_w17208_,
		_w17215_,
		_w17222_,
		_w17223_,
		_w17224_
	);
	LUT3 #(
		.INIT('h80)
	) name13177 (
		_w17190_,
		_w17207_,
		_w17224_,
		_w17225_
	);
	LUT2 #(
		.INIT('h9)
	) name13178 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w17172_,
		_w17226_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13179 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17226_,
		_w17227_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13180 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17228_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13181 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17229_
	);
	LUT2 #(
		.INIT('h8)
	) name13182 (
		_w17228_,
		_w17229_,
		_w17230_
	);
	LUT4 #(
		.INIT('h0045)
	) name13183 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17230_,
		_w17231_
	);
	LUT3 #(
		.INIT('ha8)
	) name13184 (
		_w17163_,
		_w17227_,
		_w17231_,
		_w17232_
	);
	LUT4 #(
		.INIT('h0045)
	) name13185 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w17163_,
		_w17233_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name13186 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w17171_,
		_w17234_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13187 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17234_,
		_w17235_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13188 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17236_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13189 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17237_
	);
	LUT2 #(
		.INIT('h8)
	) name13190 (
		_w17236_,
		_w17237_,
		_w17238_
	);
	LUT4 #(
		.INIT('h0045)
	) name13191 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17238_,
		_w17239_
	);
	LUT3 #(
		.INIT('ha8)
	) name13192 (
		_w17163_,
		_w17235_,
		_w17239_,
		_w17240_
	);
	LUT4 #(
		.INIT('h0045)
	) name13193 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w17163_,
		_w17241_
	);
	LUT4 #(
		.INIT('h0001)
	) name13194 (
		_w17232_,
		_w17233_,
		_w17240_,
		_w17241_,
		_w17242_
	);
	LUT3 #(
		.INIT('h63)
	) name13195 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w17171_,
		_w17243_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13196 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17243_,
		_w17244_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13197 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17245_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13198 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17246_
	);
	LUT2 #(
		.INIT('h8)
	) name13199 (
		_w17245_,
		_w17246_,
		_w17247_
	);
	LUT4 #(
		.INIT('h0045)
	) name13200 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17247_,
		_w17248_
	);
	LUT3 #(
		.INIT('ha8)
	) name13201 (
		_w17163_,
		_w17244_,
		_w17248_,
		_w17249_
	);
	LUT4 #(
		.INIT('h0045)
	) name13202 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w17163_,
		_w17250_
	);
	LUT3 #(
		.INIT('h63)
	) name13203 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w17173_,
		_w17251_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13204 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17251_,
		_w17252_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13205 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17253_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13206 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17254_
	);
	LUT2 #(
		.INIT('h8)
	) name13207 (
		_w17253_,
		_w17254_,
		_w17255_
	);
	LUT4 #(
		.INIT('h0045)
	) name13208 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17255_,
		_w17256_
	);
	LUT3 #(
		.INIT('ha8)
	) name13209 (
		_w17163_,
		_w17252_,
		_w17256_,
		_w17257_
	);
	LUT3 #(
		.INIT('h01)
	) name13210 (
		_w6263_,
		_w6362_,
		_w17163_,
		_w17258_
	);
	LUT4 #(
		.INIT('h0001)
	) name13211 (
		_w17249_,
		_w17250_,
		_w17257_,
		_w17258_,
		_w17259_
	);
	LUT2 #(
		.INIT('h8)
	) name13212 (
		_w17242_,
		_w17259_,
		_w17260_
	);
	LUT4 #(
		.INIT('h01fe)
	) name13213 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w17261_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13214 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17261_,
		_w17262_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13215 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17263_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13216 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17264_
	);
	LUT2 #(
		.INIT('h8)
	) name13217 (
		_w17263_,
		_w17264_,
		_w17265_
	);
	LUT4 #(
		.INIT('h0045)
	) name13218 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17265_,
		_w17266_
	);
	LUT3 #(
		.INIT('ha8)
	) name13219 (
		_w17163_,
		_w17262_,
		_w17266_,
		_w17267_
	);
	LUT4 #(
		.INIT('h0045)
	) name13220 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w17163_,
		_w17268_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13221 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17269_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13222 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17270_
	);
	LUT2 #(
		.INIT('h8)
	) name13223 (
		_w17269_,
		_w17270_,
		_w17271_
	);
	LUT4 #(
		.INIT('h4500)
	) name13224 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17271_,
		_w17272_
	);
	LUT2 #(
		.INIT('h9)
	) name13225 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w17174_,
		_w17273_
	);
	LUT4 #(
		.INIT('hba00)
	) name13226 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17273_,
		_w17274_
	);
	LUT4 #(
		.INIT('hddd1)
	) name13227 (
		_w5760_,
		_w17163_,
		_w17274_,
		_w17272_,
		_w17275_
	);
	LUT3 #(
		.INIT('h10)
	) name13228 (
		_w17267_,
		_w17268_,
		_w17275_,
		_w17276_
	);
	LUT3 #(
		.INIT('h1e)
	) name13229 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w17277_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13230 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17277_,
		_w17278_
	);
	LUT4 #(
		.INIT('hf35f)
	) name13231 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17279_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name13232 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17280_
	);
	LUT2 #(
		.INIT('h8)
	) name13233 (
		_w17279_,
		_w17280_,
		_w17281_
	);
	LUT4 #(
		.INIT('h0045)
	) name13234 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17281_,
		_w17282_
	);
	LUT3 #(
		.INIT('ha8)
	) name13235 (
		_w17163_,
		_w17278_,
		_w17282_,
		_w17283_
	);
	LUT4 #(
		.INIT('h0045)
	) name13236 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w17163_,
		_w17284_
	);
	LUT2 #(
		.INIT('h1)
	) name13237 (
		_w17283_,
		_w17284_,
		_w17285_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name13238 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17286_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name13239 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001 ,
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001 ,
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w17287_
	);
	LUT2 #(
		.INIT('h8)
	) name13240 (
		_w17286_,
		_w17287_,
		_w17288_
	);
	LUT4 #(
		.INIT('h0045)
	) name13241 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17288_,
		_w17289_
	);
	LUT4 #(
		.INIT('h4544)
	) name13242 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w17169_,
		_w17170_,
		_w17290_
	);
	LUT3 #(
		.INIT('h02)
	) name13243 (
		_w17163_,
		_w17290_,
		_w17289_,
		_w17291_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13244 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w17163_,
		_w17292_
	);
	LUT3 #(
		.INIT('h02)
	) name13245 (
		_w17167_,
		_w17292_,
		_w17291_,
		_w17293_
	);
	LUT3 #(
		.INIT('h80)
	) name13246 (
		_w17285_,
		_w17293_,
		_w17276_,
		_w17294_
	);
	LUT4 #(
		.INIT('heaaa)
	) name13247 (
		_w17168_,
		_w17260_,
		_w17294_,
		_w17225_,
		_w17295_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13248 (
		_w16586_,
		_w16592_,
		_w16598_,
		_w16875_,
		_w17296_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name13249 (
		\idma_ISn_reg/P0001 ,
		\idma_IWRn_reg/P0001 ,
		\idma_PM_1st_reg/NET0131 ,
		\idma_WRtrue_reg/NET0131 ,
		_w17297_
	);
	LUT2 #(
		.INIT('h2)
	) name13250 (
		_w13072_,
		_w17297_,
		_w17298_
	);
	LUT4 #(
		.INIT('h3100)
	) name13251 (
		\idma_PM_1st_reg/NET0131 ,
		_w9327_,
		_w12821_,
		_w17298_,
		_w17299_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13252 (
		\idma_DTMP_L_reg[7]/P0001 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12821_,
		_w17298_,
		_w17300_
	);
	LUT4 #(
		.INIT('hffe0)
	) name13253 (
		_w16876_,
		_w17296_,
		_w17299_,
		_w17300_,
		_w17301_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13254 (
		_w16646_,
		_w16652_,
		_w16658_,
		_w16875_,
		_w17302_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13255 (
		\idma_DTMP_L_reg[4]/P0001 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12821_,
		_w17298_,
		_w17303_
	);
	LUT4 #(
		.INIT('hffc8)
	) name13256 (
		_w16899_,
		_w17299_,
		_w17302_,
		_w17303_,
		_w17304_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13257 (
		_w16666_,
		_w16672_,
		_w16678_,
		_w16875_,
		_w17305_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13258 (
		\idma_DTMP_L_reg[3]/P0001 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12821_,
		_w17298_,
		_w17306_
	);
	LUT4 #(
		.INIT('hffc8)
	) name13259 (
		_w16907_,
		_w17299_,
		_w17305_,
		_w17306_,
		_w17307_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13260 (
		_w16606_,
		_w16612_,
		_w16618_,
		_w16875_,
		_w17308_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13261 (
		\idma_DTMP_L_reg[6]/P0001 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12821_,
		_w17298_,
		_w17309_
	);
	LUT4 #(
		.INIT('hffc8)
	) name13262 (
		_w16884_,
		_w17299_,
		_w17308_,
		_w17309_,
		_w17310_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13263 (
		_w16686_,
		_w16692_,
		_w16698_,
		_w16875_,
		_w17311_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13264 (
		\idma_DTMP_L_reg[2]/P0001 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12821_,
		_w17298_,
		_w17312_
	);
	LUT4 #(
		.INIT('hffc8)
	) name13265 (
		_w16915_,
		_w17299_,
		_w17311_,
		_w17312_,
		_w17313_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13266 (
		_w16626_,
		_w16632_,
		_w16638_,
		_w16875_,
		_w17314_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13267 (
		\idma_DTMP_L_reg[5]/P0001 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12821_,
		_w17298_,
		_w17315_
	);
	LUT4 #(
		.INIT('hffc8)
	) name13268 (
		_w16891_,
		_w17299_,
		_w17314_,
		_w17315_,
		_w17316_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13269 (
		_w16706_,
		_w16712_,
		_w16718_,
		_w16875_,
		_w17317_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13270 (
		\idma_DTMP_L_reg[1]/P0001 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12821_,
		_w17298_,
		_w17318_
	);
	LUT4 #(
		.INIT('hffc8)
	) name13271 (
		_w16923_,
		_w17299_,
		_w17317_,
		_w17318_,
		_w17319_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13272 (
		_w16726_,
		_w16732_,
		_w16738_,
		_w16875_,
		_w17320_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13273 (
		\idma_DTMP_L_reg[0]/P0001 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12821_,
		_w17298_,
		_w17321_
	);
	LUT4 #(
		.INIT('hffc8)
	) name13274 (
		_w16965_,
		_w17299_,
		_w17320_,
		_w17321_,
		_w17322_
	);
	LUT4 #(
		.INIT('h0008)
	) name13275 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w17323_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13276 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		\sice_SPC_reg[9]/P0001 ,
		_w16506_,
		_w17323_,
		_w17324_
	);
	LUT4 #(
		.INIT('h0080)
	) name13277 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17324_,
		_w17325_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13278 (
		_w13327_,
		_w16808_,
		_w16822_,
		_w17325_,
		_w17326_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13279 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\sice_SPC_reg[8]/P0001 ,
		_w16506_,
		_w17323_,
		_w17327_
	);
	LUT4 #(
		.INIT('h0080)
	) name13280 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17327_,
		_w17328_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13281 (
		_w13327_,
		_w16788_,
		_w16802_,
		_w17328_,
		_w17329_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13282 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		\sice_SPC_reg[7]/P0001 ,
		_w16506_,
		_w17323_,
		_w17330_
	);
	LUT4 #(
		.INIT('h0080)
	) name13283 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17330_,
		_w17331_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13284 (
		_w13327_,
		_w16585_,
		_w16599_,
		_w17331_,
		_w17332_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13285 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		\sice_SPC_reg[6]/P0001 ,
		_w16506_,
		_w17323_,
		_w17333_
	);
	LUT4 #(
		.INIT('h0080)
	) name13286 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17333_,
		_w17334_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13287 (
		_w13327_,
		_w16605_,
		_w16619_,
		_w17334_,
		_w17335_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13288 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\sice_SPC_reg[5]/P0001 ,
		_w16506_,
		_w17323_,
		_w17336_
	);
	LUT4 #(
		.INIT('h0080)
	) name13289 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17336_,
		_w17337_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13290 (
		_w13327_,
		_w16625_,
		_w16639_,
		_w17337_,
		_w17338_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13291 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\sice_SPC_reg[4]/P0001 ,
		_w16506_,
		_w17323_,
		_w17339_
	);
	LUT4 #(
		.INIT('h0080)
	) name13292 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17339_,
		_w17340_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13293 (
		_w13327_,
		_w16645_,
		_w16659_,
		_w17340_,
		_w17341_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13294 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		\sice_SPC_reg[3]/P0001 ,
		_w16506_,
		_w17323_,
		_w17342_
	);
	LUT4 #(
		.INIT('h0080)
	) name13295 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17342_,
		_w17343_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13296 (
		_w13327_,
		_w16665_,
		_w16679_,
		_w17343_,
		_w17344_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13297 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\sice_SPC_reg[2]/P0001 ,
		_w16506_,
		_w17323_,
		_w17345_
	);
	LUT4 #(
		.INIT('h0080)
	) name13298 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17345_,
		_w17346_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13299 (
		_w13327_,
		_w16685_,
		_w16699_,
		_w17346_,
		_w17347_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13300 (
		\core_c_dec_IR_reg[23]/NET0131 ,
		\sice_SPC_reg[23]/P0001 ,
		_w16506_,
		_w17323_,
		_w17348_
	);
	LUT4 #(
		.INIT('h0080)
	) name13301 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17348_,
		_w17349_
	);
	LUT2 #(
		.INIT('h8)
	) name13302 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[23]/P0001 ,
		_w17350_
	);
	LUT4 #(
		.INIT('h4555)
	) name13303 (
		\T_TMODE[1]_pad ,
		_w16930_,
		_w16936_,
		_w16942_,
		_w17351_
	);
	LUT4 #(
		.INIT('h3332)
	) name13304 (
		_w13327_,
		_w17349_,
		_w17350_,
		_w17351_,
		_w17352_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13305 (
		\core_c_dec_IR_reg[22]/NET0131 ,
		\sice_SPC_reg[22]/P0001 ,
		_w16506_,
		_w17323_,
		_w17353_
	);
	LUT4 #(
		.INIT('h0080)
	) name13306 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17353_,
		_w17354_
	);
	LUT2 #(
		.INIT('h8)
	) name13307 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[22]/P0001 ,
		_w17355_
	);
	LUT4 #(
		.INIT('h4555)
	) name13308 (
		\T_TMODE[1]_pad ,
		_w16947_,
		_w16953_,
		_w16959_,
		_w17356_
	);
	LUT4 #(
		.INIT('h3332)
	) name13309 (
		_w13327_,
		_w17354_,
		_w17355_,
		_w17356_,
		_w17357_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13310 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\sice_SPC_reg[21]/P0001 ,
		_w16506_,
		_w17323_,
		_w17358_
	);
	LUT4 #(
		.INIT('h0080)
	) name13311 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17358_,
		_w17359_
	);
	LUT2 #(
		.INIT('h8)
	) name13312 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[21]/P0001 ,
		_w17360_
	);
	LUT4 #(
		.INIT('h4555)
	) name13313 (
		\T_TMODE[1]_pad ,
		_w17011_,
		_w17017_,
		_w17023_,
		_w17361_
	);
	LUT4 #(
		.INIT('h3332)
	) name13314 (
		_w13327_,
		_w17359_,
		_w17360_,
		_w17361_,
		_w17362_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13315 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\sice_SPC_reg[20]/P0001 ,
		_w16506_,
		_w17323_,
		_w17363_
	);
	LUT4 #(
		.INIT('h0080)
	) name13316 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17363_,
		_w17364_
	);
	LUT2 #(
		.INIT('h8)
	) name13317 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[20]/P0001 ,
		_w17365_
	);
	LUT4 #(
		.INIT('h4555)
	) name13318 (
		\T_TMODE[1]_pad ,
		_w17029_,
		_w17035_,
		_w17041_,
		_w17366_
	);
	LUT4 #(
		.INIT('h3332)
	) name13319 (
		_w13327_,
		_w17364_,
		_w17365_,
		_w17366_,
		_w17367_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13320 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		\sice_SPC_reg[19]/P0001 ,
		_w16506_,
		_w17323_,
		_w17368_
	);
	LUT4 #(
		.INIT('h0080)
	) name13321 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17368_,
		_w17369_
	);
	LUT2 #(
		.INIT('h8)
	) name13322 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[19]/P0001 ,
		_w17370_
	);
	LUT4 #(
		.INIT('h4555)
	) name13323 (
		\T_TMODE[1]_pad ,
		_w17047_,
		_w17053_,
		_w17059_,
		_w17371_
	);
	LUT4 #(
		.INIT('h3332)
	) name13324 (
		_w13327_,
		_w17369_,
		_w17370_,
		_w17371_,
		_w17372_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13325 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\sice_SPC_reg[18]/P0001 ,
		_w16506_,
		_w17323_,
		_w17373_
	);
	LUT4 #(
		.INIT('h0080)
	) name13326 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17373_,
		_w17374_
	);
	LUT2 #(
		.INIT('h8)
	) name13327 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[18]/P0001 ,
		_w17375_
	);
	LUT4 #(
		.INIT('h4555)
	) name13328 (
		\T_TMODE[1]_pad ,
		_w17065_,
		_w17071_,
		_w17077_,
		_w17376_
	);
	LUT4 #(
		.INIT('h3332)
	) name13329 (
		_w13327_,
		_w17374_,
		_w17375_,
		_w17376_,
		_w17377_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13330 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		\sice_SPC_reg[17]/P0001 ,
		_w16506_,
		_w17323_,
		_w17378_
	);
	LUT4 #(
		.INIT('h0080)
	) name13331 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17378_,
		_w17379_
	);
	LUT2 #(
		.INIT('h8)
	) name13332 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[17]/P0001 ,
		_w17380_
	);
	LUT4 #(
		.INIT('h4555)
	) name13333 (
		\T_TMODE[1]_pad ,
		_w16975_,
		_w16981_,
		_w16987_,
		_w17381_
	);
	LUT4 #(
		.INIT('h3332)
	) name13334 (
		_w13327_,
		_w17379_,
		_w17380_,
		_w17381_,
		_w17382_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13335 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\sice_SPC_reg[16]/P0001 ,
		_w16506_,
		_w17323_,
		_w17383_
	);
	LUT4 #(
		.INIT('h0080)
	) name13336 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17383_,
		_w17384_
	);
	LUT2 #(
		.INIT('h8)
	) name13337 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[16]/P0001 ,
		_w17385_
	);
	LUT4 #(
		.INIT('h4555)
	) name13338 (
		\T_TMODE[1]_pad ,
		_w16993_,
		_w16999_,
		_w17005_,
		_w17386_
	);
	LUT4 #(
		.INIT('h3332)
	) name13339 (
		_w13327_,
		_w17384_,
		_w17385_,
		_w17386_,
		_w17387_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13340 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\sice_SPC_reg[15]/P0001 ,
		_w16506_,
		_w17323_,
		_w17388_
	);
	LUT4 #(
		.INIT('h0080)
	) name13341 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17388_,
		_w17389_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13342 (
		_w13327_,
		_w16513_,
		_w16547_,
		_w17389_,
		_w17390_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13343 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		\sice_SPC_reg[14]/P0001 ,
		_w16506_,
		_w17323_,
		_w17391_
	);
	LUT4 #(
		.INIT('h0080)
	) name13344 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17391_,
		_w17392_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13345 (
		_w13327_,
		_w16564_,
		_w16578_,
		_w17392_,
		_w17393_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13346 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\sice_SPC_reg[13]/P0001 ,
		_w16506_,
		_w17323_,
		_w17394_
	);
	LUT4 #(
		.INIT('h0080)
	) name13347 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17394_,
		_w17395_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13348 (
		_w13327_,
		_w16748_,
		_w16762_,
		_w17395_,
		_w17396_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13349 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		\sice_SPC_reg[12]/P0001 ,
		_w16506_,
		_w17323_,
		_w17397_
	);
	LUT4 #(
		.INIT('h0080)
	) name13350 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17397_,
		_w17398_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13351 (
		_w13327_,
		_w16768_,
		_w16782_,
		_w17398_,
		_w17399_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13352 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\sice_SPC_reg[11]/P0001 ,
		_w16506_,
		_w17323_,
		_w17400_
	);
	LUT4 #(
		.INIT('h0080)
	) name13353 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17400_,
		_w17401_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13354 (
		_w13327_,
		_w16828_,
		_w16842_,
		_w17401_,
		_w17402_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13355 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\sice_SPC_reg[10]/P0001 ,
		_w16506_,
		_w17323_,
		_w17403_
	);
	LUT4 #(
		.INIT('h0080)
	) name13356 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17403_,
		_w17404_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13357 (
		_w13327_,
		_w16848_,
		_w16862_,
		_w17404_,
		_w17405_
	);
	LUT3 #(
		.INIT('h80)
	) name13358 (
		\sice_SPC_reg[21]/P0001 ,
		_w16506_,
		_w16507_,
		_w17406_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13359 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w17360_,
		_w17361_,
		_w17406_,
		_w17407_
	);
	LUT3 #(
		.INIT('h80)
	) name13360 (
		\sice_SPC_reg[20]/P0001 ,
		_w16506_,
		_w16507_,
		_w17408_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13361 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w17365_,
		_w17366_,
		_w17408_,
		_w17409_
	);
	LUT3 #(
		.INIT('h80)
	) name13362 (
		\sice_SPC_reg[19]/P0001 ,
		_w16506_,
		_w16507_,
		_w17410_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13363 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w17370_,
		_w17371_,
		_w17410_,
		_w17411_
	);
	LUT3 #(
		.INIT('h80)
	) name13364 (
		\sice_SPC_reg[18]/P0001 ,
		_w16506_,
		_w16507_,
		_w17412_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13365 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w17375_,
		_w17376_,
		_w17412_,
		_w17413_
	);
	LUT3 #(
		.INIT('h80)
	) name13366 (
		\sice_SPC_reg[17]/P0001 ,
		_w16506_,
		_w16507_,
		_w17414_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13367 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w17380_,
		_w17381_,
		_w17414_,
		_w17415_
	);
	LUT3 #(
		.INIT('h80)
	) name13368 (
		\sice_SPC_reg[16]/P0001 ,
		_w16506_,
		_w16507_,
		_w17416_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13369 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w17385_,
		_w17386_,
		_w17416_,
		_w17417_
	);
	LUT3 #(
		.INIT('h80)
	) name13370 (
		\sice_SPC_reg[23]/P0001 ,
		_w16506_,
		_w16507_,
		_w17418_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13371 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w17350_,
		_w17351_,
		_w17418_,
		_w17419_
	);
	LUT3 #(
		.INIT('h80)
	) name13372 (
		\sice_SPC_reg[22]/P0001 ,
		_w16506_,
		_w16507_,
		_w17420_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13373 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w17355_,
		_w17356_,
		_w17420_,
		_w17421_
	);
	LUT4 #(
		.INIT('h2000)
	) name13374 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w4885_,
		_w4884_,
		_w9079_,
		_w17422_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13375 (
		_w16789_,
		_w16795_,
		_w16801_,
		_w17422_,
		_w17423_
	);
	LUT3 #(
		.INIT('h07)
	) name13376 (
		_w8647_,
		_w9082_,
		_w17423_,
		_w17424_
	);
	LUT4 #(
		.INIT('hfd00)
	) name13377 (
		_w5536_,
		_w7465_,
		_w7565_,
		_w17424_,
		_w17425_
	);
	LUT3 #(
		.INIT('h4e)
	) name13378 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[8]/P0001 ,
		_w17425_,
		_w17426_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13379 (
		_w16809_,
		_w16815_,
		_w16821_,
		_w17422_,
		_w17427_
	);
	LUT3 #(
		.INIT('h07)
	) name13380 (
		_w8841_,
		_w9082_,
		_w17427_,
		_w17428_
	);
	LUT4 #(
		.INIT('hfd00)
	) name13381 (
		_w5536_,
		_w7140_,
		_w7240_,
		_w17428_,
		_w17429_
	);
	LUT3 #(
		.INIT('h4e)
	) name13382 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[9]/P0001 ,
		_w17429_,
		_w17430_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13383 (
		_w16534_,
		_w16540_,
		_w16546_,
		_w17422_,
		_w17431_
	);
	LUT3 #(
		.INIT('h07)
	) name13384 (
		_w8974_,
		_w9082_,
		_w17431_,
		_w17432_
	);
	LUT4 #(
		.INIT('hfd00)
	) name13385 (
		_w5536_,
		_w8798_,
		_w8801_,
		_w17432_,
		_w17433_
	);
	LUT3 #(
		.INIT('h4e)
	) name13386 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[15]/P0001 ,
		_w17433_,
		_w17434_
	);
	LUT2 #(
		.INIT('h8)
	) name13387 (
		_w8952_,
		_w9082_,
		_w17435_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13388 (
		_w16565_,
		_w16571_,
		_w16577_,
		_w17422_,
		_w17436_
	);
	LUT4 #(
		.INIT('h00fd)
	) name13389 (
		_w5536_,
		_w8757_,
		_w8760_,
		_w17436_,
		_w17437_
	);
	LUT4 #(
		.INIT('he4ee)
	) name13390 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[14]/P0001 ,
		_w17435_,
		_w17437_,
		_w17438_
	);
	LUT2 #(
		.INIT('h4)
	) name13391 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[13]/P0001 ,
		_w17439_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13392 (
		_w16749_,
		_w16755_,
		_w16761_,
		_w17422_,
		_w17440_
	);
	LUT3 #(
		.INIT('h07)
	) name13393 (
		_w8929_,
		_w9082_,
		_w17440_,
		_w17441_
	);
	LUT4 #(
		.INIT('h80aa)
	) name13394 (
		\auctl_BSack_reg/NET0131 ,
		_w5536_,
		_w5760_,
		_w17441_,
		_w17442_
	);
	LUT2 #(
		.INIT('he)
	) name13395 (
		_w17439_,
		_w17442_,
		_w17443_
	);
	LUT2 #(
		.INIT('h4)
	) name13396 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[12]/P0001 ,
		_w17444_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13397 (
		_w16769_,
		_w16775_,
		_w16781_,
		_w17422_,
		_w17445_
	);
	LUT3 #(
		.INIT('h07)
	) name13398 (
		_w8907_,
		_w9082_,
		_w17445_,
		_w17446_
	);
	LUT4 #(
		.INIT('h80aa)
	) name13399 (
		\auctl_BSack_reg/NET0131 ,
		_w5536_,
		_w6758_,
		_w17446_,
		_w17447_
	);
	LUT2 #(
		.INIT('he)
	) name13400 (
		_w17444_,
		_w17447_,
		_w17448_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13401 (
		_w16829_,
		_w16835_,
		_w16841_,
		_w17422_,
		_w17449_
	);
	LUT3 #(
		.INIT('h07)
	) name13402 (
		_w8885_,
		_w9082_,
		_w17449_,
		_w17450_
	);
	LUT4 #(
		.INIT('hfd00)
	) name13403 (
		_w5536_,
		_w6263_,
		_w6362_,
		_w17450_,
		_w17451_
	);
	LUT3 #(
		.INIT('h4e)
	) name13404 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[11]/P0001 ,
		_w17451_,
		_w17452_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13405 (
		_w16849_,
		_w16855_,
		_w16861_,
		_w17422_,
		_w17453_
	);
	LUT3 #(
		.INIT('h07)
	) name13406 (
		_w8863_,
		_w9082_,
		_w17453_,
		_w17454_
	);
	LUT4 #(
		.INIT('hfd00)
	) name13407 (
		_w5536_,
		_w5937_,
		_w6038_,
		_w17454_,
		_w17455_
	);
	LUT3 #(
		.INIT('h4e)
	) name13408 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[10]/P0001 ,
		_w17455_,
		_w17456_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13409 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\sice_SPC_reg[1]/P0001 ,
		_w16506_,
		_w17323_,
		_w17457_
	);
	LUT4 #(
		.INIT('h0080)
	) name13410 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17457_,
		_w17458_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13411 (
		_w13327_,
		_w16705_,
		_w16719_,
		_w17458_,
		_w17459_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name13412 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\sice_SPC_reg[0]/P0001 ,
		_w16506_,
		_w17323_,
		_w17460_
	);
	LUT4 #(
		.INIT('h0080)
	) name13413 (
		_w4073_,
		_w4084_,
		_w13325_,
		_w17460_,
		_w17461_
	);
	LUT4 #(
		.INIT('h00fe)
	) name13414 (
		_w13327_,
		_w16725_,
		_w16739_,
		_w17461_,
		_w17462_
	);
	LUT4 #(
		.INIT('h2022)
	) name13415 (
		_w5536_,
		_w7793_,
		_w7903_,
		_w7905_,
		_w17463_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13416 (
		_w16586_,
		_w16592_,
		_w16598_,
		_w17422_,
		_w17464_
	);
	LUT4 #(
		.INIT('heee4)
	) name13417 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[7]/P0001 ,
		_w17463_,
		_w17464_,
		_w17465_
	);
	LUT4 #(
		.INIT('h2022)
	) name13418 (
		_w5536_,
		_w7927_,
		_w8040_,
		_w8042_,
		_w17466_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13419 (
		_w16606_,
		_w16612_,
		_w16618_,
		_w17422_,
		_w17467_
	);
	LUT4 #(
		.INIT('heee4)
	) name13420 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[6]/P0001 ,
		_w17466_,
		_w17467_,
		_w17468_
	);
	LUT4 #(
		.INIT('h2022)
	) name13421 (
		_w5536_,
		_w7592_,
		_w7707_,
		_w7709_,
		_w17469_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13422 (
		_w16626_,
		_w16632_,
		_w16638_,
		_w17422_,
		_w17470_
	);
	LUT4 #(
		.INIT('heee4)
	) name13423 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[5]/P0001 ,
		_w17469_,
		_w17470_,
		_w17471_
	);
	LUT4 #(
		.INIT('h2022)
	) name13424 (
		_w5536_,
		_w7257_,
		_w7375_,
		_w7377_,
		_w17472_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13425 (
		_w16646_,
		_w16652_,
		_w16658_,
		_w17422_,
		_w17473_
	);
	LUT4 #(
		.INIT('heee4)
	) name13426 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[4]/P0001 ,
		_w17472_,
		_w17473_,
		_w17474_
	);
	LUT4 #(
		.INIT('h2022)
	) name13427 (
		_w5536_,
		_w6054_,
		_w6173_,
		_w6175_,
		_w17475_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13428 (
		_w16666_,
		_w16672_,
		_w16678_,
		_w17422_,
		_w17476_
	);
	LUT4 #(
		.INIT('heee4)
	) name13429 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[3]/P0001 ,
		_w17475_,
		_w17476_,
		_w17477_
	);
	LUT4 #(
		.INIT('h2022)
	) name13430 (
		_w5536_,
		_w6378_,
		_w6498_,
		_w6500_,
		_w17478_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13431 (
		_w16686_,
		_w16692_,
		_w16698_,
		_w17422_,
		_w17479_
	);
	LUT4 #(
		.INIT('heee4)
	) name13432 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[2]/P0001 ,
		_w17478_,
		_w17479_,
		_w17480_
	);
	LUT2 #(
		.INIT('h4)
	) name13433 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[23]/P0001 ,
		_w17481_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13434 (
		_w16930_,
		_w16936_,
		_w16942_,
		_w17422_,
		_w17482_
	);
	LUT4 #(
		.INIT('haa80)
	) name13435 (
		\auctl_BSack_reg/NET0131 ,
		_w8821_,
		_w9082_,
		_w17482_,
		_w17483_
	);
	LUT2 #(
		.INIT('he)
	) name13436 (
		_w17481_,
		_w17483_,
		_w17484_
	);
	LUT2 #(
		.INIT('h4)
	) name13437 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[22]/P0001 ,
		_w17485_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13438 (
		_w16947_,
		_w16953_,
		_w16959_,
		_w17422_,
		_w17486_
	);
	LUT4 #(
		.INIT('haa80)
	) name13439 (
		\auctl_BSack_reg/NET0131 ,
		_w8781_,
		_w9082_,
		_w17486_,
		_w17487_
	);
	LUT2 #(
		.INIT('he)
	) name13440 (
		_w17485_,
		_w17487_,
		_w17488_
	);
	LUT2 #(
		.INIT('h4)
	) name13441 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[21]/P0001 ,
		_w17489_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13442 (
		_w17011_,
		_w17017_,
		_w17023_,
		_w17422_,
		_w17490_
	);
	LUT4 #(
		.INIT('haa80)
	) name13443 (
		\auctl_BSack_reg/NET0131 ,
		_w8740_,
		_w9082_,
		_w17490_,
		_w17491_
	);
	LUT2 #(
		.INIT('he)
	) name13444 (
		_w17489_,
		_w17491_,
		_w17492_
	);
	LUT2 #(
		.INIT('h4)
	) name13445 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[20]/P0001 ,
		_w17493_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13446 (
		_w17029_,
		_w17035_,
		_w17041_,
		_w17422_,
		_w17494_
	);
	LUT4 #(
		.INIT('haa80)
	) name13447 (
		\auctl_BSack_reg/NET0131 ,
		_w8717_,
		_w9082_,
		_w17494_,
		_w17495_
	);
	LUT2 #(
		.INIT('he)
	) name13448 (
		_w17493_,
		_w17495_,
		_w17496_
	);
	LUT4 #(
		.INIT('h2022)
	) name13449 (
		_w5536_,
		_w6774_,
		_w6894_,
		_w6896_,
		_w17497_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13450 (
		_w16706_,
		_w16712_,
		_w16718_,
		_w17422_,
		_w17498_
	);
	LUT4 #(
		.INIT('heee4)
	) name13451 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[1]/P0001 ,
		_w17497_,
		_w17498_,
		_w17499_
	);
	LUT4 #(
		.INIT('h00df)
	) name13452 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w9453_,
		_w9894_,
		_w12223_,
		_w17500_
	);
	LUT4 #(
		.INIT('h8a00)
	) name13453 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w11303_,
		_w17501_
	);
	LUT2 #(
		.INIT('h1)
	) name13454 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 ,
		_w17501_,
		_w17502_
	);
	LUT3 #(
		.INIT('h8a)
	) name13455 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11303_,
		_w11308_,
		_w17503_
	);
	LUT2 #(
		.INIT('h1)
	) name13456 (
		_w12220_,
		_w17501_,
		_w17504_
	);
	LUT2 #(
		.INIT('h2)
	) name13457 (
		_w17503_,
		_w17504_,
		_w17505_
	);
	LUT4 #(
		.INIT('hfe00)
	) name13458 (
		_w12006_,
		_w12007_,
		_w12220_,
		_w17505_,
		_w17506_
	);
	LUT4 #(
		.INIT('h1311)
	) name13459 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 ,
		_w11303_,
		_w11308_,
		_w17507_
	);
	LUT4 #(
		.INIT('h00ab)
	) name13460 (
		_w12224_,
		_w17502_,
		_w17506_,
		_w17507_,
		_w17508_
	);
	LUT2 #(
		.INIT('h2)
	) name13461 (
		_w17500_,
		_w17508_,
		_w17509_
	);
	LUT3 #(
		.INIT('h07)
	) name13462 (
		_w11624_,
		_w12239_,
		_w17509_,
		_w17510_
	);
	LUT4 #(
		.INIT('h4055)
	) name13463 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w11917_,
		_w11920_,
		_w11924_,
		_w17511_
	);
	LUT4 #(
		.INIT('h0040)
	) name13464 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w4856_,
		_w17512_
	);
	LUT2 #(
		.INIT('h1)
	) name13465 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w17513_
	);
	LUT4 #(
		.INIT('hfd20)
	) name13466 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w9470_,
		_w17513_,
		_w17514_
	);
	LUT3 #(
		.INIT('h01)
	) name13467 (
		_w17511_,
		_w17512_,
		_w17514_,
		_w17515_
	);
	LUT3 #(
		.INIT('hd0)
	) name13468 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w16289_,
		_w17516_
	);
	LUT4 #(
		.INIT('h8a00)
	) name13469 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w17516_,
		_w17517_
	);
	LUT4 #(
		.INIT('h0105)
	) name13470 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9853_,
		_w12118_,
		_w17518_
	);
	LUT3 #(
		.INIT('h02)
	) name13471 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w11313_,
		_w11314_,
		_w17519_
	);
	LUT4 #(
		.INIT('h4544)
	) name13472 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w9456_,
		_w12161_,
		_w12162_,
		_w17520_
	);
	LUT4 #(
		.INIT('h070f)
	) name13473 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17519_,
		_w17520_,
		_w17521_
	);
	LUT3 #(
		.INIT('h8a)
	) name13474 (
		_w17517_,
		_w17518_,
		_w17521_,
		_w17522_
	);
	LUT4 #(
		.INIT('h0002)
	) name13475 (
		\core_eu_em_mac_em_reg_s2_reg/P0000_reg_syn_2 ,
		_w16306_,
		_w16315_,
		_w16319_,
		_w17523_
	);
	LUT2 #(
		.INIT('h1)
	) name13476 (
		_w16314_,
		_w17523_,
		_w17524_
	);
	LUT3 #(
		.INIT('h8b)
	) name13477 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w16322_,
		_w16504_,
		_w17525_
	);
	LUT3 #(
		.INIT('h4c)
	) name13478 (
		\core_eu_em_mac_em_reg_s1_reg/P0000_reg_syn_2 ,
		_w16320_,
		_w16322_,
		_w17526_
	);
	LUT3 #(
		.INIT('h02)
	) name13479 (
		_w11318_,
		_w17525_,
		_w17526_,
		_w17527_
	);
	LUT4 #(
		.INIT('hacc0)
	) name13480 (
		_w6501_,
		_w8863_,
		_w17525_,
		_w17526_,
		_w17528_
	);
	LUT3 #(
		.INIT('ha8)
	) name13481 (
		_w17524_,
		_w17527_,
		_w17528_,
		_w17529_
	);
	LUT4 #(
		.INIT('h8088)
	) name13482 (
		_w11306_,
		_w11925_,
		_w16286_,
		_w16300_,
		_w17530_
	);
	LUT4 #(
		.INIT('h5100)
	) name13483 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w16296_,
		_w17531_
	);
	LUT3 #(
		.INIT('hd0)
	) name13484 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w16301_,
		_w17532_
	);
	LUT2 #(
		.INIT('h1)
	) name13485 (
		_w17531_,
		_w17532_,
		_w17533_
	);
	LUT3 #(
		.INIT('h08)
	) name13486 (
		_w5713_,
		_w17530_,
		_w17533_,
		_w17534_
	);
	LUT4 #(
		.INIT('h0d00)
	) name13487 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w5713_,
		_w16296_,
		_w17535_
	);
	LUT2 #(
		.INIT('h8)
	) name13488 (
		_w17530_,
		_w17535_,
		_w17536_
	);
	LUT3 #(
		.INIT('h80)
	) name13489 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w17530_,
		_w17535_,
		_w17537_
	);
	LUT2 #(
		.INIT('h1)
	) name13490 (
		_w17534_,
		_w17537_,
		_w17538_
	);
	LUT4 #(
		.INIT('h7500)
	) name13491 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w16307_,
		_w17539_
	);
	LUT3 #(
		.INIT('h20)
	) name13492 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w9463_,
		_w17540_
	);
	LUT3 #(
		.INIT('h54)
	) name13493 (
		_w6484_,
		_w17539_,
		_w17540_,
		_w17541_
	);
	LUT4 #(
		.INIT('h7500)
	) name13494 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w17531_,
		_w17542_
	);
	LUT3 #(
		.INIT('h20)
	) name13495 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w9467_,
		_w17543_
	);
	LUT3 #(
		.INIT('h54)
	) name13496 (
		_w6477_,
		_w17542_,
		_w17543_,
		_w17544_
	);
	LUT3 #(
		.INIT('h20)
	) name13497 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w9466_,
		_w17545_
	);
	LUT4 #(
		.INIT('h7500)
	) name13498 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w17532_,
		_w17546_
	);
	LUT3 #(
		.INIT('h54)
	) name13499 (
		_w6481_,
		_w17545_,
		_w17546_,
		_w17547_
	);
	LUT3 #(
		.INIT('h01)
	) name13500 (
		_w17544_,
		_w17547_,
		_w17541_,
		_w17548_
	);
	LUT2 #(
		.INIT('h8)
	) name13501 (
		_w17538_,
		_w17548_,
		_w17549_
	);
	LUT2 #(
		.INIT('h8)
	) name13502 (
		_w17525_,
		_w17549_,
		_w17550_
	);
	LUT4 #(
		.INIT('h1310)
	) name13503 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w6501_,
		_w16322_,
		_w16504_,
		_w17551_
	);
	LUT3 #(
		.INIT('h04)
	) name13504 (
		_w17524_,
		_w17526_,
		_w17551_,
		_w17552_
	);
	LUT2 #(
		.INIT('h2)
	) name13505 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w17553_
	);
	LUT3 #(
		.INIT('hd0)
	) name13506 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w16284_,
		_w17554_
	);
	LUT4 #(
		.INIT('h8a00)
	) name13507 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w17554_,
		_w17555_
	);
	LUT2 #(
		.INIT('h8)
	) name13508 (
		_w17553_,
		_w17555_,
		_w17556_
	);
	LUT2 #(
		.INIT('h4)
	) name13509 (
		_w13249_,
		_w17556_,
		_w17557_
	);
	LUT3 #(
		.INIT('h20)
	) name13510 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w9464_,
		_w17558_
	);
	LUT4 #(
		.INIT('h7500)
	) name13511 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w17516_,
		_w17559_
	);
	LUT3 #(
		.INIT('h54)
	) name13512 (
		_w6458_,
		_w17558_,
		_w17559_,
		_w17560_
	);
	LUT2 #(
		.INIT('h1)
	) name13513 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w17561_
	);
	LUT3 #(
		.INIT('he4)
	) name13514 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTSR0_E_reg/P0001 ,
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w17562_
	);
	LUT4 #(
		.INIT('h8a00)
	) name13515 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w17562_,
		_w17563_
	);
	LUT4 #(
		.INIT('hc400)
	) name13516 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		\core_c_dec_accPM_E_reg/P0001 ,
		_w4855_,
		_w16284_,
		_w17564_
	);
	LUT3 #(
		.INIT('h80)
	) name13517 (
		_w8863_,
		_w17563_,
		_w17564_,
		_w17565_
	);
	LUT4 #(
		.INIT('h3100)
	) name13518 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		\core_c_dec_accPM_E_reg/P0001 ,
		_w4855_,
		_w16284_,
		_w17566_
	);
	LUT3 #(
		.INIT('h80)
	) name13519 (
		_w6501_,
		_w17563_,
		_w17566_,
		_w17567_
	);
	LUT3 #(
		.INIT('h01)
	) name13520 (
		_w17565_,
		_w17567_,
		_w17560_,
		_w17568_
	);
	LUT2 #(
		.INIT('h8)
	) name13521 (
		_w17561_,
		_w17555_,
		_w17569_
	);
	LUT3 #(
		.INIT('h70)
	) name13522 (
		_w13270_,
		_w13282_,
		_w17569_,
		_w17570_
	);
	LUT4 #(
		.INIT('h0800)
	) name13523 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w9460_,
		_w17571_
	);
	LUT4 #(
		.INIT('h7500)
	) name13524 (
		_w11925_,
		_w16286_,
		_w16300_,
		_w17554_,
		_w17572_
	);
	LUT4 #(
		.INIT('h3230)
	) name13525 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6473_,
		_w17571_,
		_w17572_,
		_w17573_
	);
	LUT3 #(
		.INIT('h20)
	) name13526 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w17574_
	);
	LUT3 #(
		.INIT('h20)
	) name13527 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w17574_,
		_w17575_
	);
	LUT4 #(
		.INIT('h3310)
	) name13528 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6471_,
		_w17572_,
		_w17575_,
		_w17576_
	);
	LUT2 #(
		.INIT('h1)
	) name13529 (
		_w17573_,
		_w17576_,
		_w17577_
	);
	LUT3 #(
		.INIT('h40)
	) name13530 (
		_w17570_,
		_w17568_,
		_w17577_,
		_w17578_
	);
	LUT2 #(
		.INIT('h4)
	) name13531 (
		_w17557_,
		_w17578_,
		_w17579_
	);
	LUT3 #(
		.INIT('hb0)
	) name13532 (
		_w17550_,
		_w17552_,
		_w17579_,
		_w17580_
	);
	LUT2 #(
		.INIT('h4)
	) name13533 (
		_w17529_,
		_w17580_,
		_w17581_
	);
	LUT3 #(
		.INIT('h01)
	) name13534 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w17582_
	);
	LUT3 #(
		.INIT('he4)
	) name13535 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTMX0_E_reg/P0001 ,
		\core_c_dec_MTMX1_E_reg/P0001 ,
		_w17583_
	);
	LUT2 #(
		.INIT('h8)
	) name13536 (
		_w17582_,
		_w17583_,
		_w17584_
	);
	LUT3 #(
		.INIT('h40)
	) name13537 (
		_w4856_,
		_w11925_,
		_w17584_,
		_w17585_
	);
	LUT3 #(
		.INIT('h08)
	) name13538 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		\core_c_dec_MACop_E_reg/P0001 ,
		_w4855_,
		_w17586_
	);
	LUT2 #(
		.INIT('h1)
	) name13539 (
		_w11926_,
		_w17586_,
		_w17587_
	);
	LUT4 #(
		.INIT('h3353)
	) name13540 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w17588_
	);
	LUT2 #(
		.INIT('h2)
	) name13541 (
		_w6486_,
		_w17588_,
		_w17589_
	);
	LUT2 #(
		.INIT('h8)
	) name13542 (
		_w6479_,
		_w17588_,
		_w17590_
	);
	LUT3 #(
		.INIT('h01)
	) name13543 (
		_w17590_,
		_w17585_,
		_w17589_,
		_w17591_
	);
	LUT2 #(
		.INIT('h1)
	) name13544 (
		_w17587_,
		_w17591_,
		_w17592_
	);
	LUT4 #(
		.INIT('hef00)
	) name13545 (
		_w11313_,
		_w11314_,
		_w17585_,
		_w17592_,
		_w17593_
	);
	LUT3 #(
		.INIT('h01)
	) name13546 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w11926_,
		_w17586_,
		_w17594_
	);
	LUT2 #(
		.INIT('h1)
	) name13547 (
		_w17515_,
		_w17594_,
		_w17595_
	);
	LUT2 #(
		.INIT('h4)
	) name13548 (
		_w17593_,
		_w17595_,
		_w17596_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13549 (
		_w17515_,
		_w17522_,
		_w17581_,
		_w17596_,
		_w17597_
	);
	LUT2 #(
		.INIT('h4)
	) name13550 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[19]/P0001 ,
		_w17598_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13551 (
		_w17047_,
		_w17053_,
		_w17059_,
		_w17422_,
		_w17599_
	);
	LUT4 #(
		.INIT('haa80)
	) name13552 (
		\auctl_BSack_reg/NET0131 ,
		_w8694_,
		_w9082_,
		_w17599_,
		_w17600_
	);
	LUT2 #(
		.INIT('he)
	) name13553 (
		_w17598_,
		_w17600_,
		_w17601_
	);
	LUT2 #(
		.INIT('h4)
	) name13554 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[18]/P0001 ,
		_w17602_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13555 (
		_w17065_,
		_w17071_,
		_w17077_,
		_w17422_,
		_w17603_
	);
	LUT4 #(
		.INIT('haa80)
	) name13556 (
		\auctl_BSack_reg/NET0131 ,
		_w8671_,
		_w9082_,
		_w17603_,
		_w17604_
	);
	LUT2 #(
		.INIT('he)
	) name13557 (
		_w17602_,
		_w17604_,
		_w17605_
	);
	LUT2 #(
		.INIT('h4)
	) name13558 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[17]/P0001 ,
		_w17606_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13559 (
		_w16975_,
		_w16981_,
		_w16987_,
		_w17422_,
		_w17607_
	);
	LUT4 #(
		.INIT('haa80)
	) name13560 (
		\auctl_BSack_reg/NET0131 ,
		_w9021_,
		_w9082_,
		_w17607_,
		_w17608_
	);
	LUT2 #(
		.INIT('he)
	) name13561 (
		_w17606_,
		_w17608_,
		_w17609_
	);
	LUT2 #(
		.INIT('h4)
	) name13562 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[16]/P0001 ,
		_w17610_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13563 (
		_w16993_,
		_w16999_,
		_w17005_,
		_w17422_,
		_w17611_
	);
	LUT4 #(
		.INIT('haa80)
	) name13564 (
		\auctl_BSack_reg/NET0131 ,
		_w8998_,
		_w9082_,
		_w17611_,
		_w17612_
	);
	LUT2 #(
		.INIT('he)
	) name13565 (
		_w17610_,
		_w17612_,
		_w17613_
	);
	LUT4 #(
		.INIT('h2022)
	) name13566 (
		_w5536_,
		_w5784_,
		_w5911_,
		_w5913_,
		_w17614_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13567 (
		_w16726_,
		_w16732_,
		_w16738_,
		_w17422_,
		_w17615_
	);
	LUT4 #(
		.INIT('heee4)
	) name13568 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[0]/P0001 ,
		_w17614_,
		_w17615_,
		_w17616_
	);
	LUT4 #(
		.INIT('h3353)
	) name13569 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w17617_
	);
	LUT4 #(
		.INIT('h3353)
	) name13570 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4855_,
		_w17618_
	);
	LUT2 #(
		.INIT('h1)
	) name13571 (
		_w17617_,
		_w17618_,
		_w17619_
	);
	LUT2 #(
		.INIT('h2)
	) name13572 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_MTMY1_E_reg/P0001 ,
		_w17620_
	);
	LUT4 #(
		.INIT('h0504)
	) name13573 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_MTMY0_E_reg/P0001 ,
		_w17621_
	);
	LUT2 #(
		.INIT('h4)
	) name13574 (
		_w17620_,
		_w17621_,
		_w17622_
	);
	LUT3 #(
		.INIT('h70)
	) name13575 (
		_w11924_,
		_w13505_,
		_w17622_,
		_w17623_
	);
	LUT3 #(
		.INIT('h40)
	) name13576 (
		_w4856_,
		_w11925_,
		_w17623_,
		_w17624_
	);
	LUT4 #(
		.INIT('hfd08)
	) name13577 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		\core_eu_em_mac_em_reg_Sq_E_reg/P0001 ,
		_w4855_,
		_w13505_,
		_w17625_
	);
	LUT3 #(
		.INIT('h10)
	) name13578 (
		_w17619_,
		_w17624_,
		_w17625_,
		_w17626_
	);
	LUT2 #(
		.INIT('h8)
	) name13579 (
		_w17515_,
		_w17626_,
		_w17627_
	);
	LUT4 #(
		.INIT('h0100)
	) name13580 (
		_w17512_,
		_w17619_,
		_w17624_,
		_w17625_,
		_w17628_
	);
	LUT3 #(
		.INIT('h10)
	) name13581 (
		\core_c_dec_Double_E_reg/P0001 ,
		_w4104_,
		_w17624_,
		_w17629_
	);
	LUT4 #(
		.INIT('h5540)
	) name13582 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w17585_,
		_w17628_,
		_w17629_,
		_w17630_
	);
	LUT4 #(
		.INIT('h4500)
	) name13583 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w17630_,
		_w17631_
	);
	LUT3 #(
		.INIT('h10)
	) name13584 (
		_w4104_,
		_w13819_,
		_w17624_,
		_w17632_
	);
	LUT4 #(
		.INIT('h007f)
	) name13585 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w17585_,
		_w17628_,
		_w17632_,
		_w17633_
	);
	LUT3 #(
		.INIT('h02)
	) name13586 (
		_w8863_,
		_w17630_,
		_w17633_,
		_w17634_
	);
	LUT4 #(
		.INIT('h0001)
	) name13587 (
		_w17512_,
		_w17619_,
		_w17624_,
		_w17625_,
		_w17635_
	);
	LUT3 #(
		.INIT('he4)
	) name13588 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[2]/P0001 ,
		_w17636_
	);
	LUT3 #(
		.INIT('h40)
	) name13589 (
		_w17617_,
		_w17635_,
		_w17636_,
		_w17637_
	);
	LUT3 #(
		.INIT('h35)
	) name13590 (
		_w6488_,
		_w6490_,
		_w17618_,
		_w17638_
	);
	LUT3 #(
		.INIT('h80)
	) name13591 (
		_w17617_,
		_w17635_,
		_w17638_,
		_w17639_
	);
	LUT3 #(
		.INIT('h80)
	) name13592 (
		_w17514_,
		_w17591_,
		_w17628_,
		_w17640_
	);
	LUT3 #(
		.INIT('h01)
	) name13593 (
		_w17639_,
		_w17640_,
		_w17637_,
		_w17641_
	);
	LUT2 #(
		.INIT('h4)
	) name13594 (
		_w17634_,
		_w17641_,
		_w17642_
	);
	LUT3 #(
		.INIT('ha8)
	) name13595 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 ,
		_w17511_,
		_w17512_,
		_w17643_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13596 (
		_w17511_,
		_w17631_,
		_w17642_,
		_w17643_,
		_w17644_
	);
	LUT2 #(
		.INIT('h1)
	) name13597 (
		_w17627_,
		_w17644_,
		_w17645_
	);
	LUT4 #(
		.INIT('hffb0)
	) name13598 (
		_w17522_,
		_w17581_,
		_w17627_,
		_w17645_,
		_w17646_
	);
	LUT4 #(
		.INIT('h0400)
	) name13599 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[14]/NET0131 ,
		_w17647_
	);
	LUT4 #(
		.INIT('h0603)
	) name13600 (
		\tm_TCR_TMP_reg[13]/NET0131 ,
		\tm_TCR_TMP_reg[14]/NET0131 ,
		_w14103_,
		_w15996_,
		_w17648_
	);
	LUT4 #(
		.INIT('h2333)
	) name13601 (
		\tm_tpr_reg_DO_reg[14]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w17649_
	);
	LUT3 #(
		.INIT('hba)
	) name13602 (
		_w17647_,
		_w17648_,
		_w17649_,
		_w17650_
	);
	LUT3 #(
		.INIT('h13)
	) name13603 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 ,
		_w11300_,
		_w17651_
	);
	LUT4 #(
		.INIT('hccc8)
	) name13604 (
		_w11310_,
		_w11312_,
		_w12006_,
		_w12007_,
		_w17652_
	);
	LUT4 #(
		.INIT('h2322)
	) name13605 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 ,
		_w11303_,
		_w11308_,
		_w17653_
	);
	LUT4 #(
		.INIT('h00ab)
	) name13606 (
		_w11320_,
		_w17651_,
		_w17652_,
		_w17653_,
		_w17654_
	);
	LUT2 #(
		.INIT('h2)
	) name13607 (
		_w11325_,
		_w17654_,
		_w17655_
	);
	LUT3 #(
		.INIT('h07)
	) name13608 (
		_w9946_,
		_w12239_,
		_w17655_,
		_w17656_
	);
	LUT3 #(
		.INIT('hb0)
	) name13609 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w17657_
	);
	LUT3 #(
		.INIT('hd0)
	) name13610 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w13138_,
		_w17657_,
		_w17658_
	);
	LUT4 #(
		.INIT('h4500)
	) name13611 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w13161_,
		_w17659_
	);
	LUT3 #(
		.INIT('h31)
	) name13612 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13161_,
		_w17660_
	);
	LUT4 #(
		.INIT('h4544)
	) name13613 (
		_w13158_,
		_w17658_,
		_w17659_,
		_w17660_,
		_w17661_
	);
	LUT3 #(
		.INIT('h04)
	) name13614 (
		\sport0_rxctl_RXSHT_reg[0]/P0001 ,
		\sport0_rxctl_a_sync1_reg/P0001 ,
		\sport0_rxctl_a_sync2_reg/P0001 ,
		_w17662_
	);
	LUT2 #(
		.INIT('h1)
	) name13615 (
		_w17661_,
		_w17662_,
		_w17663_
	);
	LUT2 #(
		.INIT('h4)
	) name13616 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w17664_
	);
	LUT3 #(
		.INIT('h40)
	) name13617 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w17665_
	);
	LUT4 #(
		.INIT('h8000)
	) name13618 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w17666_
	);
	LUT4 #(
		.INIT('h8000)
	) name13619 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[5]/NET0131 ,
		_w17666_,
		_w17667_
	);
	LUT3 #(
		.INIT('h80)
	) name13620 (
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[7]/NET0131 ,
		_w17667_,
		_w17668_
	);
	LUT4 #(
		.INIT('h8000)
	) name13621 (
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[8]/NET0131 ,
		_w17667_,
		_w17669_
	);
	LUT2 #(
		.INIT('h8)
	) name13622 (
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w17669_,
		_w17670_
	);
	LUT3 #(
		.INIT('h80)
	) name13623 (
		\sport1_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w17669_,
		_w17671_
	);
	LUT4 #(
		.INIT('h8000)
	) name13624 (
		\sport1_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w17669_,
		_w17672_
	);
	LUT3 #(
		.INIT('h80)
	) name13625 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[13]/NET0131 ,
		_w17672_,
		_w17673_
	);
	LUT4 #(
		.INIT('h8000)
	) name13626 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[14]/NET0131 ,
		_w17672_,
		_w17674_
	);
	LUT2 #(
		.INIT('h1)
	) name13627 (
		\IRFS1_pad ,
		\ITFS1_pad ,
		_w17675_
	);
	LUT4 #(
		.INIT('hf531)
	) name13628 (
		\sport1_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[14]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w17676_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13629 (
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w17677_
	);
	LUT4 #(
		.INIT('hf531)
	) name13630 (
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w17678_
	);
	LUT4 #(
		.INIT('hf531)
	) name13631 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w17679_
	);
	LUT4 #(
		.INIT('h8000)
	) name13632 (
		_w17678_,
		_w17679_,
		_w17676_,
		_w17677_,
		_w17680_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13633 (
		\sport1_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[15]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w17681_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13634 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w17682_
	);
	LUT4 #(
		.INIT('h8caf)
	) name13635 (
		\sport1_cfg_FSi_cnt_reg[14]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w17683_
	);
	LUT4 #(
		.INIT('haf23)
	) name13636 (
		\sport1_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w17684_
	);
	LUT4 #(
		.INIT('h8000)
	) name13637 (
		_w17683_,
		_w17684_,
		_w17681_,
		_w17682_,
		_w17685_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13638 (
		\sport1_cfg_FSi_cnt_reg[5]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[8]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w17686_
	);
	LUT4 #(
		.INIT('h8caf)
	) name13639 (
		\sport1_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[5]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w17687_
	);
	LUT4 #(
		.INIT('haf23)
	) name13640 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[8]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w17688_
	);
	LUT4 #(
		.INIT('haf23)
	) name13641 (
		\sport1_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w17689_
	);
	LUT4 #(
		.INIT('h8000)
	) name13642 (
		_w17688_,
		_w17689_,
		_w17686_,
		_w17687_,
		_w17690_
	);
	LUT4 #(
		.INIT('h8caf)
	) name13643 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w17691_
	);
	LUT4 #(
		.INIT('hf531)
	) name13644 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[15]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w17692_
	);
	LUT4 #(
		.INIT('h8caf)
	) name13645 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w17693_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13646 (
		\sport1_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w17694_
	);
	LUT4 #(
		.INIT('h8000)
	) name13647 (
		_w17693_,
		_w17694_,
		_w17691_,
		_w17692_,
		_w17695_
	);
	LUT4 #(
		.INIT('h8000)
	) name13648 (
		_w17690_,
		_w17695_,
		_w17680_,
		_w17685_,
		_w17696_
	);
	LUT2 #(
		.INIT('h8)
	) name13649 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w17697_
	);
	LUT4 #(
		.INIT('h0155)
	) name13650 (
		_w17664_,
		_w17675_,
		_w17696_,
		_w17697_,
		_w17698_
	);
	LUT4 #(
		.INIT('hdcec)
	) name13651 (
		\sport1_cfg_FSi_cnt_reg[15]/NET0131 ,
		_w17665_,
		_w17698_,
		_w17674_,
		_w17699_
	);
	LUT2 #(
		.INIT('h4)
	) name13652 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w17700_
	);
	LUT3 #(
		.INIT('h40)
	) name13653 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w17701_
	);
	LUT4 #(
		.INIT('h8000)
	) name13654 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w17702_
	);
	LUT4 #(
		.INIT('h8000)
	) name13655 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[5]/NET0131 ,
		_w17702_,
		_w17703_
	);
	LUT3 #(
		.INIT('h80)
	) name13656 (
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[7]/NET0131 ,
		_w17703_,
		_w17704_
	);
	LUT4 #(
		.INIT('h8000)
	) name13657 (
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[8]/NET0131 ,
		_w17703_,
		_w17705_
	);
	LUT2 #(
		.INIT('h8)
	) name13658 (
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w17705_,
		_w17706_
	);
	LUT3 #(
		.INIT('h80)
	) name13659 (
		\sport0_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w17705_,
		_w17707_
	);
	LUT4 #(
		.INIT('h8000)
	) name13660 (
		\sport0_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w17705_,
		_w17708_
	);
	LUT3 #(
		.INIT('h80)
	) name13661 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[13]/NET0131 ,
		_w17708_,
		_w17709_
	);
	LUT4 #(
		.INIT('h8000)
	) name13662 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[14]/NET0131 ,
		_w17708_,
		_w17710_
	);
	LUT2 #(
		.INIT('h1)
	) name13663 (
		\IRFS0_pad ,
		\ITFS0_pad ,
		_w17711_
	);
	LUT4 #(
		.INIT('hf531)
	) name13664 (
		\sport0_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[14]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w17712_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13665 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w17713_
	);
	LUT4 #(
		.INIT('hf531)
	) name13666 (
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w17714_
	);
	LUT4 #(
		.INIT('hf531)
	) name13667 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w17715_
	);
	LUT4 #(
		.INIT('h8000)
	) name13668 (
		_w17714_,
		_w17715_,
		_w17712_,
		_w17713_,
		_w17716_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13669 (
		\sport0_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[15]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w17717_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13670 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w17718_
	);
	LUT4 #(
		.INIT('h8caf)
	) name13671 (
		\sport0_cfg_FSi_cnt_reg[14]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w17719_
	);
	LUT4 #(
		.INIT('haf23)
	) name13672 (
		\sport0_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w17720_
	);
	LUT4 #(
		.INIT('h8000)
	) name13673 (
		_w17719_,
		_w17720_,
		_w17717_,
		_w17718_,
		_w17721_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13674 (
		\sport0_cfg_FSi_cnt_reg[5]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[8]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w17722_
	);
	LUT4 #(
		.INIT('h8caf)
	) name13675 (
		\sport0_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[5]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w17723_
	);
	LUT4 #(
		.INIT('haf23)
	) name13676 (
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[8]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w17724_
	);
	LUT4 #(
		.INIT('haf23)
	) name13677 (
		\sport0_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w17725_
	);
	LUT4 #(
		.INIT('h8000)
	) name13678 (
		_w17724_,
		_w17725_,
		_w17722_,
		_w17723_,
		_w17726_
	);
	LUT4 #(
		.INIT('h8caf)
	) name13679 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w17727_
	);
	LUT4 #(
		.INIT('hf531)
	) name13680 (
		\sport0_cfg_FSi_cnt_reg[15]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w17728_
	);
	LUT4 #(
		.INIT('h8caf)
	) name13681 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w17729_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13682 (
		\sport0_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w17730_
	);
	LUT4 #(
		.INIT('h8000)
	) name13683 (
		_w17729_,
		_w17730_,
		_w17727_,
		_w17728_,
		_w17731_
	);
	LUT4 #(
		.INIT('h8000)
	) name13684 (
		_w17726_,
		_w17731_,
		_w17716_,
		_w17721_,
		_w17732_
	);
	LUT2 #(
		.INIT('h8)
	) name13685 (
		\memc_usysr_DO_reg[12]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w17733_
	);
	LUT4 #(
		.INIT('h0155)
	) name13686 (
		_w17700_,
		_w17711_,
		_w17732_,
		_w17733_,
		_w17734_
	);
	LUT4 #(
		.INIT('hdcec)
	) name13687 (
		\sport0_cfg_FSi_cnt_reg[15]/NET0131 ,
		_w17701_,
		_w17734_,
		_w17710_,
		_w17735_
	);
	LUT4 #(
		.INIT('h1b00)
	) name13688 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w11625_,
		_w17736_
	);
	LUT3 #(
		.INIT('h13)
	) name13689 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001 ,
		_w9894_,
		_w17737_
	);
	LUT4 #(
		.INIT('h0002)
	) name13690 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w17737_,
		_w17738_
	);
	LUT4 #(
		.INIT('h313b)
	) name13691 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001 ,
		_w11631_,
		_w11635_,
		_w17739_
	);
	LUT4 #(
		.INIT('h1055)
	) name13692 (
		_w11624_,
		_w17736_,
		_w17738_,
		_w17739_,
		_w17740_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13693 (
		_w11624_,
		_w12334_,
		_w12335_,
		_w17740_,
		_w17741_
	);
	LUT4 #(
		.INIT('he400)
	) name13694 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w11655_,
		_w17742_
	);
	LUT2 #(
		.INIT('h2)
	) name13695 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001 ,
		_w11656_,
		_w17743_
	);
	LUT3 #(
		.INIT('h01)
	) name13696 (
		_w9946_,
		_w11659_,
		_w17743_,
		_w17744_
	);
	LUT2 #(
		.INIT('h4)
	) name13697 (
		_w17742_,
		_w17744_,
		_w17745_
	);
	LUT4 #(
		.INIT('h00fd)
	) name13698 (
		_w9946_,
		_w12334_,
		_w12335_,
		_w17745_,
		_w17746_
	);
	LUT4 #(
		.INIT('hd200)
	) name13699 (
		T_IMS_pad,
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w17747_
	);
	LUT3 #(
		.INIT('hca)
	) name13700 (
		\sport1_txctl_TXSHT_reg[11]/P0001 ,
		\sport1_txctl_TX_reg[12]/P0001 ,
		_w14269_,
		_w17748_
	);
	LUT4 #(
		.INIT('h0105)
	) name13701 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9873_,
		_w12118_,
		_w17749_
	);
	LUT3 #(
		.INIT('h02)
	) name13702 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w11626_,
		_w11627_,
		_w17750_
	);
	LUT4 #(
		.INIT('h007f)
	) name13703 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w17750_,
		_w17751_
	);
	LUT3 #(
		.INIT('h8a)
	) name13704 (
		_w17517_,
		_w17749_,
		_w17751_,
		_w17752_
	);
	LUT4 #(
		.INIT('hff53)
	) name13705 (
		_w8952_,
		_w11318_,
		_w17525_,
		_w17526_,
		_w17753_
	);
	LUT2 #(
		.INIT('h2)
	) name13706 (
		_w17524_,
		_w17753_,
		_w17754_
	);
	LUT3 #(
		.INIT('h54)
	) name13707 (
		_w8026_,
		_w17539_,
		_w17540_,
		_w17755_
	);
	LUT3 #(
		.INIT('h54)
	) name13708 (
		_w8023_,
		_w17545_,
		_w17546_,
		_w17756_
	);
	LUT3 #(
		.INIT('h54)
	) name13709 (
		_w8019_,
		_w17542_,
		_w17543_,
		_w17757_
	);
	LUT3 #(
		.INIT('h01)
	) name13710 (
		_w17756_,
		_w17757_,
		_w17755_,
		_w17758_
	);
	LUT2 #(
		.INIT('h8)
	) name13711 (
		_w17538_,
		_w17758_,
		_w17759_
	);
	LUT2 #(
		.INIT('h8)
	) name13712 (
		_w17525_,
		_w17759_,
		_w17760_
	);
	LUT4 #(
		.INIT('h1310)
	) name13713 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8043_,
		_w16322_,
		_w16504_,
		_w17761_
	);
	LUT3 #(
		.INIT('h04)
	) name13714 (
		_w17524_,
		_w17526_,
		_w17761_,
		_w17762_
	);
	LUT4 #(
		.INIT('h2023)
	) name13715 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8043_,
		_w16322_,
		_w16504_,
		_w17763_
	);
	LUT4 #(
		.INIT('h1310)
	) name13716 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8952_,
		_w16322_,
		_w16504_,
		_w17764_
	);
	LUT4 #(
		.INIT('h0008)
	) name13717 (
		_w17524_,
		_w17526_,
		_w17764_,
		_w17763_,
		_w17765_
	);
	LUT4 #(
		.INIT('h3310)
	) name13718 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w8011_,
		_w17572_,
		_w17575_,
		_w17766_
	);
	LUT4 #(
		.INIT('h3230)
	) name13719 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w8015_,
		_w17571_,
		_w17572_,
		_w17767_
	);
	LUT4 #(
		.INIT('h008f)
	) name13720 (
		_w11966_,
		_w11981_,
		_w17569_,
		_w17767_,
		_w17768_
	);
	LUT2 #(
		.INIT('h4)
	) name13721 (
		_w17766_,
		_w17768_,
		_w17769_
	);
	LUT3 #(
		.INIT('h80)
	) name13722 (
		_w8952_,
		_w17563_,
		_w17564_,
		_w17770_
	);
	LUT3 #(
		.INIT('h54)
	) name13723 (
		_w7934_,
		_w17558_,
		_w17559_,
		_w17771_
	);
	LUT3 #(
		.INIT('h80)
	) name13724 (
		_w8043_,
		_w17563_,
		_w17566_,
		_w17772_
	);
	LUT3 #(
		.INIT('h01)
	) name13725 (
		_w17771_,
		_w17772_,
		_w17770_,
		_w17773_
	);
	LUT3 #(
		.INIT('hb0)
	) name13726 (
		_w11913_,
		_w17556_,
		_w17773_,
		_w17774_
	);
	LUT2 #(
		.INIT('h8)
	) name13727 (
		_w17769_,
		_w17774_,
		_w17775_
	);
	LUT4 #(
		.INIT('h4500)
	) name13728 (
		_w17765_,
		_w17760_,
		_w17762_,
		_w17775_,
		_w17776_
	);
	LUT2 #(
		.INIT('h4)
	) name13729 (
		_w17754_,
		_w17776_,
		_w17777_
	);
	LUT2 #(
		.INIT('h2)
	) name13730 (
		_w8028_,
		_w17588_,
		_w17778_
	);
	LUT2 #(
		.INIT('h8)
	) name13731 (
		_w8021_,
		_w17588_,
		_w17779_
	);
	LUT3 #(
		.INIT('h01)
	) name13732 (
		_w17585_,
		_w17779_,
		_w17778_,
		_w17780_
	);
	LUT2 #(
		.INIT('h1)
	) name13733 (
		_w17587_,
		_w17780_,
		_w17781_
	);
	LUT4 #(
		.INIT('hef00)
	) name13734 (
		_w11626_,
		_w11627_,
		_w17585_,
		_w17781_,
		_w17782_
	);
	LUT3 #(
		.INIT('h01)
	) name13735 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w11926_,
		_w17586_,
		_w17783_
	);
	LUT2 #(
		.INIT('h1)
	) name13736 (
		_w17515_,
		_w17783_,
		_w17784_
	);
	LUT2 #(
		.INIT('h4)
	) name13737 (
		_w17782_,
		_w17784_,
		_w17785_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13738 (
		_w17515_,
		_w17752_,
		_w17777_,
		_w17785_,
		_w17786_
	);
	LUT4 #(
		.INIT('h0105)
	) name13739 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9878_,
		_w12118_,
		_w17787_
	);
	LUT3 #(
		.INIT('h02)
	) name13740 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w12736_,
		_w12737_,
		_w17788_
	);
	LUT4 #(
		.INIT('h007f)
	) name13741 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w17788_,
		_w17789_
	);
	LUT3 #(
		.INIT('h8a)
	) name13742 (
		_w17517_,
		_w17787_,
		_w17789_,
		_w17790_
	);
	LUT4 #(
		.INIT('hacc0)
	) name13743 (
		_w7710_,
		_w8929_,
		_w17525_,
		_w17526_,
		_w17791_
	);
	LUT3 #(
		.INIT('ha8)
	) name13744 (
		_w17524_,
		_w17527_,
		_w17791_,
		_w17792_
	);
	LUT3 #(
		.INIT('h54)
	) name13745 (
		_w7668_,
		_w17545_,
		_w17546_,
		_w17793_
	);
	LUT3 #(
		.INIT('h54)
	) name13746 (
		_w7664_,
		_w17539_,
		_w17540_,
		_w17794_
	);
	LUT3 #(
		.INIT('h54)
	) name13747 (
		_w7671_,
		_w17542_,
		_w17543_,
		_w17795_
	);
	LUT3 #(
		.INIT('h01)
	) name13748 (
		_w17794_,
		_w17795_,
		_w17793_,
		_w17796_
	);
	LUT2 #(
		.INIT('h8)
	) name13749 (
		_w17538_,
		_w17796_,
		_w17797_
	);
	LUT2 #(
		.INIT('h8)
	) name13750 (
		_w17525_,
		_w17797_,
		_w17798_
	);
	LUT4 #(
		.INIT('h1310)
	) name13751 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w7710_,
		_w16322_,
		_w16504_,
		_w17799_
	);
	LUT3 #(
		.INIT('h04)
	) name13752 (
		_w17524_,
		_w17526_,
		_w17799_,
		_w17800_
	);
	LUT3 #(
		.INIT('h40)
	) name13753 (
		_w11430_,
		_w11871_,
		_w12629_,
		_w17801_
	);
	LUT2 #(
		.INIT('h8)
	) name13754 (
		_w11587_,
		_w11860_,
		_w17802_
	);
	LUT4 #(
		.INIT('hfca8)
	) name13755 (
		_w11534_,
		_w11492_,
		_w11512_,
		_w11454_,
		_w17803_
	);
	LUT2 #(
		.INIT('h4)
	) name13756 (
		_w17802_,
		_w17803_,
		_w17804_
	);
	LUT4 #(
		.INIT('h0080)
	) name13757 (
		_w11389_,
		_w11386_,
		_w11476_,
		_w11498_,
		_w17805_
	);
	LUT3 #(
		.INIT('h80)
	) name13758 (
		_w11389_,
		_w11541_,
		_w11445_,
		_w17806_
	);
	LUT4 #(
		.INIT('ha820)
	) name13759 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001 ,
		_w17807_
	);
	LUT4 #(
		.INIT('h007f)
	) name13760 (
		_w11473_,
		_w11389_,
		_w11341_,
		_w17807_,
		_w17808_
	);
	LUT3 #(
		.INIT('h10)
	) name13761 (
		_w17805_,
		_w17806_,
		_w17808_,
		_w17809_
	);
	LUT4 #(
		.INIT('h0f04)
	) name13762 (
		_w11444_,
		_w11428_,
		_w11489_,
		_w11455_,
		_w17810_
	);
	LUT3 #(
		.INIT('h0e)
	) name13763 (
		_w11530_,
		_w11471_,
		_w17810_,
		_w17811_
	);
	LUT3 #(
		.INIT('ha8)
	) name13764 (
		_w11532_,
		_w11973_,
		_w11974_,
		_w17812_
	);
	LUT4 #(
		.INIT('h2000)
	) name13765 (
		_w11554_,
		_w17812_,
		_w17809_,
		_w17811_,
		_w17813_
	);
	LUT2 #(
		.INIT('h8)
	) name13766 (
		_w17804_,
		_w17813_,
		_w17814_
	);
	LUT3 #(
		.INIT('hc8)
	) name13767 (
		_w11409_,
		_w11854_,
		_w11896_,
		_w17815_
	);
	LUT3 #(
		.INIT('hc8)
	) name13768 (
		_w11555_,
		_w11458_,
		_w12568_,
		_w17816_
	);
	LUT3 #(
		.INIT('h54)
	) name13769 (
		_w11514_,
		_w11522_,
		_w11523_,
		_w17817_
	);
	LUT3 #(
		.INIT('he0)
	) name13770 (
		_w11410_,
		_w11558_,
		_w11499_,
		_w17818_
	);
	LUT4 #(
		.INIT('h0001)
	) name13771 (
		_w17815_,
		_w17816_,
		_w17817_,
		_w17818_,
		_w17819_
	);
	LUT3 #(
		.INIT('ha8)
	) name13772 (
		_w11537_,
		_w11435_,
		_w12455_,
		_w17820_
	);
	LUT3 #(
		.INIT('h0d)
	) name13773 (
		_w11406_,
		_w11585_,
		_w12446_,
		_w17821_
	);
	LUT4 #(
		.INIT('h0001)
	) name13774 (
		_w11403_,
		_w11407_,
		_w11436_,
		_w11885_,
		_w17822_
	);
	LUT3 #(
		.INIT('hc8)
	) name13775 (
		_w11588_,
		_w11495_,
		_w12496_,
		_w17823_
	);
	LUT4 #(
		.INIT('h0040)
	) name13776 (
		_w17820_,
		_w17821_,
		_w17822_,
		_w17823_,
		_w17824_
	);
	LUT3 #(
		.INIT('h80)
	) name13777 (
		_w11902_,
		_w17819_,
		_w17824_,
		_w17825_
	);
	LUT4 #(
		.INIT('h8000)
	) name13778 (
		_w11837_,
		_w17801_,
		_w17814_,
		_w17825_,
		_w17826_
	);
	LUT2 #(
		.INIT('h2)
	) name13779 (
		_w17556_,
		_w17826_,
		_w17827_
	);
	LUT3 #(
		.INIT('h80)
	) name13780 (
		_w8929_,
		_w17563_,
		_w17564_,
		_w17828_
	);
	LUT3 #(
		.INIT('h54)
	) name13781 (
		_w7686_,
		_w17558_,
		_w17559_,
		_w17829_
	);
	LUT3 #(
		.INIT('h80)
	) name13782 (
		_w7710_,
		_w17563_,
		_w17566_,
		_w17830_
	);
	LUT3 #(
		.INIT('h01)
	) name13783 (
		_w17829_,
		_w17830_,
		_w17828_,
		_w17831_
	);
	LUT3 #(
		.INIT('h70)
	) name13784 (
		_w12740_,
		_w12757_,
		_w17569_,
		_w17832_
	);
	LUT4 #(
		.INIT('h3310)
	) name13785 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7695_,
		_w17572_,
		_w17575_,
		_w17833_
	);
	LUT4 #(
		.INIT('h3230)
	) name13786 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7699_,
		_w17571_,
		_w17572_,
		_w17834_
	);
	LUT2 #(
		.INIT('h1)
	) name13787 (
		_w17833_,
		_w17834_,
		_w17835_
	);
	LUT3 #(
		.INIT('h40)
	) name13788 (
		_w17832_,
		_w17831_,
		_w17835_,
		_w17836_
	);
	LUT2 #(
		.INIT('h4)
	) name13789 (
		_w17827_,
		_w17836_,
		_w17837_
	);
	LUT3 #(
		.INIT('hb0)
	) name13790 (
		_w17798_,
		_w17800_,
		_w17837_,
		_w17838_
	);
	LUT2 #(
		.INIT('h4)
	) name13791 (
		_w17792_,
		_w17838_,
		_w17839_
	);
	LUT2 #(
		.INIT('h2)
	) name13792 (
		_w7675_,
		_w17588_,
		_w17840_
	);
	LUT2 #(
		.INIT('h8)
	) name13793 (
		_w7666_,
		_w17588_,
		_w17841_
	);
	LUT3 #(
		.INIT('h01)
	) name13794 (
		_w17585_,
		_w17841_,
		_w17840_,
		_w17842_
	);
	LUT2 #(
		.INIT('h1)
	) name13795 (
		_w17587_,
		_w17842_,
		_w17843_
	);
	LUT4 #(
		.INIT('hef00)
	) name13796 (
		_w12736_,
		_w12737_,
		_w17585_,
		_w17843_,
		_w17844_
	);
	LUT3 #(
		.INIT('h01)
	) name13797 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w11926_,
		_w17586_,
		_w17845_
	);
	LUT2 #(
		.INIT('h1)
	) name13798 (
		_w17515_,
		_w17845_,
		_w17846_
	);
	LUT2 #(
		.INIT('h4)
	) name13799 (
		_w17844_,
		_w17846_,
		_w17847_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13800 (
		_w17515_,
		_w17790_,
		_w17839_,
		_w17847_,
		_w17848_
	);
	LUT4 #(
		.INIT('h0105)
	) name13801 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9860_,
		_w12118_,
		_w17849_
	);
	LUT3 #(
		.INIT('h02)
	) name13802 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w12626_,
		_w12627_,
		_w17850_
	);
	LUT4 #(
		.INIT('h007f)
	) name13803 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w17850_,
		_w17851_
	);
	LUT3 #(
		.INIT('h8a)
	) name13804 (
		_w17517_,
		_w17849_,
		_w17851_,
		_w17852_
	);
	LUT4 #(
		.INIT('hff53)
	) name13805 (
		_w8907_,
		_w11318_,
		_w17525_,
		_w17526_,
		_w17853_
	);
	LUT2 #(
		.INIT('h2)
	) name13806 (
		_w17524_,
		_w17853_,
		_w17854_
	);
	LUT3 #(
		.INIT('h54)
	) name13807 (
		_w7346_,
		_w17539_,
		_w17540_,
		_w17855_
	);
	LUT3 #(
		.INIT('h54)
	) name13808 (
		_w7349_,
		_w17542_,
		_w17543_,
		_w17856_
	);
	LUT3 #(
		.INIT('h54)
	) name13809 (
		_w7342_,
		_w17545_,
		_w17546_,
		_w17857_
	);
	LUT3 #(
		.INIT('h01)
	) name13810 (
		_w17856_,
		_w17857_,
		_w17855_,
		_w17858_
	);
	LUT2 #(
		.INIT('h8)
	) name13811 (
		_w17538_,
		_w17858_,
		_w17859_
	);
	LUT2 #(
		.INIT('h8)
	) name13812 (
		_w17525_,
		_w17859_,
		_w17860_
	);
	LUT4 #(
		.INIT('h1310)
	) name13813 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w7378_,
		_w16322_,
		_w16504_,
		_w17861_
	);
	LUT3 #(
		.INIT('h04)
	) name13814 (
		_w17524_,
		_w17526_,
		_w17861_,
		_w17862_
	);
	LUT4 #(
		.INIT('h2023)
	) name13815 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w7378_,
		_w16322_,
		_w16504_,
		_w17863_
	);
	LUT4 #(
		.INIT('h1310)
	) name13816 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8907_,
		_w16322_,
		_w16504_,
		_w17864_
	);
	LUT4 #(
		.INIT('h0008)
	) name13817 (
		_w17524_,
		_w17526_,
		_w17864_,
		_w17863_,
		_w17865_
	);
	LUT4 #(
		.INIT('h3310)
	) name13818 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7334_,
		_w17572_,
		_w17575_,
		_w17866_
	);
	LUT4 #(
		.INIT('h3230)
	) name13819 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7338_,
		_w17571_,
		_w17572_,
		_w17867_
	);
	LUT4 #(
		.INIT('h008f)
	) name13820 (
		_w12740_,
		_w14386_,
		_w17569_,
		_w17867_,
		_w17868_
	);
	LUT2 #(
		.INIT('h4)
	) name13821 (
		_w17866_,
		_w17868_,
		_w17869_
	);
	LUT3 #(
		.INIT('h80)
	) name13822 (
		_w8907_,
		_w17563_,
		_w17564_,
		_w17870_
	);
	LUT3 #(
		.INIT('h54)
	) name13823 (
		_w7365_,
		_w17558_,
		_w17559_,
		_w17871_
	);
	LUT3 #(
		.INIT('h80)
	) name13824 (
		_w7378_,
		_w17563_,
		_w17566_,
		_w17872_
	);
	LUT3 #(
		.INIT('h01)
	) name13825 (
		_w17871_,
		_w17872_,
		_w17870_,
		_w17873_
	);
	LUT3 #(
		.INIT('hb0)
	) name13826 (
		_w12668_,
		_w17556_,
		_w17873_,
		_w17874_
	);
	LUT2 #(
		.INIT('h8)
	) name13827 (
		_w17869_,
		_w17874_,
		_w17875_
	);
	LUT4 #(
		.INIT('h4500)
	) name13828 (
		_w17865_,
		_w17860_,
		_w17862_,
		_w17875_,
		_w17876_
	);
	LUT2 #(
		.INIT('h4)
	) name13829 (
		_w17854_,
		_w17876_,
		_w17877_
	);
	LUT2 #(
		.INIT('h2)
	) name13830 (
		_w7351_,
		_w17588_,
		_w17878_
	);
	LUT2 #(
		.INIT('h8)
	) name13831 (
		_w7344_,
		_w17588_,
		_w17879_
	);
	LUT3 #(
		.INIT('h01)
	) name13832 (
		_w17585_,
		_w17879_,
		_w17878_,
		_w17880_
	);
	LUT2 #(
		.INIT('h1)
	) name13833 (
		_w17587_,
		_w17880_,
		_w17881_
	);
	LUT4 #(
		.INIT('hef00)
	) name13834 (
		_w12626_,
		_w12627_,
		_w17585_,
		_w17881_,
		_w17882_
	);
	LUT3 #(
		.INIT('h01)
	) name13835 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w11926_,
		_w17586_,
		_w17883_
	);
	LUT2 #(
		.INIT('h1)
	) name13836 (
		_w17515_,
		_w17883_,
		_w17884_
	);
	LUT2 #(
		.INIT('h4)
	) name13837 (
		_w17882_,
		_w17884_,
		_w17885_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13838 (
		_w17515_,
		_w17852_,
		_w17877_,
		_w17885_,
		_w17886_
	);
	LUT4 #(
		.INIT('h1050)
	) name13839 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9847_,
		_w12118_,
		_w17887_
	);
	LUT3 #(
		.INIT('h02)
	) name13840 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w12006_,
		_w12007_,
		_w17888_
	);
	LUT4 #(
		.INIT('h007f)
	) name13841 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w17888_,
		_w17889_
	);
	LUT3 #(
		.INIT('h8a)
	) name13842 (
		_w17517_,
		_w17887_,
		_w17889_,
		_w17890_
	);
	LUT4 #(
		.INIT('hacc0)
	) name13843 (
		_w6897_,
		_w8841_,
		_w17525_,
		_w17526_,
		_w17891_
	);
	LUT3 #(
		.INIT('ha8)
	) name13844 (
		_w17524_,
		_w17527_,
		_w17891_,
		_w17892_
	);
	LUT3 #(
		.INIT('h54)
	) name13845 (
		_w6867_,
		_w17542_,
		_w17543_,
		_w17893_
	);
	LUT3 #(
		.INIT('h54)
	) name13846 (
		_w6864_,
		_w17545_,
		_w17546_,
		_w17894_
	);
	LUT3 #(
		.INIT('h54)
	) name13847 (
		_w6860_,
		_w17539_,
		_w17540_,
		_w17895_
	);
	LUT3 #(
		.INIT('h01)
	) name13848 (
		_w17894_,
		_w17895_,
		_w17893_,
		_w17896_
	);
	LUT2 #(
		.INIT('h8)
	) name13849 (
		_w17538_,
		_w17896_,
		_w17897_
	);
	LUT2 #(
		.INIT('h8)
	) name13850 (
		_w17525_,
		_w17897_,
		_w17898_
	);
	LUT4 #(
		.INIT('h1310)
	) name13851 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w6897_,
		_w16322_,
		_w16504_,
		_w17899_
	);
	LUT3 #(
		.INIT('h04)
	) name13852 (
		_w17524_,
		_w17526_,
		_w17899_,
		_w17900_
	);
	LUT2 #(
		.INIT('h4)
	) name13853 (
		_w13200_,
		_w17556_,
		_w17901_
	);
	LUT3 #(
		.INIT('h54)
	) name13854 (
		_w6848_,
		_w17558_,
		_w17559_,
		_w17902_
	);
	LUT3 #(
		.INIT('h80)
	) name13855 (
		_w8841_,
		_w17563_,
		_w17564_,
		_w17903_
	);
	LUT2 #(
		.INIT('h1)
	) name13856 (
		_w17902_,
		_w17903_,
		_w17904_
	);
	LUT3 #(
		.INIT('h80)
	) name13857 (
		_w6897_,
		_w17563_,
		_w17566_,
		_w17905_
	);
	LUT3 #(
		.INIT('h0b)
	) name13858 (
		_w12027_,
		_w17569_,
		_w17905_,
		_w17906_
	);
	LUT4 #(
		.INIT('h3230)
	) name13859 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6882_,
		_w17571_,
		_w17572_,
		_w17907_
	);
	LUT4 #(
		.INIT('h3310)
	) name13860 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6886_,
		_w17572_,
		_w17575_,
		_w17908_
	);
	LUT2 #(
		.INIT('h1)
	) name13861 (
		_w17907_,
		_w17908_,
		_w17909_
	);
	LUT3 #(
		.INIT('h80)
	) name13862 (
		_w17904_,
		_w17906_,
		_w17909_,
		_w17910_
	);
	LUT2 #(
		.INIT('h4)
	) name13863 (
		_w17901_,
		_w17910_,
		_w17911_
	);
	LUT3 #(
		.INIT('hb0)
	) name13864 (
		_w17898_,
		_w17900_,
		_w17911_,
		_w17912_
	);
	LUT2 #(
		.INIT('h4)
	) name13865 (
		_w17892_,
		_w17912_,
		_w17913_
	);
	LUT2 #(
		.INIT('h2)
	) name13866 (
		_w6871_,
		_w17588_,
		_w17914_
	);
	LUT2 #(
		.INIT('h8)
	) name13867 (
		_w6862_,
		_w17588_,
		_w17915_
	);
	LUT3 #(
		.INIT('h01)
	) name13868 (
		_w17585_,
		_w17915_,
		_w17914_,
		_w17916_
	);
	LUT2 #(
		.INIT('h1)
	) name13869 (
		_w17587_,
		_w17916_,
		_w17917_
	);
	LUT4 #(
		.INIT('hef00)
	) name13870 (
		_w12006_,
		_w12007_,
		_w17585_,
		_w17917_,
		_w17918_
	);
	LUT3 #(
		.INIT('h01)
	) name13871 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w11926_,
		_w17586_,
		_w17919_
	);
	LUT2 #(
		.INIT('h1)
	) name13872 (
		_w17515_,
		_w17919_,
		_w17920_
	);
	LUT2 #(
		.INIT('h4)
	) name13873 (
		_w17918_,
		_w17920_,
		_w17921_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13874 (
		_w17515_,
		_w17890_,
		_w17913_,
		_w17921_,
		_w17922_
	);
	LUT3 #(
		.INIT('h80)
	) name13875 (
		\sport0_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		_w12312_,
		_w17923_
	);
	LUT3 #(
		.INIT('h48)
	) name13876 (
		\sport0_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		_w12109_,
		_w17923_,
		_w17924_
	);
	LUT4 #(
		.INIT('h70f8)
	) name13877 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w12120_,
		_w12163_,
		_w17925_
	);
	LUT4 #(
		.INIT('h80d0)
	) name13878 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w11318_,
		_w17517_,
		_w17925_,
		_w17926_
	);
	LUT4 #(
		.INIT('hff53)
	) name13879 (
		_w8974_,
		_w11318_,
		_w17525_,
		_w17526_,
		_w17927_
	);
	LUT2 #(
		.INIT('h2)
	) name13880 (
		_w17524_,
		_w17927_,
		_w17928_
	);
	LUT3 #(
		.INIT('h54)
	) name13881 (
		_w8371_,
		_w17542_,
		_w17543_,
		_w17929_
	);
	LUT2 #(
		.INIT('h1)
	) name13882 (
		_w17536_,
		_w17929_,
		_w17930_
	);
	LUT3 #(
		.INIT('h54)
	) name13883 (
		_w8375_,
		_w17545_,
		_w17546_,
		_w17931_
	);
	LUT3 #(
		.INIT('h80)
	) name13884 (
		_w5713_,
		_w17532_,
		_w17530_,
		_w17932_
	);
	LUT3 #(
		.INIT('h54)
	) name13885 (
		_w5713_,
		_w17539_,
		_w17540_,
		_w17933_
	);
	LUT3 #(
		.INIT('h01)
	) name13886 (
		_w17932_,
		_w17933_,
		_w17931_,
		_w17934_
	);
	LUT2 #(
		.INIT('h8)
	) name13887 (
		_w17930_,
		_w17934_,
		_w17935_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name13888 (
		_w7906_,
		_w17525_,
		_w17526_,
		_w17935_,
		_w17936_
	);
	LUT4 #(
		.INIT('h2023)
	) name13889 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8802_,
		_w16322_,
		_w16504_,
		_w17937_
	);
	LUT4 #(
		.INIT('h1310)
	) name13890 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8821_,
		_w16322_,
		_w16504_,
		_w17938_
	);
	LUT4 #(
		.INIT('h0008)
	) name13891 (
		_w17524_,
		_w17526_,
		_w17938_,
		_w17937_,
		_w17939_
	);
	LUT3 #(
		.INIT('h80)
	) name13892 (
		_w8802_,
		_w17563_,
		_w17566_,
		_w17940_
	);
	LUT3 #(
		.INIT('h80)
	) name13893 (
		_w8821_,
		_w17563_,
		_w17564_,
		_w17941_
	);
	LUT3 #(
		.INIT('h54)
	) name13894 (
		_w8349_,
		_w17558_,
		_w17559_,
		_w17942_
	);
	LUT3 #(
		.INIT('h01)
	) name13895 (
		_w17941_,
		_w17942_,
		_w17940_,
		_w17943_
	);
	LUT4 #(
		.INIT('h3230)
	) name13896 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w8363_,
		_w17571_,
		_w17572_,
		_w17944_
	);
	LUT4 #(
		.INIT('h3310)
	) name13897 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w8365_,
		_w17572_,
		_w17575_,
		_w17945_
	);
	LUT2 #(
		.INIT('h1)
	) name13898 (
		_w17944_,
		_w17945_,
		_w17946_
	);
	LUT2 #(
		.INIT('h8)
	) name13899 (
		_w17943_,
		_w17946_,
		_w17947_
	);
	LUT4 #(
		.INIT('h54fc)
	) name13900 (
		_w11587_,
		_w11530_,
		_w11489_,
		_w11469_,
		_w17948_
	);
	LUT4 #(
		.INIT('hcf45)
	) name13901 (
		_w11496_,
		_w11510_,
		_w11522_,
		_w11953_,
		_w17949_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name13902 (
		_w11409_,
		_w11514_,
		_w11458_,
		_w11973_,
		_w17950_
	);
	LUT4 #(
		.INIT('h153f)
	) name13903 (
		_w11558_,
		_w11435_,
		_w11465_,
		_w11872_,
		_w17951_
	);
	LUT4 #(
		.INIT('h8000)
	) name13904 (
		_w17950_,
		_w17951_,
		_w17948_,
		_w17949_,
		_w17952_
	);
	LUT2 #(
		.INIT('h8)
	) name13905 (
		_w11900_,
		_w17952_,
		_w17953_
	);
	LUT4 #(
		.INIT('h4000)
	) name13906 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11386_,
		_w11358_,
		_w11476_,
		_w17954_
	);
	LUT4 #(
		.INIT('h00b1)
	) name13907 (
		_w11386_,
		_w11396_,
		_w11593_,
		_w17954_,
		_w17955_
	);
	LUT3 #(
		.INIT('hc4)
	) name13908 (
		_w11341_,
		_w11408_,
		_w17955_,
		_w17956_
	);
	LUT3 #(
		.INIT('hc8)
	) name13909 (
		_w11588_,
		_w11449_,
		_w12496_,
		_w17957_
	);
	LUT3 #(
		.INIT('hc8)
	) name13910 (
		_w11555_,
		_w11507_,
		_w11888_,
		_w17958_
	);
	LUT3 #(
		.INIT('h07)
	) name13911 (
		_w11341_,
		_w11397_,
		_w11885_,
		_w17959_
	);
	LUT3 #(
		.INIT('h04)
	) name13912 (
		_w17958_,
		_w17959_,
		_w17957_,
		_w17960_
	);
	LUT3 #(
		.INIT('h08)
	) name13913 (
		_w11386_,
		_w11415_,
		_w11510_,
		_w17961_
	);
	LUT4 #(
		.INIT('h0040)
	) name13914 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11401_,
		_w11358_,
		_w12413_,
		_w17962_
	);
	LUT4 #(
		.INIT('h1000)
	) name13915 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11542_,
		_w11358_,
		_w11491_,
		_w17963_
	);
	LUT4 #(
		.INIT('h8000)
	) name13916 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11402_,
		_w11503_,
		_w17964_
	);
	LUT4 #(
		.INIT('h0001)
	) name13917 (
		_w17961_,
		_w17962_,
		_w17963_,
		_w17964_,
		_w17965_
	);
	LUT2 #(
		.INIT('h2)
	) name13918 (
		_w11578_,
		_w12024_,
		_w17966_
	);
	LUT3 #(
		.INIT('h08)
	) name13919 (
		_w11473_,
		_w11389_,
		_w12413_,
		_w17967_
	);
	LUT3 #(
		.INIT('h80)
	) name13920 (
		_w11389_,
		_w11476_,
		_w11453_,
		_w17968_
	);
	LUT3 #(
		.INIT('h20)
	) name13921 (
		_w11389_,
		_w11542_,
		_w11392_,
		_w17969_
	);
	LUT4 #(
		.INIT('h0001)
	) name13922 (
		_w17966_,
		_w17967_,
		_w17968_,
		_w17969_,
		_w17970_
	);
	LUT4 #(
		.INIT('ha820)
	) name13923 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001 ,
		_w17971_
	);
	LUT4 #(
		.INIT('h00f7)
	) name13924 (
		_w11389_,
		_w11445_,
		_w11471_,
		_w17971_,
		_w17972_
	);
	LUT2 #(
		.INIT('h4)
	) name13925 (
		_w13293_,
		_w17972_,
		_w17973_
	);
	LUT3 #(
		.INIT('h80)
	) name13926 (
		_w17970_,
		_w17973_,
		_w17965_,
		_w17974_
	);
	LUT3 #(
		.INIT('h02)
	) name13927 (
		_w11386_,
		_w11498_,
		_w11953_,
		_w17975_
	);
	LUT2 #(
		.INIT('h2)
	) name13928 (
		_w12649_,
		_w17975_,
		_w17976_
	);
	LUT4 #(
		.INIT('h8000)
	) name13929 (
		_w17956_,
		_w17974_,
		_w17976_,
		_w17960_,
		_w17977_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name13930 (
		_w12451_,
		_w17569_,
		_w17953_,
		_w17977_,
		_w17978_
	);
	LUT3 #(
		.INIT('h0b)
	) name13931 (
		_w12435_,
		_w17556_,
		_w17978_,
		_w17979_
	);
	LUT2 #(
		.INIT('h8)
	) name13932 (
		_w17947_,
		_w17979_,
		_w17980_
	);
	LUT4 #(
		.INIT('h0e00)
	) name13933 (
		_w17524_,
		_w17936_,
		_w17939_,
		_w17980_,
		_w17981_
	);
	LUT2 #(
		.INIT('h4)
	) name13934 (
		_w17928_,
		_w17981_,
		_w17982_
	);
	LUT2 #(
		.INIT('h2)
	) name13935 (
		_w8373_,
		_w17588_,
		_w17983_
	);
	LUT2 #(
		.INIT('h8)
	) name13936 (
		_w8382_,
		_w17588_,
		_w17984_
	);
	LUT3 #(
		.INIT('h01)
	) name13937 (
		_w17585_,
		_w17984_,
		_w17983_,
		_w17985_
	);
	LUT2 #(
		.INIT('h1)
	) name13938 (
		_w17587_,
		_w17985_,
		_w17986_
	);
	LUT3 #(
		.INIT('h01)
	) name13939 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w11926_,
		_w17586_,
		_w17987_
	);
	LUT2 #(
		.INIT('h1)
	) name13940 (
		_w17515_,
		_w17987_,
		_w17988_
	);
	LUT4 #(
		.INIT('h8f00)
	) name13941 (
		_w11318_,
		_w17585_,
		_w17986_,
		_w17988_,
		_w17989_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13942 (
		_w17515_,
		_w17926_,
		_w17982_,
		_w17989_,
		_w17990_
	);
	LUT3 #(
		.INIT('hca)
	) name13943 (
		\sport0_txctl_TXSHT_reg[11]/P0001 ,
		\sport0_txctl_TX_reg[12]/P0001 ,
		_w12552_,
		_w17991_
	);
	LUT4 #(
		.INIT('h4500)
	) name13944 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w17630_,
		_w17992_
	);
	LUT3 #(
		.INIT('h02)
	) name13945 (
		_w8841_,
		_w17630_,
		_w17633_,
		_w17993_
	);
	LUT3 #(
		.INIT('he4)
	) name13946 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[1]/P0001 ,
		_w17994_
	);
	LUT3 #(
		.INIT('h40)
	) name13947 (
		_w17617_,
		_w17635_,
		_w17994_,
		_w17995_
	);
	LUT3 #(
		.INIT('h53)
	) name13948 (
		_w6869_,
		_w6873_,
		_w17618_,
		_w17996_
	);
	LUT3 #(
		.INIT('h80)
	) name13949 (
		_w17617_,
		_w17635_,
		_w17996_,
		_w17997_
	);
	LUT3 #(
		.INIT('h80)
	) name13950 (
		_w17514_,
		_w17628_,
		_w17916_,
		_w17998_
	);
	LUT3 #(
		.INIT('h01)
	) name13951 (
		_w17997_,
		_w17998_,
		_w17995_,
		_w17999_
	);
	LUT2 #(
		.INIT('h4)
	) name13952 (
		_w17993_,
		_w17999_,
		_w18000_
	);
	LUT3 #(
		.INIT('ha8)
	) name13953 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w17511_,
		_w17512_,
		_w18001_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13954 (
		_w17511_,
		_w17992_,
		_w18000_,
		_w18001_,
		_w18002_
	);
	LUT2 #(
		.INIT('h1)
	) name13955 (
		_w17627_,
		_w18002_,
		_w18003_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13956 (
		_w17627_,
		_w17890_,
		_w17913_,
		_w18003_,
		_w18004_
	);
	LUT4 #(
		.INIT('h4500)
	) name13957 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w17630_,
		_w18005_
	);
	LUT3 #(
		.INIT('h02)
	) name13958 (
		_w8907_,
		_w17630_,
		_w17633_,
		_w18006_
	);
	LUT3 #(
		.INIT('he4)
	) name13959 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[4]/P0001 ,
		_w18007_
	);
	LUT3 #(
		.INIT('h40)
	) name13960 (
		_w17617_,
		_w17635_,
		_w18007_,
		_w18008_
	);
	LUT3 #(
		.INIT('h53)
	) name13961 (
		_w7353_,
		_w7355_,
		_w17618_,
		_w18009_
	);
	LUT3 #(
		.INIT('h80)
	) name13962 (
		_w17617_,
		_w17635_,
		_w18009_,
		_w18010_
	);
	LUT3 #(
		.INIT('h80)
	) name13963 (
		_w17514_,
		_w17628_,
		_w17880_,
		_w18011_
	);
	LUT3 #(
		.INIT('h01)
	) name13964 (
		_w18010_,
		_w18011_,
		_w18008_,
		_w18012_
	);
	LUT2 #(
		.INIT('h4)
	) name13965 (
		_w18006_,
		_w18012_,
		_w18013_
	);
	LUT3 #(
		.INIT('ha8)
	) name13966 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 ,
		_w17511_,
		_w17512_,
		_w18014_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13967 (
		_w17511_,
		_w18005_,
		_w18013_,
		_w18014_,
		_w18015_
	);
	LUT2 #(
		.INIT('h1)
	) name13968 (
		_w17627_,
		_w18015_,
		_w18016_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13969 (
		_w17627_,
		_w17852_,
		_w17877_,
		_w18016_,
		_w18017_
	);
	LUT4 #(
		.INIT('h4500)
	) name13970 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w17630_,
		_w18018_
	);
	LUT3 #(
		.INIT('h02)
	) name13971 (
		_w8952_,
		_w17630_,
		_w17633_,
		_w18019_
	);
	LUT3 #(
		.INIT('he4)
	) name13972 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001 ,
		_w18020_
	);
	LUT3 #(
		.INIT('h40)
	) name13973 (
		_w17617_,
		_w17635_,
		_w18020_,
		_w18021_
	);
	LUT3 #(
		.INIT('h35)
	) name13974 (
		_w8030_,
		_w8032_,
		_w17618_,
		_w18022_
	);
	LUT3 #(
		.INIT('h80)
	) name13975 (
		_w17617_,
		_w17635_,
		_w18022_,
		_w18023_
	);
	LUT3 #(
		.INIT('h80)
	) name13976 (
		_w17514_,
		_w17628_,
		_w17780_,
		_w18024_
	);
	LUT3 #(
		.INIT('h01)
	) name13977 (
		_w18023_,
		_w18024_,
		_w18021_,
		_w18025_
	);
	LUT2 #(
		.INIT('h4)
	) name13978 (
		_w18019_,
		_w18025_,
		_w18026_
	);
	LUT3 #(
		.INIT('ha8)
	) name13979 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 ,
		_w17511_,
		_w17512_,
		_w18027_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13980 (
		_w17511_,
		_w18018_,
		_w18026_,
		_w18027_,
		_w18028_
	);
	LUT2 #(
		.INIT('h1)
	) name13981 (
		_w17627_,
		_w18028_,
		_w18029_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13982 (
		_w17627_,
		_w17752_,
		_w17777_,
		_w18029_,
		_w18030_
	);
	LUT3 #(
		.INIT('h80)
	) name13983 (
		\sport1_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		_w12733_,
		_w18031_
	);
	LUT3 #(
		.INIT('h48)
	) name13984 (
		\sport1_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		_w12087_,
		_w18031_,
		_w18032_
	);
	LUT4 #(
		.INIT('h4500)
	) name13985 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w17630_,
		_w18033_
	);
	LUT3 #(
		.INIT('h02)
	) name13986 (
		_w8929_,
		_w17630_,
		_w17633_,
		_w18034_
	);
	LUT3 #(
		.INIT('he4)
	) name13987 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001 ,
		_w18035_
	);
	LUT3 #(
		.INIT('h40)
	) name13988 (
		_w17617_,
		_w17635_,
		_w18035_,
		_w18036_
	);
	LUT3 #(
		.INIT('h53)
	) name13989 (
		_w7673_,
		_w7677_,
		_w17618_,
		_w18037_
	);
	LUT3 #(
		.INIT('h80)
	) name13990 (
		_w17617_,
		_w17635_,
		_w18037_,
		_w18038_
	);
	LUT3 #(
		.INIT('h80)
	) name13991 (
		_w17514_,
		_w17628_,
		_w17842_,
		_w18039_
	);
	LUT3 #(
		.INIT('h01)
	) name13992 (
		_w18038_,
		_w18039_,
		_w18036_,
		_w18040_
	);
	LUT2 #(
		.INIT('h4)
	) name13993 (
		_w18034_,
		_w18040_,
		_w18041_
	);
	LUT3 #(
		.INIT('ha8)
	) name13994 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w17511_,
		_w17512_,
		_w18042_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13995 (
		_w17511_,
		_w18033_,
		_w18041_,
		_w18042_,
		_w18043_
	);
	LUT2 #(
		.INIT('h1)
	) name13996 (
		_w17627_,
		_w18043_,
		_w18044_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13997 (
		_w17627_,
		_w17790_,
		_w17839_,
		_w18044_,
		_w18045_
	);
	LUT3 #(
		.INIT('h02)
	) name13998 (
		_w8821_,
		_w17630_,
		_w17633_,
		_w18046_
	);
	LUT3 #(
		.INIT('h10)
	) name13999 (
		_w8798_,
		_w8801_,
		_w17630_,
		_w18047_
	);
	LUT3 #(
		.INIT('he4)
	) name14000 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001 ,
		_w18048_
	);
	LUT3 #(
		.INIT('h40)
	) name14001 (
		_w17617_,
		_w17635_,
		_w18048_,
		_w18049_
	);
	LUT3 #(
		.INIT('h53)
	) name14002 (
		_w8378_,
		_w8380_,
		_w17618_,
		_w18050_
	);
	LUT3 #(
		.INIT('h80)
	) name14003 (
		_w17617_,
		_w17635_,
		_w18050_,
		_w18051_
	);
	LUT3 #(
		.INIT('h80)
	) name14004 (
		_w17514_,
		_w17628_,
		_w17985_,
		_w18052_
	);
	LUT3 #(
		.INIT('h01)
	) name14005 (
		_w18051_,
		_w18052_,
		_w18049_,
		_w18053_
	);
	LUT4 #(
		.INIT('h5455)
	) name14006 (
		_w17511_,
		_w18046_,
		_w18047_,
		_w18053_,
		_w18054_
	);
	LUT3 #(
		.INIT('ha8)
	) name14007 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w17511_,
		_w17512_,
		_w18055_
	);
	LUT3 #(
		.INIT('h54)
	) name14008 (
		_w17627_,
		_w18054_,
		_w18055_,
		_w18056_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14009 (
		_w17627_,
		_w17926_,
		_w17982_,
		_w18056_,
		_w18057_
	);
	LUT4 #(
		.INIT('h0060)
	) name14010 (
		_w11335_,
		_w11528_,
		_w14774_,
		_w14775_,
		_w18058_
	);
	LUT3 #(
		.INIT('h01)
	) name14011 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w14802_,
		_w18058_,
		_w18059_
	);
	LUT4 #(
		.INIT('h00fd)
	) name14012 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w12560_,
		_w12561_,
		_w18059_,
		_w18060_
	);
	LUT3 #(
		.INIT('h2e)
	) name14013 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001 ,
		_w14780_,
		_w18060_,
		_w18061_
	);
	LUT4 #(
		.INIT('h00fd)
	) name14014 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w11626_,
		_w11627_,
		_w18059_,
		_w18062_
	);
	LUT3 #(
		.INIT('h2e)
	) name14015 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001 ,
		_w14780_,
		_w18062_,
		_w18063_
	);
	LUT4 #(
		.INIT('h1b00)
	) name14016 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w11625_,
		_w18064_
	);
	LUT3 #(
		.INIT('h13)
	) name14017 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001 ,
		_w9894_,
		_w18065_
	);
	LUT4 #(
		.INIT('h0002)
	) name14018 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w18065_,
		_w18066_
	);
	LUT4 #(
		.INIT('h313b)
	) name14019 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001 ,
		_w11631_,
		_w11635_,
		_w18067_
	);
	LUT4 #(
		.INIT('h1055)
	) name14020 (
		_w11624_,
		_w18064_,
		_w18066_,
		_w18067_,
		_w18068_
	);
	LUT4 #(
		.INIT('hff02)
	) name14021 (
		_w11624_,
		_w12339_,
		_w12340_,
		_w18068_,
		_w18069_
	);
	LUT4 #(
		.INIT('h9f00)
	) name14022 (
		_w11335_,
		_w11528_,
		_w14774_,
		_w14775_,
		_w18070_
	);
	LUT4 #(
		.INIT('h3332)
	) name14023 (
		_w14802_,
		_w14803_,
		_w18058_,
		_w18070_,
		_w18071_
	);
	LUT2 #(
		.INIT('h4)
	) name14024 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w18071_,
		_w18072_
	);
	LUT4 #(
		.INIT('h0057)
	) name14025 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w12626_,
		_w12627_,
		_w18072_,
		_w18073_
	);
	LUT3 #(
		.INIT('he2)
	) name14026 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001 ,
		_w14780_,
		_w18073_,
		_w18074_
	);
	LUT4 #(
		.INIT('h00fd)
	) name14027 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w12736_,
		_w12737_,
		_w18059_,
		_w18075_
	);
	LUT3 #(
		.INIT('h2e)
	) name14028 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001 ,
		_w14780_,
		_w18075_,
		_w18076_
	);
	LUT4 #(
		.INIT('h8000)
	) name14029 (
		_w16238_,
		_w16243_,
		_w16244_,
		_w16246_,
		_w18077_
	);
	LUT3 #(
		.INIT('h51)
	) name14030 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w16247_,
		_w18077_,
		_w18078_
	);
	LUT4 #(
		.INIT('h0057)
	) name14031 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w13610_,
		_w13611_,
		_w18078_,
		_w18079_
	);
	LUT3 #(
		.INIT('he2)
	) name14032 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001 ,
		_w14780_,
		_w18079_,
		_w18080_
	);
	LUT4 #(
		.INIT('he400)
	) name14033 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w11655_,
		_w18081_
	);
	LUT2 #(
		.INIT('h2)
	) name14034 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001 ,
		_w11656_,
		_w18082_
	);
	LUT3 #(
		.INIT('h01)
	) name14035 (
		_w9946_,
		_w11659_,
		_w18082_,
		_w18083_
	);
	LUT2 #(
		.INIT('h4)
	) name14036 (
		_w18081_,
		_w18083_,
		_w18084_
	);
	LUT4 #(
		.INIT('h0057)
	) name14037 (
		_w9946_,
		_w12339_,
		_w12340_,
		_w18084_,
		_w18085_
	);
	LUT3 #(
		.INIT('h2e)
	) name14038 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001 ,
		_w14809_,
		_w18062_,
		_w18086_
	);
	LUT3 #(
		.INIT('h2e)
	) name14039 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001 ,
		_w14809_,
		_w18060_,
		_w18087_
	);
	LUT3 #(
		.INIT('h2e)
	) name14040 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001 ,
		_w14809_,
		_w18075_,
		_w18088_
	);
	LUT3 #(
		.INIT('he2)
	) name14041 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001 ,
		_w14809_,
		_w18073_,
		_w18089_
	);
	LUT3 #(
		.INIT('he2)
	) name14042 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001 ,
		_w14809_,
		_w18079_,
		_w18090_
	);
	LUT4 #(
		.INIT('h0105)
	) name14043 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9886_,
		_w12118_,
		_w18091_
	);
	LUT2 #(
		.INIT('h8)
	) name14044 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w12284_,
		_w18092_
	);
	LUT4 #(
		.INIT('h007f)
	) name14045 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18092_,
		_w18093_
	);
	LUT3 #(
		.INIT('h8a)
	) name14046 (
		_w17517_,
		_w18091_,
		_w18093_,
		_w18094_
	);
	LUT3 #(
		.INIT('h01)
	) name14047 (
		_w17534_,
		_w17537_,
		_w17933_,
		_w18095_
	);
	LUT3 #(
		.INIT('h54)
	) name14048 (
		_w7216_,
		_w17542_,
		_w17543_,
		_w18096_
	);
	LUT3 #(
		.INIT('h54)
	) name14049 (
		_w7213_,
		_w17545_,
		_w17546_,
		_w18097_
	);
	LUT2 #(
		.INIT('h1)
	) name14050 (
		_w18096_,
		_w18097_,
		_w18098_
	);
	LUT2 #(
		.INIT('h8)
	) name14051 (
		_w18095_,
		_w18098_,
		_w18099_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name14052 (
		_w7906_,
		_w17525_,
		_w17526_,
		_w18099_,
		_w18100_
	);
	LUT2 #(
		.INIT('h1)
	) name14053 (
		_w17524_,
		_w18100_,
		_w18101_
	);
	LUT4 #(
		.INIT('h1310)
	) name14054 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w9021_,
		_w16322_,
		_w16504_,
		_w18102_
	);
	LUT4 #(
		.INIT('h2023)
	) name14055 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w7241_,
		_w16322_,
		_w16504_,
		_w18103_
	);
	LUT4 #(
		.INIT('h0008)
	) name14056 (
		_w17524_,
		_w17526_,
		_w18103_,
		_w18102_,
		_w18104_
	);
	LUT3 #(
		.INIT('h80)
	) name14057 (
		_w7241_,
		_w17563_,
		_w17566_,
		_w18105_
	);
	LUT3 #(
		.INIT('h54)
	) name14058 (
		_w7228_,
		_w17558_,
		_w17559_,
		_w18106_
	);
	LUT3 #(
		.INIT('h80)
	) name14059 (
		_w9021_,
		_w17563_,
		_w17564_,
		_w18107_
	);
	LUT3 #(
		.INIT('h01)
	) name14060 (
		_w18106_,
		_w18107_,
		_w18105_,
		_w18108_
	);
	LUT4 #(
		.INIT('h3310)
	) name14061 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7203_,
		_w17572_,
		_w17575_,
		_w18109_
	);
	LUT4 #(
		.INIT('h3230)
	) name14062 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7201_,
		_w17571_,
		_w17572_,
		_w18110_
	);
	LUT2 #(
		.INIT('h1)
	) name14063 (
		_w18109_,
		_w18110_,
		_w18111_
	);
	LUT4 #(
		.INIT('h1000)
	) name14064 (
		_w11426_,
		_w11971_,
		_w12512_,
		_w12516_,
		_w18112_
	);
	LUT3 #(
		.INIT('h80)
	) name14065 (
		_w11910_,
		_w11834_,
		_w18112_,
		_w18113_
	);
	LUT2 #(
		.INIT('h4)
	) name14066 (
		_w11592_,
		_w11854_,
		_w18114_
	);
	LUT3 #(
		.INIT('he0)
	) name14067 (
		_w11552_,
		_w11474_,
		_w11874_,
		_w18115_
	);
	LUT2 #(
		.INIT('h2)
	) name14068 (
		_w11499_,
		_w11957_,
		_w18116_
	);
	LUT4 #(
		.INIT('h1113)
	) name14069 (
		_w11333_,
		_w18114_,
		_w18115_,
		_w18116_,
		_w18117_
	);
	LUT2 #(
		.INIT('h2)
	) name14070 (
		_w11385_,
		_w18117_,
		_w18118_
	);
	LUT3 #(
		.INIT('hc8)
	) name14071 (
		_w11409_,
		_w11841_,
		_w11896_,
		_w18119_
	);
	LUT3 #(
		.INIT('ha8)
	) name14072 (
		_w11537_,
		_w11547_,
		_w11976_,
		_w18120_
	);
	LUT3 #(
		.INIT('ha8)
	) name14073 (
		_w11484_,
		_w11435_,
		_w12455_,
		_w18121_
	);
	LUT3 #(
		.INIT('ha8)
	) name14074 (
		_w11507_,
		_w11973_,
		_w11974_,
		_w18122_
	);
	LUT4 #(
		.INIT('h0001)
	) name14075 (
		_w18119_,
		_w18120_,
		_w18121_,
		_w18122_,
		_w18123_
	);
	LUT3 #(
		.INIT('hc8)
	) name14076 (
		_w11552_,
		_w11459_,
		_w11474_,
		_w18124_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name14077 (
		_w11592_,
		_w11496_,
		_w11957_,
		_w12412_,
		_w18125_
	);
	LUT2 #(
		.INIT('h4)
	) name14078 (
		_w18124_,
		_w18125_,
		_w18126_
	);
	LUT4 #(
		.INIT('ha820)
	) name14079 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001 ,
		_w18127_
	);
	LUT3 #(
		.INIT('h01)
	) name14080 (
		_w11551_,
		_w11576_,
		_w18127_,
		_w18128_
	);
	LUT2 #(
		.INIT('h1)
	) name14081 (
		_w11454_,
		_w11953_,
		_w18129_
	);
	LUT3 #(
		.INIT('h0e)
	) name14082 (
		_w11393_,
		_w11589_,
		_w11471_,
		_w18130_
	);
	LUT3 #(
		.INIT('h10)
	) name14083 (
		_w18129_,
		_w18130_,
		_w18128_,
		_w18131_
	);
	LUT3 #(
		.INIT('hc8)
	) name14084 (
		_w11587_,
		_w11863_,
		_w11880_,
		_w18132_
	);
	LUT3 #(
		.INIT('he0)
	) name14085 (
		_w11420_,
		_w11421_,
		_w11860_,
		_w18133_
	);
	LUT2 #(
		.INIT('h1)
	) name14086 (
		_w18132_,
		_w18133_,
		_w18134_
	);
	LUT4 #(
		.INIT('h8000)
	) name14087 (
		_w18126_,
		_w18131_,
		_w18134_,
		_w18123_,
		_w18135_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name14088 (
		_w17569_,
		_w18113_,
		_w18118_,
		_w18135_,
		_w18136_
	);
	LUT4 #(
		.INIT('h0057)
	) name14089 (
		_w11341_,
		_w11424_,
		_w11421_,
		_w11591_,
		_w18137_
	);
	LUT2 #(
		.INIT('h4)
	) name14090 (
		_w11498_,
		_w11839_,
		_w18138_
	);
	LUT4 #(
		.INIT('h7770)
	) name14091 (
		_w11588_,
		_w11532_,
		_w11489_,
		_w11446_,
		_w18139_
	);
	LUT4 #(
		.INIT('h0800)
	) name14092 (
		_w12593_,
		_w18137_,
		_w18138_,
		_w18139_,
		_w18140_
	);
	LUT3 #(
		.INIT('ha8)
	) name14093 (
		_w11537_,
		_w11555_,
		_w12568_,
		_w18141_
	);
	LUT3 #(
		.INIT('h04)
	) name14094 (
		_w11444_,
		_w11392_,
		_w11471_,
		_w18142_
	);
	LUT3 #(
		.INIT('h04)
	) name14095 (
		_w11444_,
		_w11423_,
		_w11512_,
		_w18143_
	);
	LUT3 #(
		.INIT('h04)
	) name14096 (
		_w11444_,
		_w11428_,
		_w11454_,
		_w18144_
	);
	LUT3 #(
		.INIT('h20)
	) name14097 (
		_w11473_,
		_w11444_,
		_w11459_,
		_w18145_
	);
	LUT4 #(
		.INIT('h0001)
	) name14098 (
		_w18142_,
		_w18143_,
		_w18144_,
		_w18145_,
		_w18146_
	);
	LUT3 #(
		.INIT('ha8)
	) name14099 (
		_w11341_,
		_w11409_,
		_w11587_,
		_w18147_
	);
	LUT3 #(
		.INIT('he0)
	) name14100 (
		_w11410_,
		_w11558_,
		_w11854_,
		_w18148_
	);
	LUT4 #(
		.INIT('h0100)
	) name14101 (
		_w18141_,
		_w18147_,
		_w18148_,
		_w18146_,
		_w18149_
	);
	LUT4 #(
		.INIT('h45cf)
	) name14102 (
		_w11341_,
		_w11530_,
		_w11496_,
		_w11435_,
		_w18150_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name14103 (
		_w11534_,
		_w11515_,
		_w11522_,
		_w11860_,
		_w18151_
	);
	LUT2 #(
		.INIT('h8)
	) name14104 (
		_w18150_,
		_w18151_,
		_w18152_
	);
	LUT4 #(
		.INIT('ha820)
	) name14105 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001 ,
		_w18153_
	);
	LUT4 #(
		.INIT('h00f7)
	) name14106 (
		_w11389_,
		_w11491_,
		_w11471_,
		_w18153_,
		_w18154_
	);
	LUT2 #(
		.INIT('h2)
	) name14107 (
		_w11455_,
		_w11454_,
		_w18155_
	);
	LUT3 #(
		.INIT('h80)
	) name14108 (
		_w11401_,
		_w11389_,
		_w11459_,
		_w18156_
	);
	LUT3 #(
		.INIT('h10)
	) name14109 (
		_w18155_,
		_w18156_,
		_w18154_,
		_w18157_
	);
	LUT2 #(
		.INIT('h1)
	) name14110 (
		_w11579_,
		_w11885_,
		_w18158_
	);
	LUT4 #(
		.INIT('h7077)
	) name14111 (
		_w11529_,
		_w11500_,
		_w11512_,
		_w11462_,
		_w18159_
	);
	LUT3 #(
		.INIT('h08)
	) name14112 (
		_w11389_,
		_w11476_,
		_w12413_,
		_w18160_
	);
	LUT2 #(
		.INIT('h8)
	) name14113 (
		_w11541_,
		_w11415_,
		_w18161_
	);
	LUT3 #(
		.INIT('h10)
	) name14114 (
		_w18160_,
		_w18161_,
		_w18159_,
		_w18162_
	);
	LUT4 #(
		.INIT('h8000)
	) name14115 (
		_w11408_,
		_w18162_,
		_w18157_,
		_w18158_,
		_w18163_
	);
	LUT4 #(
		.INIT('h8000)
	) name14116 (
		_w18152_,
		_w18163_,
		_w18149_,
		_w18140_,
		_w18164_
	);
	LUT3 #(
		.INIT('h80)
	) name14117 (
		_w11902_,
		_w11905_,
		_w12629_,
		_w18165_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name14118 (
		_w11837_,
		_w17556_,
		_w18164_,
		_w18165_,
		_w18166_
	);
	LUT4 #(
		.INIT('h1000)
	) name14119 (
		_w18136_,
		_w18166_,
		_w18108_,
		_w18111_,
		_w18167_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14120 (
		_w17524_,
		_w17927_,
		_w18104_,
		_w18167_,
		_w18168_
	);
	LUT2 #(
		.INIT('h4)
	) name14121 (
		_w18101_,
		_w18168_,
		_w18169_
	);
	LUT2 #(
		.INIT('h2)
	) name14122 (
		_w9021_,
		_w17633_,
		_w18170_
	);
	LUT3 #(
		.INIT('he4)
	) name14123 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001 ,
		_w18171_
	);
	LUT3 #(
		.INIT('ha8)
	) name14124 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w17511_,
		_w17512_,
		_w18172_
	);
	LUT4 #(
		.INIT('h00bf)
	) name14125 (
		_w17617_,
		_w17635_,
		_w18171_,
		_w18172_,
		_w18173_
	);
	LUT2 #(
		.INIT('h2)
	) name14126 (
		_w7218_,
		_w17588_,
		_w18174_
	);
	LUT2 #(
		.INIT('h8)
	) name14127 (
		_w7209_,
		_w17588_,
		_w18175_
	);
	LUT3 #(
		.INIT('h01)
	) name14128 (
		_w17585_,
		_w18175_,
		_w18174_,
		_w18176_
	);
	LUT3 #(
		.INIT('h80)
	) name14129 (
		_w17514_,
		_w17628_,
		_w18176_,
		_w18177_
	);
	LUT3 #(
		.INIT('h53)
	) name14130 (
		_w7220_,
		_w7211_,
		_w17618_,
		_w18178_
	);
	LUT3 #(
		.INIT('h80)
	) name14131 (
		_w17617_,
		_w17635_,
		_w18178_,
		_w18179_
	);
	LUT4 #(
		.INIT('h0100)
	) name14132 (
		_w17630_,
		_w18177_,
		_w18179_,
		_w18173_,
		_w18180_
	);
	LUT2 #(
		.INIT('h4)
	) name14133 (
		_w18170_,
		_w18180_,
		_w18181_
	);
	LUT2 #(
		.INIT('h4)
	) name14134 (
		_w17511_,
		_w17630_,
		_w18182_
	);
	LUT2 #(
		.INIT('h4)
	) name14135 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w17511_,
		_w18183_
	);
	LUT3 #(
		.INIT('h07)
	) name14136 (
		_w17515_,
		_w17626_,
		_w18183_,
		_w18184_
	);
	LUT4 #(
		.INIT('h1f00)
	) name14137 (
		_w7140_,
		_w7240_,
		_w18182_,
		_w18184_,
		_w18185_
	);
	LUT2 #(
		.INIT('h4)
	) name14138 (
		_w18181_,
		_w18185_,
		_w18186_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14139 (
		_w17627_,
		_w18094_,
		_w18169_,
		_w18186_,
		_w18187_
	);
	LUT4 #(
		.INIT('h0105)
	) name14140 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9834_,
		_w12118_,
		_w18188_
	);
	LUT4 #(
		.INIT('ha820)
	) name14141 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w18189_
	);
	LUT4 #(
		.INIT('h007f)
	) name14142 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18189_,
		_w18190_
	);
	LUT3 #(
		.INIT('h8a)
	) name14143 (
		_w17517_,
		_w18188_,
		_w18190_,
		_w18191_
	);
	LUT3 #(
		.INIT('h54)
	) name14144 (
		_w5717_,
		_w17542_,
		_w17543_,
		_w18192_
	);
	LUT3 #(
		.INIT('h54)
	) name14145 (
		_w5720_,
		_w17545_,
		_w17546_,
		_w18193_
	);
	LUT2 #(
		.INIT('h1)
	) name14146 (
		_w18192_,
		_w18193_,
		_w18194_
	);
	LUT2 #(
		.INIT('h8)
	) name14147 (
		_w18095_,
		_w18194_,
		_w18195_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name14148 (
		_w7906_,
		_w17525_,
		_w17526_,
		_w18195_,
		_w18196_
	);
	LUT2 #(
		.INIT('h1)
	) name14149 (
		_w17524_,
		_w18196_,
		_w18197_
	);
	LUT4 #(
		.INIT('h2023)
	) name14150 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w5760_,
		_w16322_,
		_w16504_,
		_w18198_
	);
	LUT4 #(
		.INIT('h1310)
	) name14151 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8740_,
		_w16322_,
		_w16504_,
		_w18199_
	);
	LUT4 #(
		.INIT('h0008)
	) name14152 (
		_w17524_,
		_w17526_,
		_w18199_,
		_w18198_,
		_w18200_
	);
	LUT2 #(
		.INIT('h4)
	) name14153 (
		_w12481_,
		_w17569_,
		_w18201_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14154 (
		_w11433_,
		_w11546_,
		_w11597_,
		_w17556_,
		_w18202_
	);
	LUT3 #(
		.INIT('h80)
	) name14155 (
		_w5760_,
		_w17563_,
		_w17566_,
		_w18203_
	);
	LUT3 #(
		.INIT('h80)
	) name14156 (
		_w8740_,
		_w17563_,
		_w17564_,
		_w18204_
	);
	LUT3 #(
		.INIT('h54)
	) name14157 (
		_w5734_,
		_w17558_,
		_w17559_,
		_w18205_
	);
	LUT3 #(
		.INIT('h01)
	) name14158 (
		_w18204_,
		_w18205_,
		_w18203_,
		_w18206_
	);
	LUT4 #(
		.INIT('h3310)
	) name14159 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w5747_,
		_w17572_,
		_w17575_,
		_w18207_
	);
	LUT4 #(
		.INIT('h3230)
	) name14160 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w5749_,
		_w17571_,
		_w17572_,
		_w18208_
	);
	LUT2 #(
		.INIT('h1)
	) name14161 (
		_w18207_,
		_w18208_,
		_w18209_
	);
	LUT3 #(
		.INIT('h40)
	) name14162 (
		_w18202_,
		_w18206_,
		_w18209_,
		_w18210_
	);
	LUT2 #(
		.INIT('h4)
	) name14163 (
		_w18201_,
		_w18210_,
		_w18211_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14164 (
		_w17524_,
		_w17927_,
		_w18200_,
		_w18211_,
		_w18212_
	);
	LUT2 #(
		.INIT('h4)
	) name14165 (
		_w18197_,
		_w18212_,
		_w18213_
	);
	LUT2 #(
		.INIT('h8)
	) name14166 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w17512_,
		_w18214_
	);
	LUT2 #(
		.INIT('h2)
	) name14167 (
		_w5722_,
		_w17588_,
		_w18215_
	);
	LUT2 #(
		.INIT('h8)
	) name14168 (
		_w5726_,
		_w17588_,
		_w18216_
	);
	LUT3 #(
		.INIT('h01)
	) name14169 (
		_w17585_,
		_w18216_,
		_w18215_,
		_w18217_
	);
	LUT4 #(
		.INIT('h070f)
	) name14170 (
		_w17514_,
		_w17628_,
		_w18214_,
		_w18217_,
		_w18218_
	);
	LUT3 #(
		.INIT('h35)
	) name14171 (
		_w5724_,
		_w5715_,
		_w17618_,
		_w18219_
	);
	LUT3 #(
		.INIT('he4)
	) name14172 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[13]/P0001 ,
		_w18220_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14173 (
		_w17617_,
		_w17635_,
		_w18219_,
		_w18220_,
		_w18221_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name14174 (
		_w17630_,
		_w17632_,
		_w18218_,
		_w18221_,
		_w18222_
	);
	LUT4 #(
		.INIT('h3331)
	) name14175 (
		_w8740_,
		_w17511_,
		_w17630_,
		_w17633_,
		_w18223_
	);
	LUT4 #(
		.INIT('h0700)
	) name14176 (
		_w5760_,
		_w17630_,
		_w18222_,
		_w18223_,
		_w18224_
	);
	LUT2 #(
		.INIT('h4)
	) name14177 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w17511_,
		_w18225_
	);
	LUT3 #(
		.INIT('h07)
	) name14178 (
		_w17515_,
		_w17626_,
		_w18225_,
		_w18226_
	);
	LUT2 #(
		.INIT('h4)
	) name14179 (
		_w18224_,
		_w18226_,
		_w18227_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14180 (
		_w17627_,
		_w18191_,
		_w18213_,
		_w18227_,
		_w18228_
	);
	LUT4 #(
		.INIT('h0105)
	) name14181 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9768_,
		_w12118_,
		_w18229_
	);
	LUT2 #(
		.INIT('h8)
	) name14182 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w14866_,
		_w18230_
	);
	LUT4 #(
		.INIT('h007f)
	) name14183 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18230_,
		_w18231_
	);
	LUT3 #(
		.INIT('h8a)
	) name14184 (
		_w17517_,
		_w18229_,
		_w18231_,
		_w18232_
	);
	LUT3 #(
		.INIT('h54)
	) name14185 (
		_w6335_,
		_w17545_,
		_w17546_,
		_w18233_
	);
	LUT3 #(
		.INIT('h54)
	) name14186 (
		_w6331_,
		_w17542_,
		_w17543_,
		_w18234_
	);
	LUT2 #(
		.INIT('h1)
	) name14187 (
		_w18233_,
		_w18234_,
		_w18235_
	);
	LUT2 #(
		.INIT('h8)
	) name14188 (
		_w18095_,
		_w18235_,
		_w18236_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name14189 (
		_w7906_,
		_w17525_,
		_w17526_,
		_w18236_,
		_w18237_
	);
	LUT2 #(
		.INIT('h1)
	) name14190 (
		_w17524_,
		_w18237_,
		_w18238_
	);
	LUT4 #(
		.INIT('h2023)
	) name14191 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w6363_,
		_w16322_,
		_w16504_,
		_w18239_
	);
	LUT4 #(
		.INIT('h1310)
	) name14192 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8694_,
		_w16322_,
		_w16504_,
		_w18240_
	);
	LUT4 #(
		.INIT('h0008)
	) name14193 (
		_w17524_,
		_w17526_,
		_w18240_,
		_w18239_,
		_w18241_
	);
	LUT3 #(
		.INIT('h54)
	) name14194 (
		_w6349_,
		_w17558_,
		_w17559_,
		_w18242_
	);
	LUT3 #(
		.INIT('h80)
	) name14195 (
		_w8694_,
		_w17563_,
		_w17564_,
		_w18243_
	);
	LUT3 #(
		.INIT('h80)
	) name14196 (
		_w6363_,
		_w17563_,
		_w17566_,
		_w18244_
	);
	LUT3 #(
		.INIT('h01)
	) name14197 (
		_w18243_,
		_w18244_,
		_w18242_,
		_w18245_
	);
	LUT4 #(
		.INIT('h3310)
	) name14198 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6325_,
		_w17572_,
		_w17575_,
		_w18246_
	);
	LUT4 #(
		.INIT('h3230)
	) name14199 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6323_,
		_w17571_,
		_w17572_,
		_w18247_
	);
	LUT2 #(
		.INIT('h1)
	) name14200 (
		_w18246_,
		_w18247_,
		_w18248_
	);
	LUT2 #(
		.INIT('h8)
	) name14201 (
		_w18245_,
		_w18248_,
		_w18249_
	);
	LUT4 #(
		.INIT('h4000)
	) name14202 (
		_w11426_,
		_w11577_,
		_w11910_,
		_w11834_,
		_w18250_
	);
	LUT3 #(
		.INIT('h32)
	) name14203 (
		_w11552_,
		_w11501_,
		_w11474_,
		_w18251_
	);
	LUT2 #(
		.INIT('h1)
	) name14204 (
		_w11542_,
		_w11957_,
		_w18252_
	);
	LUT3 #(
		.INIT('h0e)
	) name14205 (
		_w11393_,
		_w11589_,
		_w12024_,
		_w18253_
	);
	LUT3 #(
		.INIT('h01)
	) name14206 (
		_w18252_,
		_w18253_,
		_w18251_,
		_w18254_
	);
	LUT4 #(
		.INIT('ha820)
	) name14207 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001 ,
		_w18255_
	);
	LUT3 #(
		.INIT('h0e)
	) name14208 (
		_w11471_,
		_w11953_,
		_w18255_,
		_w18256_
	);
	LUT2 #(
		.INIT('h8)
	) name14209 (
		_w12517_,
		_w18256_,
		_w18257_
	);
	LUT2 #(
		.INIT('h4)
	) name14210 (
		_w11595_,
		_w12512_,
		_w18258_
	);
	LUT3 #(
		.INIT('h80)
	) name14211 (
		_w18254_,
		_w18257_,
		_w18258_,
		_w18259_
	);
	LUT3 #(
		.INIT('hc8)
	) name14212 (
		_w11588_,
		_w11484_,
		_w12496_,
		_w18260_
	);
	LUT3 #(
		.INIT('ha8)
	) name14213 (
		_w11449_,
		_w11973_,
		_w11974_,
		_w18261_
	);
	LUT3 #(
		.INIT('hc8)
	) name14214 (
		_w11587_,
		_w11841_,
		_w11880_,
		_w18262_
	);
	LUT3 #(
		.INIT('he0)
	) name14215 (
		_w11420_,
		_w11421_,
		_w11854_,
		_w18263_
	);
	LUT4 #(
		.INIT('h0001)
	) name14216 (
		_w18260_,
		_w18261_,
		_w18262_,
		_w18263_,
		_w18264_
	);
	LUT3 #(
		.INIT('hc8)
	) name14217 (
		_w11409_,
		_w11872_,
		_w11896_,
		_w18265_
	);
	LUT3 #(
		.INIT('h32)
	) name14218 (
		_w11558_,
		_w11487_,
		_w11894_,
		_w18266_
	);
	LUT3 #(
		.INIT('hc8)
	) name14219 (
		_w11547_,
		_w11532_,
		_w11976_,
		_w18267_
	);
	LUT3 #(
		.INIT('ha8)
	) name14220 (
		_w11507_,
		_w11435_,
		_w12455_,
		_w18268_
	);
	LUT4 #(
		.INIT('h0001)
	) name14221 (
		_w18265_,
		_w18266_,
		_w18267_,
		_w18268_,
		_w18269_
	);
	LUT2 #(
		.INIT('h8)
	) name14222 (
		_w18264_,
		_w18269_,
		_w18270_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name14223 (
		_w17569_,
		_w18250_,
		_w18259_,
		_w18270_,
		_w18271_
	);
	LUT2 #(
		.INIT('h8)
	) name14224 (
		_w11910_,
		_w12409_,
		_w18272_
	);
	LUT3 #(
		.INIT('h80)
	) name14225 (
		_w11389_,
		_w11341_,
		_w11476_,
		_w18273_
	);
	LUT4 #(
		.INIT('h0010)
	) name14226 (
		_w11586_,
		_w11590_,
		_w12593_,
		_w18273_,
		_w18274_
	);
	LUT3 #(
		.INIT('h40)
	) name14227 (
		_w11444_,
		_w11423_,
		_w11449_,
		_w18275_
	);
	LUT3 #(
		.INIT('h40)
	) name14228 (
		_w11444_,
		_w11445_,
		_w11507_,
		_w18276_
	);
	LUT3 #(
		.INIT('h40)
	) name14229 (
		_w11444_,
		_w11392_,
		_w11458_,
		_w18277_
	);
	LUT3 #(
		.INIT('h20)
	) name14230 (
		_w11473_,
		_w11444_,
		_w11495_,
		_w18278_
	);
	LUT4 #(
		.INIT('h0001)
	) name14231 (
		_w18275_,
		_w18276_,
		_w18277_,
		_w18278_,
		_w18279_
	);
	LUT2 #(
		.INIT('h1)
	) name14232 (
		_w11386_,
		_w18279_,
		_w18280_
	);
	LUT2 #(
		.INIT('h4)
	) name14233 (
		_w11492_,
		_w11515_,
		_w18281_
	);
	LUT4 #(
		.INIT('hee0e)
	) name14234 (
		_w11542_,
		_w11530_,
		_w11522_,
		_w11528_,
		_w18282_
	);
	LUT3 #(
		.INIT('h20)
	) name14235 (
		_w11412_,
		_w18281_,
		_w18282_,
		_w18283_
	);
	LUT3 #(
		.INIT('h40)
	) name14236 (
		_w18280_,
		_w18274_,
		_w18283_,
		_w18284_
	);
	LUT3 #(
		.INIT('hc8)
	) name14237 (
		_w11555_,
		_w11532_,
		_w12568_,
		_w18285_
	);
	LUT3 #(
		.INIT('ha8)
	) name14238 (
		_w11341_,
		_w11557_,
		_w11558_,
		_w18286_
	);
	LUT3 #(
		.INIT('h02)
	) name14239 (
		_w11554_,
		_w18286_,
		_w18285_,
		_w18287_
	);
	LUT2 #(
		.INIT('h4)
	) name14240 (
		_w11454_,
		_w11462_,
		_w18288_
	);
	LUT3 #(
		.INIT('h80)
	) name14241 (
		_w11389_,
		_w11503_,
		_w11488_,
		_w18289_
	);
	LUT2 #(
		.INIT('h8)
	) name14242 (
		_w11455_,
		_w11470_,
		_w18290_
	);
	LUT3 #(
		.INIT('h80)
	) name14243 (
		_w11389_,
		_w11491_,
		_w11459_,
		_w18291_
	);
	LUT4 #(
		.INIT('h0001)
	) name14244 (
		_w18288_,
		_w18289_,
		_w18290_,
		_w18291_,
		_w18292_
	);
	LUT4 #(
		.INIT('ha820)
	) name14245 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001 ,
		_w18293_
	);
	LUT3 #(
		.INIT('h07)
	) name14246 (
		_w11406_,
		_w11429_,
		_w18293_,
		_w18294_
	);
	LUT3 #(
		.INIT('h08)
	) name14247 (
		_w11401_,
		_w11389_,
		_w11501_,
		_w18295_
	);
	LUT3 #(
		.INIT('h08)
	) name14248 (
		_w11389_,
		_w11434_,
		_w11512_,
		_w18296_
	);
	LUT3 #(
		.INIT('h10)
	) name14249 (
		_w18295_,
		_w18296_,
		_w18294_,
		_w18297_
	);
	LUT4 #(
		.INIT('hf400)
	) name14250 (
		_w11444_,
		_w11428_,
		_w11455_,
		_w11466_,
		_w18298_
	);
	LUT3 #(
		.INIT('h0d)
	) name14251 (
		_w11485_,
		_w11504_,
		_w18298_,
		_w18299_
	);
	LUT3 #(
		.INIT('h80)
	) name14252 (
		_w18292_,
		_w18297_,
		_w18299_,
		_w18300_
	);
	LUT3 #(
		.INIT('h40)
	) name14253 (
		_w11444_,
		_w11423_,
		_w11453_,
		_w18301_
	);
	LUT3 #(
		.INIT('h08)
	) name14254 (
		_w11386_,
		_w11415_,
		_w11528_,
		_w18302_
	);
	LUT3 #(
		.INIT('h20)
	) name14255 (
		_w11473_,
		_w11444_,
		_w11500_,
		_w18303_
	);
	LUT3 #(
		.INIT('h01)
	) name14256 (
		_w18302_,
		_w18303_,
		_w18301_,
		_w18304_
	);
	LUT3 #(
		.INIT('h40)
	) name14257 (
		_w11444_,
		_w11428_,
		_w11470_,
		_w18305_
	);
	LUT3 #(
		.INIT('h40)
	) name14258 (
		_w11444_,
		_w11445_,
		_w11511_,
		_w18306_
	);
	LUT3 #(
		.INIT('h40)
	) name14259 (
		_w11444_,
		_w11476_,
		_w11488_,
		_w18307_
	);
	LUT4 #(
		.INIT('h0001)
	) name14260 (
		_w11591_,
		_w18305_,
		_w18306_,
		_w18307_,
		_w18308_
	);
	LUT2 #(
		.INIT('h8)
	) name14261 (
		_w18304_,
		_w18308_,
		_w18309_
	);
	LUT4 #(
		.INIT('h8000)
	) name14262 (
		_w12592_,
		_w18300_,
		_w18309_,
		_w18287_,
		_w18310_
	);
	LUT4 #(
		.INIT('h8000)
	) name14263 (
		_w11836_,
		_w18272_,
		_w18310_,
		_w18284_,
		_w18311_
	);
	LUT3 #(
		.INIT('h31)
	) name14264 (
		_w17556_,
		_w18271_,
		_w18311_,
		_w18312_
	);
	LUT2 #(
		.INIT('h8)
	) name14265 (
		_w18249_,
		_w18312_,
		_w18313_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14266 (
		_w17524_,
		_w17927_,
		_w18241_,
		_w18313_,
		_w18314_
	);
	LUT2 #(
		.INIT('h4)
	) name14267 (
		_w18238_,
		_w18314_,
		_w18315_
	);
	LUT3 #(
		.INIT('h10)
	) name14268 (
		_w6263_,
		_w6362_,
		_w17630_,
		_w18316_
	);
	LUT2 #(
		.INIT('h8)
	) name14269 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		_w17512_,
		_w18317_
	);
	LUT2 #(
		.INIT('h2)
	) name14270 (
		_w6333_,
		_w17588_,
		_w18318_
	);
	LUT2 #(
		.INIT('h8)
	) name14271 (
		_w6342_,
		_w17588_,
		_w18319_
	);
	LUT3 #(
		.INIT('h01)
	) name14272 (
		_w17585_,
		_w18319_,
		_w18318_,
		_w18320_
	);
	LUT4 #(
		.INIT('h070f)
	) name14273 (
		_w17514_,
		_w17628_,
		_w18317_,
		_w18320_,
		_w18321_
	);
	LUT3 #(
		.INIT('h53)
	) name14274 (
		_w6338_,
		_w6340_,
		_w17618_,
		_w18322_
	);
	LUT3 #(
		.INIT('he4)
	) name14275 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[11]/P0001 ,
		_w18323_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14276 (
		_w17617_,
		_w17635_,
		_w18322_,
		_w18323_,
		_w18324_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name14277 (
		_w17630_,
		_w17632_,
		_w18321_,
		_w18324_,
		_w18325_
	);
	LUT4 #(
		.INIT('h3331)
	) name14278 (
		_w8694_,
		_w17511_,
		_w17630_,
		_w17633_,
		_w18326_
	);
	LUT2 #(
		.INIT('h4)
	) name14279 (
		_w18325_,
		_w18326_,
		_w18327_
	);
	LUT2 #(
		.INIT('h4)
	) name14280 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		_w17511_,
		_w18328_
	);
	LUT3 #(
		.INIT('h07)
	) name14281 (
		_w17515_,
		_w17626_,
		_w18328_,
		_w18329_
	);
	LUT3 #(
		.INIT('hb0)
	) name14282 (
		_w18316_,
		_w18327_,
		_w18329_,
		_w18330_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14283 (
		_w17627_,
		_w18232_,
		_w18315_,
		_w18330_,
		_w18331_
	);
	LUT4 #(
		.INIT('h0015)
	) name14284 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w12611_,
		_w18332_
	);
	LUT2 #(
		.INIT('h8)
	) name14285 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w12486_,
		_w18333_
	);
	LUT4 #(
		.INIT('h007f)
	) name14286 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18333_,
		_w18334_
	);
	LUT3 #(
		.INIT('h8a)
	) name14287 (
		_w17517_,
		_w18332_,
		_w18334_,
		_w18335_
	);
	LUT3 #(
		.INIT('h54)
	) name14288 (
		_w6011_,
		_w17545_,
		_w17546_,
		_w18336_
	);
	LUT3 #(
		.INIT('h54)
	) name14289 (
		_w6014_,
		_w17542_,
		_w17543_,
		_w18337_
	);
	LUT2 #(
		.INIT('h1)
	) name14290 (
		_w18336_,
		_w18337_,
		_w18338_
	);
	LUT2 #(
		.INIT('h8)
	) name14291 (
		_w18095_,
		_w18338_,
		_w18339_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name14292 (
		_w7906_,
		_w17525_,
		_w17526_,
		_w18339_,
		_w18340_
	);
	LUT2 #(
		.INIT('h1)
	) name14293 (
		_w17524_,
		_w18340_,
		_w18341_
	);
	LUT4 #(
		.INIT('h2023)
	) name14294 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w6039_,
		_w16322_,
		_w16504_,
		_w18342_
	);
	LUT4 #(
		.INIT('h1310)
	) name14295 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8671_,
		_w16322_,
		_w16504_,
		_w18343_
	);
	LUT4 #(
		.INIT('h0008)
	) name14296 (
		_w17524_,
		_w17526_,
		_w18343_,
		_w18342_,
		_w18344_
	);
	LUT3 #(
		.INIT('ha8)
	) name14297 (
		_w11341_,
		_w11409_,
		_w12496_,
		_w18345_
	);
	LUT3 #(
		.INIT('h80)
	) name14298 (
		_w11389_,
		_w11434_,
		_w11843_,
		_w18346_
	);
	LUT4 #(
		.INIT('ha820)
	) name14299 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001 ,
		_w18347_
	);
	LUT3 #(
		.INIT('h07)
	) name14300 (
		_w11529_,
		_w11962_,
		_w18347_,
		_w18348_
	);
	LUT3 #(
		.INIT('h10)
	) name14301 (
		_w11885_,
		_w18346_,
		_w18348_,
		_w18349_
	);
	LUT3 #(
		.INIT('h54)
	) name14302 (
		_w11536_,
		_w11522_,
		_w11523_,
		_w18350_
	);
	LUT3 #(
		.INIT('hc8)
	) name14303 (
		_w11555_,
		_w11854_,
		_w12568_,
		_w18351_
	);
	LUT4 #(
		.INIT('h0100)
	) name14304 (
		_w18345_,
		_w18350_,
		_w18351_,
		_w18349_,
		_w18352_
	);
	LUT2 #(
		.INIT('h1)
	) name14305 (
		_w11492_,
		_w11958_,
		_w18353_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name14306 (
		_w11534_,
		_w11504_,
		_w11864_,
		_w12506_,
		_w18354_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14307 (
		_w11444_,
		_w11428_,
		_w11455_,
		_w11950_,
		_w18355_
	);
	LUT3 #(
		.INIT('h0b)
	) name14308 (
		_w11446_,
		_w11842_,
		_w18355_,
		_w18356_
	);
	LUT4 #(
		.INIT('hf400)
	) name14309 (
		_w11444_,
		_w11423_,
		_w11462_,
		_w11873_,
		_w18357_
	);
	LUT3 #(
		.INIT('h0b)
	) name14310 (
		_w11530_,
		_w11861_,
		_w18357_,
		_w18358_
	);
	LUT4 #(
		.INIT('h4000)
	) name14311 (
		_w18353_,
		_w18356_,
		_w18358_,
		_w18354_,
		_w18359_
	);
	LUT4 #(
		.INIT('h0507)
	) name14312 (
		_w11333_,
		_w11410_,
		_w11558_,
		_w11894_,
		_w18360_
	);
	LUT4 #(
		.INIT('hc080)
	) name14313 (
		_w11335_,
		_w11408_,
		_w12593_,
		_w18360_,
		_w18361_
	);
	LUT3 #(
		.INIT('h80)
	) name14314 (
		_w18352_,
		_w18359_,
		_w18361_,
		_w18362_
	);
	LUT4 #(
		.INIT('h0f04)
	) name14315 (
		_w11444_,
		_w11423_,
		_w11506_,
		_w11462_,
		_w18363_
	);
	LUT3 #(
		.INIT('h40)
	) name14316 (
		_w11444_,
		_w11445_,
		_w11484_,
		_w18364_
	);
	LUT4 #(
		.INIT('h4000)
	) name14317 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11439_,
		_w11495_,
		_w18365_
	);
	LUT4 #(
		.INIT('haaa8)
	) name14318 (
		_w11386_,
		_w18363_,
		_w18364_,
		_w18365_,
		_w18366_
	);
	LUT4 #(
		.INIT('h0040)
	) name14319 (
		_w11549_,
		_w11554_,
		_w18137_,
		_w18366_,
		_w18367_
	);
	LUT4 #(
		.INIT('h8000)
	) name14320 (
		_w11910_,
		_w12411_,
		_w12409_,
		_w18367_,
		_w18368_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name14321 (
		_w11837_,
		_w17556_,
		_w18362_,
		_w18368_,
		_w18369_
	);
	LUT3 #(
		.INIT('h80)
	) name14322 (
		_w8671_,
		_w17563_,
		_w17564_,
		_w18370_
	);
	LUT3 #(
		.INIT('h54)
	) name14323 (
		_w6026_,
		_w17558_,
		_w17559_,
		_w18371_
	);
	LUT3 #(
		.INIT('h80)
	) name14324 (
		_w6039_,
		_w17563_,
		_w17566_,
		_w18372_
	);
	LUT3 #(
		.INIT('h01)
	) name14325 (
		_w18371_,
		_w18372_,
		_w18370_,
		_w18373_
	);
	LUT4 #(
		.INIT('h3230)
	) name14326 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w5999_,
		_w17571_,
		_w17572_,
		_w18374_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14327 (
		_w12450_,
		_w12511_,
		_w12519_,
		_w17569_,
		_w18375_
	);
	LUT4 #(
		.INIT('h3310)
	) name14328 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6001_,
		_w17572_,
		_w17575_,
		_w18376_
	);
	LUT4 #(
		.INIT('h0100)
	) name14329 (
		_w18375_,
		_w18376_,
		_w18374_,
		_w18373_,
		_w18377_
	);
	LUT2 #(
		.INIT('h4)
	) name14330 (
		_w18369_,
		_w18377_,
		_w18378_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14331 (
		_w17524_,
		_w17927_,
		_w18344_,
		_w18378_,
		_w18379_
	);
	LUT2 #(
		.INIT('h4)
	) name14332 (
		_w18341_,
		_w18379_,
		_w18380_
	);
	LUT2 #(
		.INIT('h2)
	) name14333 (
		_w8671_,
		_w17633_,
		_w18381_
	);
	LUT3 #(
		.INIT('he4)
	) name14334 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001 ,
		_w18382_
	);
	LUT3 #(
		.INIT('ha8)
	) name14335 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		_w17511_,
		_w17512_,
		_w18383_
	);
	LUT4 #(
		.INIT('h00bf)
	) name14336 (
		_w17617_,
		_w17635_,
		_w18382_,
		_w18383_,
		_w18384_
	);
	LUT2 #(
		.INIT('h2)
	) name14337 (
		_w6016_,
		_w17588_,
		_w18385_
	);
	LUT2 #(
		.INIT('h8)
	) name14338 (
		_w6007_,
		_w17588_,
		_w18386_
	);
	LUT3 #(
		.INIT('h01)
	) name14339 (
		_w17585_,
		_w18386_,
		_w18385_,
		_w18387_
	);
	LUT3 #(
		.INIT('h80)
	) name14340 (
		_w17514_,
		_w17628_,
		_w18387_,
		_w18388_
	);
	LUT3 #(
		.INIT('h53)
	) name14341 (
		_w6018_,
		_w6009_,
		_w17618_,
		_w18389_
	);
	LUT3 #(
		.INIT('h80)
	) name14342 (
		_w17617_,
		_w17635_,
		_w18389_,
		_w18390_
	);
	LUT4 #(
		.INIT('h0100)
	) name14343 (
		_w17630_,
		_w18388_,
		_w18390_,
		_w18384_,
		_w18391_
	);
	LUT2 #(
		.INIT('h4)
	) name14344 (
		_w18381_,
		_w18391_,
		_w18392_
	);
	LUT2 #(
		.INIT('h4)
	) name14345 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		_w17511_,
		_w18393_
	);
	LUT3 #(
		.INIT('h07)
	) name14346 (
		_w17515_,
		_w17626_,
		_w18393_,
		_w18394_
	);
	LUT4 #(
		.INIT('h1f00)
	) name14347 (
		_w5937_,
		_w6038_,
		_w18182_,
		_w18394_,
		_w18395_
	);
	LUT2 #(
		.INIT('h4)
	) name14348 (
		_w18392_,
		_w18395_,
		_w18396_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14349 (
		_w17627_,
		_w18335_,
		_w18380_,
		_w18396_,
		_w18397_
	);
	LUT4 #(
		.INIT('h3320)
	) name14350 (
		_w12284_,
		_w17587_,
		_w17585_,
		_w18176_,
		_w18398_
	);
	LUT3 #(
		.INIT('h02)
	) name14351 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w11926_,
		_w17586_,
		_w18399_
	);
	LUT3 #(
		.INIT('h54)
	) name14352 (
		_w17515_,
		_w18398_,
		_w18399_,
		_w18400_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14353 (
		_w17515_,
		_w18094_,
		_w18169_,
		_w18400_,
		_w18401_
	);
	LUT4 #(
		.INIT('he400)
	) name14354 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5760_,
		_w8740_,
		_w17585_,
		_w18402_
	);
	LUT4 #(
		.INIT('h4447)
	) name14355 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w17587_,
		_w18217_,
		_w18402_,
		_w18403_
	);
	LUT2 #(
		.INIT('h1)
	) name14356 (
		_w17515_,
		_w18403_,
		_w18404_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14357 (
		_w17515_,
		_w18191_,
		_w18213_,
		_w18404_,
		_w18405_
	);
	LUT4 #(
		.INIT('h3320)
	) name14358 (
		_w14866_,
		_w17587_,
		_w17585_,
		_w18320_,
		_w18406_
	);
	LUT3 #(
		.INIT('h02)
	) name14359 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w11926_,
		_w17586_,
		_w18407_
	);
	LUT3 #(
		.INIT('h54)
	) name14360 (
		_w17515_,
		_w18406_,
		_w18407_,
		_w18408_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14361 (
		_w17515_,
		_w18232_,
		_w18315_,
		_w18408_,
		_w18409_
	);
	LUT4 #(
		.INIT('h3320)
	) name14362 (
		_w12486_,
		_w17587_,
		_w17585_,
		_w18387_,
		_w18410_
	);
	LUT3 #(
		.INIT('h02)
	) name14363 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w11926_,
		_w17586_,
		_w18411_
	);
	LUT3 #(
		.INIT('h54)
	) name14364 (
		_w17515_,
		_w18410_,
		_w18411_,
		_w18412_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14365 (
		_w17515_,
		_w18335_,
		_w18380_,
		_w18412_,
		_w18413_
	);
	LUT3 #(
		.INIT('h02)
	) name14366 (
		_w8717_,
		_w17630_,
		_w17633_,
		_w18414_
	);
	LUT3 #(
		.INIT('he4)
	) name14367 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[12]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[12]/P0001 ,
		_w18415_
	);
	LUT3 #(
		.INIT('h40)
	) name14368 (
		_w17617_,
		_w17635_,
		_w18415_,
		_w18416_
	);
	LUT3 #(
		.INIT('h53)
	) name14369 (
		_w6738_,
		_w6729_,
		_w17618_,
		_w18417_
	);
	LUT3 #(
		.INIT('h80)
	) name14370 (
		_w17617_,
		_w17635_,
		_w18417_,
		_w18418_
	);
	LUT2 #(
		.INIT('h2)
	) name14371 (
		_w6736_,
		_w17588_,
		_w18419_
	);
	LUT2 #(
		.INIT('h8)
	) name14372 (
		_w6727_,
		_w17588_,
		_w18420_
	);
	LUT3 #(
		.INIT('h01)
	) name14373 (
		_w17585_,
		_w18420_,
		_w18419_,
		_w18421_
	);
	LUT3 #(
		.INIT('h80)
	) name14374 (
		_w17514_,
		_w17628_,
		_w18421_,
		_w18422_
	);
	LUT3 #(
		.INIT('h01)
	) name14375 (
		_w18418_,
		_w18422_,
		_w18416_,
		_w18423_
	);
	LUT4 #(
		.INIT('h0700)
	) name14376 (
		_w6758_,
		_w17630_,
		_w18414_,
		_w18423_,
		_w18424_
	);
	LUT3 #(
		.INIT('ha8)
	) name14377 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 ,
		_w17511_,
		_w17512_,
		_w18425_
	);
	LUT3 #(
		.INIT('h07)
	) name14378 (
		_w17515_,
		_w17626_,
		_w18425_,
		_w18426_
	);
	LUT3 #(
		.INIT('he0)
	) name14379 (
		_w17511_,
		_w18424_,
		_w18426_,
		_w18427_
	);
	LUT4 #(
		.INIT('h0105)
	) name14380 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9763_,
		_w12118_,
		_w18428_
	);
	LUT4 #(
		.INIT('ha820)
	) name14381 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w18429_
	);
	LUT4 #(
		.INIT('h007f)
	) name14382 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18429_,
		_w18430_
	);
	LUT3 #(
		.INIT('h8a)
	) name14383 (
		_w17517_,
		_w18428_,
		_w18430_,
		_w18431_
	);
	LUT3 #(
		.INIT('h54)
	) name14384 (
		_w6731_,
		_w17545_,
		_w17546_,
		_w18432_
	);
	LUT3 #(
		.INIT('h54)
	) name14385 (
		_w6734_,
		_w17542_,
		_w17543_,
		_w18433_
	);
	LUT2 #(
		.INIT('h1)
	) name14386 (
		_w18432_,
		_w18433_,
		_w18434_
	);
	LUT2 #(
		.INIT('h8)
	) name14387 (
		_w18095_,
		_w18434_,
		_w18435_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name14388 (
		_w7906_,
		_w17525_,
		_w17526_,
		_w18435_,
		_w18436_
	);
	LUT2 #(
		.INIT('h1)
	) name14389 (
		_w17524_,
		_w18436_,
		_w18437_
	);
	LUT4 #(
		.INIT('h2023)
	) name14390 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w6758_,
		_w16322_,
		_w16504_,
		_w18438_
	);
	LUT4 #(
		.INIT('h1310)
	) name14391 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8717_,
		_w16322_,
		_w16504_,
		_w18439_
	);
	LUT4 #(
		.INIT('h0008)
	) name14392 (
		_w17524_,
		_w17526_,
		_w18439_,
		_w18438_,
		_w18440_
	);
	LUT3 #(
		.INIT('h80)
	) name14393 (
		_w6758_,
		_w17563_,
		_w17566_,
		_w18441_
	);
	LUT3 #(
		.INIT('h54)
	) name14394 (
		_w6746_,
		_w17558_,
		_w17559_,
		_w18442_
	);
	LUT3 #(
		.INIT('h80)
	) name14395 (
		_w8717_,
		_w17563_,
		_w17564_,
		_w18443_
	);
	LUT3 #(
		.INIT('h01)
	) name14396 (
		_w18442_,
		_w18443_,
		_w18441_,
		_w18444_
	);
	LUT4 #(
		.INIT('h3310)
	) name14397 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6721_,
		_w17572_,
		_w17575_,
		_w18445_
	);
	LUT4 #(
		.INIT('h3230)
	) name14398 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6719_,
		_w17571_,
		_w17572_,
		_w18446_
	);
	LUT2 #(
		.INIT('h1)
	) name14399 (
		_w18445_,
		_w18446_,
		_w18447_
	);
	LUT2 #(
		.INIT('h8)
	) name14400 (
		_w18444_,
		_w18447_,
		_w18448_
	);
	LUT3 #(
		.INIT('he0)
	) name14401 (
		_w11420_,
		_w11421_,
		_w11532_,
		_w18449_
	);
	LUT3 #(
		.INIT('hc8)
	) name14402 (
		_w11409_,
		_w11449_,
		_w11896_,
		_w18450_
	);
	LUT4 #(
		.INIT('h00a8)
	) name14403 (
		_w11386_,
		_w11393_,
		_w11589_,
		_w11457_,
		_w18451_
	);
	LUT3 #(
		.INIT('h02)
	) name14404 (
		_w11386_,
		_w11464_,
		_w11953_,
		_w18452_
	);
	LUT4 #(
		.INIT('h0001)
	) name14405 (
		_w18449_,
		_w18450_,
		_w18451_,
		_w18452_,
		_w18453_
	);
	LUT4 #(
		.INIT('ha820)
	) name14406 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001 ,
		_w18454_
	);
	LUT4 #(
		.INIT('h007f)
	) name14407 (
		_w11473_,
		_w11389_,
		_w11962_,
		_w18454_,
		_w18455_
	);
	LUT3 #(
		.INIT('h08)
	) name14408 (
		_w11389_,
		_w11445_,
		_w12639_,
		_w18456_
	);
	LUT2 #(
		.INIT('h8)
	) name14409 (
		_w11415_,
		_w11864_,
		_w18457_
	);
	LUT3 #(
		.INIT('h10)
	) name14410 (
		_w18456_,
		_w18457_,
		_w18455_,
		_w18458_
	);
	LUT4 #(
		.INIT('h0040)
	) name14411 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11401_,
		_w11358_,
		_w12500_,
		_w18459_
	);
	LUT2 #(
		.INIT('h1)
	) name14412 (
		_w11427_,
		_w18459_,
		_w18460_
	);
	LUT3 #(
		.INIT('h80)
	) name14413 (
		_w11389_,
		_w11476_,
		_w11842_,
		_w18461_
	);
	LUT3 #(
		.INIT('h80)
	) name14414 (
		_w11473_,
		_w11389_,
		_w11861_,
		_w18462_
	);
	LUT2 #(
		.INIT('h8)
	) name14415 (
		_w11578_,
		_w11850_,
		_w18463_
	);
	LUT3 #(
		.INIT('h01)
	) name14416 (
		_w18462_,
		_w18463_,
		_w18461_,
		_w18464_
	);
	LUT4 #(
		.INIT('h8000)
	) name14417 (
		_w12473_,
		_w18464_,
		_w18458_,
		_w18460_,
		_w18465_
	);
	LUT3 #(
		.INIT('h04)
	) name14418 (
		_w11536_,
		_w11386_,
		_w11957_,
		_w18466_
	);
	LUT3 #(
		.INIT('hc8)
	) name14419 (
		_w11558_,
		_w11484_,
		_w11894_,
		_w18467_
	);
	LUT2 #(
		.INIT('h1)
	) name14420 (
		_w18466_,
		_w18467_,
		_w18468_
	);
	LUT4 #(
		.INIT('h0777)
	) name14421 (
		_w11587_,
		_w11507_,
		_w11469_,
		_w11973_,
		_w18469_
	);
	LUT4 #(
		.INIT('h153f)
	) name14422 (
		_w11555_,
		_w11588_,
		_w11841_,
		_w11863_,
		_w18470_
	);
	LUT2 #(
		.INIT('h8)
	) name14423 (
		_w18469_,
		_w18470_,
		_w18471_
	);
	LUT2 #(
		.INIT('h2)
	) name14424 (
		_w11855_,
		_w11957_,
		_w18472_
	);
	LUT3 #(
		.INIT('he0)
	) name14425 (
		_w11393_,
		_w11589_,
		_w12504_,
		_w18473_
	);
	LUT4 #(
		.INIT('h7707)
	) name14426 (
		_w11435_,
		_w11872_,
		_w11875_,
		_w11953_,
		_w18474_
	);
	LUT3 #(
		.INIT('h10)
	) name14427 (
		_w18472_,
		_w18473_,
		_w18474_,
		_w18475_
	);
	LUT4 #(
		.INIT('h8000)
	) name14428 (
		_w18471_,
		_w18475_,
		_w18465_,
		_w18468_,
		_w18476_
	);
	LUT4 #(
		.INIT('h8000)
	) name14429 (
		_w12449_,
		_w18250_,
		_w18453_,
		_w18476_,
		_w18477_
	);
	LUT2 #(
		.INIT('h1)
	) name14430 (
		_w11504_,
		_w11844_,
		_w18478_
	);
	LUT4 #(
		.INIT('haf8c)
	) name14431 (
		_w11530_,
		_w11446_,
		_w11855_,
		_w12639_,
		_w18479_
	);
	LUT4 #(
		.INIT('h0400)
	) name14432 (
		_w11595_,
		_w18137_,
		_w18478_,
		_w18479_,
		_w18480_
	);
	LUT4 #(
		.INIT('h8000)
	) name14433 (
		_w11560_,
		_w11584_,
		_w18274_,
		_w18480_,
		_w18481_
	);
	LUT3 #(
		.INIT('h04)
	) name14434 (
		_w11536_,
		_w11386_,
		_w11530_,
		_w18482_
	);
	LUT3 #(
		.INIT('ha8)
	) name14435 (
		_w11341_,
		_w11519_,
		_w11520_,
		_w18483_
	);
	LUT3 #(
		.INIT('h54)
	) name14436 (
		_w11335_,
		_w11522_,
		_w11523_,
		_w18484_
	);
	LUT3 #(
		.INIT('h01)
	) name14437 (
		_w18483_,
		_w18484_,
		_w18482_,
		_w18485_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14438 (
		_w11444_,
		_w11423_,
		_w11462_,
		_w11950_,
		_w18486_
	);
	LUT3 #(
		.INIT('h0e)
	) name14439 (
		_w11534_,
		_w12500_,
		_w18486_,
		_w18487_
	);
	LUT4 #(
		.INIT('hf400)
	) name14440 (
		_w11444_,
		_w11414_,
		_w11481_,
		_w11864_,
		_w18488_
	);
	LUT3 #(
		.INIT('h0b)
	) name14441 (
		_w11492_,
		_w12504_,
		_w18488_,
		_w18489_
	);
	LUT3 #(
		.INIT('h02)
	) name14442 (
		_w11386_,
		_w11492_,
		_w11457_,
		_w18490_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14443 (
		_w11444_,
		_w11428_,
		_w11455_,
		_w11958_,
		_w18491_
	);
	LUT4 #(
		.INIT('ha820)
	) name14444 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001 ,
		_w18492_
	);
	LUT2 #(
		.INIT('h1)
	) name14445 (
		_w18491_,
		_w18492_,
		_w18493_
	);
	LUT4 #(
		.INIT('h4000)
	) name14446 (
		_w18490_,
		_w18493_,
		_w18487_,
		_w18489_,
		_w18494_
	);
	LUT3 #(
		.INIT('h80)
	) name14447 (
		_w11417_,
		_w18485_,
		_w18494_,
		_w18495_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name14448 (
		_w12695_,
		_w17556_,
		_w18495_,
		_w18481_,
		_w18496_
	);
	LUT3 #(
		.INIT('h0d)
	) name14449 (
		_w17569_,
		_w18477_,
		_w18496_,
		_w18497_
	);
	LUT2 #(
		.INIT('h8)
	) name14450 (
		_w18448_,
		_w18497_,
		_w18498_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14451 (
		_w17524_,
		_w17927_,
		_w18440_,
		_w18498_,
		_w18499_
	);
	LUT2 #(
		.INIT('h4)
	) name14452 (
		_w18437_,
		_w18499_,
		_w18500_
	);
	LUT4 #(
		.INIT('h3133)
	) name14453 (
		_w17627_,
		_w18427_,
		_w18431_,
		_w18500_,
		_w18501_
	);
	LUT4 #(
		.INIT('he400)
	) name14454 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w17585_,
		_w18502_
	);
	LUT4 #(
		.INIT('h4447)
	) name14455 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w17587_,
		_w18421_,
		_w18502_,
		_w18503_
	);
	LUT2 #(
		.INIT('h1)
	) name14456 (
		_w17515_,
		_w18503_,
		_w18504_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14457 (
		_w17515_,
		_w18431_,
		_w18500_,
		_w18504_,
		_w18505_
	);
	LUT4 #(
		.INIT('h4500)
	) name14458 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w17630_,
		_w18506_
	);
	LUT3 #(
		.INIT('h02)
	) name14459 (
		_w8974_,
		_w17630_,
		_w17633_,
		_w18507_
	);
	LUT3 #(
		.INIT('he4)
	) name14460 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[7]/P0001 ,
		_w18508_
	);
	LUT3 #(
		.INIT('h40)
	) name14461 (
		_w17617_,
		_w17635_,
		_w18508_,
		_w18509_
	);
	LUT3 #(
		.INIT('h53)
	) name14462 (
		_w7891_,
		_w7893_,
		_w17618_,
		_w18510_
	);
	LUT3 #(
		.INIT('h80)
	) name14463 (
		_w17617_,
		_w17635_,
		_w18510_,
		_w18511_
	);
	LUT2 #(
		.INIT('h2)
	) name14464 (
		_w7886_,
		_w17588_,
		_w18512_
	);
	LUT2 #(
		.INIT('h8)
	) name14465 (
		_w7895_,
		_w17588_,
		_w18513_
	);
	LUT3 #(
		.INIT('h01)
	) name14466 (
		_w17585_,
		_w18513_,
		_w18512_,
		_w18514_
	);
	LUT3 #(
		.INIT('h80)
	) name14467 (
		_w17514_,
		_w17628_,
		_w18514_,
		_w18515_
	);
	LUT3 #(
		.INIT('h01)
	) name14468 (
		_w18511_,
		_w18515_,
		_w18509_,
		_w18516_
	);
	LUT2 #(
		.INIT('h4)
	) name14469 (
		_w18507_,
		_w18516_,
		_w18517_
	);
	LUT3 #(
		.INIT('ha8)
	) name14470 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w17511_,
		_w17512_,
		_w18518_
	);
	LUT3 #(
		.INIT('h07)
	) name14471 (
		_w17515_,
		_w17626_,
		_w18518_,
		_w18519_
	);
	LUT4 #(
		.INIT('hba00)
	) name14472 (
		_w17511_,
		_w18506_,
		_w18517_,
		_w18519_,
		_w18520_
	);
	LUT4 #(
		.INIT('h0015)
	) name14473 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w14583_,
		_w18521_
	);
	LUT3 #(
		.INIT('h02)
	) name14474 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w12560_,
		_w12561_,
		_w18522_
	);
	LUT4 #(
		.INIT('h007f)
	) name14475 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18522_,
		_w18523_
	);
	LUT3 #(
		.INIT('h8a)
	) name14476 (
		_w17517_,
		_w18521_,
		_w18523_,
		_w18524_
	);
	LUT3 #(
		.INIT('h54)
	) name14477 (
		_w7888_,
		_w17545_,
		_w17546_,
		_w18525_
	);
	LUT3 #(
		.INIT('h54)
	) name14478 (
		_w7884_,
		_w17542_,
		_w17543_,
		_w18526_
	);
	LUT2 #(
		.INIT('h1)
	) name14479 (
		_w18525_,
		_w18526_,
		_w18527_
	);
	LUT2 #(
		.INIT('h8)
	) name14480 (
		_w18095_,
		_w18527_,
		_w18528_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name14481 (
		_w7906_,
		_w17525_,
		_w17526_,
		_w18528_,
		_w18529_
	);
	LUT2 #(
		.INIT('h1)
	) name14482 (
		_w17524_,
		_w18529_,
		_w18530_
	);
	LUT4 #(
		.INIT('h1310)
	) name14483 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8974_,
		_w16322_,
		_w16504_,
		_w18531_
	);
	LUT4 #(
		.INIT('h2023)
	) name14484 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w7906_,
		_w16322_,
		_w16504_,
		_w18532_
	);
	LUT4 #(
		.INIT('h0008)
	) name14485 (
		_w17524_,
		_w17526_,
		_w18532_,
		_w18531_,
		_w18533_
	);
	LUT4 #(
		.INIT('h3230)
	) name14486 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7864_,
		_w17571_,
		_w17572_,
		_w18534_
	);
	LUT4 #(
		.INIT('h3310)
	) name14487 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7866_,
		_w17572_,
		_w17575_,
		_w18535_
	);
	LUT4 #(
		.INIT('ha820)
	) name14488 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001 ,
		_w18536_
	);
	LUT3 #(
		.INIT('h07)
	) name14489 (
		_w11429_,
		_w11508_,
		_w18536_,
		_w18537_
	);
	LUT3 #(
		.INIT('h80)
	) name14490 (
		_w11473_,
		_w11389_,
		_w11470_,
		_w18538_
	);
	LUT2 #(
		.INIT('h8)
	) name14491 (
		_w11578_,
		_w11488_,
		_w18539_
	);
	LUT3 #(
		.INIT('h10)
	) name14492 (
		_w18538_,
		_w18539_,
		_w18537_,
		_w18540_
	);
	LUT4 #(
		.INIT('h4000)
	) name14493 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11401_,
		_w11358_,
		_w11470_,
		_w18541_
	);
	LUT2 #(
		.INIT('h1)
	) name14494 (
		_w11570_,
		_w18541_,
		_w18542_
	);
	LUT4 #(
		.INIT('h0001)
	) name14495 (
		_w11403_,
		_w11438_,
		_w11885_,
		_w12472_,
		_w18543_
	);
	LUT3 #(
		.INIT('h80)
	) name14496 (
		_w18540_,
		_w18542_,
		_w18543_,
		_w18544_
	);
	LUT3 #(
		.INIT('hc8)
	) name14497 (
		_w11547_,
		_w11495_,
		_w11976_,
		_w18545_
	);
	LUT4 #(
		.INIT('h00a8)
	) name14498 (
		_w11386_,
		_w11393_,
		_w11589_,
		_w11452_,
		_w18546_
	);
	LUT2 #(
		.INIT('h1)
	) name14499 (
		_w18545_,
		_w18546_,
		_w18547_
	);
	LUT3 #(
		.INIT('he0)
	) name14500 (
		_w11393_,
		_w11589_,
		_w11450_,
		_w18548_
	);
	LUT3 #(
		.INIT('hc8)
	) name14501 (
		_w11552_,
		_w11466_,
		_w11474_,
		_w18549_
	);
	LUT4 #(
		.INIT('h7077)
	) name14502 (
		_w11409_,
		_w11863_,
		_w11954_,
		_w12412_,
		_w18550_
	);
	LUT3 #(
		.INIT('h10)
	) name14503 (
		_w18548_,
		_w18549_,
		_w18550_,
		_w18551_
	);
	LUT4 #(
		.INIT('heee0)
	) name14504 (
		_w11542_,
		_w11592_,
		_w11957_,
		_w12024_,
		_w18552_
	);
	LUT4 #(
		.INIT('h51f3)
	) name14505 (
		_w11507_,
		_w11511_,
		_w11953_,
		_w12468_,
		_w18553_
	);
	LUT2 #(
		.INIT('h8)
	) name14506 (
		_w18552_,
		_w18553_,
		_w18554_
	);
	LUT4 #(
		.INIT('h8000)
	) name14507 (
		_w18551_,
		_w18554_,
		_w18544_,
		_w18547_,
		_w18555_
	);
	LUT3 #(
		.INIT('he0)
	) name14508 (
		_w11420_,
		_w11421_,
		_w11499_,
		_w18556_
	);
	LUT3 #(
		.INIT('h02)
	) name14509 (
		_w11386_,
		_w11528_,
		_w11954_,
		_w18557_
	);
	LUT3 #(
		.INIT('ha8)
	) name14510 (
		_w11484_,
		_w11973_,
		_w11974_,
		_w18558_
	);
	LUT3 #(
		.INIT('h01)
	) name14511 (
		_w18557_,
		_w18558_,
		_w18556_,
		_w18559_
	);
	LUT3 #(
		.INIT('h80)
	) name14512 (
		_w11910_,
		_w11972_,
		_w18559_,
		_w18560_
	);
	LUT4 #(
		.INIT('h3111)
	) name14513 (
		_w17569_,
		_w18535_,
		_w18555_,
		_w18560_,
		_w18561_
	);
	LUT2 #(
		.INIT('h4)
	) name14514 (
		_w18534_,
		_w18561_,
		_w18562_
	);
	LUT3 #(
		.INIT('h54)
	) name14515 (
		_w7878_,
		_w17558_,
		_w17559_,
		_w18563_
	);
	LUT3 #(
		.INIT('h80)
	) name14516 (
		_w7906_,
		_w17563_,
		_w17566_,
		_w18564_
	);
	LUT3 #(
		.INIT('h80)
	) name14517 (
		_w8974_,
		_w17563_,
		_w17564_,
		_w18565_
	);
	LUT3 #(
		.INIT('h01)
	) name14518 (
		_w18564_,
		_w18565_,
		_w18563_,
		_w18566_
	);
	LUT3 #(
		.INIT('hb0)
	) name14519 (
		_w12600_,
		_w17556_,
		_w18566_,
		_w18567_
	);
	LUT2 #(
		.INIT('h8)
	) name14520 (
		_w18562_,
		_w18567_,
		_w18568_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14521 (
		_w17524_,
		_w17927_,
		_w18533_,
		_w18568_,
		_w18569_
	);
	LUT2 #(
		.INIT('h4)
	) name14522 (
		_w18530_,
		_w18569_,
		_w18570_
	);
	LUT4 #(
		.INIT('h3133)
	) name14523 (
		_w17627_,
		_w18520_,
		_w18524_,
		_w18570_,
		_w18571_
	);
	LUT3 #(
		.INIT('h40)
	) name14524 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w18572_
	);
	LUT4 #(
		.INIT('hff48)
	) name14525 (
		\sport1_cfg_FSi_cnt_reg[14]/NET0131 ,
		_w17698_,
		_w17673_,
		_w18572_,
		_w18573_
	);
	LUT3 #(
		.INIT('h02)
	) name14526 (
		_w8781_,
		_w17630_,
		_w17633_,
		_w18574_
	);
	LUT3 #(
		.INIT('h10)
	) name14527 (
		_w8757_,
		_w8760_,
		_w17630_,
		_w18575_
	);
	LUT3 #(
		.INIT('he4)
	) name14528 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[14]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[14]/P0001 ,
		_w18576_
	);
	LUT3 #(
		.INIT('h40)
	) name14529 (
		_w17617_,
		_w17635_,
		_w18576_,
		_w18577_
	);
	LUT3 #(
		.INIT('h53)
	) name14530 (
		_w8299_,
		_w8301_,
		_w17618_,
		_w18578_
	);
	LUT3 #(
		.INIT('h80)
	) name14531 (
		_w17617_,
		_w17635_,
		_w18578_,
		_w18579_
	);
	LUT2 #(
		.INIT('h2)
	) name14532 (
		_w8294_,
		_w17588_,
		_w18580_
	);
	LUT2 #(
		.INIT('h8)
	) name14533 (
		_w8303_,
		_w17588_,
		_w18581_
	);
	LUT3 #(
		.INIT('h01)
	) name14534 (
		_w17585_,
		_w18581_,
		_w18580_,
		_w18582_
	);
	LUT3 #(
		.INIT('h80)
	) name14535 (
		_w17514_,
		_w17628_,
		_w18582_,
		_w18583_
	);
	LUT3 #(
		.INIT('h01)
	) name14536 (
		_w18579_,
		_w18583_,
		_w18577_,
		_w18584_
	);
	LUT4 #(
		.INIT('h5455)
	) name14537 (
		_w17511_,
		_w18574_,
		_w18575_,
		_w18584_,
		_w18585_
	);
	LUT3 #(
		.INIT('ha8)
	) name14538 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 ,
		_w17511_,
		_w17512_,
		_w18586_
	);
	LUT3 #(
		.INIT('h07)
	) name14539 (
		_w17515_,
		_w17626_,
		_w18586_,
		_w18587_
	);
	LUT2 #(
		.INIT('h4)
	) name14540 (
		_w18585_,
		_w18587_,
		_w18588_
	);
	LUT4 #(
		.INIT('h1050)
	) name14541 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9828_,
		_w12118_,
		_w18589_
	);
	LUT2 #(
		.INIT('h8)
	) name14542 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w12673_,
		_w18590_
	);
	LUT4 #(
		.INIT('h007f)
	) name14543 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18590_,
		_w18591_
	);
	LUT3 #(
		.INIT('h8a)
	) name14544 (
		_w17517_,
		_w18589_,
		_w18591_,
		_w18592_
	);
	LUT3 #(
		.INIT('h54)
	) name14545 (
		_w8296_,
		_w17545_,
		_w17546_,
		_w18593_
	);
	LUT3 #(
		.INIT('h54)
	) name14546 (
		_w8292_,
		_w17542_,
		_w17543_,
		_w18594_
	);
	LUT2 #(
		.INIT('h1)
	) name14547 (
		_w18593_,
		_w18594_,
		_w18595_
	);
	LUT2 #(
		.INIT('h8)
	) name14548 (
		_w18095_,
		_w18595_,
		_w18596_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name14549 (
		_w7906_,
		_w17525_,
		_w17526_,
		_w18596_,
		_w18597_
	);
	LUT2 #(
		.INIT('h1)
	) name14550 (
		_w17524_,
		_w18597_,
		_w18598_
	);
	LUT4 #(
		.INIT('h2023)
	) name14551 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8761_,
		_w16322_,
		_w16504_,
		_w18599_
	);
	LUT4 #(
		.INIT('h1310)
	) name14552 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8781_,
		_w16322_,
		_w16504_,
		_w18600_
	);
	LUT4 #(
		.INIT('h0008)
	) name14553 (
		_w17524_,
		_w17526_,
		_w18600_,
		_w18599_,
		_w18601_
	);
	LUT2 #(
		.INIT('h4)
	) name14554 (
		_w13314_,
		_w17569_,
		_w18602_
	);
	LUT3 #(
		.INIT('h80)
	) name14555 (
		_w8781_,
		_w17563_,
		_w17564_,
		_w18603_
	);
	LUT3 #(
		.INIT('h54)
	) name14556 (
		_w8267_,
		_w17558_,
		_w17559_,
		_w18604_
	);
	LUT3 #(
		.INIT('h80)
	) name14557 (
		_w8761_,
		_w17563_,
		_w17566_,
		_w18605_
	);
	LUT3 #(
		.INIT('h01)
	) name14558 (
		_w18604_,
		_w18605_,
		_w18603_,
		_w18606_
	);
	LUT4 #(
		.INIT('h3230)
	) name14559 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w8284_,
		_w17571_,
		_w17572_,
		_w18607_
	);
	LUT4 #(
		.INIT('h3310)
	) name14560 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w8286_,
		_w17572_,
		_w17575_,
		_w18608_
	);
	LUT2 #(
		.INIT('h1)
	) name14561 (
		_w18607_,
		_w18608_,
		_w18609_
	);
	LUT4 #(
		.INIT('hb000)
	) name14562 (
		_w12696_,
		_w17556_,
		_w18606_,
		_w18609_,
		_w18610_
	);
	LUT2 #(
		.INIT('h4)
	) name14563 (
		_w18602_,
		_w18610_,
		_w18611_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14564 (
		_w17524_,
		_w17927_,
		_w18601_,
		_w18611_,
		_w18612_
	);
	LUT2 #(
		.INIT('h4)
	) name14565 (
		_w18598_,
		_w18612_,
		_w18613_
	);
	LUT4 #(
		.INIT('h3133)
	) name14566 (
		_w17627_,
		_w18588_,
		_w18592_,
		_w18613_,
		_w18614_
	);
	LUT3 #(
		.INIT('h40)
	) name14567 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w18615_
	);
	LUT4 #(
		.INIT('hff48)
	) name14568 (
		\sport0_cfg_FSi_cnt_reg[14]/NET0131 ,
		_w17734_,
		_w17709_,
		_w18615_,
		_w18616_
	);
	LUT4 #(
		.INIT('h00ef)
	) name14569 (
		_w12560_,
		_w12561_,
		_w17585_,
		_w18514_,
		_w18617_
	);
	LUT4 #(
		.INIT('h2023)
	) name14570 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w17515_,
		_w17587_,
		_w18617_,
		_w18618_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14571 (
		_w17515_,
		_w18524_,
		_w18570_,
		_w18618_,
		_w18619_
	);
	LUT4 #(
		.INIT('h3320)
	) name14572 (
		_w12673_,
		_w17587_,
		_w17585_,
		_w18582_,
		_w18620_
	);
	LUT3 #(
		.INIT('h02)
	) name14573 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w11926_,
		_w17586_,
		_w18621_
	);
	LUT3 #(
		.INIT('h54)
	) name14574 (
		_w17515_,
		_w18620_,
		_w18621_,
		_w18622_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14575 (
		_w17515_,
		_w18592_,
		_w18613_,
		_w18622_,
		_w18623_
	);
	LUT4 #(
		.INIT('h0105)
	) name14576 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9890_,
		_w12118_,
		_w18624_
	);
	LUT2 #(
		.INIT('h8)
	) name14577 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w14918_,
		_w18625_
	);
	LUT4 #(
		.INIT('h007f)
	) name14578 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18625_,
		_w18626_
	);
	LUT3 #(
		.INIT('h8a)
	) name14579 (
		_w17517_,
		_w18624_,
		_w18626_,
		_w18627_
	);
	LUT3 #(
		.INIT('h54)
	) name14580 (
		_w7549_,
		_w17545_,
		_w17546_,
		_w18628_
	);
	LUT3 #(
		.INIT('h54)
	) name14581 (
		_w7545_,
		_w17542_,
		_w17543_,
		_w18629_
	);
	LUT2 #(
		.INIT('h1)
	) name14582 (
		_w18628_,
		_w18629_,
		_w18630_
	);
	LUT2 #(
		.INIT('h8)
	) name14583 (
		_w18095_,
		_w18630_,
		_w18631_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name14584 (
		_w7906_,
		_w17525_,
		_w17526_,
		_w18631_,
		_w18632_
	);
	LUT2 #(
		.INIT('h1)
	) name14585 (
		_w17524_,
		_w18632_,
		_w18633_
	);
	LUT4 #(
		.INIT('h2023)
	) name14586 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w7566_,
		_w16322_,
		_w16504_,
		_w18634_
	);
	LUT4 #(
		.INIT('h1310)
	) name14587 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w8998_,
		_w16322_,
		_w16504_,
		_w18635_
	);
	LUT4 #(
		.INIT('h0008)
	) name14588 (
		_w17524_,
		_w17526_,
		_w18635_,
		_w18634_,
		_w18636_
	);
	LUT4 #(
		.INIT('h8acf)
	) name14589 (
		_w11530_,
		_w11492_,
		_w11850_,
		_w12504_,
		_w18637_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14590 (
		_w11444_,
		_w11428_,
		_w11455_,
		_w12639_,
		_w18638_
	);
	LUT3 #(
		.INIT('h07)
	) name14591 (
		_w11555_,
		_w11860_,
		_w18638_,
		_w18639_
	);
	LUT4 #(
		.INIT('h7077)
	) name14592 (
		_w11341_,
		_w11435_,
		_w11457_,
		_w11839_,
		_w18640_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14593 (
		_w11444_,
		_w11423_,
		_w11462_,
		_w11844_,
		_w18641_
	);
	LUT3 #(
		.INIT('h0b)
	) name14594 (
		_w11446_,
		_w11864_,
		_w18641_,
		_w18642_
	);
	LUT4 #(
		.INIT('h8000)
	) name14595 (
		_w18640_,
		_w18642_,
		_w18637_,
		_w18639_,
		_w18643_
	);
	LUT2 #(
		.INIT('h1)
	) name14596 (
		_w11534_,
		_w11958_,
		_w18644_
	);
	LUT4 #(
		.INIT('h45cf)
	) name14597 (
		_w11588_,
		_w11494_,
		_w11522_,
		_w11854_,
		_w18645_
	);
	LUT3 #(
		.INIT('h10)
	) name14598 (
		_w11595_,
		_w18644_,
		_w18645_,
		_w18646_
	);
	LUT2 #(
		.INIT('h8)
	) name14599 (
		_w18643_,
		_w18646_,
		_w18647_
	);
	LUT3 #(
		.INIT('h02)
	) name14600 (
		_w11386_,
		_w11492_,
		_w11448_,
		_w18648_
	);
	LUT3 #(
		.INIT('ha8)
	) name14601 (
		_w11537_,
		_w11410_,
		_w11558_,
		_w18649_
	);
	LUT3 #(
		.INIT('hc8)
	) name14602 (
		_w11587_,
		_w11532_,
		_w11880_,
		_w18650_
	);
	LUT4 #(
		.INIT('h0002)
	) name14603 (
		_w17822_,
		_w18648_,
		_w18649_,
		_w18650_,
		_w18651_
	);
	LUT4 #(
		.INIT('h2000)
	) name14604 (
		_w11389_,
		_w11536_,
		_w11386_,
		_w11476_,
		_w18652_
	);
	LUT3 #(
		.INIT('h40)
	) name14605 (
		_w11385_,
		_w11415_,
		_w11860_,
		_w18653_
	);
	LUT3 #(
		.INIT('h01)
	) name14606 (
		_w11579_,
		_w18653_,
		_w18652_,
		_w18654_
	);
	LUT4 #(
		.INIT('ha820)
	) name14607 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001 ,
		_w18655_
	);
	LUT3 #(
		.INIT('h07)
	) name14608 (
		_w11529_,
		_w12505_,
		_w18655_,
		_w18656_
	);
	LUT2 #(
		.INIT('h8)
	) name14609 (
		_w11415_,
		_w11962_,
		_w18657_
	);
	LUT3 #(
		.INIT('h80)
	) name14610 (
		_w11389_,
		_w11476_,
		_w11855_,
		_w18658_
	);
	LUT3 #(
		.INIT('h10)
	) name14611 (
		_w18657_,
		_w18658_,
		_w18656_,
		_w18659_
	);
	LUT3 #(
		.INIT('h40)
	) name14612 (
		_w11586_,
		_w18659_,
		_w18654_,
		_w18660_
	);
	LUT2 #(
		.INIT('h2)
	) name14613 (
		_w11554_,
		_w12597_,
		_w18661_
	);
	LUT4 #(
		.INIT('h8000)
	) name14614 (
		_w11902_,
		_w18660_,
		_w18661_,
		_w18651_,
		_w18662_
	);
	LUT4 #(
		.INIT('h8000)
	) name14615 (
		_w12591_,
		_w17801_,
		_w18647_,
		_w18662_,
		_w18663_
	);
	LUT2 #(
		.INIT('h2)
	) name14616 (
		_w17556_,
		_w18663_,
		_w18664_
	);
	LUT3 #(
		.INIT('h54)
	) name14617 (
		_w7538_,
		_w17558_,
		_w17559_,
		_w18665_
	);
	LUT3 #(
		.INIT('h80)
	) name14618 (
		_w7566_,
		_w17563_,
		_w17566_,
		_w18666_
	);
	LUT3 #(
		.INIT('h80)
	) name14619 (
		_w8998_,
		_w17563_,
		_w17564_,
		_w18667_
	);
	LUT3 #(
		.INIT('h01)
	) name14620 (
		_w18666_,
		_w18667_,
		_w18665_,
		_w18668_
	);
	LUT4 #(
		.INIT('h3310)
	) name14621 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7528_,
		_w17572_,
		_w17575_,
		_w18669_
	);
	LUT3 #(
		.INIT('h32)
	) name14622 (
		_w11409_,
		_w11483_,
		_w11896_,
		_w18670_
	);
	LUT3 #(
		.INIT('hc8)
	) name14623 (
		_w11435_,
		_w11863_,
		_w12455_,
		_w18671_
	);
	LUT3 #(
		.INIT('h02)
	) name14624 (
		_w11386_,
		_w11457_,
		_w11957_,
		_w18672_
	);
	LUT4 #(
		.INIT('h0a08)
	) name14625 (
		_w11386_,
		_w11552_,
		_w11464_,
		_w11474_,
		_w18673_
	);
	LUT4 #(
		.INIT('h0001)
	) name14626 (
		_w18670_,
		_w18671_,
		_w18672_,
		_w18673_,
		_w18674_
	);
	LUT2 #(
		.INIT('h2)
	) name14627 (
		_w11852_,
		_w11953_,
		_w18675_
	);
	LUT3 #(
		.INIT('h0e)
	) name14628 (
		_w11393_,
		_w11589_,
		_w11950_,
		_w18676_
	);
	LUT4 #(
		.INIT('h4000)
	) name14629 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11382_,
		_w11873_,
		_w18677_
	);
	LUT4 #(
		.INIT('ha820)
	) name14630 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001 ,
		_w18678_
	);
	LUT2 #(
		.INIT('h1)
	) name14631 (
		_w18677_,
		_w18678_,
		_w18679_
	);
	LUT3 #(
		.INIT('h10)
	) name14632 (
		_w18676_,
		_w18675_,
		_w18679_,
		_w18680_
	);
	LUT3 #(
		.INIT('hc8)
	) name14633 (
		_w11547_,
		_w11860_,
		_w11976_,
		_w18681_
	);
	LUT3 #(
		.INIT('ha8)
	) name14634 (
		_w11841_,
		_w11973_,
		_w11974_,
		_w18682_
	);
	LUT2 #(
		.INIT('h1)
	) name14635 (
		_w18681_,
		_w18682_,
		_w18683_
	);
	LUT3 #(
		.INIT('h80)
	) name14636 (
		_w18680_,
		_w18683_,
		_w18674_,
		_w18684_
	);
	LUT2 #(
		.INIT('h8)
	) name14637 (
		_w11429_,
		_w11872_,
		_w18685_
	);
	LUT4 #(
		.INIT('h0045)
	) name14638 (
		_w11551_,
		_w11592_,
		_w11854_,
		_w18685_,
		_w18686_
	);
	LUT4 #(
		.INIT('h5455)
	) name14639 (
		_w11386_,
		_w18115_,
		_w18116_,
		_w18686_,
		_w18687_
	);
	LUT3 #(
		.INIT('h04)
	) name14640 (
		_w11536_,
		_w11386_,
		_w11592_,
		_w18688_
	);
	LUT3 #(
		.INIT('h02)
	) name14641 (
		_w11386_,
		_w11335_,
		_w11954_,
		_w18689_
	);
	LUT3 #(
		.INIT('he0)
	) name14642 (
		_w11420_,
		_w11421_,
		_w11495_,
		_w18690_
	);
	LUT3 #(
		.INIT('h01)
	) name14643 (
		_w18689_,
		_w18690_,
		_w18688_,
		_w18691_
	);
	LUT2 #(
		.INIT('h4)
	) name14644 (
		_w18687_,
		_w18691_,
		_w18692_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name14645 (
		_w17569_,
		_w18113_,
		_w18684_,
		_w18692_,
		_w18693_
	);
	LUT4 #(
		.INIT('h3230)
	) name14646 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w7526_,
		_w17571_,
		_w17572_,
		_w18694_
	);
	LUT4 #(
		.INIT('h0100)
	) name14647 (
		_w18693_,
		_w18694_,
		_w18669_,
		_w18668_,
		_w18695_
	);
	LUT2 #(
		.INIT('h4)
	) name14648 (
		_w18664_,
		_w18695_,
		_w18696_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14649 (
		_w17524_,
		_w17927_,
		_w18636_,
		_w18696_,
		_w18697_
	);
	LUT2 #(
		.INIT('h4)
	) name14650 (
		_w18633_,
		_w18697_,
		_w18698_
	);
	LUT3 #(
		.INIT('h10)
	) name14651 (
		_w7465_,
		_w7565_,
		_w17630_,
		_w18699_
	);
	LUT2 #(
		.INIT('h8)
	) name14652 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		_w17512_,
		_w18700_
	);
	LUT2 #(
		.INIT('h2)
	) name14653 (
		_w7547_,
		_w17588_,
		_w18701_
	);
	LUT2 #(
		.INIT('h8)
	) name14654 (
		_w7556_,
		_w17588_,
		_w18702_
	);
	LUT3 #(
		.INIT('h01)
	) name14655 (
		_w17585_,
		_w18702_,
		_w18701_,
		_w18703_
	);
	LUT4 #(
		.INIT('h070f)
	) name14656 (
		_w17514_,
		_w17628_,
		_w18700_,
		_w18703_,
		_w18704_
	);
	LUT3 #(
		.INIT('h53)
	) name14657 (
		_w7552_,
		_w7554_,
		_w17618_,
		_w18705_
	);
	LUT3 #(
		.INIT('he4)
	) name14658 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[8]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[8]/P0001 ,
		_w18706_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14659 (
		_w17617_,
		_w17635_,
		_w18705_,
		_w18706_,
		_w18707_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name14660 (
		_w17630_,
		_w17632_,
		_w18704_,
		_w18707_,
		_w18708_
	);
	LUT4 #(
		.INIT('h3331)
	) name14661 (
		_w8998_,
		_w17511_,
		_w17630_,
		_w17633_,
		_w18709_
	);
	LUT2 #(
		.INIT('h4)
	) name14662 (
		_w18708_,
		_w18709_,
		_w18710_
	);
	LUT2 #(
		.INIT('h4)
	) name14663 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		_w17511_,
		_w18711_
	);
	LUT3 #(
		.INIT('h07)
	) name14664 (
		_w17515_,
		_w17626_,
		_w18711_,
		_w18712_
	);
	LUT3 #(
		.INIT('hb0)
	) name14665 (
		_w18699_,
		_w18710_,
		_w18712_,
		_w18713_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14666 (
		_w17627_,
		_w18627_,
		_w18698_,
		_w18713_,
		_w18714_
	);
	LUT4 #(
		.INIT('h3320)
	) name14667 (
		_w14918_,
		_w17587_,
		_w17585_,
		_w18703_,
		_w18715_
	);
	LUT3 #(
		.INIT('h02)
	) name14668 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w11926_,
		_w17586_,
		_w18716_
	);
	LUT3 #(
		.INIT('h54)
	) name14669 (
		_w17515_,
		_w18715_,
		_w18716_,
		_w18717_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14670 (
		_w17515_,
		_w18627_,
		_w18698_,
		_w18717_,
		_w18718_
	);
	LUT4 #(
		.INIT('h0105)
	) name14671 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9866_,
		_w12118_,
		_w18719_
	);
	LUT3 #(
		.INIT('h02)
	) name14672 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w13610_,
		_w13611_,
		_w18720_
	);
	LUT4 #(
		.INIT('h007f)
	) name14673 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18720_,
		_w18721_
	);
	LUT3 #(
		.INIT('h8a)
	) name14674 (
		_w17517_,
		_w18719_,
		_w18721_,
		_w18722_
	);
	LUT4 #(
		.INIT('hacc0)
	) name14675 (
		_w6176_,
		_w8885_,
		_w17525_,
		_w17526_,
		_w18723_
	);
	LUT3 #(
		.INIT('ha8)
	) name14676 (
		_w17524_,
		_w17527_,
		_w18723_,
		_w18724_
	);
	LUT3 #(
		.INIT('h54)
	) name14677 (
		_w6148_,
		_w17542_,
		_w17543_,
		_w18725_
	);
	LUT3 #(
		.INIT('h54)
	) name14678 (
		_w6145_,
		_w17539_,
		_w17540_,
		_w18726_
	);
	LUT3 #(
		.INIT('h54)
	) name14679 (
		_w6141_,
		_w17545_,
		_w17546_,
		_w18727_
	);
	LUT3 #(
		.INIT('h01)
	) name14680 (
		_w18726_,
		_w18727_,
		_w18725_,
		_w18728_
	);
	LUT2 #(
		.INIT('h8)
	) name14681 (
		_w17538_,
		_w18728_,
		_w18729_
	);
	LUT2 #(
		.INIT('h8)
	) name14682 (
		_w17525_,
		_w18729_,
		_w18730_
	);
	LUT4 #(
		.INIT('h1310)
	) name14683 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w6176_,
		_w16322_,
		_w16504_,
		_w18731_
	);
	LUT3 #(
		.INIT('h04)
	) name14684 (
		_w17524_,
		_w17526_,
		_w18731_,
		_w18732_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14685 (
		_w12451_,
		_w13224_,
		_w13631_,
		_w17556_,
		_w18733_
	);
	LUT3 #(
		.INIT('h80)
	) name14686 (
		_w6176_,
		_w17563_,
		_w17566_,
		_w18734_
	);
	LUT4 #(
		.INIT('h008f)
	) name14687 (
		_w13793_,
		_w13805_,
		_w17569_,
		_w18734_,
		_w18735_
	);
	LUT3 #(
		.INIT('h54)
	) name14688 (
		_w6163_,
		_w17558_,
		_w17559_,
		_w18736_
	);
	LUT3 #(
		.INIT('h80)
	) name14689 (
		_w8885_,
		_w17563_,
		_w17564_,
		_w18737_
	);
	LUT2 #(
		.INIT('h1)
	) name14690 (
		_w18736_,
		_w18737_,
		_w18738_
	);
	LUT4 #(
		.INIT('h3310)
	) name14691 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6135_,
		_w17572_,
		_w17575_,
		_w18739_
	);
	LUT4 #(
		.INIT('h3230)
	) name14692 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6137_,
		_w17571_,
		_w17572_,
		_w18740_
	);
	LUT2 #(
		.INIT('h1)
	) name14693 (
		_w18739_,
		_w18740_,
		_w18741_
	);
	LUT4 #(
		.INIT('h4000)
	) name14694 (
		_w18733_,
		_w18735_,
		_w18738_,
		_w18741_,
		_w18742_
	);
	LUT3 #(
		.INIT('hb0)
	) name14695 (
		_w18730_,
		_w18732_,
		_w18742_,
		_w18743_
	);
	LUT2 #(
		.INIT('h4)
	) name14696 (
		_w18724_,
		_w18743_,
		_w18744_
	);
	LUT2 #(
		.INIT('h2)
	) name14697 (
		_w6143_,
		_w17588_,
		_w18745_
	);
	LUT2 #(
		.INIT('h8)
	) name14698 (
		_w6150_,
		_w17588_,
		_w18746_
	);
	LUT3 #(
		.INIT('h01)
	) name14699 (
		_w17585_,
		_w18746_,
		_w18745_,
		_w18747_
	);
	LUT2 #(
		.INIT('h1)
	) name14700 (
		_w17587_,
		_w18747_,
		_w18748_
	);
	LUT4 #(
		.INIT('hef00)
	) name14701 (
		_w13610_,
		_w13611_,
		_w17585_,
		_w18748_,
		_w18749_
	);
	LUT3 #(
		.INIT('h01)
	) name14702 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w11926_,
		_w17586_,
		_w18750_
	);
	LUT2 #(
		.INIT('h1)
	) name14703 (
		_w17515_,
		_w18750_,
		_w18751_
	);
	LUT2 #(
		.INIT('h4)
	) name14704 (
		_w18749_,
		_w18751_,
		_w18752_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14705 (
		_w17515_,
		_w18722_,
		_w18744_,
		_w18752_,
		_w18753_
	);
	LUT4 #(
		.INIT('h0105)
	) name14706 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w9841_,
		_w12118_,
		_w18754_
	);
	LUT3 #(
		.INIT('h02)
	) name14707 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w12315_,
		_w12316_,
		_w18755_
	);
	LUT4 #(
		.INIT('h007f)
	) name14708 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w12118_,
		_w17520_,
		_w18755_,
		_w18756_
	);
	LUT3 #(
		.INIT('h8a)
	) name14709 (
		_w17517_,
		_w18754_,
		_w18756_,
		_w18757_
	);
	LUT4 #(
		.INIT('hacc0)
	) name14710 (
		_w5914_,
		_w8647_,
		_w17525_,
		_w17526_,
		_w18758_
	);
	LUT3 #(
		.INIT('ha8)
	) name14711 (
		_w17524_,
		_w17527_,
		_w18758_,
		_w18759_
	);
	LUT3 #(
		.INIT('h54)
	) name14712 (
		_w5872_,
		_w17542_,
		_w17543_,
		_w18760_
	);
	LUT3 #(
		.INIT('h54)
	) name14713 (
		_w5865_,
		_w17539_,
		_w17540_,
		_w18761_
	);
	LUT3 #(
		.INIT('h54)
	) name14714 (
		_w5869_,
		_w17545_,
		_w17546_,
		_w18762_
	);
	LUT3 #(
		.INIT('h01)
	) name14715 (
		_w18761_,
		_w18762_,
		_w18760_,
		_w18763_
	);
	LUT2 #(
		.INIT('h8)
	) name14716 (
		_w17538_,
		_w18763_,
		_w18764_
	);
	LUT2 #(
		.INIT('h8)
	) name14717 (
		_w17525_,
		_w18764_,
		_w18765_
	);
	LUT4 #(
		.INIT('h1310)
	) name14718 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w5914_,
		_w16322_,
		_w16504_,
		_w18766_
	);
	LUT3 #(
		.INIT('h04)
	) name14719 (
		_w17524_,
		_w17526_,
		_w18766_,
		_w18767_
	);
	LUT3 #(
		.INIT('he0)
	) name14720 (
		_w11393_,
		_w11589_,
		_w11855_,
		_w18768_
	);
	LUT2 #(
		.INIT('h8)
	) name14721 (
		_w11507_,
		_w11522_,
		_w18769_
	);
	LUT3 #(
		.INIT('he0)
	) name14722 (
		_w11552_,
		_w11474_,
		_w12767_,
		_w18770_
	);
	LUT3 #(
		.INIT('h01)
	) name14723 (
		_w18769_,
		_w18770_,
		_w18768_,
		_w18771_
	);
	LUT3 #(
		.INIT('h80)
	) name14724 (
		_w11900_,
		_w11833_,
		_w18771_,
		_w18772_
	);
	LUT4 #(
		.INIT('h4000)
	) name14725 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11358_,
		_w11382_,
		_w11861_,
		_w18773_
	);
	LUT3 #(
		.INIT('h08)
	) name14726 (
		_w11386_,
		_w11415_,
		_w11506_,
		_w18774_
	);
	LUT4 #(
		.INIT('h0001)
	) name14727 (
		_w11570_,
		_w17964_,
		_w18773_,
		_w18774_,
		_w18775_
	);
	LUT3 #(
		.INIT('h80)
	) name14728 (
		_w11401_,
		_w11389_,
		_w11864_,
		_w18776_
	);
	LUT4 #(
		.INIT('h777f)
	) name14729 (
		_w11389_,
		_w11445_,
		_w11848_,
		_w11875_,
		_w18777_
	);
	LUT2 #(
		.INIT('h4)
	) name14730 (
		_w18776_,
		_w18777_,
		_w18778_
	);
	LUT4 #(
		.INIT('ha820)
	) name14731 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001 ,
		_w18779_
	);
	LUT3 #(
		.INIT('h07)
	) name14732 (
		_w11578_,
		_w12504_,
		_w18779_,
		_w18780_
	);
	LUT3 #(
		.INIT('h08)
	) name14733 (
		_w11389_,
		_w11476_,
		_w11950_,
		_w18781_
	);
	LUT2 #(
		.INIT('h8)
	) name14734 (
		_w11429_,
		_w11861_,
		_w18782_
	);
	LUT3 #(
		.INIT('h10)
	) name14735 (
		_w18781_,
		_w18782_,
		_w18780_,
		_w18783_
	);
	LUT3 #(
		.INIT('h80)
	) name14736 (
		_w18778_,
		_w18783_,
		_w18775_,
		_w18784_
	);
	LUT2 #(
		.INIT('h8)
	) name14737 (
		_w17821_,
		_w17959_,
		_w18785_
	);
	LUT4 #(
		.INIT('h135f)
	) name14738 (
		_w11588_,
		_w11435_,
		_w11469_,
		_w11874_,
		_w18786_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name14739 (
		_w11558_,
		_w11530_,
		_w11449_,
		_w11844_,
		_w18787_
	);
	LUT4 #(
		.INIT('h0111)
	) name14740 (
		_w11550_,
		_w11551_,
		_w11587_,
		_w11465_,
		_w18788_
	);
	LUT4 #(
		.INIT('h7707)
	) name14741 (
		_w11499_,
		_w11973_,
		_w11962_,
		_w11953_,
		_w18789_
	);
	LUT4 #(
		.INIT('h8000)
	) name14742 (
		_w18788_,
		_w18789_,
		_w18786_,
		_w18787_,
		_w18790_
	);
	LUT3 #(
		.INIT('h80)
	) name14743 (
		_w18784_,
		_w18785_,
		_w18790_,
		_w18791_
	);
	LUT3 #(
		.INIT('hc8)
	) name14744 (
		_w11409_,
		_w11458_,
		_w11896_,
		_w18792_
	);
	LUT4 #(
		.INIT('h4440)
	) name14745 (
		_w11536_,
		_w11386_,
		_w11393_,
		_w11589_,
		_w18793_
	);
	LUT3 #(
		.INIT('hc8)
	) name14746 (
		_w11555_,
		_w11872_,
		_w11888_,
		_w18794_
	);
	LUT3 #(
		.INIT('h20)
	) name14747 (
		_w11473_,
		_w11444_,
		_w11863_,
		_w18795_
	);
	LUT3 #(
		.INIT('h54)
	) name14748 (
		_w11385_,
		_w11475_,
		_w18795_,
		_w18796_
	);
	LUT4 #(
		.INIT('h0001)
	) name14749 (
		_w18792_,
		_w18793_,
		_w18794_,
		_w18796_,
		_w18797_
	);
	LUT2 #(
		.INIT('h8)
	) name14750 (
		_w17956_,
		_w18797_,
		_w18798_
	);
	LUT4 #(
		.INIT('h8000)
	) name14751 (
		_w12630_,
		_w18772_,
		_w18791_,
		_w18798_,
		_w18799_
	);
	LUT2 #(
		.INIT('h2)
	) name14752 (
		_w17556_,
		_w18799_,
		_w18800_
	);
	LUT3 #(
		.INIT('h80)
	) name14753 (
		_w5914_,
		_w17563_,
		_w17566_,
		_w18801_
	);
	LUT3 #(
		.INIT('h54)
	) name14754 (
		_w5901_,
		_w17558_,
		_w17559_,
		_w18802_
	);
	LUT2 #(
		.INIT('h1)
	) name14755 (
		_w18801_,
		_w18802_,
		_w18803_
	);
	LUT3 #(
		.INIT('h80)
	) name14756 (
		_w8647_,
		_w17563_,
		_w17564_,
		_w18804_
	);
	LUT3 #(
		.INIT('h0b)
	) name14757 (
		_w12779_,
		_w17569_,
		_w18804_,
		_w18805_
	);
	LUT4 #(
		.INIT('h3230)
	) name14758 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w5891_,
		_w17571_,
		_w17572_,
		_w18806_
	);
	LUT4 #(
		.INIT('h3310)
	) name14759 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w5887_,
		_w17572_,
		_w17575_,
		_w18807_
	);
	LUT2 #(
		.INIT('h1)
	) name14760 (
		_w18806_,
		_w18807_,
		_w18808_
	);
	LUT3 #(
		.INIT('h80)
	) name14761 (
		_w18803_,
		_w18805_,
		_w18808_,
		_w18809_
	);
	LUT2 #(
		.INIT('h4)
	) name14762 (
		_w18800_,
		_w18809_,
		_w18810_
	);
	LUT3 #(
		.INIT('hb0)
	) name14763 (
		_w18765_,
		_w18767_,
		_w18810_,
		_w18811_
	);
	LUT2 #(
		.INIT('h4)
	) name14764 (
		_w18759_,
		_w18811_,
		_w18812_
	);
	LUT2 #(
		.INIT('h2)
	) name14765 (
		_w5876_,
		_w17588_,
		_w18813_
	);
	LUT2 #(
		.INIT('h8)
	) name14766 (
		_w5867_,
		_w17588_,
		_w18814_
	);
	LUT3 #(
		.INIT('h01)
	) name14767 (
		_w17585_,
		_w18814_,
		_w18813_,
		_w18815_
	);
	LUT2 #(
		.INIT('h1)
	) name14768 (
		_w17587_,
		_w18815_,
		_w18816_
	);
	LUT4 #(
		.INIT('hef00)
	) name14769 (
		_w12315_,
		_w12316_,
		_w17585_,
		_w18816_,
		_w18817_
	);
	LUT3 #(
		.INIT('h01)
	) name14770 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w11926_,
		_w17586_,
		_w18818_
	);
	LUT2 #(
		.INIT('h1)
	) name14771 (
		_w17515_,
		_w18818_,
		_w18819_
	);
	LUT2 #(
		.INIT('h4)
	) name14772 (
		_w18817_,
		_w18819_,
		_w18820_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14773 (
		_w17515_,
		_w18757_,
		_w18812_,
		_w18820_,
		_w18821_
	);
	LUT4 #(
		.INIT('h4500)
	) name14774 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w17630_,
		_w18822_
	);
	LUT3 #(
		.INIT('h02)
	) name14775 (
		_w8647_,
		_w17630_,
		_w17633_,
		_w18823_
	);
	LUT3 #(
		.INIT('he4)
	) name14776 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001 ,
		_w18824_
	);
	LUT3 #(
		.INIT('h40)
	) name14777 (
		_w17617_,
		_w17635_,
		_w18824_,
		_w18825_
	);
	LUT3 #(
		.INIT('h53)
	) name14778 (
		_w5874_,
		_w5878_,
		_w17618_,
		_w18826_
	);
	LUT3 #(
		.INIT('h80)
	) name14779 (
		_w17617_,
		_w17635_,
		_w18826_,
		_w18827_
	);
	LUT3 #(
		.INIT('h80)
	) name14780 (
		_w17514_,
		_w17628_,
		_w18815_,
		_w18828_
	);
	LUT3 #(
		.INIT('h01)
	) name14781 (
		_w18827_,
		_w18828_,
		_w18825_,
		_w18829_
	);
	LUT2 #(
		.INIT('h4)
	) name14782 (
		_w18823_,
		_w18829_,
		_w18830_
	);
	LUT3 #(
		.INIT('ha8)
	) name14783 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		_w17511_,
		_w17512_,
		_w18831_
	);
	LUT4 #(
		.INIT('h00ba)
	) name14784 (
		_w17511_,
		_w18822_,
		_w18830_,
		_w18831_,
		_w18832_
	);
	LUT2 #(
		.INIT('h1)
	) name14785 (
		_w17627_,
		_w18832_,
		_w18833_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14786 (
		_w17627_,
		_w18757_,
		_w18812_,
		_w18833_,
		_w18834_
	);
	LUT4 #(
		.INIT('h4500)
	) name14787 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w17630_,
		_w18835_
	);
	LUT3 #(
		.INIT('h02)
	) name14788 (
		_w8885_,
		_w17630_,
		_w17633_,
		_w18836_
	);
	LUT3 #(
		.INIT('he4)
	) name14789 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[3]/P0001 ,
		_w18837_
	);
	LUT3 #(
		.INIT('h40)
	) name14790 (
		_w17617_,
		_w17635_,
		_w18837_,
		_w18838_
	);
	LUT3 #(
		.INIT('h35)
	) name14791 (
		_w6152_,
		_w6154_,
		_w17618_,
		_w18839_
	);
	LUT3 #(
		.INIT('h80)
	) name14792 (
		_w17617_,
		_w17635_,
		_w18839_,
		_w18840_
	);
	LUT3 #(
		.INIT('h80)
	) name14793 (
		_w17514_,
		_w17628_,
		_w18747_,
		_w18841_
	);
	LUT3 #(
		.INIT('h01)
	) name14794 (
		_w18840_,
		_w18841_,
		_w18838_,
		_w18842_
	);
	LUT2 #(
		.INIT('h4)
	) name14795 (
		_w18836_,
		_w18842_,
		_w18843_
	);
	LUT3 #(
		.INIT('ha8)
	) name14796 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w17511_,
		_w17512_,
		_w18844_
	);
	LUT4 #(
		.INIT('h00ba)
	) name14797 (
		_w17511_,
		_w18835_,
		_w18843_,
		_w18844_,
		_w18845_
	);
	LUT2 #(
		.INIT('h1)
	) name14798 (
		_w17627_,
		_w18845_,
		_w18846_
	);
	LUT4 #(
		.INIT('hff8a)
	) name14799 (
		_w17627_,
		_w18722_,
		_w18744_,
		_w18846_,
		_w18847_
	);
	LUT4 #(
		.INIT('hab00)
	) name14800 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w11305_,
		_w17501_,
		_w18848_
	);
	LUT4 #(
		.INIT('h5455)
	) name14801 (
		_w12224_,
		_w12560_,
		_w12561_,
		_w18848_,
		_w18849_
	);
	LUT4 #(
		.INIT('haa8a)
	) name14802 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 ,
		_w11632_,
		_w17503_,
		_w17504_,
		_w18850_
	);
	LUT4 #(
		.INIT('h5504)
	) name14803 (
		_w11624_,
		_w17503_,
		_w18849_,
		_w18850_,
		_w18851_
	);
	LUT4 #(
		.INIT('h4c08)
	) name14804 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w14365_,
		_w14367_,
		_w18852_
	);
	LUT2 #(
		.INIT('he)
	) name14805 (
		_w18851_,
		_w18852_,
		_w18853_
	);
	LUT4 #(
		.INIT('h0400)
	) name14806 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[1]/NET0131 ,
		_w18854_
	);
	LUT3 #(
		.INIT('h01)
	) name14807 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TCR_TMP_reg[0]/NET0131 ,
		_w14107_,
		_w18855_
	);
	LUT4 #(
		.INIT('h0001)
	) name14808 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TCR_TMP_reg[0]/NET0131 ,
		\tm_TCR_TMP_reg[1]/NET0131 ,
		_w14107_,
		_w18856_
	);
	LUT4 #(
		.INIT('h2333)
	) name14809 (
		\tm_tpr_reg_DO_reg[1]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w18857_
	);
	LUT4 #(
		.INIT('hde00)
	) name14810 (
		\tm_TCR_TMP_reg[1]/NET0131 ,
		_w14103_,
		_w18855_,
		_w18857_,
		_w18858_
	);
	LUT2 #(
		.INIT('he)
	) name14811 (
		_w18854_,
		_w18858_,
		_w18859_
	);
	LUT4 #(
		.INIT('h0400)
	) name14812 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[2]/NET0131 ,
		_w18860_
	);
	LUT4 #(
		.INIT('h2333)
	) name14813 (
		\tm_tpr_reg_DO_reg[2]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w18861_
	);
	LUT4 #(
		.INIT('hde00)
	) name14814 (
		\tm_TCR_TMP_reg[2]/NET0131 ,
		_w14103_,
		_w18856_,
		_w18861_,
		_w18862_
	);
	LUT2 #(
		.INIT('he)
	) name14815 (
		_w18860_,
		_w18862_,
		_w18863_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name14816 (
		\tm_TCR_TMP_reg[6]/NET0131 ,
		\tm_tpr_reg_DO_reg[6]/NET0131 ,
		_w14103_,
		_w17151_,
		_w18864_
	);
	LUT3 #(
		.INIT('hb8)
	) name14817 (
		\tm_tcr_reg_DO_reg[6]/NET0131 ,
		_w12803_,
		_w18864_,
		_w18865_
	);
	LUT4 #(
		.INIT('h0400)
	) name14818 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[5]/NET0131 ,
		_w18866_
	);
	LUT3 #(
		.INIT('hc9)
	) name14819 (
		\T_TMODE[0]_pad ,
		\tm_TCR_TMP_reg[4]/NET0131 ,
		_w12797_,
		_w18867_
	);
	LUT3 #(
		.INIT('h01)
	) name14820 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w14107_,
		_w18867_,
		_w18868_
	);
	LUT4 #(
		.INIT('hccc8)
	) name14821 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TCR_TMP_reg[5]/NET0131 ,
		_w14107_,
		_w18867_,
		_w18869_
	);
	LUT4 #(
		.INIT('hfcbd)
	) name14822 (
		\T_TMODE[0]_pad ,
		\tm_TCR_TMP_reg[4]/NET0131 ,
		\tm_TCR_TMP_reg[5]/NET0131 ,
		_w12797_,
		_w18870_
	);
	LUT3 #(
		.INIT('h01)
	) name14823 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w14107_,
		_w18870_,
		_w18871_
	);
	LUT4 #(
		.INIT('h2333)
	) name14824 (
		\tm_tpr_reg_DO_reg[5]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w18872_
	);
	LUT4 #(
		.INIT('hfe00)
	) name14825 (
		_w14103_,
		_w18871_,
		_w18869_,
		_w18872_,
		_w18873_
	);
	LUT2 #(
		.INIT('he)
	) name14826 (
		_w18866_,
		_w18873_,
		_w18874_
	);
	LUT3 #(
		.INIT('h04)
	) name14827 (
		\sport1_cfg_RFSg_d1_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w18875_
	);
	LUT4 #(
		.INIT('h3500)
	) name14828 (
		\sport1_cfg_RFSg_d2_reg/NET0131 ,
		\sport1_cfg_RFSg_d3_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w18876_
	);
	LUT2 #(
		.INIT('h1)
	) name14829 (
		_w18875_,
		_w18876_,
		_w18877_
	);
	LUT4 #(
		.INIT('h8f00)
	) name14830 (
		_w13425_,
		_w13426_,
		_w14257_,
		_w18877_,
		_w18878_
	);
	LUT4 #(
		.INIT('h0001)
	) name14831 (
		\sport1_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[1]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[2]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[3]/NET0131 ,
		_w18879_
	);
	LUT2 #(
		.INIT('h4)
	) name14832 (
		\sport1_rxctl_LMcnt_reg[4]/NET0131 ,
		_w18879_,
		_w18880_
	);
	LUT3 #(
		.INIT('h0d)
	) name14833 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		_w18878_,
		_w18880_,
		_w18881_
	);
	LUT4 #(
		.INIT('h00c4)
	) name14834 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[0]/P0001 ,
		_w18878_,
		_w18880_,
		_w18882_
	);
	LUT3 #(
		.INIT('he0)
	) name14835 (
		\sport1_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport1_rxctl_sht2nd_reg/P0001 ,
		_w18883_
	);
	LUT2 #(
		.INIT('h8)
	) name14836 (
		_w18882_,
		_w18883_,
		_w18884_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14837 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[15]/P0001 ,
		_w18878_,
		_w18880_,
		_w18885_
	);
	LUT4 #(
		.INIT('h0031)
	) name14838 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_sht2nd_reg/P0001 ,
		_w18878_,
		_w18880_,
		_w18886_
	);
	LUT3 #(
		.INIT('h13)
	) name14839 (
		\sport1_rxctl_RXSHT_reg[14]/P0001 ,
		_w18885_,
		_w18886_,
		_w18887_
	);
	LUT2 #(
		.INIT('hb)
	) name14840 (
		_w18884_,
		_w18887_,
		_w18888_
	);
	LUT3 #(
		.INIT('h04)
	) name14841 (
		\sport0_cfg_RFSg_d1_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w18889_
	);
	LUT4 #(
		.INIT('h3500)
	) name14842 (
		\sport0_cfg_RFSg_d2_reg/NET0131 ,
		\sport0_cfg_RFSg_d3_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w18890_
	);
	LUT2 #(
		.INIT('h1)
	) name14843 (
		_w18889_,
		_w18890_,
		_w18891_
	);
	LUT4 #(
		.INIT('hd500)
	) name14844 (
		_w12540_,
		_w13428_,
		_w13429_,
		_w18891_,
		_w18892_
	);
	LUT4 #(
		.INIT('h0001)
	) name14845 (
		\sport0_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[1]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[2]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[3]/NET0131 ,
		_w18893_
	);
	LUT2 #(
		.INIT('h4)
	) name14846 (
		\sport0_rxctl_LMcnt_reg[4]/NET0131 ,
		_w18893_,
		_w18894_
	);
	LUT3 #(
		.INIT('h0d)
	) name14847 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		_w18892_,
		_w18894_,
		_w18895_
	);
	LUT4 #(
		.INIT('h00c4)
	) name14848 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[0]/P0001 ,
		_w18892_,
		_w18894_,
		_w18896_
	);
	LUT3 #(
		.INIT('he0)
	) name14849 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_sht2nd_reg/P0001 ,
		_w18897_
	);
	LUT2 #(
		.INIT('h8)
	) name14850 (
		_w18896_,
		_w18897_,
		_w18898_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14851 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[10]/P0001 ,
		_w18892_,
		_w18894_,
		_w18899_
	);
	LUT4 #(
		.INIT('h0031)
	) name14852 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_sht2nd_reg/P0001 ,
		_w18892_,
		_w18894_,
		_w18900_
	);
	LUT3 #(
		.INIT('h13)
	) name14853 (
		\sport0_rxctl_RXSHT_reg[9]/P0001 ,
		_w18899_,
		_w18900_,
		_w18901_
	);
	LUT2 #(
		.INIT('hb)
	) name14854 (
		_w18898_,
		_w18901_,
		_w18902_
	);
	LUT2 #(
		.INIT('h8)
	) name14855 (
		\sport1_rxctl_RXSHT_reg[9]/P0001 ,
		_w18886_,
		_w18903_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14856 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[10]/P0001 ,
		_w18878_,
		_w18880_,
		_w18904_
	);
	LUT3 #(
		.INIT('h07)
	) name14857 (
		_w18882_,
		_w18883_,
		_w18904_,
		_w18905_
	);
	LUT2 #(
		.INIT('hb)
	) name14858 (
		_w18903_,
		_w18905_,
		_w18906_
	);
	LUT2 #(
		.INIT('h8)
	) name14859 (
		\sport1_rxctl_RXSHT_reg[10]/P0001 ,
		_w18886_,
		_w18907_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14860 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[11]/P0001 ,
		_w18878_,
		_w18880_,
		_w18908_
	);
	LUT3 #(
		.INIT('h07)
	) name14861 (
		_w18882_,
		_w18883_,
		_w18908_,
		_w18909_
	);
	LUT2 #(
		.INIT('hb)
	) name14862 (
		_w18907_,
		_w18909_,
		_w18910_
	);
	LUT4 #(
		.INIT('h084c)
	) name14863 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w14367_,
		_w14391_,
		_w18911_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name14864 (
		_w11626_,
		_w11627_,
		_w12224_,
		_w18848_,
		_w18912_
	);
	LUT4 #(
		.INIT('h44c4)
	) name14865 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001 ,
		_w17500_,
		_w17503_,
		_w17504_,
		_w18913_
	);
	LUT3 #(
		.INIT('hd0)
	) name14866 (
		_w17503_,
		_w18912_,
		_w18913_,
		_w18914_
	);
	LUT2 #(
		.INIT('h1)
	) name14867 (
		_w18911_,
		_w18914_,
		_w18915_
	);
	LUT2 #(
		.INIT('h8)
	) name14868 (
		\sport1_rxctl_RXSHT_reg[11]/P0001 ,
		_w18886_,
		_w18916_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14869 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[12]/P0001 ,
		_w18878_,
		_w18880_,
		_w18917_
	);
	LUT3 #(
		.INIT('h07)
	) name14870 (
		_w18882_,
		_w18883_,
		_w18917_,
		_w18918_
	);
	LUT2 #(
		.INIT('hb)
	) name14871 (
		_w18916_,
		_w18918_,
		_w18919_
	);
	LUT2 #(
		.INIT('h8)
	) name14872 (
		\sport1_rxctl_RXSHT_reg[12]/P0001 ,
		_w18886_,
		_w18920_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14873 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[13]/P0001 ,
		_w18878_,
		_w18880_,
		_w18921_
	);
	LUT3 #(
		.INIT('h07)
	) name14874 (
		_w18882_,
		_w18883_,
		_w18921_,
		_w18922_
	);
	LUT2 #(
		.INIT('hb)
	) name14875 (
		_w18920_,
		_w18922_,
		_w18923_
	);
	LUT2 #(
		.INIT('h8)
	) name14876 (
		\sport1_rxctl_RXSHT_reg[13]/P0001 ,
		_w18886_,
		_w18924_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14877 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[14]/P0001 ,
		_w18878_,
		_w18880_,
		_w18925_
	);
	LUT3 #(
		.INIT('h07)
	) name14878 (
		_w18882_,
		_w18883_,
		_w18925_,
		_w18926_
	);
	LUT2 #(
		.INIT('hb)
	) name14879 (
		_w18924_,
		_w18926_,
		_w18927_
	);
	LUT2 #(
		.INIT('h8)
	) name14880 (
		\sport1_rxctl_RXSHT_reg[1]/P0001 ,
		_w18886_,
		_w18928_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14881 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[2]/P0001 ,
		_w18878_,
		_w18880_,
		_w18929_
	);
	LUT3 #(
		.INIT('h07)
	) name14882 (
		_w18882_,
		_w18883_,
		_w18929_,
		_w18930_
	);
	LUT2 #(
		.INIT('hb)
	) name14883 (
		_w18928_,
		_w18930_,
		_w18931_
	);
	LUT2 #(
		.INIT('h8)
	) name14884 (
		\sport1_rxctl_RXSHT_reg[2]/P0001 ,
		_w18886_,
		_w18932_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14885 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[3]/P0001 ,
		_w18878_,
		_w18880_,
		_w18933_
	);
	LUT3 #(
		.INIT('h07)
	) name14886 (
		_w18882_,
		_w18883_,
		_w18933_,
		_w18934_
	);
	LUT2 #(
		.INIT('hb)
	) name14887 (
		_w18932_,
		_w18934_,
		_w18935_
	);
	LUT2 #(
		.INIT('h8)
	) name14888 (
		\sport1_rxctl_RXSHT_reg[3]/P0001 ,
		_w18886_,
		_w18936_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14889 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[4]/P0001 ,
		_w18878_,
		_w18880_,
		_w18937_
	);
	LUT3 #(
		.INIT('h07)
	) name14890 (
		_w18882_,
		_w18883_,
		_w18937_,
		_w18938_
	);
	LUT2 #(
		.INIT('hb)
	) name14891 (
		_w18936_,
		_w18938_,
		_w18939_
	);
	LUT2 #(
		.INIT('h8)
	) name14892 (
		\sport1_rxctl_RXSHT_reg[4]/P0001 ,
		_w18886_,
		_w18940_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14893 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[5]/P0001 ,
		_w18878_,
		_w18880_,
		_w18941_
	);
	LUT3 #(
		.INIT('h07)
	) name14894 (
		_w18882_,
		_w18883_,
		_w18941_,
		_w18942_
	);
	LUT2 #(
		.INIT('hb)
	) name14895 (
		_w18940_,
		_w18942_,
		_w18943_
	);
	LUT2 #(
		.INIT('h8)
	) name14896 (
		\sport1_rxctl_RXSHT_reg[5]/P0001 ,
		_w18886_,
		_w18944_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14897 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[6]/P0001 ,
		_w18878_,
		_w18880_,
		_w18945_
	);
	LUT3 #(
		.INIT('h07)
	) name14898 (
		_w18882_,
		_w18883_,
		_w18945_,
		_w18946_
	);
	LUT2 #(
		.INIT('hb)
	) name14899 (
		_w18944_,
		_w18946_,
		_w18947_
	);
	LUT2 #(
		.INIT('h8)
	) name14900 (
		\sport1_rxctl_RXSHT_reg[7]/P0001 ,
		_w18886_,
		_w18948_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14901 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[8]/P0001 ,
		_w18878_,
		_w18880_,
		_w18949_
	);
	LUT3 #(
		.INIT('h07)
	) name14902 (
		_w18882_,
		_w18883_,
		_w18949_,
		_w18950_
	);
	LUT2 #(
		.INIT('hb)
	) name14903 (
		_w18948_,
		_w18950_,
		_w18951_
	);
	LUT2 #(
		.INIT('h8)
	) name14904 (
		\sport1_rxctl_RXSHT_reg[8]/P0001 ,
		_w18886_,
		_w18952_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14905 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[9]/P0001 ,
		_w18878_,
		_w18880_,
		_w18953_
	);
	LUT3 #(
		.INIT('h07)
	) name14906 (
		_w18882_,
		_w18883_,
		_w18953_,
		_w18954_
	);
	LUT2 #(
		.INIT('hb)
	) name14907 (
		_w18952_,
		_w18954_,
		_w18955_
	);
	LUT2 #(
		.INIT('h8)
	) name14908 (
		\sport0_rxctl_RXSHT_reg[10]/P0001 ,
		_w18900_,
		_w18956_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14909 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[11]/P0001 ,
		_w18892_,
		_w18894_,
		_w18957_
	);
	LUT3 #(
		.INIT('h07)
	) name14910 (
		_w18896_,
		_w18897_,
		_w18957_,
		_w18958_
	);
	LUT2 #(
		.INIT('hb)
	) name14911 (
		_w18956_,
		_w18958_,
		_w18959_
	);
	LUT2 #(
		.INIT('h8)
	) name14912 (
		\sport0_rxctl_RXSHT_reg[13]/P0001 ,
		_w18900_,
		_w18960_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14913 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[14]/P0001 ,
		_w18892_,
		_w18894_,
		_w18961_
	);
	LUT3 #(
		.INIT('h07)
	) name14914 (
		_w18896_,
		_w18897_,
		_w18961_,
		_w18962_
	);
	LUT2 #(
		.INIT('hb)
	) name14915 (
		_w18960_,
		_w18962_,
		_w18963_
	);
	LUT2 #(
		.INIT('h8)
	) name14916 (
		\sport0_rxctl_RXSHT_reg[14]/P0001 ,
		_w18900_,
		_w18964_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14917 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[15]/P0001 ,
		_w18892_,
		_w18894_,
		_w18965_
	);
	LUT3 #(
		.INIT('h07)
	) name14918 (
		_w18896_,
		_w18897_,
		_w18965_,
		_w18966_
	);
	LUT2 #(
		.INIT('hb)
	) name14919 (
		_w18964_,
		_w18966_,
		_w18967_
	);
	LUT2 #(
		.INIT('h8)
	) name14920 (
		\sport0_rxctl_RXSHT_reg[1]/P0001 ,
		_w18900_,
		_w18968_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14921 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[2]/P0001 ,
		_w18892_,
		_w18894_,
		_w18969_
	);
	LUT3 #(
		.INIT('h07)
	) name14922 (
		_w18896_,
		_w18897_,
		_w18969_,
		_w18970_
	);
	LUT2 #(
		.INIT('hb)
	) name14923 (
		_w18968_,
		_w18970_,
		_w18971_
	);
	LUT2 #(
		.INIT('h8)
	) name14924 (
		\sport0_rxctl_RXSHT_reg[2]/P0001 ,
		_w18900_,
		_w18972_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14925 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[3]/P0001 ,
		_w18892_,
		_w18894_,
		_w18973_
	);
	LUT3 #(
		.INIT('h07)
	) name14926 (
		_w18896_,
		_w18897_,
		_w18973_,
		_w18974_
	);
	LUT2 #(
		.INIT('hb)
	) name14927 (
		_w18972_,
		_w18974_,
		_w18975_
	);
	LUT2 #(
		.INIT('h8)
	) name14928 (
		\sport0_rxctl_RXSHT_reg[3]/P0001 ,
		_w18900_,
		_w18976_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14929 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[4]/P0001 ,
		_w18892_,
		_w18894_,
		_w18977_
	);
	LUT3 #(
		.INIT('h07)
	) name14930 (
		_w18896_,
		_w18897_,
		_w18977_,
		_w18978_
	);
	LUT2 #(
		.INIT('hb)
	) name14931 (
		_w18976_,
		_w18978_,
		_w18979_
	);
	LUT2 #(
		.INIT('h8)
	) name14932 (
		\sport0_rxctl_RXSHT_reg[4]/P0001 ,
		_w18900_,
		_w18980_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14933 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[5]/P0001 ,
		_w18892_,
		_w18894_,
		_w18981_
	);
	LUT3 #(
		.INIT('h07)
	) name14934 (
		_w18896_,
		_w18897_,
		_w18981_,
		_w18982_
	);
	LUT2 #(
		.INIT('hb)
	) name14935 (
		_w18980_,
		_w18982_,
		_w18983_
	);
	LUT2 #(
		.INIT('h8)
	) name14936 (
		\sport0_rxctl_RXSHT_reg[5]/P0001 ,
		_w18900_,
		_w18984_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14937 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[6]/P0001 ,
		_w18892_,
		_w18894_,
		_w18985_
	);
	LUT3 #(
		.INIT('h07)
	) name14938 (
		_w18896_,
		_w18897_,
		_w18985_,
		_w18986_
	);
	LUT2 #(
		.INIT('hb)
	) name14939 (
		_w18984_,
		_w18986_,
		_w18987_
	);
	LUT2 #(
		.INIT('h8)
	) name14940 (
		\sport0_rxctl_RXSHT_reg[6]/P0001 ,
		_w18900_,
		_w18988_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14941 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[7]/P0001 ,
		_w18892_,
		_w18894_,
		_w18989_
	);
	LUT3 #(
		.INIT('h07)
	) name14942 (
		_w18896_,
		_w18897_,
		_w18989_,
		_w18990_
	);
	LUT2 #(
		.INIT('hb)
	) name14943 (
		_w18988_,
		_w18990_,
		_w18991_
	);
	LUT2 #(
		.INIT('h8)
	) name14944 (
		\sport0_rxctl_RXSHT_reg[7]/P0001 ,
		_w18900_,
		_w18992_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14945 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[8]/P0001 ,
		_w18892_,
		_w18894_,
		_w18993_
	);
	LUT3 #(
		.INIT('h07)
	) name14946 (
		_w18896_,
		_w18897_,
		_w18993_,
		_w18994_
	);
	LUT2 #(
		.INIT('hb)
	) name14947 (
		_w18992_,
		_w18994_,
		_w18995_
	);
	LUT2 #(
		.INIT('h8)
	) name14948 (
		\sport0_rxctl_RXSHT_reg[8]/P0001 ,
		_w18900_,
		_w18996_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14949 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[9]/P0001 ,
		_w18892_,
		_w18894_,
		_w18997_
	);
	LUT3 #(
		.INIT('h07)
	) name14950 (
		_w18896_,
		_w18897_,
		_w18997_,
		_w18998_
	);
	LUT2 #(
		.INIT('hb)
	) name14951 (
		_w18996_,
		_w18998_,
		_w18999_
	);
	LUT2 #(
		.INIT('h8)
	) name14952 (
		\sport1_rxctl_RXSHT_reg[6]/P0001 ,
		_w18886_,
		_w19000_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14953 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[7]/P0001 ,
		_w18878_,
		_w18880_,
		_w19001_
	);
	LUT3 #(
		.INIT('h07)
	) name14954 (
		_w18882_,
		_w18883_,
		_w19001_,
		_w19002_
	);
	LUT2 #(
		.INIT('hb)
	) name14955 (
		_w19000_,
		_w19002_,
		_w19003_
	);
	LUT2 #(
		.INIT('h8)
	) name14956 (
		\sport0_rxctl_RXSHT_reg[12]/P0001 ,
		_w18900_,
		_w19004_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14957 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[13]/P0001 ,
		_w18892_,
		_w18894_,
		_w19005_
	);
	LUT3 #(
		.INIT('h07)
	) name14958 (
		_w18896_,
		_w18897_,
		_w19005_,
		_w19006_
	);
	LUT2 #(
		.INIT('hb)
	) name14959 (
		_w19004_,
		_w19006_,
		_w19007_
	);
	LUT2 #(
		.INIT('h8)
	) name14960 (
		\sport0_rxctl_RXSHT_reg[11]/P0001 ,
		_w18900_,
		_w19008_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14961 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[12]/P0001 ,
		_w18892_,
		_w18894_,
		_w19009_
	);
	LUT3 #(
		.INIT('h07)
	) name14962 (
		_w18896_,
		_w18897_,
		_w19009_,
		_w19010_
	);
	LUT2 #(
		.INIT('hb)
	) name14963 (
		_w19008_,
		_w19010_,
		_w19011_
	);
	LUT3 #(
		.INIT('h8c)
	) name14964 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w4142_,
		_w12114_,
		_w19012_
	);
	LUT4 #(
		.INIT('hef00)
	) name14965 (
		_w12114_,
		_w12121_,
		_w12134_,
		_w19012_,
		_w19013_
	);
	LUT2 #(
		.INIT('h8)
	) name14966 (
		_w11301_,
		_w11307_,
		_w19014_
	);
	LUT4 #(
		.INIT('h5455)
	) name14967 (
		_w11320_,
		_w12560_,
		_w12561_,
		_w19014_,
		_w19015_
	);
	LUT4 #(
		.INIT('haaa2)
	) name14968 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 ,
		_w11309_,
		_w11311_,
		_w11323_,
		_w19016_
	);
	LUT4 #(
		.INIT('h5504)
	) name14969 (
		_w9946_,
		_w11309_,
		_w19015_,
		_w19016_,
		_w19017_
	);
	LUT4 #(
		.INIT('h4c08)
	) name14970 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w14365_,
		_w14367_,
		_w19018_
	);
	LUT2 #(
		.INIT('he)
	) name14971 (
		_w19017_,
		_w19018_,
		_w19019_
	);
	LUT4 #(
		.INIT('h0400)
	) name14972 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[13]/NET0131 ,
		_w19020_
	);
	LUT4 #(
		.INIT('h2333)
	) name14973 (
		\tm_tpr_reg_DO_reg[13]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w19021_
	);
	LUT4 #(
		.INIT('hde00)
	) name14974 (
		\tm_TCR_TMP_reg[13]/NET0131 ,
		_w14103_,
		_w15996_,
		_w19021_,
		_w19022_
	);
	LUT2 #(
		.INIT('he)
	) name14975 (
		_w19020_,
		_w19022_,
		_w19023_
	);
	LUT4 #(
		.INIT('h084c)
	) name14976 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w14367_,
		_w14391_,
		_w19024_
	);
	LUT3 #(
		.INIT('h13)
	) name14977 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001 ,
		_w11300_,
		_w19025_
	);
	LUT4 #(
		.INIT('hccc8)
	) name14978 (
		_w11310_,
		_w11312_,
		_w11626_,
		_w11627_,
		_w19026_
	);
	LUT4 #(
		.INIT('h2322)
	) name14979 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001 ,
		_w11303_,
		_w11308_,
		_w19027_
	);
	LUT4 #(
		.INIT('h00ab)
	) name14980 (
		_w11320_,
		_w19025_,
		_w19026_,
		_w19027_,
		_w19028_
	);
	LUT2 #(
		.INIT('h2)
	) name14981 (
		_w11325_,
		_w19028_,
		_w19029_
	);
	LUT2 #(
		.INIT('h1)
	) name14982 (
		_w19024_,
		_w19029_,
		_w19030_
	);
	LUT4 #(
		.INIT('h2000)
	) name14983 (
		\core_c_dec_pMFMAC_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19031_
	);
	LUT4 #(
		.INIT('h00bf)
	) name14984 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w12389_,
		_w19032_
	);
	LUT2 #(
		.INIT('h4)
	) name14985 (
		_w5045_,
		_w5564_,
		_w19033_
	);
	LUT3 #(
		.INIT('h80)
	) name14986 (
		_w5027_,
		_w5028_,
		_w12392_,
		_w19034_
	);
	LUT4 #(
		.INIT('h0080)
	) name14987 (
		_w5027_,
		_w5028_,
		_w12392_,
		_w16302_,
		_w19035_
	);
	LUT2 #(
		.INIT('h1)
	) name14988 (
		_w19033_,
		_w19035_,
		_w19036_
	);
	LUT3 #(
		.INIT('h80)
	) name14989 (
		_w5027_,
		_w5028_,
		_w13333_,
		_w19037_
	);
	LUT3 #(
		.INIT('h07)
	) name14990 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w9323_,
		_w11918_,
		_w19038_
	);
	LUT3 #(
		.INIT('h10)
	) name14991 (
		_w15324_,
		_w19037_,
		_w19038_,
		_w19039_
	);
	LUT4 #(
		.INIT('h007f)
	) name14992 (
		_w5027_,
		_w5028_,
		_w12392_,
		_w15325_,
		_w19040_
	);
	LUT3 #(
		.INIT('h40)
	) name14993 (
		_w5026_,
		_w5045_,
		_w5046_,
		_w19041_
	);
	LUT4 #(
		.INIT('h2000)
	) name14994 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w5026_,
		_w5045_,
		_w5046_,
		_w19042_
	);
	LUT2 #(
		.INIT('h2)
	) name14995 (
		_w19040_,
		_w19042_,
		_w19043_
	);
	LUT3 #(
		.INIT('h80)
	) name14996 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w5027_,
		_w5028_,
		_w19044_
	);
	LUT4 #(
		.INIT('hff37)
	) name14997 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w19045_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14998 (
		_w5028_,
		_w5045_,
		_w15564_,
		_w19045_,
		_w19046_
	);
	LUT4 #(
		.INIT('h5355)
	) name14999 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w19044_,
		_w19046_,
		_w19047_
	);
	LUT3 #(
		.INIT('h70)
	) name15000 (
		_w19039_,
		_w19043_,
		_w19047_,
		_w19048_
	);
	LUT4 #(
		.INIT('h7000)
	) name15001 (
		_w19039_,
		_w19043_,
		_w19047_,
		_w19036_,
		_w19049_
	);
	LUT4 #(
		.INIT('h5355)
	) name15002 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w19044_,
		_w19046_,
		_w19050_
	);
	LUT4 #(
		.INIT('h5355)
	) name15003 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w19044_,
		_w19046_,
		_w19051_
	);
	LUT4 #(
		.INIT('h5355)
	) name15004 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w19044_,
		_w19046_,
		_w19052_
	);
	LUT2 #(
		.INIT('h4)
	) name15005 (
		_w19051_,
		_w19052_,
		_w19053_
	);
	LUT3 #(
		.INIT('h04)
	) name15006 (
		_w19051_,
		_w19052_,
		_w19050_,
		_w19054_
	);
	LUT2 #(
		.INIT('h8)
	) name15007 (
		_w19049_,
		_w19054_,
		_w19055_
	);
	LUT3 #(
		.INIT('h07)
	) name15008 (
		_w19039_,
		_w19043_,
		_w19047_,
		_w19056_
	);
	LUT4 #(
		.INIT('h0700)
	) name15009 (
		_w19039_,
		_w19043_,
		_w19047_,
		_w19036_,
		_w19057_
	);
	LUT2 #(
		.INIT('h2)
	) name15010 (
		_w19051_,
		_w19052_,
		_w19058_
	);
	LUT3 #(
		.INIT('h08)
	) name15011 (
		_w19036_,
		_w19051_,
		_w19052_,
		_w19059_
	);
	LUT3 #(
		.INIT('h70)
	) name15012 (
		_w19039_,
		_w19043_,
		_w19050_,
		_w19060_
	);
	LUT4 #(
		.INIT('h153f)
	) name15013 (
		_w19059_,
		_w19057_,
		_w19054_,
		_w19060_,
		_w19061_
	);
	LUT2 #(
		.INIT('h4)
	) name15014 (
		_w19055_,
		_w19061_,
		_w19062_
	);
	LUT2 #(
		.INIT('h1)
	) name15015 (
		_w19051_,
		_w19052_,
		_w19063_
	);
	LUT3 #(
		.INIT('h80)
	) name15016 (
		_w19050_,
		_w19063_,
		_w19049_,
		_w19064_
	);
	LUT4 #(
		.INIT('h0008)
	) name15017 (
		_w19036_,
		_w19051_,
		_w19052_,
		_w19050_,
		_w19065_
	);
	LUT2 #(
		.INIT('h8)
	) name15018 (
		_w19056_,
		_w19065_,
		_w19066_
	);
	LUT3 #(
		.INIT('h80)
	) name15019 (
		_w19050_,
		_w19063_,
		_w19057_,
		_w19067_
	);
	LUT3 #(
		.INIT('h01)
	) name15020 (
		_w19066_,
		_w19067_,
		_w19064_,
		_w19068_
	);
	LUT4 #(
		.INIT('haeee)
	) name15021 (
		_w19031_,
		_w19032_,
		_w19062_,
		_w19068_,
		_w19069_
	);
	LUT4 #(
		.INIT('h2000)
	) name15022 (
		\core_c_dec_MFMAC_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19070_
	);
	LUT4 #(
		.INIT('hff2a)
	) name15023 (
		_w15539_,
		_w19062_,
		_w19068_,
		_w19070_,
		_w19071_
	);
	LUT3 #(
		.INIT('h40)
	) name15024 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w19072_
	);
	LUT4 #(
		.INIT('hff48)
	) name15025 (
		\sport1_cfg_FSi_cnt_reg[11]/NET0131 ,
		_w17698_,
		_w17671_,
		_w19072_,
		_w19073_
	);
	LUT3 #(
		.INIT('h40)
	) name15026 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w19074_
	);
	LUT4 #(
		.INIT('hff48)
	) name15027 (
		\sport0_cfg_FSi_cnt_reg[11]/NET0131 ,
		_w17734_,
		_w17707_,
		_w19074_,
		_w19075_
	);
	LUT4 #(
		.INIT('h0400)
	) name15028 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[0]/NET0131 ,
		_w19076_
	);
	LUT4 #(
		.INIT('h2333)
	) name15029 (
		\tm_tpr_reg_DO_reg[0]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w19077_
	);
	LUT4 #(
		.INIT('hde00)
	) name15030 (
		\tm_TCR_TMP_reg[0]/NET0131 ,
		_w14103_,
		_w14108_,
		_w19077_,
		_w19078_
	);
	LUT2 #(
		.INIT('he)
	) name15031 (
		_w19076_,
		_w19078_,
		_w19079_
	);
	LUT4 #(
		.INIT('h0400)
	) name15032 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[3]/NET0131 ,
		_w19080_
	);
	LUT3 #(
		.INIT('h8c)
	) name15033 (
		\tm_TCR_TMP_reg[2]/NET0131 ,
		\tm_TCR_TMP_reg[3]/NET0131 ,
		_w18856_,
		_w19081_
	);
	LUT4 #(
		.INIT('h0010)
	) name15034 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TCR_TMP_reg[0]/NET0131 ,
		_w12796_,
		_w14107_,
		_w19082_
	);
	LUT2 #(
		.INIT('h1)
	) name15035 (
		_w14103_,
		_w19082_,
		_w19083_
	);
	LUT4 #(
		.INIT('h2333)
	) name15036 (
		\tm_tpr_reg_DO_reg[3]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w19084_
	);
	LUT4 #(
		.INIT('hefaa)
	) name15037 (
		_w19080_,
		_w19081_,
		_w19083_,
		_w19084_,
		_w19085_
	);
	LUT4 #(
		.INIT('h0400)
	) name15038 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[4]/NET0131 ,
		_w19086_
	);
	LUT3 #(
		.INIT('hc8)
	) name15039 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TCR_TMP_reg[4]/NET0131 ,
		_w14107_,
		_w19087_
	);
	LUT4 #(
		.INIT('h2333)
	) name15040 (
		\tm_tpr_reg_DO_reg[4]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w19088_
	);
	LUT4 #(
		.INIT('hfe00)
	) name15041 (
		_w14103_,
		_w18868_,
		_w19087_,
		_w19088_,
		_w19089_
	);
	LUT2 #(
		.INIT('he)
	) name15042 (
		_w19086_,
		_w19089_,
		_w19090_
	);
	LUT4 #(
		.INIT('h0008)
	) name15043 (
		_w13136_,
		_w13140_,
		_w13148_,
		_w13153_,
		_w19091_
	);
	LUT4 #(
		.INIT('ha851)
	) name15044 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w19092_
	);
	LUT2 #(
		.INIT('h2)
	) name15045 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w19092_,
		_w19093_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15046 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13103_,
		_w13100_,
		_w13101_,
		_w19094_
	);
	LUT2 #(
		.INIT('h4)
	) name15047 (
		_w19093_,
		_w19094_,
		_w19095_
	);
	LUT4 #(
		.INIT('h41cb)
	) name15048 (
		_w13098_,
		_w13147_,
		_w13152_,
		_w19095_,
		_w19096_
	);
	LUT3 #(
		.INIT('h21)
	) name15049 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w19097_
	);
	LUT4 #(
		.INIT('h0021)
	) name15050 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w19098_
	);
	LUT4 #(
		.INIT('h5540)
	) name15051 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w19091_,
		_w19096_,
		_w19098_,
		_w19099_
	);
	LUT4 #(
		.INIT('h0001)
	) name15052 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w19100_
	);
	LUT4 #(
		.INIT('hea00)
	) name15053 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w19091_,
		_w19096_,
		_w19100_,
		_w19101_
	);
	LUT4 #(
		.INIT('h0a08)
	) name15054 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w19101_,
		_w19099_,
		_w19102_
	);
	LUT3 #(
		.INIT('he0)
	) name15055 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[12]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w19103_
	);
	LUT2 #(
		.INIT('h4)
	) name15056 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13161_,
		_w19104_
	);
	LUT2 #(
		.INIT('h8)
	) name15057 (
		_w6758_,
		_w19104_,
		_w19105_
	);
	LUT4 #(
		.INIT('h5510)
	) name15058 (
		_w13158_,
		_w19102_,
		_w19103_,
		_w19105_,
		_w19106_
	);
	LUT4 #(
		.INIT('h0002)
	) name15059 (
		\sport0_rxctl_RX_reg[12]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w19107_
	);
	LUT3 #(
		.INIT('h08)
	) name15060 (
		\sport0_rxctl_RXSHT_reg[12]/P0001 ,
		\sport0_rxctl_a_sync1_reg/P0001 ,
		\sport0_rxctl_a_sync2_reg/P0001 ,
		_w19108_
	);
	LUT2 #(
		.INIT('h1)
	) name15061 (
		_w19107_,
		_w19108_,
		_w19109_
	);
	LUT2 #(
		.INIT('hb)
	) name15062 (
		_w19106_,
		_w19109_,
		_w19110_
	);
	LUT2 #(
		.INIT('h1)
	) name15063 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_dec_updAR_E_reg/P0001 ,
		_w19111_
	);
	LUT3 #(
		.INIT('h04)
	) name15064 (
		_w9453_,
		_w9894_,
		_w19111_,
		_w19112_
	);
	LUT4 #(
		.INIT('h8d00)
	) name15065 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w11318_,
		_w17925_,
		_w19112_,
		_w19113_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15066 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001 ,
		_w9453_,
		_w9894_,
		_w19111_,
		_w19114_
	);
	LUT2 #(
		.INIT('he)
	) name15067 (
		_w19113_,
		_w19114_,
		_w19115_
	);
	LUT4 #(
		.INIT('h00e0)
	) name15068 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w19116_
	);
	LUT3 #(
		.INIT('h07)
	) name15069 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w9931_,
		_w19116_,
		_w19117_
	);
	LUT4 #(
		.INIT('h5355)
	) name15070 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w15565_,
		_w19117_,
		_w19118_
	);
	LUT4 #(
		.INIT('h5355)
	) name15071 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w15565_,
		_w19117_,
		_w19119_
	);
	LUT2 #(
		.INIT('h1)
	) name15072 (
		_w19118_,
		_w19119_,
		_w19120_
	);
	LUT3 #(
		.INIT('h54)
	) name15073 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w15565_,
		_w19041_,
		_w19121_
	);
	LUT4 #(
		.INIT('hffd7)
	) name15074 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w19122_
	);
	LUT3 #(
		.INIT('hb0)
	) name15075 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w9323_,
		_w19122_,
		_w19123_
	);
	LUT3 #(
		.INIT('h13)
	) name15076 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w8177_,
		_w9931_,
		_w19124_
	);
	LUT4 #(
		.INIT('h1000)
	) name15077 (
		_w8176_,
		_w19044_,
		_w19124_,
		_w19123_,
		_w19125_
	);
	LUT4 #(
		.INIT('h8000)
	) name15078 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19126_
	);
	LUT4 #(
		.INIT('h8000)
	) name15079 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19127_
	);
	LUT4 #(
		.INIT('h131f)
	) name15080 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w5564_,
		_w9931_,
		_w19128_
	);
	LUT3 #(
		.INIT('h10)
	) name15081 (
		_w19127_,
		_w19126_,
		_w19128_,
		_w19129_
	);
	LUT4 #(
		.INIT('h5355)
	) name15082 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w15565_,
		_w19117_,
		_w19130_
	);
	LUT4 #(
		.INIT('h00b0)
	) name15083 (
		_w19121_,
		_w19125_,
		_w19129_,
		_w19130_,
		_w19131_
	);
	LUT4 #(
		.INIT('h5355)
	) name15084 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w15565_,
		_w19117_,
		_w19132_
	);
	LUT4 #(
		.INIT('h0800)
	) name15085 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w19133_
	);
	LUT4 #(
		.INIT('h00bf)
	) name15086 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19133_,
		_w19134_
	);
	LUT4 #(
		.INIT('h7f00)
	) name15087 (
		_w19120_,
		_w19131_,
		_w19132_,
		_w19134_,
		_w19135_
	);
	LUT4 #(
		.INIT('h1000)
	) name15088 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19136_
	);
	LUT2 #(
		.INIT('h2)
	) name15089 (
		_w4102_,
		_w19136_,
		_w19137_
	);
	LUT2 #(
		.INIT('h4)
	) name15090 (
		_w19135_,
		_w19137_,
		_w19138_
	);
	LUT4 #(
		.INIT('hb000)
	) name15091 (
		_w19121_,
		_w19125_,
		_w19129_,
		_w19130_,
		_w19139_
	);
	LUT4 #(
		.INIT('h0400)
	) name15092 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w19140_
	);
	LUT4 #(
		.INIT('h00bf)
	) name15093 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19140_,
		_w19141_
	);
	LUT4 #(
		.INIT('h7f00)
	) name15094 (
		_w19120_,
		_w19132_,
		_w19139_,
		_w19141_,
		_w19142_
	);
	LUT4 #(
		.INIT('h1000)
	) name15095 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19143_
	);
	LUT2 #(
		.INIT('h2)
	) name15096 (
		_w4102_,
		_w19143_,
		_w19144_
	);
	LUT2 #(
		.INIT('h4)
	) name15097 (
		_w19142_,
		_w19144_,
		_w19145_
	);
	LUT3 #(
		.INIT('h20)
	) name15098 (
		_w19118_,
		_w19119_,
		_w19132_,
		_w19146_
	);
	LUT4 #(
		.INIT('h4777)
	) name15099 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		_w4104_,
		_w19131_,
		_w19146_,
		_w19147_
	);
	LUT2 #(
		.INIT('h2)
	) name15100 (
		_w4102_,
		_w19147_,
		_w19148_
	);
	LUT4 #(
		.INIT('h4777)
	) name15101 (
		\core_c_dec_MTAY0_E_reg/P0001 ,
		_w4104_,
		_w19139_,
		_w19146_,
		_w19149_
	);
	LUT2 #(
		.INIT('h2)
	) name15102 (
		_w4102_,
		_w19149_,
		_w19150_
	);
	LUT3 #(
		.INIT('h48)
	) name15103 (
		\sport0_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		_w12109_,
		_w12310_,
		_w19151_
	);
	LUT4 #(
		.INIT('h0004)
	) name15104 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9452_,
		_w9453_,
		_w19111_,
		_w19152_
	);
	LUT4 #(
		.INIT('h8d00)
	) name15105 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w11318_,
		_w17925_,
		_w19152_,
		_w19153_
	);
	LUT2 #(
		.INIT('h2)
	) name15106 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001 ,
		_w19152_,
		_w19154_
	);
	LUT2 #(
		.INIT('he)
	) name15107 (
		_w19153_,
		_w19154_,
		_w19155_
	);
	LUT3 #(
		.INIT('h13)
	) name15108 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001 ,
		_w9894_,
		_w19156_
	);
	LUT4 #(
		.INIT('h0002)
	) name15109 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w19156_,
		_w19157_
	);
	LUT4 #(
		.INIT('h313b)
	) name15110 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001 ,
		_w11631_,
		_w11635_,
		_w19158_
	);
	LUT4 #(
		.INIT('h2f00)
	) name15111 (
		_w11625_,
		_w14866_,
		_w19157_,
		_w19158_,
		_w19159_
	);
	LUT2 #(
		.INIT('h1)
	) name15112 (
		_w11624_,
		_w19159_,
		_w19160_
	);
	LUT4 #(
		.INIT('hc480)
	) name15113 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w12338_,
		_w12343_,
		_w19161_
	);
	LUT2 #(
		.INIT('he)
	) name15114 (
		_w19160_,
		_w19161_,
		_w19162_
	);
	LUT4 #(
		.INIT('h084c)
	) name15115 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w12338_,
		_w12343_,
		_w19163_
	);
	LUT2 #(
		.INIT('h2)
	) name15116 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001 ,
		_w11656_,
		_w19164_
	);
	LUT3 #(
		.INIT('h01)
	) name15117 (
		_w9946_,
		_w11659_,
		_w19164_,
		_w19165_
	);
	LUT3 #(
		.INIT('h70)
	) name15118 (
		_w11655_,
		_w14866_,
		_w19165_,
		_w19166_
	);
	LUT2 #(
		.INIT('h1)
	) name15119 (
		_w19163_,
		_w19166_,
		_w19167_
	);
	LUT4 #(
		.INIT('h3b38)
	) name15120 (
		IACKn_pad,
		\sice_RCS_reg[0]/NET0131 ,
		\sice_RCS_reg[1]/NET0131 ,
		\sice_RST_req_reg/NET0131 ,
		_w19168_
	);
	LUT3 #(
		.INIT('h13)
	) name15121 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 ,
		_w9894_,
		_w19169_
	);
	LUT4 #(
		.INIT('h0002)
	) name15122 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w19169_,
		_w19170_
	);
	LUT4 #(
		.INIT('h313b)
	) name15123 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 ,
		_w11308_,
		_w11635_,
		_w19171_
	);
	LUT4 #(
		.INIT('h2f00)
	) name15124 (
		_w12282_,
		_w14866_,
		_w19170_,
		_w19171_,
		_w19172_
	);
	LUT2 #(
		.INIT('h1)
	) name15125 (
		_w11624_,
		_w19172_,
		_w19173_
	);
	LUT4 #(
		.INIT('h4c08)
	) name15126 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w12243_,
		_w12248_,
		_w19174_
	);
	LUT2 #(
		.INIT('he)
	) name15127 (
		_w19173_,
		_w19174_,
		_w19175_
	);
	LUT3 #(
		.INIT('h54)
	) name15128 (
		_w9455_,
		_w15254_,
		_w15255_,
		_w19176_
	);
	LUT4 #(
		.INIT('haa20)
	) name15129 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w9797_,
		_w9800_,
		_w9801_,
		_w19177_
	);
	LUT4 #(
		.INIT('h0154)
	) name15130 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w9456_,
		_w12116_,
		_w12119_,
		_w19178_
	);
	LUT3 #(
		.INIT('h56)
	) name15131 (
		_w9473_,
		_w19177_,
		_w19178_,
		_w19179_
	);
	LUT4 #(
		.INIT('h0b07)
	) name15132 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w9455_,
		_w19176_,
		_w19179_,
		_w19180_
	);
	LUT3 #(
		.INIT('he2)
	) name15133 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001 ,
		_w13818_,
		_w19180_,
		_w19181_
	);
	LUT3 #(
		.INIT('he2)
	) name15134 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001 ,
		_w13902_,
		_w19180_,
		_w19182_
	);
	LUT3 #(
		.INIT('h48)
	) name15135 (
		\sport1_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		_w12087_,
		_w12731_,
		_w19183_
	);
	LUT4 #(
		.INIT('h2800)
	) name15136 (
		_w9841_,
		_w9843_,
		_w9846_,
		_w12115_,
		_w19184_
	);
	LUT4 #(
		.INIT('h8200)
	) name15137 (
		_w9853_,
		_w9862_,
		_w9865_,
		_w19184_,
		_w19185_
	);
	LUT3 #(
		.INIT('h80)
	) name15138 (
		_w9860_,
		_w9878_,
		_w19185_,
		_w19186_
	);
	LUT4 #(
		.INIT('h8000)
	) name15139 (
		_w9873_,
		_w9890_,
		_w14583_,
		_w19186_,
		_w19187_
	);
	LUT4 #(
		.INIT('h8000)
	) name15140 (
		_w9768_,
		_w9886_,
		_w12611_,
		_w19187_,
		_w19188_
	);
	LUT4 #(
		.INIT('h2000)
	) name15141 (
		_w9763_,
		_w9828_,
		_w9834_,
		_w19188_,
		_w19189_
	);
	LUT4 #(
		.INIT('h2000)
	) name15142 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001 ,
		_w19190_
	);
	LUT4 #(
		.INIT('h0800)
	) name15143 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001 ,
		_w19191_
	);
	LUT4 #(
		.INIT('h4000)
	) name15144 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001 ,
		_w19192_
	);
	LUT3 #(
		.INIT('h01)
	) name15145 (
		_w19191_,
		_w19192_,
		_w19190_,
		_w19193_
	);
	LUT4 #(
		.INIT('h0400)
	) name15146 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001 ,
		_w19194_
	);
	LUT4 #(
		.INIT('h0100)
	) name15147 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001 ,
		_w19195_
	);
	LUT4 #(
		.INIT('h0200)
	) name15148 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001 ,
		_w19196_
	);
	LUT4 #(
		.INIT('h1000)
	) name15149 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001 ,
		_w19197_
	);
	LUT4 #(
		.INIT('h0001)
	) name15150 (
		_w19194_,
		_w19195_,
		_w19196_,
		_w19197_,
		_w19198_
	);
	LUT2 #(
		.INIT('h8)
	) name15151 (
		_w19193_,
		_w19198_,
		_w19199_
	);
	LUT2 #(
		.INIT('h2)
	) name15152 (
		_w9911_,
		_w19199_,
		_w19200_
	);
	LUT4 #(
		.INIT('h2022)
	) name15153 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w5784_,
		_w5911_,
		_w5913_,
		_w19201_
	);
	LUT3 #(
		.INIT('h01)
	) name15154 (
		_w12114_,
		_w19200_,
		_w19201_,
		_w19202_
	);
	LUT3 #(
		.INIT('h8c)
	) name15155 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w4142_,
		_w12114_,
		_w19203_
	);
	LUT4 #(
		.INIT('h8f00)
	) name15156 (
		_w12120_,
		_w19189_,
		_w19202_,
		_w19203_,
		_w19204_
	);
	LUT4 #(
		.INIT('h80c4)
	) name15157 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w12243_,
		_w12248_,
		_w19205_
	);
	LUT2 #(
		.INIT('h2)
	) name15158 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001 ,
		_w11310_,
		_w19206_
	);
	LUT3 #(
		.INIT('h01)
	) name15159 (
		_w9946_,
		_w12442_,
		_w19206_,
		_w19207_
	);
	LUT3 #(
		.INIT('h70)
	) name15160 (
		_w12440_,
		_w14866_,
		_w19207_,
		_w19208_
	);
	LUT2 #(
		.INIT('h1)
	) name15161 (
		_w19205_,
		_w19208_,
		_w19209_
	);
	LUT4 #(
		.INIT('h2228)
	) name15162 (
		_w9455_,
		_w9473_,
		_w19177_,
		_w19178_,
		_w19210_
	);
	LUT3 #(
		.INIT('hb0)
	) name15163 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9455_,
		_w19211_
	);
	LUT4 #(
		.INIT('h0007)
	) name15164 (
		_w9910_,
		_w11802_,
		_w12111_,
		_w19211_,
		_w19212_
	);
	LUT4 #(
		.INIT('h2022)
	) name15165 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w7592_,
		_w7707_,
		_w7709_,
		_w19213_
	);
	LUT4 #(
		.INIT('h4000)
	) name15166 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001 ,
		_w19214_
	);
	LUT4 #(
		.INIT('h0800)
	) name15167 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001 ,
		_w19215_
	);
	LUT4 #(
		.INIT('h2000)
	) name15168 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001 ,
		_w19216_
	);
	LUT3 #(
		.INIT('h01)
	) name15169 (
		_w19215_,
		_w19216_,
		_w19214_,
		_w19217_
	);
	LUT4 #(
		.INIT('h0400)
	) name15170 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001 ,
		_w19218_
	);
	LUT4 #(
		.INIT('h0100)
	) name15171 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001 ,
		_w19219_
	);
	LUT4 #(
		.INIT('h1000)
	) name15172 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001 ,
		_w19220_
	);
	LUT4 #(
		.INIT('h0200)
	) name15173 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001 ,
		_w19221_
	);
	LUT4 #(
		.INIT('h0001)
	) name15174 (
		_w19218_,
		_w19219_,
		_w19220_,
		_w19221_,
		_w19222_
	);
	LUT2 #(
		.INIT('h8)
	) name15175 (
		_w19217_,
		_w19222_,
		_w19223_
	);
	LUT2 #(
		.INIT('h2)
	) name15176 (
		_w9911_,
		_w19223_,
		_w19224_
	);
	LUT3 #(
		.INIT('h01)
	) name15177 (
		_w19212_,
		_w19213_,
		_w19224_,
		_w19225_
	);
	LUT3 #(
		.INIT('h8c)
	) name15178 (
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w4142_,
		_w19212_,
		_w19226_
	);
	LUT3 #(
		.INIT('hb0)
	) name15179 (
		_w19210_,
		_w19225_,
		_w19226_,
		_w19227_
	);
	LUT4 #(
		.INIT('h2000)
	) name15180 (
		\core_c_dec_pMFALU_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19228_
	);
	LUT2 #(
		.INIT('h8)
	) name15181 (
		_w19065_,
		_w19048_,
		_w19229_
	);
	LUT2 #(
		.INIT('h8)
	) name15182 (
		_w19036_,
		_w19052_,
		_w19230_
	);
	LUT4 #(
		.INIT('h8000)
	) name15183 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19231_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15184 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w5028_,
		_w12392_,
		_w19232_
	);
	LUT3 #(
		.INIT('h54)
	) name15185 (
		_w19040_,
		_w19231_,
		_w19232_,
		_w19233_
	);
	LUT2 #(
		.INIT('h1)
	) name15186 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w19234_
	);
	LUT4 #(
		.INIT('h5400)
	) name15187 (
		_w19040_,
		_w19231_,
		_w19232_,
		_w19234_,
		_w19235_
	);
	LUT4 #(
		.INIT('h8000)
	) name15188 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19236_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name15189 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w5028_,
		_w12392_,
		_w19237_
	);
	LUT2 #(
		.INIT('h1)
	) name15190 (
		_w19236_,
		_w19237_,
		_w19238_
	);
	LUT3 #(
		.INIT('h54)
	) name15191 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w19236_,
		_w19237_,
		_w19239_
	);
	LUT4 #(
		.INIT('h1110)
	) name15192 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w19236_,
		_w19237_,
		_w19240_
	);
	LUT2 #(
		.INIT('h8)
	) name15193 (
		_w19235_,
		_w19240_,
		_w19241_
	);
	LUT3 #(
		.INIT('h07)
	) name15194 (
		_w19060_,
		_w19230_,
		_w19241_,
		_w19242_
	);
	LUT4 #(
		.INIT('hecee)
	) name15195 (
		_w19032_,
		_w19228_,
		_w19229_,
		_w19242_,
		_w19243_
	);
	LUT4 #(
		.INIT('h2000)
	) name15196 (
		\core_c_dec_MFALU_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19244_
	);
	LUT4 #(
		.INIT('hff8a)
	) name15197 (
		_w15539_,
		_w19229_,
		_w19242_,
		_w19244_,
		_w19245_
	);
	LUT3 #(
		.INIT('hca)
	) name15198 (
		\sport1_txctl_TXSHT_reg[6]/P0001 ,
		\sport1_txctl_TX_reg[7]/P0001 ,
		_w14269_,
		_w19246_
	);
	LUT3 #(
		.INIT('h40)
	) name15199 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w19247_
	);
	LUT4 #(
		.INIT('hff48)
	) name15200 (
		\sport1_cfg_FSi_cnt_reg[10]/NET0131 ,
		_w17698_,
		_w17670_,
		_w19247_,
		_w19248_
	);
	LUT3 #(
		.INIT('h40)
	) name15201 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w19249_
	);
	LUT4 #(
		.INIT('hff48)
	) name15202 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		_w17698_,
		_w17672_,
		_w19249_,
		_w19250_
	);
	LUT3 #(
		.INIT('h40)
	) name15203 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w19251_
	);
	LUT4 #(
		.INIT('hff48)
	) name15204 (
		\sport0_cfg_FSi_cnt_reg[10]/NET0131 ,
		_w17734_,
		_w17706_,
		_w19251_,
		_w19252_
	);
	LUT3 #(
		.INIT('hca)
	) name15205 (
		\sport0_txctl_TXSHT_reg[6]/P0001 ,
		\sport0_txctl_TX_reg[7]/P0001 ,
		_w12552_,
		_w19253_
	);
	LUT3 #(
		.INIT('h40)
	) name15206 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w19254_
	);
	LUT4 #(
		.INIT('hff48)
	) name15207 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		_w17734_,
		_w17708_,
		_w19254_,
		_w19255_
	);
	LUT2 #(
		.INIT('h2)
	) name15208 (
		\core_dag_ilm2reg_M_E_reg[1]/NET0131 ,
		_w4857_,
		_w19256_
	);
	LUT4 #(
		.INIT('h4440)
	) name15209 (
		_w4061_,
		_w4062_,
		_w15895_,
		_w15896_,
		_w19257_
	);
	LUT3 #(
		.INIT('h80)
	) name15210 (
		\sport1_regs_AUTOreg_DO_reg[3]/NET0131 ,
		_w4061_,
		_w4062_,
		_w19258_
	);
	LUT4 #(
		.INIT('h0040)
	) name15211 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[3]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w19259_
	);
	LUT3 #(
		.INIT('h40)
	) name15212 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[8]/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w19260_
	);
	LUT4 #(
		.INIT('h0007)
	) name15213 (
		\sport1_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w4982_,
		_w19259_,
		_w19260_,
		_w19261_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15214 (
		_w4857_,
		_w19257_,
		_w19258_,
		_w19261_,
		_w19262_
	);
	LUT2 #(
		.INIT('h1)
	) name15215 (
		_w19256_,
		_w19262_,
		_w19263_
	);
	LUT2 #(
		.INIT('h2)
	) name15216 (
		\core_dag_ilm2reg_M_E_reg[0]/NET0131 ,
		_w4857_,
		_w19264_
	);
	LUT4 #(
		.INIT('h4440)
	) name15217 (
		_w4061_,
		_w4062_,
		_w15901_,
		_w15902_,
		_w19265_
	);
	LUT3 #(
		.INIT('h80)
	) name15218 (
		\sport1_regs_AUTOreg_DO_reg[2]/NET0131 ,
		_w4061_,
		_w4062_,
		_w19266_
	);
	LUT3 #(
		.INIT('h40)
	) name15219 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[7]/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w19267_
	);
	LUT4 #(
		.INIT('h0040)
	) name15220 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[2]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w19268_
	);
	LUT4 #(
		.INIT('h0007)
	) name15221 (
		\sport1_regs_AUTOreg_DO_reg[7]/NET0131 ,
		_w4982_,
		_w19267_,
		_w19268_,
		_w19269_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15222 (
		_w4857_,
		_w19265_,
		_w19266_,
		_w19269_,
		_w19270_
	);
	LUT2 #(
		.INIT('h1)
	) name15223 (
		_w19264_,
		_w19270_,
		_w19271_
	);
	LUT4 #(
		.INIT('h3050)
	) name15224 (
		_w16130_,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19272_
	);
	LUT4 #(
		.INIT('h000e)
	) name15225 (
		_w19256_,
		_w19262_,
		_w19264_,
		_w19270_,
		_w19273_
	);
	LUT4 #(
		.INIT('heee0)
	) name15226 (
		_w19256_,
		_w19262_,
		_w19264_,
		_w19270_,
		_w19274_
	);
	LUT4 #(
		.INIT('hfafc)
	) name15227 (
		_w16129_,
		_w16140_,
		_w19263_,
		_w19271_,
		_w19275_
	);
	LUT2 #(
		.INIT('h4)
	) name15228 (
		_w19272_,
		_w19275_,
		_w19276_
	);
	LUT3 #(
		.INIT('h20)
	) name15229 (
		\core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19277_
	);
	LUT3 #(
		.INIT('h20)
	) name15230 (
		\core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19278_
	);
	LUT4 #(
		.INIT('h000b)
	) name15231 (
		_w12398_,
		_w13536_,
		_w19277_,
		_w19278_,
		_w19279_
	);
	LUT4 #(
		.INIT('h0020)
	) name15232 (
		\core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19280_
	);
	LUT4 #(
		.INIT('h2000)
	) name15233 (
		\core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19281_
	);
	LUT2 #(
		.INIT('h1)
	) name15234 (
		_w19280_,
		_w19281_,
		_w19282_
	);
	LUT2 #(
		.INIT('h8)
	) name15235 (
		_w19279_,
		_w19282_,
		_w19283_
	);
	LUT4 #(
		.INIT('hef00)
	) name15236 (
		_w7140_,
		_w7240_,
		_w19276_,
		_w19283_,
		_w19284_
	);
	LUT3 #(
		.INIT('h10)
	) name15237 (
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w12398_,
		_w13536_,
		_w19285_
	);
	LUT2 #(
		.INIT('h1)
	) name15238 (
		_w19284_,
		_w19285_,
		_w19286_
	);
	LUT3 #(
		.INIT('h20)
	) name15239 (
		\core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19287_
	);
	LUT3 #(
		.INIT('h20)
	) name15240 (
		\core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19288_
	);
	LUT4 #(
		.INIT('h000b)
	) name15241 (
		_w12398_,
		_w13536_,
		_w19287_,
		_w19288_,
		_w19289_
	);
	LUT4 #(
		.INIT('h0020)
	) name15242 (
		\core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19290_
	);
	LUT4 #(
		.INIT('h2000)
	) name15243 (
		\core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19291_
	);
	LUT2 #(
		.INIT('h1)
	) name15244 (
		_w19290_,
		_w19291_,
		_w19292_
	);
	LUT2 #(
		.INIT('h8)
	) name15245 (
		_w19289_,
		_w19292_,
		_w19293_
	);
	LUT3 #(
		.INIT('h10)
	) name15246 (
		\core_dag_ilm2reg_M_reg[12]/NET0131 ,
		_w12398_,
		_w13536_,
		_w19294_
	);
	LUT4 #(
		.INIT('h008f)
	) name15247 (
		_w6758_,
		_w19276_,
		_w19293_,
		_w19294_,
		_w19295_
	);
	LUT3 #(
		.INIT('h20)
	) name15248 (
		\core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19296_
	);
	LUT3 #(
		.INIT('h20)
	) name15249 (
		\core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19297_
	);
	LUT4 #(
		.INIT('h000b)
	) name15250 (
		_w12398_,
		_w13536_,
		_w19296_,
		_w19297_,
		_w19298_
	);
	LUT4 #(
		.INIT('h0020)
	) name15251 (
		\core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19299_
	);
	LUT4 #(
		.INIT('h2000)
	) name15252 (
		\core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19300_
	);
	LUT2 #(
		.INIT('h1)
	) name15253 (
		_w19299_,
		_w19300_,
		_w19301_
	);
	LUT2 #(
		.INIT('h8)
	) name15254 (
		_w19298_,
		_w19301_,
		_w19302_
	);
	LUT4 #(
		.INIT('hef00)
	) name15255 (
		_w6263_,
		_w6362_,
		_w19276_,
		_w19302_,
		_w19303_
	);
	LUT3 #(
		.INIT('h10)
	) name15256 (
		\core_dag_ilm2reg_M_reg[11]/NET0131 ,
		_w12398_,
		_w13536_,
		_w19304_
	);
	LUT2 #(
		.INIT('h1)
	) name15257 (
		_w19303_,
		_w19304_,
		_w19305_
	);
	LUT3 #(
		.INIT('h20)
	) name15258 (
		\core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19306_
	);
	LUT3 #(
		.INIT('h20)
	) name15259 (
		\core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19307_
	);
	LUT4 #(
		.INIT('h000b)
	) name15260 (
		_w12398_,
		_w13536_,
		_w19306_,
		_w19307_,
		_w19308_
	);
	LUT4 #(
		.INIT('h0020)
	) name15261 (
		\core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19309_
	);
	LUT4 #(
		.INIT('h2000)
	) name15262 (
		\core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19310_
	);
	LUT2 #(
		.INIT('h1)
	) name15263 (
		_w19309_,
		_w19310_,
		_w19311_
	);
	LUT2 #(
		.INIT('h8)
	) name15264 (
		_w19308_,
		_w19311_,
		_w19312_
	);
	LUT4 #(
		.INIT('hef00)
	) name15265 (
		_w5937_,
		_w6038_,
		_w19276_,
		_w19312_,
		_w19313_
	);
	LUT3 #(
		.INIT('h10)
	) name15266 (
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w12398_,
		_w13536_,
		_w19314_
	);
	LUT2 #(
		.INIT('h1)
	) name15267 (
		_w19313_,
		_w19314_,
		_w19315_
	);
	LUT2 #(
		.INIT('h2)
	) name15268 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w4857_,
		_w19316_
	);
	LUT3 #(
		.INIT('h20)
	) name15269 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w4061_,
		_w4062_,
		_w19317_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15270 (
		_w4857_,
		_w19258_,
		_w19261_,
		_w19317_,
		_w19318_
	);
	LUT2 #(
		.INIT('h1)
	) name15271 (
		_w19316_,
		_w19318_,
		_w19319_
	);
	LUT2 #(
		.INIT('h2)
	) name15272 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w4857_,
		_w19320_
	);
	LUT3 #(
		.INIT('h20)
	) name15273 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w4061_,
		_w4062_,
		_w19321_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15274 (
		_w4857_,
		_w19266_,
		_w19269_,
		_w19321_,
		_w19322_
	);
	LUT2 #(
		.INIT('h1)
	) name15275 (
		_w19320_,
		_w19322_,
		_w19323_
	);
	LUT4 #(
		.INIT('h3050)
	) name15276 (
		_w16142_,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19324_
	);
	LUT4 #(
		.INIT('h000e)
	) name15277 (
		_w19316_,
		_w19318_,
		_w19320_,
		_w19322_,
		_w19325_
	);
	LUT4 #(
		.INIT('heee0)
	) name15278 (
		_w19316_,
		_w19318_,
		_w19320_,
		_w19322_,
		_w19326_
	);
	LUT4 #(
		.INIT('hfcfa)
	) name15279 (
		_w16143_,
		_w16145_,
		_w19319_,
		_w19323_,
		_w19327_
	);
	LUT2 #(
		.INIT('h4)
	) name15280 (
		_w19324_,
		_w19327_,
		_w19328_
	);
	LUT3 #(
		.INIT('h20)
	) name15281 (
		\core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19329_
	);
	LUT3 #(
		.INIT('h20)
	) name15282 (
		\core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19330_
	);
	LUT3 #(
		.INIT('h01)
	) name15283 (
		_w13546_,
		_w19329_,
		_w19330_,
		_w19331_
	);
	LUT4 #(
		.INIT('h2000)
	) name15284 (
		\core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19332_
	);
	LUT4 #(
		.INIT('h0020)
	) name15285 (
		\core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19333_
	);
	LUT2 #(
		.INIT('h1)
	) name15286 (
		_w19332_,
		_w19333_,
		_w19334_
	);
	LUT2 #(
		.INIT('h8)
	) name15287 (
		_w19331_,
		_w19334_,
		_w19335_
	);
	LUT4 #(
		.INIT('hef00)
	) name15288 (
		_w7140_,
		_w7240_,
		_w19328_,
		_w19335_,
		_w19336_
	);
	LUT2 #(
		.INIT('h4)
	) name15289 (
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w13546_,
		_w19337_
	);
	LUT2 #(
		.INIT('h1)
	) name15290 (
		_w19336_,
		_w19337_,
		_w19338_
	);
	LUT3 #(
		.INIT('h20)
	) name15291 (
		\core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19339_
	);
	LUT3 #(
		.INIT('h20)
	) name15292 (
		\core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19340_
	);
	LUT3 #(
		.INIT('h01)
	) name15293 (
		_w13546_,
		_w19339_,
		_w19340_,
		_w19341_
	);
	LUT4 #(
		.INIT('h2000)
	) name15294 (
		\core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19342_
	);
	LUT4 #(
		.INIT('h0020)
	) name15295 (
		\core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19343_
	);
	LUT2 #(
		.INIT('h1)
	) name15296 (
		_w19342_,
		_w19343_,
		_w19344_
	);
	LUT2 #(
		.INIT('h8)
	) name15297 (
		_w19341_,
		_w19344_,
		_w19345_
	);
	LUT4 #(
		.INIT('hef00)
	) name15298 (
		_w7465_,
		_w7565_,
		_w19328_,
		_w19345_,
		_w19346_
	);
	LUT2 #(
		.INIT('h4)
	) name15299 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w13546_,
		_w19347_
	);
	LUT2 #(
		.INIT('h1)
	) name15300 (
		_w19346_,
		_w19347_,
		_w19348_
	);
	LUT3 #(
		.INIT('h20)
	) name15301 (
		\core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19349_
	);
	LUT3 #(
		.INIT('h20)
	) name15302 (
		\core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19350_
	);
	LUT3 #(
		.INIT('h01)
	) name15303 (
		_w13546_,
		_w19349_,
		_w19350_,
		_w19351_
	);
	LUT4 #(
		.INIT('h2000)
	) name15304 (
		\core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19352_
	);
	LUT4 #(
		.INIT('h0020)
	) name15305 (
		\core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19353_
	);
	LUT2 #(
		.INIT('h1)
	) name15306 (
		_w19352_,
		_w19353_,
		_w19354_
	);
	LUT2 #(
		.INIT('h8)
	) name15307 (
		_w19351_,
		_w19354_,
		_w19355_
	);
	LUT2 #(
		.INIT('h4)
	) name15308 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w13546_,
		_w19356_
	);
	LUT4 #(
		.INIT('h008f)
	) name15309 (
		_w5760_,
		_w19328_,
		_w19355_,
		_w19356_,
		_w19357_
	);
	LUT3 #(
		.INIT('h20)
	) name15310 (
		\core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19358_
	);
	LUT3 #(
		.INIT('h20)
	) name15311 (
		\core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19359_
	);
	LUT3 #(
		.INIT('h01)
	) name15312 (
		_w13546_,
		_w19358_,
		_w19359_,
		_w19360_
	);
	LUT4 #(
		.INIT('h2000)
	) name15313 (
		\core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19361_
	);
	LUT4 #(
		.INIT('h0020)
	) name15314 (
		\core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19362_
	);
	LUT2 #(
		.INIT('h1)
	) name15315 (
		_w19361_,
		_w19362_,
		_w19363_
	);
	LUT2 #(
		.INIT('h8)
	) name15316 (
		_w19360_,
		_w19363_,
		_w19364_
	);
	LUT4 #(
		.INIT('hef00)
	) name15317 (
		_w6263_,
		_w6362_,
		_w19328_,
		_w19364_,
		_w19365_
	);
	LUT2 #(
		.INIT('h4)
	) name15318 (
		\core_dag_ilm1reg_M_reg[11]/NET0131 ,
		_w13546_,
		_w19366_
	);
	LUT2 #(
		.INIT('h1)
	) name15319 (
		_w19365_,
		_w19366_,
		_w19367_
	);
	LUT3 #(
		.INIT('h20)
	) name15320 (
		\core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19368_
	);
	LUT3 #(
		.INIT('h20)
	) name15321 (
		\core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19369_
	);
	LUT3 #(
		.INIT('h01)
	) name15322 (
		_w13546_,
		_w19368_,
		_w19369_,
		_w19370_
	);
	LUT4 #(
		.INIT('h2000)
	) name15323 (
		\core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19371_
	);
	LUT4 #(
		.INIT('h0020)
	) name15324 (
		\core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19372_
	);
	LUT2 #(
		.INIT('h1)
	) name15325 (
		_w19371_,
		_w19372_,
		_w19373_
	);
	LUT2 #(
		.INIT('h8)
	) name15326 (
		_w19370_,
		_w19373_,
		_w19374_
	);
	LUT4 #(
		.INIT('hef00)
	) name15327 (
		_w5937_,
		_w6038_,
		_w19328_,
		_w19374_,
		_w19375_
	);
	LUT2 #(
		.INIT('h4)
	) name15328 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		_w13546_,
		_w19376_
	);
	LUT2 #(
		.INIT('h1)
	) name15329 (
		_w19375_,
		_w19376_,
		_w19377_
	);
	LUT3 #(
		.INIT('h13)
	) name15330 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 ,
		_w9894_,
		_w19378_
	);
	LUT4 #(
		.INIT('h0002)
	) name15331 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11308_,
		_w11632_,
		_w19378_,
		_w19379_
	);
	LUT4 #(
		.INIT('h313b)
	) name15332 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 ,
		_w11308_,
		_w11635_,
		_w19380_
	);
	LUT4 #(
		.INIT('h2f00)
	) name15333 (
		_w12282_,
		_w12486_,
		_w19379_,
		_w19380_,
		_w19381_
	);
	LUT2 #(
		.INIT('h1)
	) name15334 (
		_w11624_,
		_w19381_,
		_w19382_
	);
	LUT4 #(
		.INIT('h80c4)
	) name15335 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w12248_,
		_w12291_,
		_w19383_
	);
	LUT2 #(
		.INIT('he)
	) name15336 (
		_w19382_,
		_w19383_,
		_w19384_
	);
	LUT4 #(
		.INIT('h4c08)
	) name15337 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w12248_,
		_w12291_,
		_w19385_
	);
	LUT2 #(
		.INIT('h2)
	) name15338 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001 ,
		_w11310_,
		_w19386_
	);
	LUT3 #(
		.INIT('h01)
	) name15339 (
		_w9946_,
		_w12442_,
		_w19386_,
		_w19387_
	);
	LUT3 #(
		.INIT('h70)
	) name15340 (
		_w12440_,
		_w12486_,
		_w19387_,
		_w19388_
	);
	LUT2 #(
		.INIT('h1)
	) name15341 (
		_w19385_,
		_w19388_,
		_w19389_
	);
	LUT4 #(
		.INIT('h8000)
	) name15342 (
		\clkc_STDcnt_reg[0]/NET0131 ,
		\clkc_STDcnt_reg[1]/NET0131 ,
		\clkc_STDcnt_reg[2]/NET0131 ,
		\clkc_STDcnt_reg[3]/NET0131 ,
		_w19390_
	);
	LUT2 #(
		.INIT('h8)
	) name15343 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		_w19390_,
		_w19391_
	);
	LUT3 #(
		.INIT('h80)
	) name15344 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		\clkc_STDcnt_reg[5]/NET0131 ,
		_w19390_,
		_w19392_
	);
	LUT4 #(
		.INIT('h8000)
	) name15345 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		\clkc_STDcnt_reg[5]/NET0131 ,
		\clkc_STDcnt_reg[6]/NET0131 ,
		_w19390_,
		_w19393_
	);
	LUT2 #(
		.INIT('h8)
	) name15346 (
		\clkc_STDcnt_reg[7]/NET0131 ,
		_w19393_,
		_w19394_
	);
	LUT3 #(
		.INIT('h80)
	) name15347 (
		\clkc_STDcnt_reg[7]/NET0131 ,
		\clkc_STDcnt_reg[8]/NET0131 ,
		_w19393_,
		_w19395_
	);
	LUT4 #(
		.INIT('h8000)
	) name15348 (
		\clkc_STDcnt_reg[7]/NET0131 ,
		\clkc_STDcnt_reg[8]/NET0131 ,
		\clkc_STDcnt_reg[9]/NET0131 ,
		_w19393_,
		_w19396_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name15349 (
		\clkc_STDcnt_reg[7]/NET0131 ,
		\clkc_STDcnt_reg[8]/NET0131 ,
		\clkc_ckr_reg_DO_reg[4]/NET0131 ,
		\clkc_ckr_reg_DO_reg[5]/NET0131 ,
		_w19397_
	);
	LUT4 #(
		.INIT('h8caf)
	) name15350 (
		\clkc_STDcnt_reg[5]/NET0131 ,
		\clkc_STDcnt_reg[7]/NET0131 ,
		\clkc_ckr_reg_DO_reg[2]/NET0131 ,
		\clkc_ckr_reg_DO_reg[4]/NET0131 ,
		_w19398_
	);
	LUT4 #(
		.INIT('h8241)
	) name15351 (
		\clkc_STDcnt_reg[10]/NET0131 ,
		\clkc_STDcnt_reg[9]/NET0131 ,
		\clkc_ckr_reg_DO_reg[6]/NET0131 ,
		\clkc_ckr_reg_DO_reg[7]/NET0131 ,
		_w19399_
	);
	LUT3 #(
		.INIT('h80)
	) name15352 (
		_w19397_,
		_w19398_,
		_w19399_,
		_w19400_
	);
	LUT4 #(
		.INIT('hf531)
	) name15353 (
		\clkc_STDcnt_reg[3]/NET0131 ,
		\clkc_STDcnt_reg[6]/NET0131 ,
		\clkc_ckr_reg_DO_reg[0]/NET0131 ,
		\clkc_ckr_reg_DO_reg[3]/NET0131 ,
		_w19401_
	);
	LUT4 #(
		.INIT('haf23)
	) name15354 (
		\clkc_STDcnt_reg[3]/NET0131 ,
		\clkc_STDcnt_reg[8]/NET0131 ,
		\clkc_ckr_reg_DO_reg[0]/NET0131 ,
		\clkc_ckr_reg_DO_reg[5]/NET0131 ,
		_w19402_
	);
	LUT4 #(
		.INIT('hf531)
	) name15355 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		\clkc_STDcnt_reg[5]/NET0131 ,
		\clkc_ckr_reg_DO_reg[1]/NET0131 ,
		\clkc_ckr_reg_DO_reg[2]/NET0131 ,
		_w19403_
	);
	LUT4 #(
		.INIT('h8caf)
	) name15356 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		\clkc_STDcnt_reg[6]/NET0131 ,
		\clkc_ckr_reg_DO_reg[1]/NET0131 ,
		\clkc_ckr_reg_DO_reg[3]/NET0131 ,
		_w19404_
	);
	LUT4 #(
		.INIT('h8000)
	) name15357 (
		_w19403_,
		_w19404_,
		_w19401_,
		_w19402_,
		_w19405_
	);
	LUT2 #(
		.INIT('h8)
	) name15358 (
		_w19400_,
		_w19405_,
		_w19406_
	);
	LUT3 #(
		.INIT('h12)
	) name15359 (
		\clkc_STDcnt_reg[10]/NET0131 ,
		_w19406_,
		_w19396_,
		_w19407_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15360 (
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w19408_
	);
	LUT3 #(
		.INIT('h04)
	) name15361 (
		\sport0_regs_AUTOreg_DO_reg[1]/NET0131 ,
		\sport0_txctl_c_sync1_reg/P0001 ,
		\sport0_txctl_c_sync2_reg/P0001 ,
		_w19409_
	);
	LUT4 #(
		.INIT('h0111)
	) name15362 (
		\core_c_psq_IFC_reg[14]/NET0131 ,
		\core_c_psq_Iflag_reg[6]/NET0131 ,
		\core_dag_modulo1_T0wrap_reg/P0001 ,
		\sport0_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w19410_
	);
	LUT3 #(
		.INIT('h45)
	) name15363 (
		\core_c_psq_IFC_reg[6]/NET0131 ,
		_w19409_,
		_w19410_,
		_w19411_
	);
	LUT2 #(
		.INIT('h4)
	) name15364 (
		_w19408_,
		_w19411_,
		_w19412_
	);
	LUT2 #(
		.INIT('h4)
	) name15365 (
		_w19118_,
		_w19119_,
		_w19413_
	);
	LUT2 #(
		.INIT('h8)
	) name15366 (
		_w4967_,
		_w5027_,
		_w19414_
	);
	LUT4 #(
		.INIT('h00bf)
	) name15367 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19414_,
		_w19415_
	);
	LUT4 #(
		.INIT('h7f00)
	) name15368 (
		_w19131_,
		_w19132_,
		_w19413_,
		_w19415_,
		_w19416_
	);
	LUT4 #(
		.INIT('h1000)
	) name15369 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19417_
	);
	LUT2 #(
		.INIT('h2)
	) name15370 (
		_w4102_,
		_w19417_,
		_w19418_
	);
	LUT2 #(
		.INIT('h4)
	) name15371 (
		_w19416_,
		_w19418_,
		_w19419_
	);
	LUT2 #(
		.INIT('h8)
	) name15372 (
		_w4967_,
		_w12393_,
		_w19420_
	);
	LUT4 #(
		.INIT('h00bf)
	) name15373 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19420_,
		_w19421_
	);
	LUT4 #(
		.INIT('h7f00)
	) name15374 (
		_w19132_,
		_w19139_,
		_w19413_,
		_w19421_,
		_w19422_
	);
	LUT4 #(
		.INIT('h1000)
	) name15375 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19423_
	);
	LUT2 #(
		.INIT('h2)
	) name15376 (
		_w4102_,
		_w19423_,
		_w19424_
	);
	LUT2 #(
		.INIT('h4)
	) name15377 (
		_w19422_,
		_w19424_,
		_w19425_
	);
	LUT3 #(
		.INIT('h80)
	) name15378 (
		_w19118_,
		_w19129_,
		_w19132_,
		_w19426_
	);
	LUT4 #(
		.INIT('h008a)
	) name15379 (
		_w19119_,
		_w19121_,
		_w19125_,
		_w19130_,
		_w19427_
	);
	LUT2 #(
		.INIT('h8)
	) name15380 (
		_w4967_,
		_w12916_,
		_w19428_
	);
	LUT4 #(
		.INIT('h00bf)
	) name15381 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19428_,
		_w19429_
	);
	LUT3 #(
		.INIT('h70)
	) name15382 (
		_w19426_,
		_w19427_,
		_w19429_,
		_w19430_
	);
	LUT4 #(
		.INIT('h1000)
	) name15383 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19431_
	);
	LUT2 #(
		.INIT('h2)
	) name15384 (
		_w4102_,
		_w19431_,
		_w19432_
	);
	LUT2 #(
		.INIT('h4)
	) name15385 (
		_w19430_,
		_w19432_,
		_w19433_
	);
	LUT4 #(
		.INIT('h60c0)
	) name15386 (
		\sport0_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		_w12109_,
		_w12312_,
		_w19434_
	);
	LUT4 #(
		.INIT('h208a)
	) name15387 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14289_,
		_w14292_,
		_w15551_,
		_w19435_
	);
	LUT3 #(
		.INIT('hf4)
	) name15388 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11294_,
		_w19435_,
		_w19436_
	);
	LUT4 #(
		.INIT('h60c0)
	) name15389 (
		\sport1_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		_w12087_,
		_w12733_,
		_w19437_
	);
	LUT4 #(
		.INIT('h8a00)
	) name15390 (
		_w19119_,
		_w19121_,
		_w19125_,
		_w19130_,
		_w19438_
	);
	LUT3 #(
		.INIT('h40)
	) name15391 (
		_w4104_,
		_w19426_,
		_w19438_,
		_w19439_
	);
	LUT4 #(
		.INIT('h2000)
	) name15392 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19440_
	);
	LUT3 #(
		.INIT('h07)
	) name15393 (
		_w5045_,
		_w15929_,
		_w19440_,
		_w19441_
	);
	LUT3 #(
		.INIT('h8a)
	) name15394 (
		_w4102_,
		_w19439_,
		_w19441_,
		_w19442_
	);
	LUT4 #(
		.INIT('h0155)
	) name15395 (
		\sport1_cfg_FSi_reg/NET0131 ,
		_w17675_,
		_w17696_,
		_w17697_,
		_w19443_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name15396 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w19444_
	);
	LUT2 #(
		.INIT('h9)
	) name15397 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w19445_
	);
	LUT2 #(
		.INIT('h8)
	) name15398 (
		_w19444_,
		_w19445_,
		_w19446_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name15399 (
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w19447_
	);
	LUT4 #(
		.INIT('hcf45)
	) name15400 (
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w19448_
	);
	LUT4 #(
		.INIT('haf23)
	) name15401 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w19449_
	);
	LUT3 #(
		.INIT('h80)
	) name15402 (
		_w19447_,
		_w19448_,
		_w19449_,
		_w19450_
	);
	LUT2 #(
		.INIT('h8)
	) name15403 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		_w19451_
	);
	LUT4 #(
		.INIT('h0800)
	) name15404 (
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w19452_
	);
	LUT2 #(
		.INIT('h8)
	) name15405 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w19453_
	);
	LUT3 #(
		.INIT('h70)
	) name15406 (
		_w19451_,
		_w19452_,
		_w19453_,
		_w19454_
	);
	LUT4 #(
		.INIT('h80aa)
	) name15407 (
		\sport1_cfg_FSi_reg/NET0131 ,
		_w19446_,
		_w19450_,
		_w19454_,
		_w19455_
	);
	LUT2 #(
		.INIT('h1)
	) name15408 (
		_w19443_,
		_w19455_,
		_w19456_
	);
	LUT4 #(
		.INIT('h0155)
	) name15409 (
		\sport0_cfg_FSi_reg/NET0131 ,
		_w17711_,
		_w17732_,
		_w17733_,
		_w19457_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name15410 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w19458_
	);
	LUT2 #(
		.INIT('h9)
	) name15411 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w19459_
	);
	LUT2 #(
		.INIT('h8)
	) name15412 (
		_w19458_,
		_w19459_,
		_w19460_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name15413 (
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w19461_
	);
	LUT4 #(
		.INIT('hcf45)
	) name15414 (
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w19462_
	);
	LUT4 #(
		.INIT('haf23)
	) name15415 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w19463_
	);
	LUT3 #(
		.INIT('h80)
	) name15416 (
		_w19461_,
		_w19462_,
		_w19463_,
		_w19464_
	);
	LUT2 #(
		.INIT('h8)
	) name15417 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		_w19465_
	);
	LUT4 #(
		.INIT('h0800)
	) name15418 (
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w19466_
	);
	LUT2 #(
		.INIT('h8)
	) name15419 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w19467_
	);
	LUT3 #(
		.INIT('h70)
	) name15420 (
		_w19465_,
		_w19466_,
		_w19467_,
		_w19468_
	);
	LUT4 #(
		.INIT('h80aa)
	) name15421 (
		\sport0_cfg_FSi_reg/NET0131 ,
		_w19460_,
		_w19464_,
		_w19468_,
		_w19469_
	);
	LUT2 #(
		.INIT('h1)
	) name15422 (
		_w19457_,
		_w19469_,
		_w19470_
	);
	LUT4 #(
		.INIT('h2000)
	) name15423 (
		\core_c_dec_pMFSHT_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19471_
	);
	LUT3 #(
		.INIT('h01)
	) name15424 (
		_w19051_,
		_w19052_,
		_w19050_,
		_w19472_
	);
	LUT2 #(
		.INIT('h8)
	) name15425 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w19473_
	);
	LUT4 #(
		.INIT('h5400)
	) name15426 (
		_w19040_,
		_w19231_,
		_w19232_,
		_w19473_,
		_w19474_
	);
	LUT2 #(
		.INIT('h8)
	) name15427 (
		_w19240_,
		_w19474_,
		_w19475_
	);
	LUT3 #(
		.INIT('h07)
	) name15428 (
		_w19057_,
		_w19472_,
		_w19475_,
		_w19476_
	);
	LUT2 #(
		.INIT('h8)
	) name15429 (
		_w19051_,
		_w19052_,
		_w19477_
	);
	LUT3 #(
		.INIT('h08)
	) name15430 (
		_w19051_,
		_w19052_,
		_w19050_,
		_w19478_
	);
	LUT4 #(
		.INIT('h113f)
	) name15431 (
		_w19057_,
		_w19049_,
		_w19472_,
		_w19478_,
		_w19479_
	);
	LUT4 #(
		.INIT('hceee)
	) name15432 (
		_w19032_,
		_w19471_,
		_w19476_,
		_w19479_,
		_w19480_
	);
	LUT4 #(
		.INIT('h2000)
	) name15433 (
		\core_c_dec_MFSHT_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19481_
	);
	LUT4 #(
		.INIT('hff2a)
	) name15434 (
		_w15539_,
		_w19476_,
		_w19479_,
		_w19481_,
		_w19482_
	);
	LUT4 #(
		.INIT('h3c2d)
	) name15435 (
		\T_TMODE[0]_pad ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TSR_TMP_reg[4]/NET0131 ,
		_w14105_,
		_w19483_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name15436 (
		\tm_tsr_reg_DO_reg[4]/NET0131 ,
		_w12802_,
		_w15792_,
		_w19483_,
		_w19484_
	);
	LUT3 #(
		.INIT('h40)
	) name15437 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w19485_
	);
	LUT3 #(
		.INIT('h6c)
	) name15438 (
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[7]/NET0131 ,
		_w17703_,
		_w19486_
	);
	LUT3 #(
		.INIT('hec)
	) name15439 (
		_w17734_,
		_w19485_,
		_w19486_,
		_w19487_
	);
	LUT3 #(
		.INIT('h40)
	) name15440 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w19488_
	);
	LUT3 #(
		.INIT('h6c)
	) name15441 (
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[7]/NET0131 ,
		_w17667_,
		_w19489_
	);
	LUT3 #(
		.INIT('hec)
	) name15442 (
		_w17698_,
		_w19488_,
		_w19489_,
		_w19490_
	);
	LUT3 #(
		.INIT('h40)
	) name15443 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w19491_
	);
	LUT4 #(
		.INIT('hff48)
	) name15444 (
		\sport1_cfg_FSi_cnt_reg[8]/NET0131 ,
		_w17698_,
		_w17668_,
		_w19491_,
		_w19492_
	);
	LUT3 #(
		.INIT('h40)
	) name15445 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w19493_
	);
	LUT4 #(
		.INIT('hff48)
	) name15446 (
		\sport0_cfg_FSi_cnt_reg[8]/NET0131 ,
		_w17734_,
		_w17704_,
		_w19493_,
		_w19494_
	);
	LUT3 #(
		.INIT('h04)
	) name15447 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RCS_reg[1]/NET0131 ,
		\sport1_rxctl_RCS_reg[2]/NET0131 ,
		_w19495_
	);
	LUT3 #(
		.INIT('h12)
	) name15448 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RCS_reg[1]/NET0131 ,
		\sport1_rxctl_RCS_reg[2]/NET0131 ,
		_w19496_
	);
	LUT3 #(
		.INIT('hd0)
	) name15449 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		_w18878_,
		_w19496_,
		_w19497_
	);
	LUT4 #(
		.INIT('he9eb)
	) name15450 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RCS_reg[1]/NET0131 ,
		\sport1_rxctl_RCS_reg[2]/NET0131 ,
		_w18878_,
		_w19498_
	);
	LUT4 #(
		.INIT('h0001)
	) name15451 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[2]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[3]/NET0131 ,
		_w19499_
	);
	LUT2 #(
		.INIT('h4)
	) name15452 (
		\sport1_rxctl_Bcnt_reg[4]/NET0131 ,
		_w19499_,
		_w19500_
	);
	LUT4 #(
		.INIT('h2f00)
	) name15453 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		_w18878_,
		_w19496_,
		_w19500_,
		_w19501_
	);
	LUT2 #(
		.INIT('h1)
	) name15454 (
		_w19498_,
		_w19501_,
		_w19502_
	);
	LUT3 #(
		.INIT('ha8)
	) name15455 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w19498_,
		_w19501_,
		_w19503_
	);
	LUT4 #(
		.INIT('h01fe)
	) name15456 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[2]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[3]/NET0131 ,
		_w19504_
	);
	LUT4 #(
		.INIT('h5554)
	) name15457 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w19504_,
		_w19498_,
		_w19501_,
		_w19505_
	);
	LUT2 #(
		.INIT('hb)
	) name15458 (
		_w19503_,
		_w19505_,
		_w19506_
	);
	LUT3 #(
		.INIT('h1e)
	) name15459 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[2]/NET0131 ,
		_w19507_
	);
	LUT3 #(
		.INIT('h01)
	) name15460 (
		_w19498_,
		_w19501_,
		_w19507_,
		_w19508_
	);
	LUT4 #(
		.INIT('h1113)
	) name15461 (
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w19498_,
		_w19501_,
		_w19509_
	);
	LUT2 #(
		.INIT('hb)
	) name15462 (
		_w19508_,
		_w19509_,
		_w19510_
	);
	LUT2 #(
		.INIT('h6)
	) name15463 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[1]/NET0131 ,
		_w19511_
	);
	LUT3 #(
		.INIT('h01)
	) name15464 (
		_w19498_,
		_w19501_,
		_w19511_,
		_w19512_
	);
	LUT4 #(
		.INIT('h1113)
	) name15465 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w19498_,
		_w19501_,
		_w19513_
	);
	LUT2 #(
		.INIT('hb)
	) name15466 (
		_w19512_,
		_w19513_,
		_w19514_
	);
	LUT3 #(
		.INIT('ha8)
	) name15467 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w19498_,
		_w19501_,
		_w19515_
	);
	LUT4 #(
		.INIT('h3332)
	) name15468 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w19498_,
		_w19501_,
		_w19516_
	);
	LUT2 #(
		.INIT('hb)
	) name15469 (
		_w19515_,
		_w19516_,
		_w19517_
	);
	LUT4 #(
		.INIT('h4500)
	) name15470 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w19276_,
		_w19518_
	);
	LUT4 #(
		.INIT('h2000)
	) name15471 (
		\core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19519_
	);
	LUT4 #(
		.INIT('h0020)
	) name15472 (
		\core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19520_
	);
	LUT3 #(
		.INIT('h20)
	) name15473 (
		\core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19521_
	);
	LUT3 #(
		.INIT('h20)
	) name15474 (
		\core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19522_
	);
	LUT4 #(
		.INIT('h0001)
	) name15475 (
		_w19520_,
		_w19521_,
		_w19519_,
		_w19522_,
		_w19523_
	);
	LUT2 #(
		.INIT('hb)
	) name15476 (
		_w19518_,
		_w19523_,
		_w19524_
	);
	LUT4 #(
		.INIT('h4500)
	) name15477 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w19276_,
		_w19525_
	);
	LUT4 #(
		.INIT('h2000)
	) name15478 (
		\core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19526_
	);
	LUT4 #(
		.INIT('h0020)
	) name15479 (
		\core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19527_
	);
	LUT3 #(
		.INIT('h20)
	) name15480 (
		\core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19528_
	);
	LUT3 #(
		.INIT('h20)
	) name15481 (
		\core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19529_
	);
	LUT4 #(
		.INIT('h0001)
	) name15482 (
		_w19527_,
		_w19528_,
		_w19526_,
		_w19529_,
		_w19530_
	);
	LUT2 #(
		.INIT('hb)
	) name15483 (
		_w19525_,
		_w19530_,
		_w19531_
	);
	LUT4 #(
		.INIT('h4500)
	) name15484 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w19276_,
		_w19532_
	);
	LUT4 #(
		.INIT('h0020)
	) name15485 (
		\core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19533_
	);
	LUT4 #(
		.INIT('h2000)
	) name15486 (
		\core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19534_
	);
	LUT3 #(
		.INIT('h20)
	) name15487 (
		\core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19535_
	);
	LUT3 #(
		.INIT('h20)
	) name15488 (
		\core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19536_
	);
	LUT4 #(
		.INIT('h0001)
	) name15489 (
		_w19534_,
		_w19535_,
		_w19533_,
		_w19536_,
		_w19537_
	);
	LUT2 #(
		.INIT('hb)
	) name15490 (
		_w19532_,
		_w19537_,
		_w19538_
	);
	LUT4 #(
		.INIT('h4500)
	) name15491 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w19276_,
		_w19539_
	);
	LUT4 #(
		.INIT('h0020)
	) name15492 (
		\core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19540_
	);
	LUT4 #(
		.INIT('h2000)
	) name15493 (
		\core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19541_
	);
	LUT3 #(
		.INIT('h20)
	) name15494 (
		\core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19542_
	);
	LUT3 #(
		.INIT('h20)
	) name15495 (
		\core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19543_
	);
	LUT4 #(
		.INIT('h0001)
	) name15496 (
		_w19541_,
		_w19542_,
		_w19540_,
		_w19543_,
		_w19544_
	);
	LUT2 #(
		.INIT('hb)
	) name15497 (
		_w19539_,
		_w19544_,
		_w19545_
	);
	LUT4 #(
		.INIT('h4500)
	) name15498 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w19276_,
		_w19546_
	);
	LUT4 #(
		.INIT('h0020)
	) name15499 (
		\core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19547_
	);
	LUT4 #(
		.INIT('h2000)
	) name15500 (
		\core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19548_
	);
	LUT3 #(
		.INIT('h20)
	) name15501 (
		\core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19549_
	);
	LUT3 #(
		.INIT('h20)
	) name15502 (
		\core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19550_
	);
	LUT4 #(
		.INIT('h0001)
	) name15503 (
		_w19548_,
		_w19549_,
		_w19547_,
		_w19550_,
		_w19551_
	);
	LUT2 #(
		.INIT('hb)
	) name15504 (
		_w19546_,
		_w19551_,
		_w19552_
	);
	LUT4 #(
		.INIT('h4500)
	) name15505 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w19276_,
		_w19553_
	);
	LUT4 #(
		.INIT('h0020)
	) name15506 (
		\core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19554_
	);
	LUT4 #(
		.INIT('h2000)
	) name15507 (
		\core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19555_
	);
	LUT3 #(
		.INIT('h20)
	) name15508 (
		\core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19556_
	);
	LUT3 #(
		.INIT('h20)
	) name15509 (
		\core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19557_
	);
	LUT4 #(
		.INIT('h0001)
	) name15510 (
		_w19555_,
		_w19556_,
		_w19554_,
		_w19557_,
		_w19558_
	);
	LUT2 #(
		.INIT('hb)
	) name15511 (
		_w19553_,
		_w19558_,
		_w19559_
	);
	LUT4 #(
		.INIT('h4500)
	) name15512 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w19328_,
		_w19560_
	);
	LUT4 #(
		.INIT('h0020)
	) name15513 (
		\core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19561_
	);
	LUT4 #(
		.INIT('h2000)
	) name15514 (
		\core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19562_
	);
	LUT3 #(
		.INIT('h20)
	) name15515 (
		\core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19563_
	);
	LUT3 #(
		.INIT('h20)
	) name15516 (
		\core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19564_
	);
	LUT4 #(
		.INIT('h0001)
	) name15517 (
		_w19562_,
		_w19563_,
		_w19561_,
		_w19564_,
		_w19565_
	);
	LUT2 #(
		.INIT('hb)
	) name15518 (
		_w19560_,
		_w19565_,
		_w19566_
	);
	LUT4 #(
		.INIT('h4500)
	) name15519 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w19328_,
		_w19567_
	);
	LUT4 #(
		.INIT('h0020)
	) name15520 (
		\core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19568_
	);
	LUT4 #(
		.INIT('h2000)
	) name15521 (
		\core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19569_
	);
	LUT3 #(
		.INIT('h20)
	) name15522 (
		\core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19570_
	);
	LUT3 #(
		.INIT('h20)
	) name15523 (
		\core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19571_
	);
	LUT4 #(
		.INIT('h0001)
	) name15524 (
		_w19569_,
		_w19570_,
		_w19568_,
		_w19571_,
		_w19572_
	);
	LUT2 #(
		.INIT('hb)
	) name15525 (
		_w19567_,
		_w19572_,
		_w19573_
	);
	LUT4 #(
		.INIT('h4500)
	) name15526 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w19328_,
		_w19574_
	);
	LUT4 #(
		.INIT('h0020)
	) name15527 (
		\core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19575_
	);
	LUT4 #(
		.INIT('h2000)
	) name15528 (
		\core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19576_
	);
	LUT3 #(
		.INIT('h20)
	) name15529 (
		\core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19577_
	);
	LUT3 #(
		.INIT('h20)
	) name15530 (
		\core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19578_
	);
	LUT4 #(
		.INIT('h0001)
	) name15531 (
		_w19576_,
		_w19577_,
		_w19575_,
		_w19578_,
		_w19579_
	);
	LUT2 #(
		.INIT('hb)
	) name15532 (
		_w19574_,
		_w19579_,
		_w19580_
	);
	LUT4 #(
		.INIT('h4500)
	) name15533 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w19328_,
		_w19581_
	);
	LUT4 #(
		.INIT('h2000)
	) name15534 (
		\core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19582_
	);
	LUT4 #(
		.INIT('h0020)
	) name15535 (
		\core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19583_
	);
	LUT3 #(
		.INIT('h20)
	) name15536 (
		\core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19584_
	);
	LUT3 #(
		.INIT('h20)
	) name15537 (
		\core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19585_
	);
	LUT4 #(
		.INIT('h0001)
	) name15538 (
		_w19583_,
		_w19584_,
		_w19582_,
		_w19585_,
		_w19586_
	);
	LUT2 #(
		.INIT('hb)
	) name15539 (
		_w19581_,
		_w19586_,
		_w19587_
	);
	LUT4 #(
		.INIT('h4500)
	) name15540 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w19328_,
		_w19588_
	);
	LUT4 #(
		.INIT('h2000)
	) name15541 (
		\core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19589_
	);
	LUT4 #(
		.INIT('h0020)
	) name15542 (
		\core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19590_
	);
	LUT3 #(
		.INIT('h20)
	) name15543 (
		\core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19591_
	);
	LUT3 #(
		.INIT('h20)
	) name15544 (
		\core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19592_
	);
	LUT4 #(
		.INIT('h0001)
	) name15545 (
		_w19590_,
		_w19591_,
		_w19589_,
		_w19592_,
		_w19593_
	);
	LUT2 #(
		.INIT('hb)
	) name15546 (
		_w19588_,
		_w19593_,
		_w19594_
	);
	LUT4 #(
		.INIT('h4500)
	) name15547 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w19328_,
		_w19595_
	);
	LUT4 #(
		.INIT('h2000)
	) name15548 (
		\core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19596_
	);
	LUT4 #(
		.INIT('h0020)
	) name15549 (
		\core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19597_
	);
	LUT3 #(
		.INIT('h20)
	) name15550 (
		\core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19598_
	);
	LUT3 #(
		.INIT('h20)
	) name15551 (
		\core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19599_
	);
	LUT4 #(
		.INIT('h0001)
	) name15552 (
		_w19597_,
		_w19598_,
		_w19596_,
		_w19599_,
		_w19600_
	);
	LUT2 #(
		.INIT('hb)
	) name15553 (
		_w19595_,
		_w19600_,
		_w19601_
	);
	LUT4 #(
		.INIT('h0408)
	) name15554 (
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12306_,
		_w19602_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name15555 (
		\core_c_dec_updMF_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001 ,
		_w9453_,
		_w9894_,
		_w19603_
	);
	LUT4 #(
		.INIT('h8d00)
	) name15556 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12248_,
		_w12291_,
		_w13091_,
		_w19604_
	);
	LUT2 #(
		.INIT('he)
	) name15557 (
		_w19603_,
		_w19604_,
		_w19605_
	);
	LUT4 #(
		.INIT('h2000)
	) name15558 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19606_
	);
	LUT4 #(
		.INIT('h4a00)
	) name15559 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		\core_c_dec_updMR_E_reg/P0001 ,
		_w19607_
	);
	LUT3 #(
		.INIT('h40)
	) name15560 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_updMF_E_reg/P0001 ,
		_w19608_
	);
	LUT4 #(
		.INIT('h080f)
	) name15561 (
		_w11924_,
		_w13505_,
		_w19607_,
		_w19608_,
		_w19609_
	);
	LUT2 #(
		.INIT('h2)
	) name15562 (
		_w11926_,
		_w19609_,
		_w19610_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name15563 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9453_,
		_w19606_,
		_w19610_,
		_w19611_
	);
	LUT2 #(
		.INIT('h2)
	) name15564 (
		_w4102_,
		_w19611_,
		_w19612_
	);
	LUT2 #(
		.INIT('h9)
	) name15565 (
		\sport1_rxctl_Bcnt_reg[4]/NET0131 ,
		_w19499_,
		_w19613_
	);
	LUT3 #(
		.INIT('h10)
	) name15566 (
		_w19498_,
		_w19501_,
		_w19613_,
		_w19614_
	);
	LUT4 #(
		.INIT('h2223)
	) name15567 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w19498_,
		_w19501_,
		_w19615_
	);
	LUT2 #(
		.INIT('h4)
	) name15568 (
		_w19614_,
		_w19615_,
		_w19616_
	);
	LUT3 #(
		.INIT('h04)
	) name15569 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RCS_reg[1]/NET0131 ,
		\sport0_rxctl_RCS_reg[2]/NET0131 ,
		_w19617_
	);
	LUT3 #(
		.INIT('h12)
	) name15570 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RCS_reg[1]/NET0131 ,
		\sport0_rxctl_RCS_reg[2]/NET0131 ,
		_w19618_
	);
	LUT3 #(
		.INIT('hd0)
	) name15571 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		_w18892_,
		_w19618_,
		_w19619_
	);
	LUT4 #(
		.INIT('he9eb)
	) name15572 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RCS_reg[1]/NET0131 ,
		\sport0_rxctl_RCS_reg[2]/NET0131 ,
		_w18892_,
		_w19620_
	);
	LUT4 #(
		.INIT('h0001)
	) name15573 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[2]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[3]/NET0131 ,
		_w19621_
	);
	LUT2 #(
		.INIT('h4)
	) name15574 (
		\sport0_rxctl_Bcnt_reg[4]/NET0131 ,
		_w19621_,
		_w19622_
	);
	LUT4 #(
		.INIT('h2f00)
	) name15575 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		_w18892_,
		_w19618_,
		_w19622_,
		_w19623_
	);
	LUT2 #(
		.INIT('h1)
	) name15576 (
		_w19620_,
		_w19623_,
		_w19624_
	);
	LUT2 #(
		.INIT('h9)
	) name15577 (
		\sport0_rxctl_Bcnt_reg[4]/NET0131 ,
		_w19621_,
		_w19625_
	);
	LUT3 #(
		.INIT('h10)
	) name15578 (
		_w19620_,
		_w19623_,
		_w19625_,
		_w19626_
	);
	LUT4 #(
		.INIT('h2223)
	) name15579 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w19620_,
		_w19623_,
		_w19627_
	);
	LUT2 #(
		.INIT('h4)
	) name15580 (
		_w19626_,
		_w19627_,
		_w19628_
	);
	LUT4 #(
		.INIT('h01fe)
	) name15581 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[2]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[3]/NET0131 ,
		_w19629_
	);
	LUT3 #(
		.INIT('h01)
	) name15582 (
		_w19620_,
		_w19623_,
		_w19629_,
		_w19630_
	);
	LUT4 #(
		.INIT('h1113)
	) name15583 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w19620_,
		_w19623_,
		_w19631_
	);
	LUT2 #(
		.INIT('hb)
	) name15584 (
		_w19630_,
		_w19631_,
		_w19632_
	);
	LUT3 #(
		.INIT('h1e)
	) name15585 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[2]/NET0131 ,
		_w19633_
	);
	LUT3 #(
		.INIT('h01)
	) name15586 (
		_w19620_,
		_w19623_,
		_w19633_,
		_w19634_
	);
	LUT4 #(
		.INIT('h1113)
	) name15587 (
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w19620_,
		_w19623_,
		_w19635_
	);
	LUT2 #(
		.INIT('hb)
	) name15588 (
		_w19634_,
		_w19635_,
		_w19636_
	);
	LUT2 #(
		.INIT('h6)
	) name15589 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[1]/NET0131 ,
		_w19637_
	);
	LUT3 #(
		.INIT('h01)
	) name15590 (
		_w19620_,
		_w19623_,
		_w19637_,
		_w19638_
	);
	LUT4 #(
		.INIT('h1113)
	) name15591 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w19620_,
		_w19623_,
		_w19639_
	);
	LUT2 #(
		.INIT('hb)
	) name15592 (
		_w19638_,
		_w19639_,
		_w19640_
	);
	LUT3 #(
		.INIT('ha8)
	) name15593 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w19620_,
		_w19623_,
		_w19641_
	);
	LUT4 #(
		.INIT('h3332)
	) name15594 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w19620_,
		_w19623_,
		_w19642_
	);
	LUT2 #(
		.INIT('hb)
	) name15595 (
		_w19641_,
		_w19642_,
		_w19643_
	);
	LUT4 #(
		.INIT('h0408)
	) name15596 (
		\sport1_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12722_,
		_w19644_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15597 (
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w19645_
	);
	LUT2 #(
		.INIT('h8)
	) name15598 (
		\core_dag_modulo1_R0wrap_reg/P0001 ,
		\sport0_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w19646_
	);
	LUT4 #(
		.INIT('h1011)
	) name15599 (
		\core_c_psq_IFC_reg[13]/NET0131 ,
		\core_c_psq_Iflag_reg[5]/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[0]/NET0131 ,
		\sport0_rxctl_ISRa_reg/P0001 ,
		_w19647_
	);
	LUT3 #(
		.INIT('h45)
	) name15600 (
		\core_c_psq_IFC_reg[5]/NET0131 ,
		_w19646_,
		_w19647_,
		_w19648_
	);
	LUT2 #(
		.INIT('h4)
	) name15601 (
		_w19645_,
		_w19648_,
		_w19649_
	);
	LUT4 #(
		.INIT('h0001)
	) name15602 (
		\clkc_oscntr_reg_DO_reg[10]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[11]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		_w19650_
	);
	LUT2 #(
		.INIT('h2)
	) name15603 (
		\T_TMODE[0]_pad ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		_w19651_
	);
	LUT3 #(
		.INIT('h40)
	) name15604 (
		\T_TMODE[0]_pad ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		_w19652_
	);
	LUT3 #(
		.INIT('h80)
	) name15605 (
		\clkc_oscntr_reg_DO_reg[11]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		_w19653_
	);
	LUT4 #(
		.INIT('h0777)
	) name15606 (
		_w19650_,
		_w19651_,
		_w19652_,
		_w19653_,
		_w19654_
	);
	LUT2 #(
		.INIT('h4)
	) name15607 (
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		_w19655_
	);
	LUT4 #(
		.INIT('hb000)
	) name15608 (
		\clkc_oscntr_reg_DO_reg[10]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		\sport0_regs_AUTO_a_reg[14]/NET0131 ,
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w19656_
	);
	LUT4 #(
		.INIT('h0800)
	) name15609 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		_w14698_,
		_w19655_,
		_w19656_,
		_w19657_
	);
	LUT4 #(
		.INIT('h3111)
	) name15610 (
		\clkc_Cnt128_reg/NET0131 ,
		\clkc_Cnt4096_reg/NET0131 ,
		\sport0_regs_AUTO_a_reg[14]/NET0131 ,
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w19658_
	);
	LUT4 #(
		.INIT('h1055)
	) name15611 (
		\clkc_Awake_reg/NET0131 ,
		_w19654_,
		_w19657_,
		_w19658_,
		_w19659_
	);
	LUT3 #(
		.INIT('h2e)
	) name15612 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w17167_,
		_w17275_,
		_w19660_
	);
	LUT2 #(
		.INIT('h6)
	) name15613 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TSR_TMP_reg[0]/NET0131 ,
		_w19661_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name15614 (
		\tm_tsr_reg_DO_reg[0]/NET0131 ,
		_w12802_,
		_w15792_,
		_w19661_,
		_w19662_
	);
	LUT3 #(
		.INIT('h13)
	) name15615 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001 ,
		_w9894_,
		_w19663_
	);
	LUT4 #(
		.INIT('h0002)
	) name15616 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w19663_,
		_w19664_
	);
	LUT4 #(
		.INIT('h5700)
	) name15617 (
		_w11625_,
		_w12006_,
		_w12007_,
		_w19664_,
		_w19665_
	);
	LUT4 #(
		.INIT('h313b)
	) name15618 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001 ,
		_w11631_,
		_w11635_,
		_w19666_
	);
	LUT4 #(
		.INIT('h2000)
	) name15619 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w9453_,
		_w9894_,
		_w12367_,
		_w19667_
	);
	LUT4 #(
		.INIT('hff45)
	) name15620 (
		_w11624_,
		_w19665_,
		_w19666_,
		_w19667_,
		_w19668_
	);
	LUT2 #(
		.INIT('h2)
	) name15621 (
		_w9946_,
		_w12367_,
		_w19669_
	);
	LUT2 #(
		.INIT('h2)
	) name15622 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001 ,
		_w11656_,
		_w19670_
	);
	LUT3 #(
		.INIT('h01)
	) name15623 (
		_w9946_,
		_w11659_,
		_w19670_,
		_w19671_
	);
	LUT4 #(
		.INIT('hfd00)
	) name15624 (
		_w11655_,
		_w12006_,
		_w12007_,
		_w19671_,
		_w19672_
	);
	LUT2 #(
		.INIT('h1)
	) name15625 (
		_w19669_,
		_w19672_,
		_w19673_
	);
	LUT2 #(
		.INIT('h2)
	) name15626 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001 ,
		_w13168_,
		_w19674_
	);
	LUT4 #(
		.INIT('h8d00)
	) name15627 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w12248_,
		_w12291_,
		_w13168_,
		_w19675_
	);
	LUT2 #(
		.INIT('he)
	) name15628 (
		_w19674_,
		_w19675_,
		_w19676_
	);
	LUT4 #(
		.INIT('h1015)
	) name15629 (
		\core_c_psq_IFC_reg[9]/NET0131 ,
		\core_dag_modulo1_R1wrap_reg/P0001 ,
		\sport1_regs_AUTOreg_DO_reg[0]/NET0131 ,
		\sport1_rxctl_ISRa_reg/P0001 ,
		_w19677_
	);
	LUT3 #(
		.INIT('h51)
	) name15630 (
		\core_c_psq_Iflag_reg[1]/NET0131 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w19677_,
		_w19678_
	);
	LUT3 #(
		.INIT('h01)
	) name15631 (
		\core_c_psq_IFC_reg[1]/NET0131 ,
		_w13442_,
		_w19678_,
		_w19679_
	);
	LUT4 #(
		.INIT('h1000)
	) name15632 (
		\core_c_dec_MFDAG1_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19680_
	);
	LUT3 #(
		.INIT('h01)
	) name15633 (
		_w19040_,
		_w19236_,
		_w19237_,
		_w19681_
	);
	LUT4 #(
		.INIT('h0001)
	) name15634 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w19040_,
		_w19236_,
		_w19237_,
		_w19682_
	);
	LUT4 #(
		.INIT('h8880)
	) name15635 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12156_,
		_w19231_,
		_w19232_,
		_w19683_
	);
	LUT2 #(
		.INIT('h8)
	) name15636 (
		_w19682_,
		_w19683_,
		_w19684_
	);
	LUT4 #(
		.INIT('h8880)
	) name15637 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12153_,
		_w19231_,
		_w19232_,
		_w19685_
	);
	LUT2 #(
		.INIT('h8)
	) name15638 (
		_w19682_,
		_w19685_,
		_w19686_
	);
	LUT3 #(
		.INIT('h54)
	) name15639 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w19236_,
		_w19237_,
		_w19687_
	);
	LUT4 #(
		.INIT('h2220)
	) name15640 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w19236_,
		_w19237_,
		_w19688_
	);
	LUT4 #(
		.INIT('h153f)
	) name15641 (
		_w19474_,
		_w19682_,
		_w19685_,
		_w19688_,
		_w19689_
	);
	LUT2 #(
		.INIT('h4)
	) name15642 (
		_w19684_,
		_w19689_,
		_w19690_
	);
	LUT4 #(
		.INIT('h8880)
	) name15643 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12150_,
		_w19231_,
		_w19232_,
		_w19691_
	);
	LUT2 #(
		.INIT('h8)
	) name15644 (
		_w19682_,
		_w19691_,
		_w19692_
	);
	LUT3 #(
		.INIT('h54)
	) name15645 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w19231_,
		_w19232_,
		_w19693_
	);
	LUT4 #(
		.INIT('h8880)
	) name15646 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w12158_,
		_w19231_,
		_w19232_,
		_w19694_
	);
	LUT2 #(
		.INIT('h8)
	) name15647 (
		_w19682_,
		_w19694_,
		_w19695_
	);
	LUT4 #(
		.INIT('h3b3f)
	) name15648 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w19681_,
		_w19693_,
		_w19694_,
		_w19696_
	);
	LUT3 #(
		.INIT('h10)
	) name15649 (
		_w4104_,
		_w19692_,
		_w19696_,
		_w19697_
	);
	LUT3 #(
		.INIT('h15)
	) name15650 (
		_w19680_,
		_w19690_,
		_w19697_,
		_w19698_
	);
	LUT2 #(
		.INIT('h8)
	) name15651 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4106_,
		_w19699_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name15652 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[18]/NET0131 ,
		_w19034_,
		_w19124_,
		_w19700_
	);
	LUT2 #(
		.INIT('h1)
	) name15653 (
		_w19126_,
		_w19237_,
		_w19701_
	);
	LUT2 #(
		.INIT('h2)
	) name15654 (
		_w19700_,
		_w19701_,
		_w19702_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15655 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19703_
	);
	LUT4 #(
		.INIT('h8000)
	) name15656 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19704_
	);
	LUT2 #(
		.INIT('h1)
	) name15657 (
		_w19703_,
		_w19704_,
		_w19705_
	);
	LUT3 #(
		.INIT('h02)
	) name15658 (
		_w19700_,
		_w19701_,
		_w19705_,
		_w19706_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15659 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19707_
	);
	LUT4 #(
		.INIT('h8000)
	) name15660 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19708_
	);
	LUT2 #(
		.INIT('h1)
	) name15661 (
		_w19707_,
		_w19708_,
		_w19709_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15662 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19710_
	);
	LUT4 #(
		.INIT('h8000)
	) name15663 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19711_
	);
	LUT2 #(
		.INIT('h1)
	) name15664 (
		_w19710_,
		_w19711_,
		_w19712_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15665 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19713_
	);
	LUT4 #(
		.INIT('h8000)
	) name15666 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w5027_,
		_w5028_,
		_w12392_,
		_w19714_
	);
	LUT2 #(
		.INIT('h1)
	) name15667 (
		_w19713_,
		_w19714_,
		_w19715_
	);
	LUT4 #(
		.INIT('heee0)
	) name15668 (
		_w19710_,
		_w19711_,
		_w19713_,
		_w19714_,
		_w19716_
	);
	LUT2 #(
		.INIT('h4)
	) name15669 (
		_w19709_,
		_w19716_,
		_w19717_
	);
	LUT2 #(
		.INIT('h8)
	) name15670 (
		_w19706_,
		_w19717_,
		_w19718_
	);
	LUT3 #(
		.INIT('ha8)
	) name15671 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w19236_,
		_w19237_,
		_w19719_
	);
	LUT4 #(
		.INIT('h8880)
	) name15672 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w19236_,
		_w19237_,
		_w19720_
	);
	LUT2 #(
		.INIT('h8)
	) name15673 (
		_w19474_,
		_w19720_,
		_w19721_
	);
	LUT3 #(
		.INIT('h01)
	) name15674 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w19722_
	);
	LUT4 #(
		.INIT('h0080)
	) name15675 (
		_w5028_,
		_w12393_,
		_w13333_,
		_w19722_,
		_w19723_
	);
	LUT3 #(
		.INIT('h01)
	) name15676 (
		_w13334_,
		_w15673_,
		_w19723_,
		_w19724_
	);
	LUT3 #(
		.INIT('h70)
	) name15677 (
		_w19474_,
		_w19720_,
		_w19724_,
		_w19725_
	);
	LUT3 #(
		.INIT('h70)
	) name15678 (
		_w19706_,
		_w19717_,
		_w19725_,
		_w19726_
	);
	LUT4 #(
		.INIT('h0001)
	) name15679 (
		_w19707_,
		_w19708_,
		_w19710_,
		_w19711_,
		_w19727_
	);
	LUT4 #(
		.INIT('h0200)
	) name15680 (
		_w19700_,
		_w19701_,
		_w19705_,
		_w19727_,
		_w19728_
	);
	LUT4 #(
		.INIT('h0001)
	) name15681 (
		_w19710_,
		_w19711_,
		_w19713_,
		_w19714_,
		_w19729_
	);
	LUT2 #(
		.INIT('h8)
	) name15682 (
		_w19705_,
		_w19729_,
		_w19730_
	);
	LUT3 #(
		.INIT('h08)
	) name15683 (
		_w19709_,
		_w19700_,
		_w19701_,
		_w19731_
	);
	LUT2 #(
		.INIT('h4)
	) name15684 (
		_w19709_,
		_w19700_,
		_w19732_
	);
	LUT3 #(
		.INIT('h40)
	) name15685 (
		_w19709_,
		_w19700_,
		_w19701_,
		_w19733_
	);
	LUT4 #(
		.INIT('h4000)
	) name15686 (
		_w19709_,
		_w19716_,
		_w19700_,
		_w19701_,
		_w19734_
	);
	LUT4 #(
		.INIT('h0007)
	) name15687 (
		_w19730_,
		_w19731_,
		_w19734_,
		_w19728_,
		_w19735_
	);
	LUT2 #(
		.INIT('h8)
	) name15688 (
		_w19726_,
		_w19735_,
		_w19736_
	);
	LUT3 #(
		.INIT('hce)
	) name15689 (
		_w14570_,
		_w19699_,
		_w19736_,
		_w19737_
	);
	LUT4 #(
		.INIT('h1555)
	) name15690 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sice_ICYC_reg[22]/NET0131 ,
		\sice_ICYC_reg[23]/NET0131 ,
		_w13019_,
		_w19738_
	);
	LUT2 #(
		.INIT('h1)
	) name15691 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w4084_,
		_w19739_
	);
	LUT2 #(
		.INIT('h8)
	) name15692 (
		_w19738_,
		_w19739_,
		_w19740_
	);
	LUT4 #(
		.INIT('h8000)
	) name15693 (
		\sice_IIRC_reg[18]/NET0131 ,
		_w14202_,
		_w19738_,
		_w19739_,
		_w19741_
	);
	LUT3 #(
		.INIT('h6c)
	) name15694 (
		\sice_IIRC_reg[19]/NET0131 ,
		\sice_IIRC_reg[20]/NET0131 ,
		_w19741_,
		_w19742_
	);
	LUT3 #(
		.INIT('h01)
	) name15695 (
		_w4967_,
		_w4969_,
		_w5327_,
		_w19743_
	);
	LUT2 #(
		.INIT('h4)
	) name15696 (
		_w5049_,
		_w19743_,
		_w19744_
	);
	LUT3 #(
		.INIT('h23)
	) name15697 (
		_w5041_,
		_w5108_,
		_w19744_,
		_w19745_
	);
	LUT3 #(
		.INIT('h23)
	) name15698 (
		_w5104_,
		_w4970_,
		_w5049_,
		_w19746_
	);
	LUT3 #(
		.INIT('h8c)
	) name15699 (
		_w5041_,
		_w4970_,
		_w5328_,
		_w19747_
	);
	LUT2 #(
		.INIT('h1)
	) name15700 (
		_w19746_,
		_w19747_,
		_w19748_
	);
	LUT4 #(
		.INIT('hbf00)
	) name15701 (
		_w5312_,
		_w5315_,
		_w19745_,
		_w19748_,
		_w19749_
	);
	LUT3 #(
		.INIT('hd0)
	) name15702 (
		_w5771_,
		_w19745_,
		_w19749_,
		_w19750_
	);
	LUT4 #(
		.INIT('h0001)
	) name15703 (
		_w6909_,
		_w6910_,
		_w6911_,
		_w19745_,
		_w19751_
	);
	LUT3 #(
		.INIT('h02)
	) name15704 (
		_w5041_,
		_w5049_,
		_w6918_,
		_w19752_
	);
	LUT4 #(
		.INIT('h0203)
	) name15705 (
		_w5041_,
		_w5108_,
		_w6926_,
		_w19744_,
		_w19753_
	);
	LUT4 #(
		.INIT('he0ee)
	) name15706 (
		_w19746_,
		_w19747_,
		_w19752_,
		_w19753_,
		_w19754_
	);
	LUT3 #(
		.INIT('h32)
	) name15707 (
		_w4967_,
		_w5107_,
		_w4969_,
		_w19755_
	);
	LUT2 #(
		.INIT('h4)
	) name15708 (
		_w5104_,
		_w19755_,
		_w19756_
	);
	LUT2 #(
		.INIT('h1)
	) name15709 (
		_w19747_,
		_w19756_,
		_w19757_
	);
	LUT4 #(
		.INIT('h00ba)
	) name15710 (
		_w19750_,
		_w19751_,
		_w19754_,
		_w19757_,
		_w19758_
	);
	LUT2 #(
		.INIT('h4)
	) name15711 (
		_w5760_,
		_w19745_,
		_w19759_
	);
	LUT4 #(
		.INIT('h00ba)
	) name15712 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w19745_,
		_w19760_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name15713 (
		_w5041_,
		_w5108_,
		_w5562_,
		_w19744_,
		_w19761_
	);
	LUT4 #(
		.INIT('h2030)
	) name15714 (
		_w5041_,
		_w5108_,
		_w5325_,
		_w19744_,
		_w19762_
	);
	LUT4 #(
		.INIT('h000e)
	) name15715 (
		_w19746_,
		_w19747_,
		_w19762_,
		_w19761_,
		_w19763_
	);
	LUT4 #(
		.INIT('h00fd)
	) name15716 (
		_w19748_,
		_w19760_,
		_w19759_,
		_w19763_,
		_w19764_
	);
	LUT2 #(
		.INIT('h2)
	) name15717 (
		_w19757_,
		_w19764_,
		_w19765_
	);
	LUT3 #(
		.INIT('h2a)
	) name15718 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		_w11917_,
		_w15505_,
		_w19766_
	);
	LUT3 #(
		.INIT('h10)
	) name15719 (
		_w19758_,
		_w19765_,
		_w19766_,
		_w19767_
	);
	LUT4 #(
		.INIT('h5040)
	) name15720 (
		PM_bdry_sel_pad,
		_w5041_,
		_w6608_,
		_w12984_,
		_w19768_
	);
	LUT3 #(
		.INIT('h8a)
	) name15721 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w4967_,
		_w12389_,
		_w19769_
	);
	LUT4 #(
		.INIT('h3233)
	) name15722 (
		_w12978_,
		_w15565_,
		_w19768_,
		_w19769_,
		_w19770_
	);
	LUT2 #(
		.INIT('hb)
	) name15723 (
		_w19767_,
		_w19770_,
		_w19771_
	);
	LUT4 #(
		.INIT('h4555)
	) name15724 (
		\T_TMODE[1]_pad ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19772_
	);
	LUT4 #(
		.INIT('h7500)
	) name15725 (
		_w8173_,
		_w19767_,
		_w19770_,
		_w19772_,
		_w19773_
	);
	LUT4 #(
		.INIT('h4000)
	) name15726 (
		\sice_GO_NX_reg/NET0131 ,
		_w4069_,
		_w4073_,
		_w4084_,
		_w19774_
	);
	LUT2 #(
		.INIT('h1)
	) name15727 (
		_w19773_,
		_w19774_,
		_w19775_
	);
	LUT3 #(
		.INIT('h20)
	) name15728 (
		\core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19776_
	);
	LUT3 #(
		.INIT('h20)
	) name15729 (
		\core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19777_
	);
	LUT4 #(
		.INIT('h000b)
	) name15730 (
		_w12398_,
		_w13536_,
		_w19776_,
		_w19777_,
		_w19778_
	);
	LUT4 #(
		.INIT('h0020)
	) name15731 (
		\core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19779_
	);
	LUT4 #(
		.INIT('h2000)
	) name15732 (
		\core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19780_
	);
	LUT2 #(
		.INIT('h1)
	) name15733 (
		_w19779_,
		_w19780_,
		_w19781_
	);
	LUT2 #(
		.INIT('h8)
	) name15734 (
		_w19778_,
		_w19781_,
		_w19782_
	);
	LUT4 #(
		.INIT('hef00)
	) name15735 (
		_w7465_,
		_w7565_,
		_w19276_,
		_w19782_,
		_w19783_
	);
	LUT3 #(
		.INIT('h10)
	) name15736 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		_w12398_,
		_w13536_,
		_w19784_
	);
	LUT2 #(
		.INIT('h1)
	) name15737 (
		_w19783_,
		_w19784_,
		_w19785_
	);
	LUT3 #(
		.INIT('h20)
	) name15738 (
		\core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19786_
	);
	LUT3 #(
		.INIT('h20)
	) name15739 (
		\core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19787_
	);
	LUT4 #(
		.INIT('h000b)
	) name15740 (
		_w12398_,
		_w13536_,
		_w19786_,
		_w19787_,
		_w19788_
	);
	LUT4 #(
		.INIT('h2000)
	) name15741 (
		\core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19789_
	);
	LUT4 #(
		.INIT('h0020)
	) name15742 (
		\core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19790_
	);
	LUT2 #(
		.INIT('h1)
	) name15743 (
		_w19789_,
		_w19790_,
		_w19791_
	);
	LUT2 #(
		.INIT('h8)
	) name15744 (
		_w19788_,
		_w19791_,
		_w19792_
	);
	LUT3 #(
		.INIT('h10)
	) name15745 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w12398_,
		_w13536_,
		_w19793_
	);
	LUT4 #(
		.INIT('h008f)
	) name15746 (
		_w5760_,
		_w19276_,
		_w19792_,
		_w19793_,
		_w19794_
	);
	LUT3 #(
		.INIT('h20)
	) name15747 (
		\core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19795_
	);
	LUT3 #(
		.INIT('h20)
	) name15748 (
		\core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19796_
	);
	LUT3 #(
		.INIT('h01)
	) name15749 (
		_w13546_,
		_w19795_,
		_w19796_,
		_w19797_
	);
	LUT4 #(
		.INIT('h0020)
	) name15750 (
		\core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19798_
	);
	LUT4 #(
		.INIT('h2000)
	) name15751 (
		\core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19799_
	);
	LUT2 #(
		.INIT('h1)
	) name15752 (
		_w19798_,
		_w19799_,
		_w19800_
	);
	LUT2 #(
		.INIT('h8)
	) name15753 (
		_w19797_,
		_w19800_,
		_w19801_
	);
	LUT2 #(
		.INIT('h4)
	) name15754 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w13546_,
		_w19802_
	);
	LUT4 #(
		.INIT('h008f)
	) name15755 (
		_w6758_,
		_w19328_,
		_w19801_,
		_w19802_,
		_w19803_
	);
	LUT4 #(
		.INIT('h4500)
	) name15756 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w19276_,
		_w19804_
	);
	LUT3 #(
		.INIT('h20)
	) name15757 (
		\core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19805_
	);
	LUT3 #(
		.INIT('h20)
	) name15758 (
		\core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19806_
	);
	LUT4 #(
		.INIT('h000b)
	) name15759 (
		_w12398_,
		_w13536_,
		_w19805_,
		_w19806_,
		_w19807_
	);
	LUT4 #(
		.INIT('h2000)
	) name15760 (
		\core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19808_
	);
	LUT4 #(
		.INIT('h0020)
	) name15761 (
		\core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19809_
	);
	LUT2 #(
		.INIT('h1)
	) name15762 (
		_w19808_,
		_w19809_,
		_w19810_
	);
	LUT2 #(
		.INIT('h8)
	) name15763 (
		_w19807_,
		_w19810_,
		_w19811_
	);
	LUT3 #(
		.INIT('h10)
	) name15764 (
		\core_dag_ilm2reg_M_reg[7]/NET0131 ,
		_w12398_,
		_w13536_,
		_w19812_
	);
	LUT3 #(
		.INIT('h0b)
	) name15765 (
		_w19804_,
		_w19811_,
		_w19812_,
		_w19813_
	);
	LUT4 #(
		.INIT('h4500)
	) name15766 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w19276_,
		_w19814_
	);
	LUT3 #(
		.INIT('h20)
	) name15767 (
		\core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131 ,
		_w16140_,
		_w19274_,
		_w19815_
	);
	LUT3 #(
		.INIT('h20)
	) name15768 (
		\core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131 ,
		_w16129_,
		_w19273_,
		_w19816_
	);
	LUT4 #(
		.INIT('h000b)
	) name15769 (
		_w12398_,
		_w13536_,
		_w19815_,
		_w19816_,
		_w19817_
	);
	LUT4 #(
		.INIT('h2000)
	) name15770 (
		\core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131 ,
		_w16141_,
		_w19263_,
		_w19271_,
		_w19818_
	);
	LUT4 #(
		.INIT('h0020)
	) name15771 (
		\core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131 ,
		_w16130_,
		_w19263_,
		_w19271_,
		_w19819_
	);
	LUT2 #(
		.INIT('h1)
	) name15772 (
		_w19818_,
		_w19819_,
		_w19820_
	);
	LUT2 #(
		.INIT('h8)
	) name15773 (
		_w19817_,
		_w19820_,
		_w19821_
	);
	LUT3 #(
		.INIT('h10)
	) name15774 (
		\core_dag_ilm2reg_M_reg[0]/NET0131 ,
		_w12398_,
		_w13536_,
		_w19822_
	);
	LUT3 #(
		.INIT('h0b)
	) name15775 (
		_w19814_,
		_w19821_,
		_w19822_,
		_w19823_
	);
	LUT4 #(
		.INIT('h4500)
	) name15776 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w19328_,
		_w19824_
	);
	LUT3 #(
		.INIT('h20)
	) name15777 (
		\core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19825_
	);
	LUT3 #(
		.INIT('h20)
	) name15778 (
		\core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19826_
	);
	LUT3 #(
		.INIT('h01)
	) name15779 (
		_w13546_,
		_w19825_,
		_w19826_,
		_w19827_
	);
	LUT4 #(
		.INIT('h0020)
	) name15780 (
		\core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19828_
	);
	LUT4 #(
		.INIT('h2000)
	) name15781 (
		\core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19829_
	);
	LUT2 #(
		.INIT('h1)
	) name15782 (
		_w19828_,
		_w19829_,
		_w19830_
	);
	LUT2 #(
		.INIT('h8)
	) name15783 (
		_w19827_,
		_w19830_,
		_w19831_
	);
	LUT2 #(
		.INIT('h4)
	) name15784 (
		\core_dag_ilm1reg_M_reg[7]/NET0131 ,
		_w13546_,
		_w19832_
	);
	LUT3 #(
		.INIT('h0b)
	) name15785 (
		_w19824_,
		_w19831_,
		_w19832_,
		_w19833_
	);
	LUT4 #(
		.INIT('h4500)
	) name15786 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w19328_,
		_w19834_
	);
	LUT3 #(
		.INIT('h20)
	) name15787 (
		\core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131 ,
		_w16145_,
		_w19325_,
		_w19835_
	);
	LUT3 #(
		.INIT('h20)
	) name15788 (
		\core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131 ,
		_w16143_,
		_w19326_,
		_w19836_
	);
	LUT3 #(
		.INIT('h01)
	) name15789 (
		_w13546_,
		_w19835_,
		_w19836_,
		_w19837_
	);
	LUT4 #(
		.INIT('h2000)
	) name15790 (
		\core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131 ,
		_w16146_,
		_w19319_,
		_w19323_,
		_w19838_
	);
	LUT4 #(
		.INIT('h0020)
	) name15791 (
		\core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131 ,
		_w16142_,
		_w19319_,
		_w19323_,
		_w19839_
	);
	LUT2 #(
		.INIT('h1)
	) name15792 (
		_w19838_,
		_w19839_,
		_w19840_
	);
	LUT2 #(
		.INIT('h8)
	) name15793 (
		_w19837_,
		_w19840_,
		_w19841_
	);
	LUT2 #(
		.INIT('h4)
	) name15794 (
		\core_dag_ilm1reg_M_reg[3]/NET0131 ,
		_w13546_,
		_w19842_
	);
	LUT3 #(
		.INIT('h0b)
	) name15795 (
		_w19834_,
		_w19841_,
		_w19842_,
		_w19843_
	);
	LUT3 #(
		.INIT('h40)
	) name15796 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w19844_
	);
	LUT3 #(
		.INIT('h6c)
	) name15797 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		_w17666_,
		_w19845_
	);
	LUT3 #(
		.INIT('hec)
	) name15798 (
		_w17698_,
		_w19844_,
		_w19845_,
		_w19846_
	);
	LUT3 #(
		.INIT('h40)
	) name15799 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w19847_
	);
	LUT3 #(
		.INIT('h6c)
	) name15800 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		_w17702_,
		_w19848_
	);
	LUT3 #(
		.INIT('hec)
	) name15801 (
		_w17734_,
		_w19847_,
		_w19848_,
		_w19849_
	);
	LUT3 #(
		.INIT('h40)
	) name15802 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w19850_
	);
	LUT2 #(
		.INIT('h6)
	) name15803 (
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		_w17667_,
		_w19851_
	);
	LUT3 #(
		.INIT('hec)
	) name15804 (
		_w17698_,
		_w19850_,
		_w19851_,
		_w19852_
	);
	LUT3 #(
		.INIT('h40)
	) name15805 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w19853_
	);
	LUT2 #(
		.INIT('h6)
	) name15806 (
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		_w17703_,
		_w19854_
	);
	LUT3 #(
		.INIT('hec)
	) name15807 (
		_w17734_,
		_w19853_,
		_w19854_,
		_w19855_
	);
	LUT3 #(
		.INIT('h1e)
	) name15808 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TSR_TMP_reg[0]/NET0131 ,
		\tm_TSR_TMP_reg[1]/NET0131 ,
		_w19856_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name15809 (
		\tm_tsr_reg_DO_reg[1]/NET0131 ,
		_w12802_,
		_w15792_,
		_w19856_,
		_w19857_
	);
	LUT4 #(
		.INIT('h01fe)
	) name15810 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TSR_TMP_reg[0]/NET0131 ,
		\tm_TSR_TMP_reg[1]/NET0131 ,
		\tm_TSR_TMP_reg[2]/NET0131 ,
		_w19858_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name15811 (
		\tm_tsr_reg_DO_reg[2]/NET0131 ,
		_w12802_,
		_w15792_,
		_w19858_,
		_w19859_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name15812 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TSR_TMP_reg[0]/NET0131 ,
		\tm_TSR_TMP_reg[3]/NET0131 ,
		_w14104_,
		_w19860_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name15813 (
		\tm_tsr_reg_DO_reg[3]/NET0131 ,
		_w12802_,
		_w15792_,
		_w19860_,
		_w19861_
	);
	LUT3 #(
		.INIT('h04)
	) name15814 (
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		\sport1_txctl_c_sync1_reg/P0001 ,
		\sport1_txctl_c_sync2_reg/P0001 ,
		_w19862_
	);
	LUT3 #(
		.INIT('h15)
	) name15815 (
		\core_c_psq_IFC_reg[10]/NET0131 ,
		\core_dag_modulo1_T1wrap_reg/P0001 ,
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w19863_
	);
	LUT4 #(
		.INIT('h1511)
	) name15816 (
		\core_c_psq_Iflag_reg[2]/NET0131 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w19862_,
		_w19863_,
		_w19864_
	);
	LUT3 #(
		.INIT('h01)
	) name15817 (
		\core_c_psq_IFC_reg[2]/NET0131 ,
		_w13437_,
		_w19864_,
		_w19865_
	);
	LUT4 #(
		.INIT('h0100)
	) name15818 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w4971_,
		_w9453_,
		_w14777_,
		_w19866_
	);
	LUT4 #(
		.INIT('h0007)
	) name15819 (
		_w9910_,
		_w11802_,
		_w12111_,
		_w19866_,
		_w19867_
	);
	LUT4 #(
		.INIT('h0400)
	) name15820 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001 ,
		_w19868_
	);
	LUT4 #(
		.INIT('h1000)
	) name15821 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001 ,
		_w19869_
	);
	LUT4 #(
		.INIT('h0100)
	) name15822 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001 ,
		_w19870_
	);
	LUT3 #(
		.INIT('h01)
	) name15823 (
		_w19869_,
		_w19870_,
		_w19868_,
		_w19871_
	);
	LUT4 #(
		.INIT('h0200)
	) name15824 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001 ,
		_w19872_
	);
	LUT4 #(
		.INIT('h2000)
	) name15825 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001 ,
		_w19873_
	);
	LUT4 #(
		.INIT('h4000)
	) name15826 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001 ,
		_w19874_
	);
	LUT4 #(
		.INIT('h0800)
	) name15827 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001 ,
		_w19875_
	);
	LUT4 #(
		.INIT('h0001)
	) name15828 (
		_w19872_,
		_w19873_,
		_w19874_,
		_w19875_,
		_w19876_
	);
	LUT2 #(
		.INIT('h8)
	) name15829 (
		_w19871_,
		_w19876_,
		_w19877_
	);
	LUT2 #(
		.INIT('h2)
	) name15830 (
		_w9911_,
		_w19877_,
		_w19878_
	);
	LUT4 #(
		.INIT('h2022)
	) name15831 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w7793_,
		_w7903_,
		_w7905_,
		_w19879_
	);
	LUT3 #(
		.INIT('h84)
	) name15832 (
		_w11335_,
		_w14777_,
		_w14801_,
		_w19880_
	);
	LUT3 #(
		.INIT('h10)
	) name15833 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9453_,
		_w19880_,
		_w19881_
	);
	LUT4 #(
		.INIT('h0001)
	) name15834 (
		_w19867_,
		_w19879_,
		_w19878_,
		_w19881_,
		_w19882_
	);
	LUT3 #(
		.INIT('h8c)
	) name15835 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w4142_,
		_w19867_,
		_w19883_
	);
	LUT2 #(
		.INIT('h4)
	) name15836 (
		_w19882_,
		_w19883_,
		_w19884_
	);
	LUT3 #(
		.INIT('h8c)
	) name15837 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w4142_,
		_w12114_,
		_w19885_
	);
	LUT3 #(
		.INIT('hb0)
	) name15838 (
		_w12114_,
		_w12149_,
		_w19885_,
		_w19886_
	);
	LUT3 #(
		.INIT('h48)
	) name15839 (
		\sport0_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		_w12109_,
		_w12311_,
		_w19887_
	);
	LUT4 #(
		.INIT('h0408)
	) name15840 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12309_,
		_w19888_
	);
	LUT3 #(
		.INIT('h1e)
	) name15841 (
		\sport1_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[1]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[2]/NET0131 ,
		_w19889_
	);
	LUT4 #(
		.INIT('h0001)
	) name15842 (
		_w18880_,
		_w19498_,
		_w19501_,
		_w19889_,
		_w19890_
	);
	LUT3 #(
		.INIT('h01)
	) name15843 (
		_w19118_,
		_w19119_,
		_w19132_,
		_w19891_
	);
	LUT4 #(
		.INIT('h4777)
	) name15844 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w4104_,
		_w19131_,
		_w19891_,
		_w19892_
	);
	LUT2 #(
		.INIT('h2)
	) name15845 (
		_w4102_,
		_w19892_,
		_w19893_
	);
	LUT4 #(
		.INIT('h4777)
	) name15846 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w4104_,
		_w19139_,
		_w19891_,
		_w19894_
	);
	LUT2 #(
		.INIT('h2)
	) name15847 (
		_w4102_,
		_w19894_,
		_w19895_
	);
	LUT3 #(
		.INIT('h08)
	) name15848 (
		_w19118_,
		_w19119_,
		_w19132_,
		_w19896_
	);
	LUT4 #(
		.INIT('h4777)
	) name15849 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		_w4104_,
		_w19139_,
		_w19896_,
		_w19897_
	);
	LUT2 #(
		.INIT('h2)
	) name15850 (
		_w4102_,
		_w19897_,
		_w19898_
	);
	LUT4 #(
		.INIT('h4777)
	) name15851 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w4104_,
		_w19131_,
		_w19896_,
		_w19899_
	);
	LUT2 #(
		.INIT('h2)
	) name15852 (
		_w4102_,
		_w19899_,
		_w19900_
	);
	LUT3 #(
		.INIT('h02)
	) name15853 (
		_w19118_,
		_w19119_,
		_w19132_,
		_w19901_
	);
	LUT4 #(
		.INIT('h4777)
	) name15854 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		_w4104_,
		_w19131_,
		_w19901_,
		_w19902_
	);
	LUT2 #(
		.INIT('h2)
	) name15855 (
		_w4102_,
		_w19902_,
		_w19903_
	);
	LUT4 #(
		.INIT('h4777)
	) name15856 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w4104_,
		_w19139_,
		_w19901_,
		_w19904_
	);
	LUT2 #(
		.INIT('h2)
	) name15857 (
		_w4102_,
		_w19904_,
		_w19905_
	);
	LUT3 #(
		.INIT('h04)
	) name15858 (
		_w19118_,
		_w19119_,
		_w19132_,
		_w19906_
	);
	LUT4 #(
		.INIT('h4777)
	) name15859 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		_w4104_,
		_w19131_,
		_w19906_,
		_w19907_
	);
	LUT2 #(
		.INIT('h2)
	) name15860 (
		_w4102_,
		_w19907_,
		_w19908_
	);
	LUT4 #(
		.INIT('h4777)
	) name15861 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w4104_,
		_w19139_,
		_w19906_,
		_w19909_
	);
	LUT2 #(
		.INIT('h2)
	) name15862 (
		_w4102_,
		_w19909_,
		_w19910_
	);
	LUT4 #(
		.INIT('h01fe)
	) name15863 (
		\sport1_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[1]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[2]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[3]/NET0131 ,
		_w19911_
	);
	LUT4 #(
		.INIT('h0001)
	) name15864 (
		_w18880_,
		_w19498_,
		_w19501_,
		_w19911_,
		_w19912_
	);
	LUT2 #(
		.INIT('h6)
	) name15865 (
		\sport1_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[1]/NET0131 ,
		_w19913_
	);
	LUT4 #(
		.INIT('h0001)
	) name15866 (
		_w18880_,
		_w19498_,
		_w19501_,
		_w19913_,
		_w19914_
	);
	LUT4 #(
		.INIT('h01fe)
	) name15867 (
		\sport0_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[1]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[2]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[3]/NET0131 ,
		_w19915_
	);
	LUT4 #(
		.INIT('h0001)
	) name15868 (
		_w18894_,
		_w19620_,
		_w19623_,
		_w19915_,
		_w19916_
	);
	LUT3 #(
		.INIT('h1e)
	) name15869 (
		\sport0_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[1]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[2]/NET0131 ,
		_w19917_
	);
	LUT4 #(
		.INIT('h0001)
	) name15870 (
		_w18894_,
		_w19620_,
		_w19623_,
		_w19917_,
		_w19918_
	);
	LUT2 #(
		.INIT('h6)
	) name15871 (
		\sport0_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[1]/NET0131 ,
		_w19919_
	);
	LUT4 #(
		.INIT('h0001)
	) name15872 (
		_w18894_,
		_w19620_,
		_w19623_,
		_w19919_,
		_w19920_
	);
	LUT4 #(
		.INIT('h0001)
	) name15873 (
		\sport0_rxctl_LMcnt_reg[0]/NET0131 ,
		_w18894_,
		_w19620_,
		_w19623_,
		_w19921_
	);
	LUT2 #(
		.INIT('h1)
	) name15874 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		_w19922_
	);
	LUT4 #(
		.INIT('hbffd)
	) name15875 (
		\T_TMODE[0]_pad ,
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		_w19923_
	);
	LUT3 #(
		.INIT('ha2)
	) name15876 (
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w14698_,
		_w19923_,
		_w19924_
	);
	LUT4 #(
		.INIT('h0001)
	) name15877 (
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[1]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[2]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[3]/NET0131 ,
		_w19925_
	);
	LUT3 #(
		.INIT('h01)
	) name15878 (
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w19926_
	);
	LUT4 #(
		.INIT('h8000)
	) name15879 (
		_w19650_,
		_w19922_,
		_w19926_,
		_w19925_,
		_w19927_
	);
	LUT4 #(
		.INIT('h4445)
	) name15880 (
		\clkc_Awake_reg/NET0131 ,
		\clkc_Cnt128_reg/NET0131 ,
		_w19924_,
		_w19927_,
		_w19928_
	);
	LUT3 #(
		.INIT('h48)
	) name15881 (
		\sport1_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		_w12087_,
		_w12732_,
		_w19929_
	);
	LUT4 #(
		.INIT('h0408)
	) name15882 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12725_,
		_w19930_
	);
	LUT4 #(
		.INIT('h0001)
	) name15883 (
		\sport1_rxctl_LMcnt_reg[0]/NET0131 ,
		_w18880_,
		_w19498_,
		_w19501_,
		_w19931_
	);
	LUT2 #(
		.INIT('h2)
	) name15884 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w12284_,
		_w19932_
	);
	LUT4 #(
		.INIT('h4000)
	) name15885 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11837_,
		_w18164_,
		_w18165_,
		_w19933_
	);
	LUT4 #(
		.INIT('h222e)
	) name15886 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001 ,
		_w11830_,
		_w19932_,
		_w19933_,
		_w19934_
	);
	LUT4 #(
		.INIT('ha800)
	) name15887 (
		_w4067_,
		_w9414_,
		_w9415_,
		_w9423_,
		_w19935_
	);
	LUT4 #(
		.INIT('h1101)
	) name15888 (
		\core_c_psq_IFC_reg[11]/NET0131 ,
		\core_c_psq_Iflag_reg[3]/NET0131 ,
		\core_c_psq_T_IRQE0_reg/P0001 ,
		\core_c_psq_T_IRQE0_s1_reg/P0001 ,
		_w19936_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15889 (
		\core_c_psq_Iact_E_reg[3]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w19937_
	);
	LUT2 #(
		.INIT('h1)
	) name15890 (
		\core_c_psq_IFC_reg[3]/NET0131 ,
		_w19937_,
		_w19938_
	);
	LUT3 #(
		.INIT('hb0)
	) name15891 (
		_w19935_,
		_w19936_,
		_w19938_,
		_w19939_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15892 (
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		_w4094_,
		_w4097_,
		_w4101_,
		_w19940_
	);
	LUT3 #(
		.INIT('h10)
	) name15893 (
		\T_TMODE[0]_pad ,
		\tm_TINT_GEN1_reg/NET0131 ,
		\tm_TINT_GEN2_reg/NET0131 ,
		_w19941_
	);
	LUT2 #(
		.INIT('h1)
	) name15894 (
		\core_c_psq_IFC_reg[8]/NET0131 ,
		\core_c_psq_Iflag_reg[0]/NET0131 ,
		_w19942_
	);
	LUT3 #(
		.INIT('h45)
	) name15895 (
		\core_c_psq_IFC_reg[0]/NET0131 ,
		_w19941_,
		_w19942_,
		_w19943_
	);
	LUT2 #(
		.INIT('h4)
	) name15896 (
		_w19940_,
		_w19943_,
		_w19944_
	);
	LUT3 #(
		.INIT('h45)
	) name15897 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4094_,
		_w4097_,
		_w19945_
	);
	LUT3 #(
		.INIT('h32)
	) name15898 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w4971_,
		_w9911_,
		_w19946_
	);
	LUT4 #(
		.INIT('h0032)
	) name15899 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w4971_,
		_w9911_,
		_w19945_,
		_w19947_
	);
	LUT4 #(
		.INIT('h8a88)
	) name15900 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w6054_,
		_w6173_,
		_w6175_,
		_w19948_
	);
	LUT4 #(
		.INIT('h2000)
	) name15901 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001 ,
		_w19949_
	);
	LUT4 #(
		.INIT('h0800)
	) name15902 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001 ,
		_w19950_
	);
	LUT4 #(
		.INIT('h0100)
	) name15903 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001 ,
		_w19951_
	);
	LUT4 #(
		.INIT('h1000)
	) name15904 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001 ,
		_w19952_
	);
	LUT4 #(
		.INIT('h0001)
	) name15905 (
		_w19949_,
		_w19950_,
		_w19951_,
		_w19952_,
		_w19953_
	);
	LUT4 #(
		.INIT('h0200)
	) name15906 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001 ,
		_w19954_
	);
	LUT4 #(
		.INIT('h0400)
	) name15907 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001 ,
		_w19955_
	);
	LUT4 #(
		.INIT('h4000)
	) name15908 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001 ,
		_w19956_
	);
	LUT4 #(
		.INIT('h0001)
	) name15909 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w19954_,
		_w19955_,
		_w19956_,
		_w19957_
	);
	LUT2 #(
		.INIT('h8)
	) name15910 (
		_w19953_,
		_w19957_,
		_w19958_
	);
	LUT4 #(
		.INIT('haaa8)
	) name15911 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		_w19959_
	);
	LUT4 #(
		.INIT('h0045)
	) name15912 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4094_,
		_w4097_,
		_w19959_,
		_w19960_
	);
	LUT2 #(
		.INIT('h2)
	) name15913 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w19960_,
		_w19961_
	);
	LUT2 #(
		.INIT('h4)
	) name15914 (
		_w19947_,
		_w19961_,
		_w19962_
	);
	LUT4 #(
		.INIT('hff02)
	) name15915 (
		_w19947_,
		_w19948_,
		_w19958_,
		_w19962_,
		_w19963_
	);
	LUT4 #(
		.INIT('h222e)
	) name15916 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001 ,
		_w11329_,
		_w19932_,
		_w19933_,
		_w19964_
	);
	LUT4 #(
		.INIT('h4000)
	) name15917 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		_w19965_
	);
	LUT3 #(
		.INIT('h20)
	) name15918 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[7]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w19966_
	);
	LUT4 #(
		.INIT('hdf00)
	) name15919 (
		_w13097_,
		_w13099_,
		_w19965_,
		_w19966_,
		_w19967_
	);
	LUT3 #(
		.INIT('h40)
	) name15920 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[14]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w19968_
	);
	LUT2 #(
		.INIT('h1)
	) name15921 (
		_w13158_,
		_w19968_,
		_w19969_
	);
	LUT2 #(
		.INIT('h4)
	) name15922 (
		_w19967_,
		_w19969_,
		_w19970_
	);
	LUT4 #(
		.INIT('hfe00)
	) name15923 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w8757_,
		_w8760_,
		_w19970_,
		_w19971_
	);
	LUT4 #(
		.INIT('hafac)
	) name15924 (
		\sport0_rxctl_RXSHT_reg[14]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w19972_
	);
	LUT4 #(
		.INIT('h0002)
	) name15925 (
		\sport0_rxctl_RX_reg[14]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w19973_
	);
	LUT3 #(
		.INIT('hf4)
	) name15926 (
		_w19971_,
		_w19972_,
		_w19973_,
		_w19974_
	);
	LUT3 #(
		.INIT('h40)
	) name15927 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[15]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w19975_
	);
	LUT2 #(
		.INIT('h1)
	) name15928 (
		_w13158_,
		_w19975_,
		_w19976_
	);
	LUT2 #(
		.INIT('h4)
	) name15929 (
		_w19967_,
		_w19976_,
		_w19977_
	);
	LUT4 #(
		.INIT('hfe00)
	) name15930 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w8798_,
		_w8801_,
		_w19977_,
		_w19978_
	);
	LUT4 #(
		.INIT('hafac)
	) name15931 (
		\sport0_rxctl_RXSHT_reg[15]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w19979_
	);
	LUT4 #(
		.INIT('h0002)
	) name15932 (
		\sport0_rxctl_RX_reg[15]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w19980_
	);
	LUT3 #(
		.INIT('hf4)
	) name15933 (
		_w19978_,
		_w19979_,
		_w19980_,
		_w19981_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name15934 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001 ,
		_w18091_,
		_w18093_,
		_w19112_,
		_w19982_
	);
	LUT4 #(
		.INIT('heee2)
	) name15935 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w17167_,
		_w17222_,
		_w17223_,
		_w19983_
	);
	LUT4 #(
		.INIT('heee2)
	) name15936 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w17167_,
		_w17197_,
		_w17198_,
		_w19984_
	);
	LUT4 #(
		.INIT('heee2)
	) name15937 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w17167_,
		_w17205_,
		_w17206_,
		_w19985_
	);
	LUT4 #(
		.INIT('heee2)
	) name15938 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w17167_,
		_w17267_,
		_w17268_,
		_w19986_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name15939 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001 ,
		_w18624_,
		_w18626_,
		_w19112_,
		_w19987_
	);
	LUT4 #(
		.INIT('heee2)
	) name15940 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w17167_,
		_w17283_,
		_w17284_,
		_w19988_
	);
	LUT3 #(
		.INIT('h2e)
	) name15941 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w17167_,
		_w17181_,
		_w19989_
	);
	LUT4 #(
		.INIT('heee2)
	) name15942 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w17167_,
		_w17257_,
		_w17258_,
		_w19990_
	);
	LUT4 #(
		.INIT('heee2)
	) name15943 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w17167_,
		_w17188_,
		_w17189_,
		_w19991_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name15944 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001 ,
		_w18521_,
		_w18523_,
		_w19112_,
		_w19992_
	);
	LUT3 #(
		.INIT('h10)
	) name15945 (
		IACKn_pad,
		\idma_IAL_reg/P0001 ,
		\memc_MMR_web_reg/NET0131 ,
		_w19993_
	);
	LUT2 #(
		.INIT('h1)
	) name15946 (
		_w12623_,
		_w19993_,
		_w19994_
	);
	LUT4 #(
		.INIT('h888b)
	) name15947 (
		\idma_IADi_reg[8]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w7465_,
		_w7565_,
		_w19995_
	);
	LUT2 #(
		.INIT('h4)
	) name15948 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		_w19996_
	);
	LUT4 #(
		.INIT('hc088)
	) name15949 (
		\auctl_DSack_reg/NET0131 ,
		\idma_WRcyc_reg/NET0131 ,
		_w12812_,
		_w19996_,
		_w19997_
	);
	LUT2 #(
		.INIT('h1)
	) name15950 (
		_w19993_,
		_w19996_,
		_w19998_
	);
	LUT4 #(
		.INIT('ha800)
	) name15951 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w12821_,
		_w19997_,
		_w19998_,
		_w19999_
	);
	LUT4 #(
		.INIT('h8000)
	) name15952 (
		\idma_DCTL_reg[1]/NET0131 ,
		\idma_DCTL_reg[2]/NET0131 ,
		\idma_DCTL_reg[3]/NET0131 ,
		_w19999_,
		_w20000_
	);
	LUT3 #(
		.INIT('h80)
	) name15953 (
		\idma_DCTL_reg[4]/NET0131 ,
		\idma_DCTL_reg[5]/NET0131 ,
		_w20000_,
		_w20001_
	);
	LUT4 #(
		.INIT('h8000)
	) name15954 (
		\idma_DCTL_reg[4]/NET0131 ,
		\idma_DCTL_reg[5]/NET0131 ,
		\idma_DCTL_reg[6]/NET0131 ,
		_w20000_,
		_w20002_
	);
	LUT2 #(
		.INIT('h8)
	) name15955 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w20002_,
		_w20003_
	);
	LUT3 #(
		.INIT('h80)
	) name15956 (
		\idma_DCTL_reg[7]/NET0131 ,
		\idma_DCTL_reg[8]/NET0131 ,
		_w20002_,
		_w20004_
	);
	LUT3 #(
		.INIT('h12)
	) name15957 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w19994_,
		_w20003_,
		_w20005_
	);
	LUT3 #(
		.INIT('hf8)
	) name15958 (
		_w19994_,
		_w19995_,
		_w20005_,
		_w20006_
	);
	LUT4 #(
		.INIT('h888b)
	) name15959 (
		\idma_IADi_reg[9]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w7140_,
		_w7240_,
		_w20007_
	);
	LUT4 #(
		.INIT('h8000)
	) name15960 (
		\idma_DCTL_reg[7]/NET0131 ,
		\idma_DCTL_reg[8]/NET0131 ,
		\idma_DCTL_reg[9]/NET0131 ,
		_w20002_,
		_w20008_
	);
	LUT3 #(
		.INIT('h12)
	) name15961 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w19994_,
		_w20004_,
		_w20009_
	);
	LUT3 #(
		.INIT('hf8)
	) name15962 (
		_w19994_,
		_w20007_,
		_w20009_,
		_w20010_
	);
	LUT2 #(
		.INIT('h4)
	) name15963 (
		\idma_IADi_reg[13]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20011_
	);
	LUT3 #(
		.INIT('h01)
	) name15964 (
		_w12623_,
		_w19993_,
		_w20011_,
		_w20012_
	);
	LUT3 #(
		.INIT('he0)
	) name15965 (
		\idma_IAL_reg/P0001 ,
		_w5760_,
		_w20012_,
		_w20013_
	);
	LUT4 #(
		.INIT('h8000)
	) name15966 (
		\idma_DCTL_reg[10]/NET0131 ,
		\idma_DCTL_reg[11]/NET0131 ,
		\idma_DCTL_reg[12]/NET0131 ,
		_w20008_,
		_w20014_
	);
	LUT3 #(
		.INIT('h12)
	) name15967 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w19994_,
		_w20014_,
		_w20015_
	);
	LUT2 #(
		.INIT('he)
	) name15968 (
		_w20013_,
		_w20015_,
		_w20016_
	);
	LUT4 #(
		.INIT('h78f0)
	) name15969 (
		\idma_DCTL_reg[10]/NET0131 ,
		\idma_DCTL_reg[11]/NET0131 ,
		\idma_DCTL_reg[12]/NET0131 ,
		_w20008_,
		_w20017_
	);
	LUT2 #(
		.INIT('h1)
	) name15970 (
		_w19994_,
		_w20017_,
		_w20018_
	);
	LUT2 #(
		.INIT('h8)
	) name15971 (
		\idma_IADi_reg[12]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20019_
	);
	LUT3 #(
		.INIT('h01)
	) name15972 (
		_w12623_,
		_w19993_,
		_w20019_,
		_w20020_
	);
	LUT3 #(
		.INIT('hb0)
	) name15973 (
		\idma_IAL_reg/P0001 ,
		_w6758_,
		_w20020_,
		_w20021_
	);
	LUT2 #(
		.INIT('h1)
	) name15974 (
		_w20018_,
		_w20021_,
		_w20022_
	);
	LUT4 #(
		.INIT('h888b)
	) name15975 (
		\idma_IADi_reg[11]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w6263_,
		_w6362_,
		_w20023_
	);
	LUT4 #(
		.INIT('h060c)
	) name15976 (
		\idma_DCTL_reg[10]/NET0131 ,
		\idma_DCTL_reg[11]/NET0131 ,
		_w19994_,
		_w20008_,
		_w20024_
	);
	LUT3 #(
		.INIT('hf8)
	) name15977 (
		_w19994_,
		_w20023_,
		_w20024_,
		_w20025_
	);
	LUT4 #(
		.INIT('h888b)
	) name15978 (
		\idma_IADi_reg[10]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w5937_,
		_w6038_,
		_w20026_
	);
	LUT3 #(
		.INIT('h12)
	) name15979 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w19994_,
		_w20008_,
		_w20027_
	);
	LUT3 #(
		.INIT('hf8)
	) name15980 (
		_w19994_,
		_w20026_,
		_w20027_,
		_w20028_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name15981 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001 ,
		_w17749_,
		_w17751_,
		_w19112_,
		_w20029_
	);
	LUT3 #(
		.INIT('h40)
	) name15982 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[13]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w20030_
	);
	LUT2 #(
		.INIT('h1)
	) name15983 (
		_w13158_,
		_w20030_,
		_w20031_
	);
	LUT2 #(
		.INIT('h4)
	) name15984 (
		_w19967_,
		_w20031_,
		_w20032_
	);
	LUT4 #(
		.INIT('hafac)
	) name15985 (
		\sport0_rxctl_RXSHT_reg[13]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w20033_
	);
	LUT4 #(
		.INIT('h4f00)
	) name15986 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w5760_,
		_w20032_,
		_w20033_,
		_w20034_
	);
	LUT4 #(
		.INIT('h0002)
	) name15987 (
		\sport0_rxctl_RX_reg[13]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w20035_
	);
	LUT2 #(
		.INIT('he)
	) name15988 (
		_w20034_,
		_w20035_,
		_w20036_
	);
	LUT4 #(
		.INIT('h4544)
	) name15989 (
		\idma_IAL_reg/P0001 ,
		_w7793_,
		_w7903_,
		_w7905_,
		_w20037_
	);
	LUT2 #(
		.INIT('h4)
	) name15990 (
		\idma_IADi_reg[7]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20038_
	);
	LUT4 #(
		.INIT('h54a8)
	) name15991 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w12623_,
		_w19993_,
		_w20002_,
		_w20039_
	);
	LUT4 #(
		.INIT('hff02)
	) name15992 (
		_w19994_,
		_w20037_,
		_w20038_,
		_w20039_,
		_w20040_
	);
	LUT4 #(
		.INIT('h4544)
	) name15993 (
		\idma_IAL_reg/P0001 ,
		_w7592_,
		_w7707_,
		_w7709_,
		_w20041_
	);
	LUT2 #(
		.INIT('h4)
	) name15994 (
		\idma_IADi_reg[5]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20042_
	);
	LUT3 #(
		.INIT('h6c)
	) name15995 (
		\idma_DCTL_reg[4]/NET0131 ,
		\idma_DCTL_reg[5]/NET0131 ,
		_w20000_,
		_w20043_
	);
	LUT3 #(
		.INIT('he0)
	) name15996 (
		_w12623_,
		_w19993_,
		_w20043_,
		_w20044_
	);
	LUT4 #(
		.INIT('hff02)
	) name15997 (
		_w19994_,
		_w20041_,
		_w20042_,
		_w20044_,
		_w20045_
	);
	LUT4 #(
		.INIT('h4544)
	) name15998 (
		\idma_IAL_reg/P0001 ,
		_w7927_,
		_w8040_,
		_w8042_,
		_w20046_
	);
	LUT2 #(
		.INIT('h4)
	) name15999 (
		\idma_IADi_reg[6]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20047_
	);
	LUT4 #(
		.INIT('h54a8)
	) name16000 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w12623_,
		_w19993_,
		_w20001_,
		_w20048_
	);
	LUT4 #(
		.INIT('hff02)
	) name16001 (
		_w19994_,
		_w20046_,
		_w20047_,
		_w20048_,
		_w20049_
	);
	LUT4 #(
		.INIT('h4544)
	) name16002 (
		\idma_IAL_reg/P0001 ,
		_w7257_,
		_w7375_,
		_w7377_,
		_w20050_
	);
	LUT2 #(
		.INIT('h4)
	) name16003 (
		\idma_IADi_reg[4]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20051_
	);
	LUT2 #(
		.INIT('h6)
	) name16004 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w20000_,
		_w20052_
	);
	LUT3 #(
		.INIT('he0)
	) name16005 (
		_w12623_,
		_w19993_,
		_w20052_,
		_w20053_
	);
	LUT4 #(
		.INIT('hff02)
	) name16006 (
		_w19994_,
		_w20050_,
		_w20051_,
		_w20053_,
		_w20054_
	);
	LUT4 #(
		.INIT('h4544)
	) name16007 (
		\idma_IAL_reg/P0001 ,
		_w6054_,
		_w6173_,
		_w6175_,
		_w20055_
	);
	LUT2 #(
		.INIT('h4)
	) name16008 (
		\idma_IADi_reg[3]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20056_
	);
	LUT4 #(
		.INIT('h78f0)
	) name16009 (
		\idma_DCTL_reg[1]/NET0131 ,
		\idma_DCTL_reg[2]/NET0131 ,
		\idma_DCTL_reg[3]/NET0131 ,
		_w19999_,
		_w20057_
	);
	LUT3 #(
		.INIT('he0)
	) name16010 (
		_w12623_,
		_w19993_,
		_w20057_,
		_w20058_
	);
	LUT4 #(
		.INIT('hff02)
	) name16011 (
		_w19994_,
		_w20055_,
		_w20056_,
		_w20058_,
		_w20059_
	);
	LUT4 #(
		.INIT('h4544)
	) name16012 (
		\idma_IAL_reg/P0001 ,
		_w6378_,
		_w6498_,
		_w6500_,
		_w20060_
	);
	LUT2 #(
		.INIT('h4)
	) name16013 (
		\idma_IADi_reg[2]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20061_
	);
	LUT3 #(
		.INIT('h6c)
	) name16014 (
		\idma_DCTL_reg[1]/NET0131 ,
		\idma_DCTL_reg[2]/NET0131 ,
		_w19999_,
		_w20062_
	);
	LUT3 #(
		.INIT('he0)
	) name16015 (
		_w12623_,
		_w19993_,
		_w20062_,
		_w20063_
	);
	LUT4 #(
		.INIT('hff02)
	) name16016 (
		_w19994_,
		_w20060_,
		_w20061_,
		_w20063_,
		_w20064_
	);
	LUT4 #(
		.INIT('h4544)
	) name16017 (
		\idma_IAL_reg/P0001 ,
		_w5784_,
		_w5911_,
		_w5913_,
		_w20065_
	);
	LUT2 #(
		.INIT('h4)
	) name16018 (
		\idma_IADi_reg[0]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20066_
	);
	LUT4 #(
		.INIT('h56aa)
	) name16019 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w12821_,
		_w19997_,
		_w19998_,
		_w20067_
	);
	LUT3 #(
		.INIT('he0)
	) name16020 (
		_w12623_,
		_w19993_,
		_w20067_,
		_w20068_
	);
	LUT4 #(
		.INIT('hff02)
	) name16021 (
		_w19994_,
		_w20065_,
		_w20066_,
		_w20068_,
		_w20069_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16022 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001 ,
		_w17787_,
		_w17789_,
		_w19112_,
		_w20070_
	);
	LUT4 #(
		.INIT('heee2)
	) name16023 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w17167_,
		_w17232_,
		_w17233_,
		_w20071_
	);
	LUT4 #(
		.INIT('heee2)
	) name16024 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w17167_,
		_w17240_,
		_w17241_,
		_w20072_
	);
	LUT4 #(
		.INIT('h222e)
	) name16025 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		_w17167_,
		_w17292_,
		_w17291_,
		_w20073_
	);
	LUT3 #(
		.INIT('h40)
	) name16026 (
		\sport1_rxctl_Bcnt_reg[4]/NET0131 ,
		_w19499_,
		_w19495_,
		_w20074_
	);
	LUT2 #(
		.INIT('h1)
	) name16027 (
		\sport1_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[1]/NET0131 ,
		_w20075_
	);
	LUT4 #(
		.INIT('h0001)
	) name16028 (
		\sport1_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[1]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[2]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		_w20076_
	);
	LUT2 #(
		.INIT('h8)
	) name16029 (
		_w12829_,
		_w20076_,
		_w20077_
	);
	LUT2 #(
		.INIT('h8)
	) name16030 (
		_w20074_,
		_w20077_,
		_w20078_
	);
	LUT2 #(
		.INIT('h1)
	) name16031 (
		_w19498_,
		_w20078_,
		_w20079_
	);
	LUT2 #(
		.INIT('he)
	) name16032 (
		_w19498_,
		_w20078_,
		_w20080_
	);
	LUT2 #(
		.INIT('h2)
	) name16033 (
		_w20074_,
		_w20077_,
		_w20081_
	);
	LUT4 #(
		.INIT('h0040)
	) name16034 (
		\sport1_rxctl_Wcnt_reg[2]/NET0131 ,
		_w20074_,
		_w20075_,
		_w20077_,
		_w20082_
	);
	LUT3 #(
		.INIT('h63)
	) name16035 (
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[4]/NET0131 ,
		_w20082_,
		_w20083_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16036 (
		\sport1_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w19498_,
		_w20078_,
		_w20083_,
		_w20084_
	);
	LUT4 #(
		.INIT('heee2)
	) name16037 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w17167_,
		_w17249_,
		_w17250_,
		_w20085_
	);
	LUT4 #(
		.INIT('heee2)
	) name16038 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w17167_,
		_w17208_,
		_w17215_,
		_w20086_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16039 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001 ,
		_w17849_,
		_w17851_,
		_w19112_,
		_w20087_
	);
	LUT4 #(
		.INIT('h2000)
	) name16040 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20088_
	);
	LUT4 #(
		.INIT('h4000)
	) name16041 (
		_w4104_,
		_w19050_,
		_w19063_,
		_w19057_,
		_w20089_
	);
	LUT2 #(
		.INIT('he)
	) name16042 (
		_w20088_,
		_w20089_,
		_w20090_
	);
	LUT4 #(
		.INIT('h2000)
	) name16043 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20091_
	);
	LUT4 #(
		.INIT('h4000)
	) name16044 (
		_w4104_,
		_w19050_,
		_w19063_,
		_w19049_,
		_w20092_
	);
	LUT2 #(
		.INIT('he)
	) name16045 (
		_w20091_,
		_w20092_,
		_w20093_
	);
	LUT4 #(
		.INIT('h2000)
	) name16046 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20094_
	);
	LUT4 #(
		.INIT('h4000)
	) name16047 (
		_w4104_,
		_w19058_,
		_w19050_,
		_w19049_,
		_w20095_
	);
	LUT2 #(
		.INIT('he)
	) name16048 (
		_w20094_,
		_w20095_,
		_w20096_
	);
	LUT4 #(
		.INIT('h2000)
	) name16049 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20097_
	);
	LUT4 #(
		.INIT('h4000)
	) name16050 (
		_w4104_,
		_w19050_,
		_w19057_,
		_w19053_,
		_w20098_
	);
	LUT2 #(
		.INIT('he)
	) name16051 (
		_w20097_,
		_w20098_,
		_w20099_
	);
	LUT4 #(
		.INIT('h2000)
	) name16052 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20100_
	);
	LUT4 #(
		.INIT('h4000)
	) name16053 (
		_w4104_,
		_w19050_,
		_w19049_,
		_w19053_,
		_w20101_
	);
	LUT2 #(
		.INIT('he)
	) name16054 (
		_w20100_,
		_w20101_,
		_w20102_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16055 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001 ,
		_w18719_,
		_w18721_,
		_w19112_,
		_w20103_
	);
	LUT3 #(
		.INIT('h40)
	) name16056 (
		\sport0_rxctl_Bcnt_reg[4]/NET0131 ,
		_w19617_,
		_w19621_,
		_w20104_
	);
	LUT2 #(
		.INIT('h1)
	) name16057 (
		\sport0_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[1]/NET0131 ,
		_w20105_
	);
	LUT4 #(
		.INIT('h0001)
	) name16058 (
		\sport0_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[1]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[2]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		_w20106_
	);
	LUT2 #(
		.INIT('h8)
	) name16059 (
		_w12841_,
		_w20106_,
		_w20107_
	);
	LUT2 #(
		.INIT('h8)
	) name16060 (
		_w20104_,
		_w20107_,
		_w20108_
	);
	LUT2 #(
		.INIT('h1)
	) name16061 (
		_w19620_,
		_w20108_,
		_w20109_
	);
	LUT2 #(
		.INIT('he)
	) name16062 (
		_w19620_,
		_w20108_,
		_w20110_
	);
	LUT2 #(
		.INIT('h2)
	) name16063 (
		_w20104_,
		_w20107_,
		_w20111_
	);
	LUT4 #(
		.INIT('h0040)
	) name16064 (
		\sport0_rxctl_Wcnt_reg[2]/NET0131 ,
		_w20104_,
		_w20105_,
		_w20107_,
		_w20112_
	);
	LUT3 #(
		.INIT('h63)
	) name16065 (
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[4]/NET0131 ,
		_w20112_,
		_w20113_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16066 (
		\sport0_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w19620_,
		_w20108_,
		_w20113_,
		_w20114_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16067 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001 ,
		_w17518_,
		_w17521_,
		_w19112_,
		_w20115_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16068 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001 ,
		_w17887_,
		_w17889_,
		_w19112_,
		_w20116_
	);
	LUT4 #(
		.INIT('h4544)
	) name16069 (
		\idma_IAL_reg/P0001 ,
		_w6774_,
		_w6894_,
		_w6896_,
		_w20117_
	);
	LUT2 #(
		.INIT('h4)
	) name16070 (
		\idma_IADi_reg[1]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w20118_
	);
	LUT2 #(
		.INIT('h6)
	) name16071 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w19999_,
		_w20119_
	);
	LUT3 #(
		.INIT('he0)
	) name16072 (
		_w12623_,
		_w19993_,
		_w20119_,
		_w20120_
	);
	LUT4 #(
		.INIT('hff02)
	) name16073 (
		_w19994_,
		_w20117_,
		_w20118_,
		_w20120_,
		_w20121_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16074 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001 ,
		_w18589_,
		_w18591_,
		_w19112_,
		_w20122_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16075 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001 ,
		_w18188_,
		_w18190_,
		_w19112_,
		_w20123_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16076 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001 ,
		_w18428_,
		_w18430_,
		_w19112_,
		_w20124_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16077 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001 ,
		_w18229_,
		_w18231_,
		_w19112_,
		_w20125_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16078 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001 ,
		_w18332_,
		_w18334_,
		_w19112_,
		_w20126_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16079 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001 ,
		_w18754_,
		_w18756_,
		_w19112_,
		_w20127_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16080 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001 ,
		_w18091_,
		_w18093_,
		_w19152_,
		_w20128_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16081 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001 ,
		_w18624_,
		_w18626_,
		_w19152_,
		_w20129_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16082 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001 ,
		_w18521_,
		_w18523_,
		_w19152_,
		_w20130_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16083 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001 ,
		_w17749_,
		_w17751_,
		_w19152_,
		_w20131_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16084 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001 ,
		_w17849_,
		_w17851_,
		_w19152_,
		_w20132_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16085 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001 ,
		_w18719_,
		_w18721_,
		_w19152_,
		_w20133_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16086 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001 ,
		_w17787_,
		_w17789_,
		_w19152_,
		_w20134_
	);
	LUT3 #(
		.INIT('h12)
	) name16087 (
		\clkc_STDcnt_reg[8]/NET0131 ,
		_w19406_,
		_w19394_,
		_w20135_
	);
	LUT4 #(
		.INIT('h152a)
	) name16088 (
		\clkc_STDcnt_reg[6]/NET0131 ,
		_w19400_,
		_w19405_,
		_w19392_,
		_w20136_
	);
	LUT4 #(
		.INIT('h0408)
	) name16089 (
		\sport0_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w12307_,
		_w20137_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16090 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001 ,
		_w17518_,
		_w17521_,
		_w19152_,
		_w20138_
	);
	LUT4 #(
		.INIT('h0408)
	) name16091 (
		\sport1_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w12723_,
		_w20139_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16092 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001 ,
		_w17887_,
		_w17889_,
		_w19152_,
		_w20140_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16093 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001 ,
		_w18589_,
		_w18591_,
		_w19152_,
		_w20141_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16094 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001 ,
		_w18188_,
		_w18190_,
		_w19152_,
		_w20142_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16095 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001 ,
		_w18428_,
		_w18430_,
		_w19152_,
		_w20143_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16096 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001 ,
		_w18229_,
		_w18231_,
		_w19152_,
		_w20144_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16097 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001 ,
		_w18332_,
		_w18334_,
		_w19152_,
		_w20145_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name16098 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001 ,
		_w18754_,
		_w18756_,
		_w19152_,
		_w20146_
	);
	LUT4 #(
		.INIT('ha800)
	) name16099 (
		\bdma_BCTL_reg[3]/NET0131 ,
		_w9414_,
		_w9415_,
		_w9423_,
		_w20147_
	);
	LUT2 #(
		.INIT('h1)
	) name16100 (
		\bdma_BRST_s2_reg/NET0131 ,
		\sice_IRST_syn_reg/P0001 ,
		_w20148_
	);
	LUT2 #(
		.INIT('hb)
	) name16101 (
		_w20147_,
		_w20148_,
		_w20149_
	);
	LUT4 #(
		.INIT('h4500)
	) name16102 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w19745_,
		_w20150_
	);
	LUT4 #(
		.INIT('h0045)
	) name16103 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w19745_,
		_w20151_
	);
	LUT3 #(
		.INIT('h02)
	) name16104 (
		_w19757_,
		_w20150_,
		_w20151_,
		_w20152_
	);
	LUT3 #(
		.INIT('hb0)
	) name16105 (
		_w7911_,
		_w7914_,
		_w19745_,
		_w20153_
	);
	LUT4 #(
		.INIT('h000e)
	) name16106 (
		_w7731_,
		_w19745_,
		_w19757_,
		_w20153_,
		_w20154_
	);
	LUT3 #(
		.INIT('ha8)
	) name16107 (
		_w19748_,
		_w20152_,
		_w20154_,
		_w20155_
	);
	LUT4 #(
		.INIT('h00fd)
	) name16108 (
		_w5041_,
		_w5049_,
		_w7748_,
		_w7756_,
		_w20156_
	);
	LUT4 #(
		.INIT('hfc54)
	) name16109 (
		_w19745_,
		_w19747_,
		_w19756_,
		_w20156_,
		_w20157_
	);
	LUT4 #(
		.INIT('hf100)
	) name16110 (
		_w7715_,
		_w7720_,
		_w19745_,
		_w20157_,
		_w20158_
	);
	LUT4 #(
		.INIT('h0203)
	) name16111 (
		_w5041_,
		_w5108_,
		_w7742_,
		_w19744_,
		_w20159_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name16112 (
		_w5041_,
		_w5108_,
		_w7776_,
		_w19744_,
		_w20160_
	);
	LUT4 #(
		.INIT('h0001)
	) name16113 (
		_w19747_,
		_w19756_,
		_w20160_,
		_w20159_,
		_w20161_
	);
	LUT3 #(
		.INIT('h54)
	) name16114 (
		_w19748_,
		_w20158_,
		_w20161_,
		_w20162_
	);
	LUT4 #(
		.INIT('h0045)
	) name16115 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w19745_,
		_w20163_
	);
	LUT3 #(
		.INIT('h10)
	) name16116 (
		_w7465_,
		_w7565_,
		_w19745_,
		_w20164_
	);
	LUT3 #(
		.INIT('h02)
	) name16117 (
		_w19757_,
		_w20164_,
		_w20163_,
		_w20165_
	);
	LUT4 #(
		.INIT('h00ac)
	) name16118 (
		_w7400_,
		_w7579_,
		_w19745_,
		_w19757_,
		_w20166_
	);
	LUT3 #(
		.INIT('ha8)
	) name16119 (
		_w19748_,
		_w20165_,
		_w20166_,
		_w20167_
	);
	LUT4 #(
		.INIT('h00fd)
	) name16120 (
		_w5041_,
		_w5049_,
		_w8093_,
		_w8101_,
		_w20168_
	);
	LUT4 #(
		.INIT('hfc54)
	) name16121 (
		_w19745_,
		_w19747_,
		_w19756_,
		_w20168_,
		_w20169_
	);
	LUT4 #(
		.INIT('hf400)
	) name16122 (
		_w8118_,
		_w8121_,
		_w19745_,
		_w20169_,
		_w20170_
	);
	LUT4 #(
		.INIT('h0203)
	) name16123 (
		_w5041_,
		_w5108_,
		_w7448_,
		_w19744_,
		_w20171_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name16124 (
		_w5041_,
		_w5108_,
		_w7413_,
		_w19744_,
		_w20172_
	);
	LUT4 #(
		.INIT('h0001)
	) name16125 (
		_w19747_,
		_w19756_,
		_w20172_,
		_w20171_,
		_w20173_
	);
	LUT3 #(
		.INIT('h54)
	) name16126 (
		_w19748_,
		_w20170_,
		_w20173_,
		_w20174_
	);
	LUT4 #(
		.INIT('h0001)
	) name16127 (
		_w20155_,
		_w20162_,
		_w20167_,
		_w20174_,
		_w20175_
	);
	LUT4 #(
		.INIT('h0045)
	) name16128 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w19745_,
		_w20176_
	);
	LUT4 #(
		.INIT('h0007)
	) name16129 (
		_w6758_,
		_w19745_,
		_w19747_,
		_w19756_,
		_w20177_
	);
	LUT2 #(
		.INIT('h4)
	) name16130 (
		_w20176_,
		_w20177_,
		_w20178_
	);
	LUT3 #(
		.INIT('hb0)
	) name16131 (
		_w6643_,
		_w6646_,
		_w19745_,
		_w20179_
	);
	LUT4 #(
		.INIT('h000e)
	) name16132 (
		_w6591_,
		_w19745_,
		_w19757_,
		_w20179_,
		_w20180_
	);
	LUT3 #(
		.INIT('ha8)
	) name16133 (
		_w19748_,
		_w20178_,
		_w20180_,
		_w20181_
	);
	LUT4 #(
		.INIT('h00fd)
	) name16134 (
		_w5041_,
		_w5049_,
		_w6608_,
		_w6616_,
		_w20182_
	);
	LUT4 #(
		.INIT('hfc54)
	) name16135 (
		_w19745_,
		_w19747_,
		_w19756_,
		_w20182_,
		_w20183_
	);
	LUT4 #(
		.INIT('hf400)
	) name16136 (
		_w6576_,
		_w6580_,
		_w19745_,
		_w20183_,
		_w20184_
	);
	LUT4 #(
		.INIT('h0203)
	) name16137 (
		_w5041_,
		_w5108_,
		_w6602_,
		_w19744_,
		_w20185_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name16138 (
		_w5041_,
		_w5108_,
		_w6637_,
		_w19744_,
		_w20186_
	);
	LUT4 #(
		.INIT('h0001)
	) name16139 (
		_w19747_,
		_w19756_,
		_w20186_,
		_w20185_,
		_w20187_
	);
	LUT3 #(
		.INIT('h54)
	) name16140 (
		_w19748_,
		_w20184_,
		_w20187_,
		_w20188_
	);
	LUT4 #(
		.INIT('h0045)
	) name16141 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w19745_,
		_w20189_
	);
	LUT3 #(
		.INIT('h10)
	) name16142 (
		_w6263_,
		_w6362_,
		_w19745_,
		_w20190_
	);
	LUT3 #(
		.INIT('h02)
	) name16143 (
		_w19757_,
		_w20190_,
		_w20189_,
		_w20191_
	);
	LUT3 #(
		.INIT('hb0)
	) name16144 (
		_w6245_,
		_w6250_,
		_w19745_,
		_w20192_
	);
	LUT4 #(
		.INIT('h000e)
	) name16145 (
		_w6555_,
		_w19745_,
		_w19757_,
		_w20192_,
		_w20193_
	);
	LUT3 #(
		.INIT('ha8)
	) name16146 (
		_w19748_,
		_w20191_,
		_w20193_,
		_w20194_
	);
	LUT4 #(
		.INIT('h00fd)
	) name16147 (
		_w5041_,
		_w5049_,
		_w6506_,
		_w6535_,
		_w20195_
	);
	LUT4 #(
		.INIT('hfc54)
	) name16148 (
		_w19745_,
		_w19747_,
		_w19756_,
		_w20195_,
		_w20196_
	);
	LUT4 #(
		.INIT('hf400)
	) name16149 (
		_w6529_,
		_w6533_,
		_w19745_,
		_w20196_,
		_w20197_
	);
	LUT4 #(
		.INIT('h0203)
	) name16150 (
		_w5041_,
		_w5108_,
		_w6522_,
		_w19744_,
		_w20198_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name16151 (
		_w5041_,
		_w5108_,
		_w6566_,
		_w19744_,
		_w20199_
	);
	LUT4 #(
		.INIT('h0001)
	) name16152 (
		_w19747_,
		_w19756_,
		_w20199_,
		_w20198_,
		_w20200_
	);
	LUT3 #(
		.INIT('h54)
	) name16153 (
		_w19748_,
		_w20197_,
		_w20200_,
		_w20201_
	);
	LUT4 #(
		.INIT('h0001)
	) name16154 (
		_w20181_,
		_w20188_,
		_w20194_,
		_w20201_,
		_w20202_
	);
	LUT2 #(
		.INIT('h8)
	) name16155 (
		_w20175_,
		_w20202_,
		_w20203_
	);
	LUT3 #(
		.INIT('h54)
	) name16156 (
		_w15328_,
		_w19758_,
		_w19765_,
		_w20204_
	);
	LUT3 #(
		.INIT('h01)
	) name16157 (
		_w7465_,
		_w7565_,
		_w19745_,
		_w20205_
	);
	LUT4 #(
		.INIT('h4500)
	) name16158 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w19745_,
		_w20206_
	);
	LUT3 #(
		.INIT('h02)
	) name16159 (
		_w19757_,
		_w20206_,
		_w20205_,
		_w20207_
	);
	LUT4 #(
		.INIT('h00ca)
	) name16160 (
		_w7400_,
		_w7579_,
		_w19745_,
		_w19757_,
		_w20208_
	);
	LUT3 #(
		.INIT('ha8)
	) name16161 (
		_w19748_,
		_w20207_,
		_w20208_,
		_w20209_
	);
	LUT4 #(
		.INIT('h00fd)
	) name16162 (
		_w5041_,
		_w5049_,
		_w7419_,
		_w7427_,
		_w20210_
	);
	LUT4 #(
		.INIT('hfc54)
	) name16163 (
		_w19745_,
		_w19747_,
		_w19756_,
		_w20210_,
		_w20211_
	);
	LUT4 #(
		.INIT('hf400)
	) name16164 (
		_w7386_,
		_w7390_,
		_w19745_,
		_w20211_,
		_w20212_
	);
	LUT4 #(
		.INIT('h0203)
	) name16165 (
		_w5041_,
		_w5108_,
		_w7413_,
		_w19744_,
		_w20213_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name16166 (
		_w5041_,
		_w5108_,
		_w7448_,
		_w19744_,
		_w20214_
	);
	LUT4 #(
		.INIT('h0001)
	) name16167 (
		_w19747_,
		_w19756_,
		_w20214_,
		_w20213_,
		_w20215_
	);
	LUT3 #(
		.INIT('h54)
	) name16168 (
		_w19748_,
		_w20212_,
		_w20215_,
		_w20216_
	);
	LUT4 #(
		.INIT('h0045)
	) name16169 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w19745_,
		_w20217_
	);
	LUT4 #(
		.INIT('h4500)
	) name16170 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w19745_,
		_w20218_
	);
	LUT3 #(
		.INIT('h02)
	) name16171 (
		_w19757_,
		_w20218_,
		_w20217_,
		_w20219_
	);
	LUT3 #(
		.INIT('h0b)
	) name16172 (
		_w7911_,
		_w7914_,
		_w19745_,
		_w20220_
	);
	LUT4 #(
		.INIT('h000b)
	) name16173 (
		_w7731_,
		_w19745_,
		_w19757_,
		_w20220_,
		_w20221_
	);
	LUT3 #(
		.INIT('ha8)
	) name16174 (
		_w19748_,
		_w20219_,
		_w20221_,
		_w20222_
	);
	LUT4 #(
		.INIT('h00fd)
	) name16175 (
		_w5041_,
		_w5049_,
		_w8061_,
		_w8069_,
		_w20223_
	);
	LUT4 #(
		.INIT('hfc54)
	) name16176 (
		_w19745_,
		_w19747_,
		_w19756_,
		_w20223_,
		_w20224_
	);
	LUT4 #(
		.INIT('hf400)
	) name16177 (
		_w8052_,
		_w8055_,
		_w19745_,
		_w20224_,
		_w20225_
	);
	LUT4 #(
		.INIT('h0203)
	) name16178 (
		_w5041_,
		_w5108_,
		_w7776_,
		_w19744_,
		_w20226_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name16179 (
		_w5041_,
		_w5108_,
		_w7742_,
		_w19744_,
		_w20227_
	);
	LUT4 #(
		.INIT('h0001)
	) name16180 (
		_w19747_,
		_w19756_,
		_w20227_,
		_w20226_,
		_w20228_
	);
	LUT3 #(
		.INIT('h54)
	) name16181 (
		_w19748_,
		_w20225_,
		_w20228_,
		_w20229_
	);
	LUT4 #(
		.INIT('h0001)
	) name16182 (
		_w20209_,
		_w20216_,
		_w20222_,
		_w20229_,
		_w20230_
	);
	LUT4 #(
		.INIT('h0045)
	) name16183 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w19745_,
		_w20231_
	);
	LUT3 #(
		.INIT('h10)
	) name16184 (
		_w7140_,
		_w7240_,
		_w19745_,
		_w20232_
	);
	LUT3 #(
		.INIT('h02)
	) name16185 (
		_w19757_,
		_w20232_,
		_w20231_,
		_w20233_
	);
	LUT3 #(
		.INIT('h0b)
	) name16186 (
		_w7122_,
		_w7126_,
		_w19745_,
		_w20234_
	);
	LUT4 #(
		.INIT('h001f)
	) name16187 (
		_w7062_,
		_w7067_,
		_w19745_,
		_w19757_,
		_w20235_
	);
	LUT4 #(
		.INIT('h8a88)
	) name16188 (
		_w19748_,
		_w20233_,
		_w20234_,
		_w20235_,
		_w20236_
	);
	LUT4 #(
		.INIT('h00fd)
	) name16189 (
		_w5041_,
		_w5049_,
		_w8132_,
		_w8143_,
		_w20237_
	);
	LUT4 #(
		.INIT('hfc54)
	) name16190 (
		_w19745_,
		_w19747_,
		_w19756_,
		_w20237_,
		_w20238_
	);
	LUT4 #(
		.INIT('hf400)
	) name16191 (
		_w8157_,
		_w8162_,
		_w19745_,
		_w20238_,
		_w20239_
	);
	LUT4 #(
		.INIT('h0203)
	) name16192 (
		_w5041_,
		_w5108_,
		_w7077_,
		_w19744_,
		_w20240_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name16193 (
		_w5041_,
		_w5108_,
		_w7108_,
		_w19744_,
		_w20241_
	);
	LUT4 #(
		.INIT('h0001)
	) name16194 (
		_w19747_,
		_w19756_,
		_w20241_,
		_w20240_,
		_w20242_
	);
	LUT4 #(
		.INIT('h2223)
	) name16195 (
		_w19748_,
		_w20236_,
		_w20239_,
		_w20242_,
		_w20243_
	);
	LUT4 #(
		.INIT('h0045)
	) name16196 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w19745_,
		_w20244_
	);
	LUT3 #(
		.INIT('h10)
	) name16197 (
		_w5937_,
		_w6038_,
		_w19745_,
		_w20245_
	);
	LUT3 #(
		.INIT('h02)
	) name16198 (
		_w19757_,
		_w20245_,
		_w20244_,
		_w20246_
	);
	LUT3 #(
		.INIT('h0b)
	) name16199 (
		_w6204_,
		_w6207_,
		_w19745_,
		_w20247_
	);
	LUT4 #(
		.INIT('h004f)
	) name16200 (
		_w5920_,
		_w5924_,
		_w19745_,
		_w19757_,
		_w20248_
	);
	LUT4 #(
		.INIT('h8a88)
	) name16201 (
		_w19748_,
		_w20246_,
		_w20247_,
		_w20248_,
		_w20249_
	);
	LUT4 #(
		.INIT('h00fd)
	) name16202 (
		_w5041_,
		_w5049_,
		_w6181_,
		_w6218_,
		_w20250_
	);
	LUT4 #(
		.INIT('hfc54)
	) name16203 (
		_w19745_,
		_w19747_,
		_w19756_,
		_w20250_,
		_w20251_
	);
	LUT4 #(
		.INIT('hf100)
	) name16204 (
		_w6209_,
		_w6215_,
		_w19745_,
		_w20251_,
		_w20252_
	);
	LUT4 #(
		.INIT('h0203)
	) name16205 (
		_w5041_,
		_w5108_,
		_w6197_,
		_w19744_,
		_w20253_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name16206 (
		_w5041_,
		_w5108_,
		_w6237_,
		_w19744_,
		_w20254_
	);
	LUT4 #(
		.INIT('h0001)
	) name16207 (
		_w19747_,
		_w19756_,
		_w20254_,
		_w20253_,
		_w20255_
	);
	LUT4 #(
		.INIT('h2223)
	) name16208 (
		_w19748_,
		_w20249_,
		_w20252_,
		_w20255_,
		_w20256_
	);
	LUT2 #(
		.INIT('h8)
	) name16209 (
		_w20243_,
		_w20256_,
		_w20257_
	);
	LUT3 #(
		.INIT('h80)
	) name16210 (
		_w20204_,
		_w20230_,
		_w20257_,
		_w20258_
	);
	LUT2 #(
		.INIT('h7)
	) name16211 (
		_w20203_,
		_w20258_,
		_w20259_
	);
	LUT4 #(
		.INIT('h6663)
	) name16212 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		_w12821_,
		_w19997_,
		_w20260_
	);
	LUT3 #(
		.INIT('h7f)
	) name16213 (
		_w12619_,
		_w12623_,
		_w20260_,
		_w20261_
	);
	LUT3 #(
		.INIT('ha8)
	) name16214 (
		_w4142_,
		_w15960_,
		_w15961_,
		_w20262_
	);
	LUT4 #(
		.INIT('h0400)
	) name16215 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[12]/NET0131 ,
		_w20263_
	);
	LUT4 #(
		.INIT('h2333)
	) name16216 (
		\tm_tpr_reg_DO_reg[12]/NET0131 ,
		_w12803_,
		_w12801_,
		_w14102_,
		_w20264_
	);
	LUT4 #(
		.INIT('hde00)
	) name16217 (
		\tm_TCR_TMP_reg[12]/NET0131 ,
		_w14103_,
		_w15995_,
		_w20264_,
		_w20265_
	);
	LUT2 #(
		.INIT('he)
	) name16218 (
		_w20263_,
		_w20265_,
		_w20266_
	);
	LUT2 #(
		.INIT('h2)
	) name16219 (
		\sport1_rxctl_LMcnt_reg[4]/NET0131 ,
		_w18879_,
		_w20267_
	);
	LUT3 #(
		.INIT('hfe)
	) name16220 (
		_w19498_,
		_w19501_,
		_w20267_,
		_w20268_
	);
	LUT2 #(
		.INIT('h2)
	) name16221 (
		\sport0_rxctl_LMcnt_reg[4]/NET0131 ,
		_w18893_,
		_w20269_
	);
	LUT3 #(
		.INIT('hfe)
	) name16222 (
		_w19620_,
		_w19623_,
		_w20269_,
		_w20270_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name16223 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w4063_,
		_w5030_,
		_w20271_
	);
	LUT3 #(
		.INIT('h20)
	) name16224 (
		_w4857_,
		_w4981_,
		_w4986_,
		_w20272_
	);
	LUT2 #(
		.INIT('h1)
	) name16225 (
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		_w4857_,
		_w20273_
	);
	LUT3 #(
		.INIT('h0b)
	) name16226 (
		_w20271_,
		_w20272_,
		_w20273_,
		_w20274_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name16227 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w4063_,
		_w5030_,
		_w20275_
	);
	LUT3 #(
		.INIT('h20)
	) name16228 (
		_w4857_,
		_w4994_,
		_w4997_,
		_w20276_
	);
	LUT2 #(
		.INIT('h1)
	) name16229 (
		\core_dag_ilm2reg_IL_E_reg[0]/P0001 ,
		_w4857_,
		_w20277_
	);
	LUT3 #(
		.INIT('h0b)
	) name16230 (
		_w20275_,
		_w20276_,
		_w20277_,
		_w20278_
	);
	LUT4 #(
		.INIT('hf53f)
	) name16231 (
		_w16061_,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20279_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name16232 (
		_w16060_,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20280_
	);
	LUT2 #(
		.INIT('h8)
	) name16233 (
		_w20279_,
		_w20280_,
		_w20281_
	);
	LUT4 #(
		.INIT('h0045)
	) name16234 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w20281_,
		_w20282_
	);
	LUT4 #(
		.INIT('h0020)
	) name16235 (
		\core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20283_
	);
	LUT3 #(
		.INIT('h0b)
	) name16236 (
		_w12398_,
		_w13536_,
		_w20283_,
		_w20284_
	);
	LUT4 #(
		.INIT('h0200)
	) name16237 (
		\core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20285_
	);
	LUT4 #(
		.INIT('h0002)
	) name16238 (
		\core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20286_
	);
	LUT4 #(
		.INIT('h2000)
	) name16239 (
		\core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20287_
	);
	LUT3 #(
		.INIT('h01)
	) name16240 (
		_w20286_,
		_w20287_,
		_w20285_,
		_w20288_
	);
	LUT2 #(
		.INIT('h8)
	) name16241 (
		_w20284_,
		_w20288_,
		_w20289_
	);
	LUT3 #(
		.INIT('h10)
	) name16242 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20290_
	);
	LUT3 #(
		.INIT('h0b)
	) name16243 (
		_w20282_,
		_w20289_,
		_w20290_,
		_w20291_
	);
	LUT4 #(
		.INIT('h0045)
	) name16244 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w20281_,
		_w20292_
	);
	LUT4 #(
		.INIT('h0020)
	) name16245 (
		\core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20293_
	);
	LUT3 #(
		.INIT('h0b)
	) name16246 (
		_w12398_,
		_w13536_,
		_w20293_,
		_w20294_
	);
	LUT4 #(
		.INIT('h0200)
	) name16247 (
		\core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20295_
	);
	LUT4 #(
		.INIT('h0002)
	) name16248 (
		\core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20296_
	);
	LUT4 #(
		.INIT('h2000)
	) name16249 (
		\core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20297_
	);
	LUT3 #(
		.INIT('h01)
	) name16250 (
		_w20296_,
		_w20297_,
		_w20295_,
		_w20298_
	);
	LUT2 #(
		.INIT('h8)
	) name16251 (
		_w20294_,
		_w20298_,
		_w20299_
	);
	LUT3 #(
		.INIT('h10)
	) name16252 (
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20300_
	);
	LUT3 #(
		.INIT('h0b)
	) name16253 (
		_w20292_,
		_w20299_,
		_w20300_,
		_w20301_
	);
	LUT4 #(
		.INIT('h0045)
	) name16254 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w20281_,
		_w20302_
	);
	LUT4 #(
		.INIT('h0002)
	) name16255 (
		\core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20303_
	);
	LUT3 #(
		.INIT('h0b)
	) name16256 (
		_w12398_,
		_w13536_,
		_w20303_,
		_w20304_
	);
	LUT4 #(
		.INIT('h2000)
	) name16257 (
		\core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20305_
	);
	LUT4 #(
		.INIT('h0020)
	) name16258 (
		\core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20306_
	);
	LUT4 #(
		.INIT('h0200)
	) name16259 (
		\core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20307_
	);
	LUT3 #(
		.INIT('h01)
	) name16260 (
		_w20306_,
		_w20307_,
		_w20305_,
		_w20308_
	);
	LUT2 #(
		.INIT('h8)
	) name16261 (
		_w20304_,
		_w20308_,
		_w20309_
	);
	LUT3 #(
		.INIT('h10)
	) name16262 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20310_
	);
	LUT3 #(
		.INIT('h0b)
	) name16263 (
		_w20302_,
		_w20309_,
		_w20310_,
		_w20311_
	);
	LUT4 #(
		.INIT('h0045)
	) name16264 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w20281_,
		_w20312_
	);
	LUT4 #(
		.INIT('h0020)
	) name16265 (
		\core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20313_
	);
	LUT3 #(
		.INIT('h0b)
	) name16266 (
		_w12398_,
		_w13536_,
		_w20313_,
		_w20314_
	);
	LUT4 #(
		.INIT('h0200)
	) name16267 (
		\core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20315_
	);
	LUT4 #(
		.INIT('h0002)
	) name16268 (
		\core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20316_
	);
	LUT4 #(
		.INIT('h2000)
	) name16269 (
		\core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20317_
	);
	LUT3 #(
		.INIT('h01)
	) name16270 (
		_w20316_,
		_w20317_,
		_w20315_,
		_w20318_
	);
	LUT2 #(
		.INIT('h8)
	) name16271 (
		_w20314_,
		_w20318_,
		_w20319_
	);
	LUT3 #(
		.INIT('h10)
	) name16272 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20320_
	);
	LUT3 #(
		.INIT('h0b)
	) name16273 (
		_w20312_,
		_w20319_,
		_w20320_,
		_w20321_
	);
	LUT4 #(
		.INIT('h0045)
	) name16274 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w20281_,
		_w20322_
	);
	LUT4 #(
		.INIT('h0020)
	) name16275 (
		\core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20323_
	);
	LUT3 #(
		.INIT('h0b)
	) name16276 (
		_w12398_,
		_w13536_,
		_w20323_,
		_w20324_
	);
	LUT4 #(
		.INIT('h0200)
	) name16277 (
		\core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20325_
	);
	LUT4 #(
		.INIT('h0002)
	) name16278 (
		\core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20326_
	);
	LUT4 #(
		.INIT('h2000)
	) name16279 (
		\core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20327_
	);
	LUT3 #(
		.INIT('h01)
	) name16280 (
		_w20326_,
		_w20327_,
		_w20325_,
		_w20328_
	);
	LUT2 #(
		.INIT('h8)
	) name16281 (
		_w20324_,
		_w20328_,
		_w20329_
	);
	LUT3 #(
		.INIT('h10)
	) name16282 (
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20330_
	);
	LUT3 #(
		.INIT('h0b)
	) name16283 (
		_w20322_,
		_w20329_,
		_w20330_,
		_w20331_
	);
	LUT4 #(
		.INIT('h0045)
	) name16284 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w20281_,
		_w20332_
	);
	LUT4 #(
		.INIT('h0002)
	) name16285 (
		\core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20333_
	);
	LUT3 #(
		.INIT('h0b)
	) name16286 (
		_w12398_,
		_w13536_,
		_w20333_,
		_w20334_
	);
	LUT4 #(
		.INIT('h2000)
	) name16287 (
		\core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20335_
	);
	LUT4 #(
		.INIT('h0020)
	) name16288 (
		\core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20336_
	);
	LUT4 #(
		.INIT('h0200)
	) name16289 (
		\core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20337_
	);
	LUT3 #(
		.INIT('h01)
	) name16290 (
		_w20336_,
		_w20337_,
		_w20335_,
		_w20338_
	);
	LUT2 #(
		.INIT('h8)
	) name16291 (
		_w20334_,
		_w20338_,
		_w20339_
	);
	LUT3 #(
		.INIT('h10)
	) name16292 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20340_
	);
	LUT3 #(
		.INIT('h0b)
	) name16293 (
		_w20332_,
		_w20339_,
		_w20340_,
		_w20341_
	);
	LUT4 #(
		.INIT('h0045)
	) name16294 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w20281_,
		_w20342_
	);
	LUT4 #(
		.INIT('h0020)
	) name16295 (
		\core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20343_
	);
	LUT3 #(
		.INIT('h0b)
	) name16296 (
		_w12398_,
		_w13536_,
		_w20343_,
		_w20344_
	);
	LUT4 #(
		.INIT('h0200)
	) name16297 (
		\core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20345_
	);
	LUT4 #(
		.INIT('h0002)
	) name16298 (
		\core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20346_
	);
	LUT4 #(
		.INIT('h2000)
	) name16299 (
		\core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20347_
	);
	LUT3 #(
		.INIT('h01)
	) name16300 (
		_w20346_,
		_w20347_,
		_w20345_,
		_w20348_
	);
	LUT2 #(
		.INIT('h8)
	) name16301 (
		_w20344_,
		_w20348_,
		_w20349_
	);
	LUT3 #(
		.INIT('h10)
	) name16302 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20350_
	);
	LUT3 #(
		.INIT('h0b)
	) name16303 (
		_w20342_,
		_w20349_,
		_w20350_,
		_w20351_
	);
	LUT2 #(
		.INIT('h1)
	) name16304 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w4857_,
		_w20352_
	);
	LUT3 #(
		.INIT('h20)
	) name16305 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w4061_,
		_w4062_,
		_w20353_
	);
	LUT4 #(
		.INIT('h0020)
	) name16306 (
		_w4857_,
		_w4981_,
		_w4986_,
		_w20353_,
		_w20354_
	);
	LUT2 #(
		.INIT('h1)
	) name16307 (
		_w20352_,
		_w20354_,
		_w20355_
	);
	LUT2 #(
		.INIT('h1)
	) name16308 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w4857_,
		_w20356_
	);
	LUT3 #(
		.INIT('h20)
	) name16309 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w4061_,
		_w4062_,
		_w20357_
	);
	LUT4 #(
		.INIT('h0020)
	) name16310 (
		_w4857_,
		_w4994_,
		_w4997_,
		_w20357_,
		_w20358_
	);
	LUT2 #(
		.INIT('h1)
	) name16311 (
		_w20356_,
		_w20358_,
		_w20359_
	);
	LUT4 #(
		.INIT('h0001)
	) name16312 (
		_w20352_,
		_w20354_,
		_w20356_,
		_w20358_,
		_w20360_
	);
	LUT4 #(
		.INIT('heee0)
	) name16313 (
		_w20352_,
		_w20354_,
		_w20356_,
		_w20358_,
		_w20361_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name16314 (
		_w16073_,
		_w16074_,
		_w20355_,
		_w20359_,
		_w20362_
	);
	LUT4 #(
		.INIT('h1110)
	) name16315 (
		_w20352_,
		_w20354_,
		_w20356_,
		_w20358_,
		_w20363_
	);
	LUT4 #(
		.INIT('h000e)
	) name16316 (
		_w20352_,
		_w20354_,
		_w20356_,
		_w20358_,
		_w20364_
	);
	LUT4 #(
		.INIT('hf35f)
	) name16317 (
		_w16071_,
		_w16072_,
		_w20355_,
		_w20359_,
		_w20365_
	);
	LUT2 #(
		.INIT('h8)
	) name16318 (
		_w20362_,
		_w20365_,
		_w20366_
	);
	LUT4 #(
		.INIT('h0045)
	) name16319 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w20366_,
		_w20367_
	);
	LUT3 #(
		.INIT('h20)
	) name16320 (
		\core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20368_
	);
	LUT3 #(
		.INIT('h20)
	) name16321 (
		\core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20369_
	);
	LUT3 #(
		.INIT('h20)
	) name16322 (
		\core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20370_
	);
	LUT3 #(
		.INIT('h20)
	) name16323 (
		\core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20371_
	);
	LUT4 #(
		.INIT('h0001)
	) name16324 (
		_w20368_,
		_w20369_,
		_w20370_,
		_w20371_,
		_w20372_
	);
	LUT2 #(
		.INIT('h4)
	) name16325 (
		_w13546_,
		_w20372_,
		_w20373_
	);
	LUT2 #(
		.INIT('h4)
	) name16326 (
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		_w13546_,
		_w20374_
	);
	LUT3 #(
		.INIT('h0b)
	) name16327 (
		_w20367_,
		_w20373_,
		_w20374_,
		_w20375_
	);
	LUT4 #(
		.INIT('h0045)
	) name16328 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w20366_,
		_w20376_
	);
	LUT3 #(
		.INIT('h20)
	) name16329 (
		\core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20377_
	);
	LUT3 #(
		.INIT('h20)
	) name16330 (
		\core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20378_
	);
	LUT3 #(
		.INIT('h20)
	) name16331 (
		\core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20379_
	);
	LUT3 #(
		.INIT('h20)
	) name16332 (
		\core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20380_
	);
	LUT4 #(
		.INIT('h0001)
	) name16333 (
		_w20377_,
		_w20378_,
		_w20379_,
		_w20380_,
		_w20381_
	);
	LUT2 #(
		.INIT('h4)
	) name16334 (
		_w13546_,
		_w20381_,
		_w20382_
	);
	LUT2 #(
		.INIT('h4)
	) name16335 (
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		_w13546_,
		_w20383_
	);
	LUT3 #(
		.INIT('h0b)
	) name16336 (
		_w20376_,
		_w20382_,
		_w20383_,
		_w20384_
	);
	LUT4 #(
		.INIT('h0045)
	) name16337 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w20366_,
		_w20385_
	);
	LUT3 #(
		.INIT('h20)
	) name16338 (
		\core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20386_
	);
	LUT3 #(
		.INIT('h20)
	) name16339 (
		\core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20387_
	);
	LUT3 #(
		.INIT('h20)
	) name16340 (
		\core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20388_
	);
	LUT3 #(
		.INIT('h20)
	) name16341 (
		\core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20389_
	);
	LUT4 #(
		.INIT('h0001)
	) name16342 (
		_w20386_,
		_w20387_,
		_w20388_,
		_w20389_,
		_w20390_
	);
	LUT2 #(
		.INIT('h4)
	) name16343 (
		_w13546_,
		_w20390_,
		_w20391_
	);
	LUT2 #(
		.INIT('h4)
	) name16344 (
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w13546_,
		_w20392_
	);
	LUT3 #(
		.INIT('h0b)
	) name16345 (
		_w20385_,
		_w20391_,
		_w20392_,
		_w20393_
	);
	LUT4 #(
		.INIT('h0045)
	) name16346 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w20366_,
		_w20394_
	);
	LUT3 #(
		.INIT('h20)
	) name16347 (
		\core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20395_
	);
	LUT3 #(
		.INIT('h20)
	) name16348 (
		\core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20396_
	);
	LUT3 #(
		.INIT('h20)
	) name16349 (
		\core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20397_
	);
	LUT3 #(
		.INIT('h20)
	) name16350 (
		\core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20398_
	);
	LUT4 #(
		.INIT('h0001)
	) name16351 (
		_w20395_,
		_w20396_,
		_w20397_,
		_w20398_,
		_w20399_
	);
	LUT2 #(
		.INIT('h4)
	) name16352 (
		_w13546_,
		_w20399_,
		_w20400_
	);
	LUT2 #(
		.INIT('h4)
	) name16353 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		_w13546_,
		_w20401_
	);
	LUT3 #(
		.INIT('h0b)
	) name16354 (
		_w20394_,
		_w20400_,
		_w20401_,
		_w20402_
	);
	LUT4 #(
		.INIT('h0045)
	) name16355 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w20366_,
		_w20403_
	);
	LUT3 #(
		.INIT('h20)
	) name16356 (
		\core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20404_
	);
	LUT3 #(
		.INIT('h20)
	) name16357 (
		\core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20405_
	);
	LUT3 #(
		.INIT('h20)
	) name16358 (
		\core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20406_
	);
	LUT3 #(
		.INIT('h20)
	) name16359 (
		\core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20407_
	);
	LUT4 #(
		.INIT('h0001)
	) name16360 (
		_w20404_,
		_w20405_,
		_w20406_,
		_w20407_,
		_w20408_
	);
	LUT2 #(
		.INIT('h4)
	) name16361 (
		_w13546_,
		_w20408_,
		_w20409_
	);
	LUT2 #(
		.INIT('h4)
	) name16362 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		_w13546_,
		_w20410_
	);
	LUT3 #(
		.INIT('h0b)
	) name16363 (
		_w20403_,
		_w20409_,
		_w20410_,
		_w20411_
	);
	LUT4 #(
		.INIT('h0045)
	) name16364 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w20366_,
		_w20412_
	);
	LUT3 #(
		.INIT('h20)
	) name16365 (
		\core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20413_
	);
	LUT3 #(
		.INIT('h20)
	) name16366 (
		\core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20414_
	);
	LUT3 #(
		.INIT('h20)
	) name16367 (
		\core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20415_
	);
	LUT3 #(
		.INIT('h20)
	) name16368 (
		\core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20416_
	);
	LUT4 #(
		.INIT('h0001)
	) name16369 (
		_w20413_,
		_w20414_,
		_w20415_,
		_w20416_,
		_w20417_
	);
	LUT2 #(
		.INIT('h4)
	) name16370 (
		_w13546_,
		_w20417_,
		_w20418_
	);
	LUT2 #(
		.INIT('h4)
	) name16371 (
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w13546_,
		_w20419_
	);
	LUT3 #(
		.INIT('h0b)
	) name16372 (
		_w20412_,
		_w20418_,
		_w20419_,
		_w20420_
	);
	LUT4 #(
		.INIT('h0045)
	) name16373 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w20366_,
		_w20421_
	);
	LUT3 #(
		.INIT('h20)
	) name16374 (
		\core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20422_
	);
	LUT3 #(
		.INIT('h20)
	) name16375 (
		\core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20423_
	);
	LUT3 #(
		.INIT('h20)
	) name16376 (
		\core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20424_
	);
	LUT3 #(
		.INIT('h20)
	) name16377 (
		\core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20425_
	);
	LUT4 #(
		.INIT('h0001)
	) name16378 (
		_w20422_,
		_w20423_,
		_w20424_,
		_w20425_,
		_w20426_
	);
	LUT2 #(
		.INIT('h4)
	) name16379 (
		_w13546_,
		_w20426_,
		_w20427_
	);
	LUT2 #(
		.INIT('h4)
	) name16380 (
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		_w13546_,
		_w20428_
	);
	LUT3 #(
		.INIT('h0b)
	) name16381 (
		_w20421_,
		_w20427_,
		_w20428_,
		_w20429_
	);
	LUT4 #(
		.INIT('h0045)
	) name16382 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w20366_,
		_w20430_
	);
	LUT3 #(
		.INIT('h20)
	) name16383 (
		\core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20431_
	);
	LUT3 #(
		.INIT('h20)
	) name16384 (
		\core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20432_
	);
	LUT3 #(
		.INIT('h20)
	) name16385 (
		\core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20433_
	);
	LUT3 #(
		.INIT('h20)
	) name16386 (
		\core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20434_
	);
	LUT4 #(
		.INIT('h0001)
	) name16387 (
		_w20431_,
		_w20432_,
		_w20433_,
		_w20434_,
		_w20435_
	);
	LUT2 #(
		.INIT('h4)
	) name16388 (
		_w13546_,
		_w20435_,
		_w20436_
	);
	LUT2 #(
		.INIT('h4)
	) name16389 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		_w13546_,
		_w20437_
	);
	LUT3 #(
		.INIT('h0b)
	) name16390 (
		_w20430_,
		_w20436_,
		_w20437_,
		_w20438_
	);
	LUT4 #(
		.INIT('hc444)
	) name16391 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20439_
	);
	LUT2 #(
		.INIT('h1)
	) name16392 (
		_w12273_,
		_w12272_,
		_w20440_
	);
	LUT3 #(
		.INIT('h40)
	) name16393 (
		_w12270_,
		_w12279_,
		_w20440_,
		_w20441_
	);
	LUT4 #(
		.INIT('ha088)
	) name16394 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		\core_c_psq_Iflag_reg[12]/NET0131 ,
		\core_c_psq_Iflag_reg[2]/NET0131 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w20442_
	);
	LUT2 #(
		.INIT('h4)
	) name16395 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w20442_,
		_w20443_
	);
	LUT2 #(
		.INIT('h1)
	) name16396 (
		\core_c_psq_Iflag_reg[11]/NET0131 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w20444_
	);
	LUT4 #(
		.INIT('h080a)
	) name16397 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		\core_c_psq_Iflag_reg[1]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w20445_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16398 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w20442_,
		_w20444_,
		_w20445_,
		_w20446_
	);
	LUT3 #(
		.INIT('h08)
	) name16399 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_Iflag_reg[0]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w20447_
	);
	LUT3 #(
		.INIT('h08)
	) name16400 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_Iflag_reg[3]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w20448_
	);
	LUT2 #(
		.INIT('h1)
	) name16401 (
		_w20447_,
		_w20448_,
		_w20449_
	);
	LUT2 #(
		.INIT('h8)
	) name16402 (
		_w20446_,
		_w20449_,
		_w20450_
	);
	LUT4 #(
		.INIT('h8ddd)
	) name16403 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_c_psq_TRAP_R_L_reg/NET0131 ,
		_w20441_,
		_w20450_,
		_w20451_
	);
	LUT2 #(
		.INIT('h8)
	) name16404 (
		_w12267_,
		_w20451_,
		_w20452_
	);
	LUT4 #(
		.INIT('h1000)
	) name16405 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4428_,
		_w8172_,
		_w20452_,
		_w20453_
	);
	LUT2 #(
		.INIT('he)
	) name16406 (
		_w20439_,
		_w20453_,
		_w20454_
	);
	LUT4 #(
		.INIT('h8a88)
	) name16407 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w7927_,
		_w8040_,
		_w8042_,
		_w20455_
	);
	LUT4 #(
		.INIT('h0800)
	) name16408 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001 ,
		_w20456_
	);
	LUT4 #(
		.INIT('h0200)
	) name16409 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001 ,
		_w20457_
	);
	LUT4 #(
		.INIT('h0400)
	) name16410 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001 ,
		_w20458_
	);
	LUT4 #(
		.INIT('h0100)
	) name16411 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001 ,
		_w20459_
	);
	LUT4 #(
		.INIT('h0001)
	) name16412 (
		_w20456_,
		_w20457_,
		_w20458_,
		_w20459_,
		_w20460_
	);
	LUT4 #(
		.INIT('h4000)
	) name16413 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001 ,
		_w20461_
	);
	LUT4 #(
		.INIT('h1000)
	) name16414 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001 ,
		_w20462_
	);
	LUT4 #(
		.INIT('h2000)
	) name16415 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001 ,
		_w20463_
	);
	LUT4 #(
		.INIT('h0001)
	) name16416 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w20461_,
		_w20462_,
		_w20463_,
		_w20464_
	);
	LUT2 #(
		.INIT('h8)
	) name16417 (
		_w20460_,
		_w20464_,
		_w20465_
	);
	LUT4 #(
		.INIT('h0001)
	) name16418 (
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		\core_c_psq_Iact_E_reg[3]/NET0131 ,
		_w20466_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name16419 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		_w20466_,
		_w20467_
	);
	LUT4 #(
		.INIT('h0045)
	) name16420 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4094_,
		_w4097_,
		_w20467_,
		_w20468_
	);
	LUT2 #(
		.INIT('h2)
	) name16421 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w20468_,
		_w20469_
	);
	LUT2 #(
		.INIT('h4)
	) name16422 (
		_w19947_,
		_w20469_,
		_w20470_
	);
	LUT4 #(
		.INIT('hff02)
	) name16423 (
		_w19947_,
		_w20455_,
		_w20465_,
		_w20470_,
		_w20471_
	);
	LUT4 #(
		.INIT('h8a88)
	) name16424 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w7592_,
		_w7707_,
		_w7709_,
		_w20472_
	);
	LUT4 #(
		.INIT('h0800)
	) name16425 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001 ,
		_w20473_
	);
	LUT4 #(
		.INIT('h2000)
	) name16426 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001 ,
		_w20474_
	);
	LUT4 #(
		.INIT('h4000)
	) name16427 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001 ,
		_w20475_
	);
	LUT4 #(
		.INIT('h0100)
	) name16428 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001 ,
		_w20476_
	);
	LUT4 #(
		.INIT('h0001)
	) name16429 (
		_w20473_,
		_w20474_,
		_w20475_,
		_w20476_,
		_w20477_
	);
	LUT4 #(
		.INIT('h0400)
	) name16430 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001 ,
		_w20478_
	);
	LUT4 #(
		.INIT('h1000)
	) name16431 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001 ,
		_w20479_
	);
	LUT4 #(
		.INIT('h0200)
	) name16432 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001 ,
		_w20480_
	);
	LUT4 #(
		.INIT('h0001)
	) name16433 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w20478_,
		_w20479_,
		_w20480_,
		_w20481_
	);
	LUT2 #(
		.INIT('h8)
	) name16434 (
		_w20477_,
		_w20481_,
		_w20482_
	);
	LUT3 #(
		.INIT('h8a)
	) name16435 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		_w20466_,
		_w20483_
	);
	LUT4 #(
		.INIT('h0045)
	) name16436 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4094_,
		_w4097_,
		_w20483_,
		_w20484_
	);
	LUT2 #(
		.INIT('h2)
	) name16437 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w20484_,
		_w20485_
	);
	LUT2 #(
		.INIT('h4)
	) name16438 (
		_w19947_,
		_w20485_,
		_w20486_
	);
	LUT4 #(
		.INIT('hff02)
	) name16439 (
		_w19947_,
		_w20472_,
		_w20482_,
		_w20486_,
		_w20487_
	);
	LUT4 #(
		.INIT('h1000)
	) name16440 (
		\core_c_dec_MFPSQ_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20488_
	);
	LUT3 #(
		.INIT('h3e)
	) name16441 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w20489_
	);
	LUT4 #(
		.INIT('h5400)
	) name16442 (
		_w19040_,
		_w19231_,
		_w19232_,
		_w20489_,
		_w20490_
	);
	LUT2 #(
		.INIT('h8)
	) name16443 (
		_w19687_,
		_w20490_,
		_w20491_
	);
	LUT4 #(
		.INIT('h0002)
	) name16444 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w19040_,
		_w19236_,
		_w19237_,
		_w20492_
	);
	LUT2 #(
		.INIT('h8)
	) name16445 (
		_w19694_,
		_w20492_,
		_w20493_
	);
	LUT2 #(
		.INIT('h8)
	) name16446 (
		_w19691_,
		_w20492_,
		_w20494_
	);
	LUT3 #(
		.INIT('h1f)
	) name16447 (
		_w19691_,
		_w19694_,
		_w20492_,
		_w20495_
	);
	LUT2 #(
		.INIT('h4)
	) name16448 (
		_w20491_,
		_w20495_,
		_w20496_
	);
	LUT2 #(
		.INIT('h8)
	) name16449 (
		_w19683_,
		_w20492_,
		_w20497_
	);
	LUT3 #(
		.INIT('h70)
	) name16450 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w9931_,
		_w15227_,
		_w20498_
	);
	LUT3 #(
		.INIT('h70)
	) name16451 (
		_w19474_,
		_w19720_,
		_w20498_,
		_w20499_
	);
	LUT3 #(
		.INIT('h10)
	) name16452 (
		_w4104_,
		_w20497_,
		_w20499_,
		_w20500_
	);
	LUT3 #(
		.INIT('h15)
	) name16453 (
		_w20488_,
		_w20496_,
		_w20500_,
		_w20501_
	);
	LUT4 #(
		.INIT('h4440)
	) name16454 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		_w9418_,
		_w9414_,
		_w9415_,
		_w20502_
	);
	LUT3 #(
		.INIT('h10)
	) name16455 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		\bdma_BWCOUNT_reg[8]/NET0131 ,
		_w20502_,
		_w20503_
	);
	LUT4 #(
		.INIT('h0100)
	) name16456 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		\bdma_BWCOUNT_reg[8]/NET0131 ,
		\bdma_BWCOUNT_reg[9]/NET0131 ,
		_w20502_,
		_w20504_
	);
	LUT3 #(
		.INIT('h10)
	) name16457 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		\bdma_BWCOUNT_reg[11]/NET0131 ,
		_w20504_,
		_w20505_
	);
	LUT4 #(
		.INIT('h0100)
	) name16458 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		\bdma_BWCOUNT_reg[11]/NET0131 ,
		\bdma_BWCOUNT_reg[12]/NET0131 ,
		_w20504_,
		_w20506_
	);
	LUT2 #(
		.INIT('h4)
	) name16459 (
		_w5760_,
		_w9432_,
		_w20507_
	);
	LUT4 #(
		.INIT('h00de)
	) name16460 (
		\bdma_BWCOUNT_reg[13]/NET0131 ,
		_w9432_,
		_w20506_,
		_w20507_,
		_w20508_
	);
	LUT3 #(
		.INIT('h80)
	) name16461 (
		\bdma_BEAD_reg[2]/NET0131 ,
		\bdma_BEAD_reg[3]/NET0131 ,
		_w13031_,
		_w20509_
	);
	LUT4 #(
		.INIT('h8000)
	) name16462 (
		\bdma_BEAD_reg[2]/NET0131 ,
		\bdma_BEAD_reg[3]/NET0131 ,
		\bdma_BEAD_reg[4]/NET0131 ,
		_w13031_,
		_w20510_
	);
	LUT3 #(
		.INIT('h80)
	) name16463 (
		\bdma_BEAD_reg[5]/NET0131 ,
		\bdma_BEAD_reg[6]/NET0131 ,
		_w20510_,
		_w20511_
	);
	LUT4 #(
		.INIT('h8000)
	) name16464 (
		\bdma_BEAD_reg[5]/NET0131 ,
		\bdma_BEAD_reg[6]/NET0131 ,
		\bdma_BEAD_reg[7]/NET0131 ,
		_w20510_,
		_w20512_
	);
	LUT3 #(
		.INIT('h80)
	) name16465 (
		\bdma_BEAD_reg[8]/NET0131 ,
		\bdma_BEAD_reg[9]/NET0131 ,
		_w20512_,
		_w20513_
	);
	LUT4 #(
		.INIT('h8000)
	) name16466 (
		\bdma_BEAD_reg[10]/NET0131 ,
		\bdma_BEAD_reg[8]/NET0131 ,
		\bdma_BEAD_reg[9]/NET0131 ,
		_w20512_,
		_w20514_
	);
	LUT4 #(
		.INIT('h060c)
	) name16467 (
		\bdma_BEAD_reg[11]/NET0131 ,
		\bdma_BEAD_reg[12]/NET0131 ,
		_w13032_,
		_w20514_,
		_w20515_
	);
	LUT2 #(
		.INIT('h8)
	) name16468 (
		_w6758_,
		_w13032_,
		_w20516_
	);
	LUT2 #(
		.INIT('he)
	) name16469 (
		_w20515_,
		_w20516_,
		_w20517_
	);
	LUT3 #(
		.INIT('h13)
	) name16470 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001 ,
		_w9894_,
		_w20518_
	);
	LUT4 #(
		.INIT('h0002)
	) name16471 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w20518_,
		_w20519_
	);
	LUT4 #(
		.INIT('h5700)
	) name16472 (
		_w11625_,
		_w12315_,
		_w12316_,
		_w20519_,
		_w20520_
	);
	LUT4 #(
		.INIT('h313b)
	) name16473 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001 ,
		_w11631_,
		_w11635_,
		_w20521_
	);
	LUT4 #(
		.INIT('h0020)
	) name16474 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w9453_,
		_w9894_,
		_w12370_,
		_w20522_
	);
	LUT4 #(
		.INIT('hff45)
	) name16475 (
		_w11624_,
		_w20520_,
		_w20521_,
		_w20522_,
		_w20523_
	);
	LUT2 #(
		.INIT('h8)
	) name16476 (
		_w9946_,
		_w12370_,
		_w20524_
	);
	LUT2 #(
		.INIT('h2)
	) name16477 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001 ,
		_w11656_,
		_w20525_
	);
	LUT3 #(
		.INIT('h01)
	) name16478 (
		_w9946_,
		_w11659_,
		_w20525_,
		_w20526_
	);
	LUT4 #(
		.INIT('hfd00)
	) name16479 (
		_w11655_,
		_w12315_,
		_w12316_,
		_w20526_,
		_w20527_
	);
	LUT2 #(
		.INIT('h1)
	) name16480 (
		_w20524_,
		_w20527_,
		_w20528_
	);
	LUT4 #(
		.INIT('h20aa)
	) name16481 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9438_,
		_w20529_
	);
	LUT3 #(
		.INIT('h07)
	) name16482 (
		\core_c_dec_MTCNTR_Eg_reg/P0001 ,
		\core_c_psq_CNTRval_reg/NET0131 ,
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		_w20530_
	);
	LUT4 #(
		.INIT('h1300)
	) name16483 (
		_w5088_,
		_w17162_,
		_w17161_,
		_w20530_,
		_w20531_
	);
	LUT2 #(
		.INIT('h1)
	) name16484 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w20531_,
		_w20532_
	);
	LUT4 #(
		.INIT('h4500)
	) name16485 (
		_w4971_,
		_w17169_,
		_w17170_,
		_w20532_,
		_w20533_
	);
	LUT2 #(
		.INIT('he)
	) name16486 (
		_w9440_,
		_w20533_,
		_w20534_
	);
	LUT4 #(
		.INIT('h4500)
	) name16487 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9438_,
		_w20535_
	);
	LUT3 #(
		.INIT('h0e)
	) name16488 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w20536_
	);
	LUT3 #(
		.INIT('h71)
	) name16489 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w20537_
	);
	LUT2 #(
		.INIT('h4)
	) name16490 (
		_w20535_,
		_w20537_,
		_w20538_
	);
	LUT4 #(
		.INIT('hfecc)
	) name16491 (
		_w9440_,
		_w20529_,
		_w20533_,
		_w20538_,
		_w20539_
	);
	LUT3 #(
		.INIT('h56)
	) name16492 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		_w9440_,
		_w20533_,
		_w20540_
	);
	LUT4 #(
		.INIT('h0100)
	) name16493 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001 ,
		_w20541_
	);
	LUT4 #(
		.INIT('h2000)
	) name16494 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001 ,
		_w20542_
	);
	LUT4 #(
		.INIT('h1000)
	) name16495 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001 ,
		_w20543_
	);
	LUT4 #(
		.INIT('h0400)
	) name16496 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001 ,
		_w20544_
	);
	LUT4 #(
		.INIT('h0001)
	) name16497 (
		_w20541_,
		_w20542_,
		_w20543_,
		_w20544_,
		_w20545_
	);
	LUT4 #(
		.INIT('h4000)
	) name16498 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001 ,
		_w20546_
	);
	LUT4 #(
		.INIT('h0800)
	) name16499 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001 ,
		_w20547_
	);
	LUT4 #(
		.INIT('h0200)
	) name16500 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001 ,
		_w20548_
	);
	LUT4 #(
		.INIT('h0001)
	) name16501 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w20546_,
		_w20547_,
		_w20548_,
		_w20549_
	);
	LUT4 #(
		.INIT('h4070)
	) name16502 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w20550_
	);
	LUT2 #(
		.INIT('h1)
	) name16503 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w20550_,
		_w20551_
	);
	LUT3 #(
		.INIT('h70)
	) name16504 (
		_w20545_,
		_w20549_,
		_w20551_,
		_w20552_
	);
	LUT4 #(
		.INIT('h2022)
	) name16505 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w7927_,
		_w8040_,
		_w8042_,
		_w20553_
	);
	LUT4 #(
		.INIT('heee2)
	) name16506 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w14577_,
		_w20552_,
		_w20553_,
		_w20554_
	);
	LUT4 #(
		.INIT('h0400)
	) name16507 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001 ,
		_w20555_
	);
	LUT4 #(
		.INIT('h2000)
	) name16508 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001 ,
		_w20556_
	);
	LUT4 #(
		.INIT('h0200)
	) name16509 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001 ,
		_w20557_
	);
	LUT4 #(
		.INIT('h0800)
	) name16510 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001 ,
		_w20558_
	);
	LUT4 #(
		.INIT('h0001)
	) name16511 (
		_w20555_,
		_w20556_,
		_w20557_,
		_w20558_,
		_w20559_
	);
	LUT4 #(
		.INIT('h0100)
	) name16512 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001 ,
		_w20560_
	);
	LUT4 #(
		.INIT('h1000)
	) name16513 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001 ,
		_w20561_
	);
	LUT4 #(
		.INIT('h4000)
	) name16514 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001 ,
		_w20562_
	);
	LUT4 #(
		.INIT('h0001)
	) name16515 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w20560_,
		_w20561_,
		_w20562_,
		_w20563_
	);
	LUT4 #(
		.INIT('h4070)
	) name16516 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_IRE_reg[15]/NET0131 ,
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w20564_
	);
	LUT2 #(
		.INIT('h1)
	) name16517 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w20564_,
		_w20565_
	);
	LUT3 #(
		.INIT('h70)
	) name16518 (
		_w20559_,
		_w20563_,
		_w20565_,
		_w20566_
	);
	LUT4 #(
		.INIT('h2022)
	) name16519 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w7592_,
		_w7707_,
		_w7709_,
		_w20567_
	);
	LUT4 #(
		.INIT('heee2)
	) name16520 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w14577_,
		_w20566_,
		_w20567_,
		_w20568_
	);
	LUT4 #(
		.INIT('h4000)
	) name16521 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001 ,
		_w20569_
	);
	LUT4 #(
		.INIT('h0200)
	) name16522 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001 ,
		_w20570_
	);
	LUT4 #(
		.INIT('h2000)
	) name16523 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001 ,
		_w20571_
	);
	LUT4 #(
		.INIT('h0800)
	) name16524 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001 ,
		_w20572_
	);
	LUT4 #(
		.INIT('h0001)
	) name16525 (
		_w20569_,
		_w20570_,
		_w20571_,
		_w20572_,
		_w20573_
	);
	LUT4 #(
		.INIT('h0100)
	) name16526 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001 ,
		_w20574_
	);
	LUT4 #(
		.INIT('h1000)
	) name16527 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001 ,
		_w20575_
	);
	LUT4 #(
		.INIT('h0400)
	) name16528 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001 ,
		_w20576_
	);
	LUT4 #(
		.INIT('h0001)
	) name16529 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w20574_,
		_w20575_,
		_w20576_,
		_w20577_
	);
	LUT4 #(
		.INIT('h4070)
	) name16530 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w20578_
	);
	LUT2 #(
		.INIT('h1)
	) name16531 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w20578_,
		_w20579_
	);
	LUT3 #(
		.INIT('h70)
	) name16532 (
		_w20573_,
		_w20577_,
		_w20579_,
		_w20580_
	);
	LUT4 #(
		.INIT('h2022)
	) name16533 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w6054_,
		_w6173_,
		_w6175_,
		_w20581_
	);
	LUT4 #(
		.INIT('heee2)
	) name16534 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w14577_,
		_w20580_,
		_w20581_,
		_w20582_
	);
	LUT4 #(
		.INIT('h1000)
	) name16535 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001 ,
		_w20583_
	);
	LUT4 #(
		.INIT('h0200)
	) name16536 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001 ,
		_w20584_
	);
	LUT4 #(
		.INIT('h0800)
	) name16537 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001 ,
		_w20585_
	);
	LUT4 #(
		.INIT('h4000)
	) name16538 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001 ,
		_w20586_
	);
	LUT4 #(
		.INIT('h0001)
	) name16539 (
		_w20583_,
		_w20584_,
		_w20585_,
		_w20586_,
		_w20587_
	);
	LUT4 #(
		.INIT('h2000)
	) name16540 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001 ,
		_w20588_
	);
	LUT4 #(
		.INIT('h0400)
	) name16541 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001 ,
		_w20589_
	);
	LUT4 #(
		.INIT('h0100)
	) name16542 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001 ,
		_w20590_
	);
	LUT4 #(
		.INIT('h0001)
	) name16543 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w20588_,
		_w20589_,
		_w20590_,
		_w20591_
	);
	LUT4 #(
		.INIT('h4070)
	) name16544 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w20592_
	);
	LUT2 #(
		.INIT('h1)
	) name16545 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w20592_,
		_w20593_
	);
	LUT3 #(
		.INIT('h70)
	) name16546 (
		_w20587_,
		_w20591_,
		_w20593_,
		_w20594_
	);
	LUT4 #(
		.INIT('h2022)
	) name16547 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w6378_,
		_w6498_,
		_w6500_,
		_w20595_
	);
	LUT4 #(
		.INIT('heee2)
	) name16548 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w14577_,
		_w20594_,
		_w20595_,
		_w20596_
	);
	LUT4 #(
		.INIT('h0400)
	) name16549 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001 ,
		_w20597_
	);
	LUT4 #(
		.INIT('h2000)
	) name16550 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001 ,
		_w20598_
	);
	LUT4 #(
		.INIT('h0200)
	) name16551 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001 ,
		_w20599_
	);
	LUT4 #(
		.INIT('h0800)
	) name16552 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001 ,
		_w20600_
	);
	LUT4 #(
		.INIT('h0001)
	) name16553 (
		_w20597_,
		_w20598_,
		_w20599_,
		_w20600_,
		_w20601_
	);
	LUT4 #(
		.INIT('h0100)
	) name16554 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001 ,
		_w20602_
	);
	LUT4 #(
		.INIT('h1000)
	) name16555 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001 ,
		_w20603_
	);
	LUT4 #(
		.INIT('h4000)
	) name16556 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001 ,
		_w20604_
	);
	LUT4 #(
		.INIT('h0001)
	) name16557 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w20602_,
		_w20603_,
		_w20604_,
		_w20605_
	);
	LUT4 #(
		.INIT('h2070)
	) name16558 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w20606_
	);
	LUT2 #(
		.INIT('h1)
	) name16559 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w20606_,
		_w20607_
	);
	LUT3 #(
		.INIT('h70)
	) name16560 (
		_w20601_,
		_w20605_,
		_w20607_,
		_w20608_
	);
	LUT4 #(
		.INIT('h2022)
	) name16561 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w6774_,
		_w6894_,
		_w6896_,
		_w20609_
	);
	LUT4 #(
		.INIT('heee2)
	) name16562 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w14577_,
		_w20608_,
		_w20609_,
		_w20610_
	);
	LUT4 #(
		.INIT('h0800)
	) name16563 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001 ,
		_w20611_
	);
	LUT4 #(
		.INIT('h2000)
	) name16564 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001 ,
		_w20612_
	);
	LUT4 #(
		.INIT('h4000)
	) name16565 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001 ,
		_w20613_
	);
	LUT4 #(
		.INIT('h0100)
	) name16566 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001 ,
		_w20614_
	);
	LUT4 #(
		.INIT('h0001)
	) name16567 (
		_w20611_,
		_w20612_,
		_w20613_,
		_w20614_,
		_w20615_
	);
	LUT4 #(
		.INIT('h0400)
	) name16568 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001 ,
		_w20616_
	);
	LUT4 #(
		.INIT('h1000)
	) name16569 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001 ,
		_w20617_
	);
	LUT4 #(
		.INIT('h0200)
	) name16570 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001 ,
		_w20618_
	);
	LUT4 #(
		.INIT('h0001)
	) name16571 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w20616_,
		_w20617_,
		_w20618_,
		_w20619_
	);
	LUT2 #(
		.INIT('h8)
	) name16572 (
		_w20615_,
		_w20619_,
		_w20620_
	);
	LUT4 #(
		.INIT('h0057)
	) name16573 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w7140_,
		_w7240_,
		_w20620_,
		_w20621_
	);
	LUT4 #(
		.INIT('h0100)
	) name16574 (
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		_w20466_,
		_w20622_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name16575 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[7]/NET0131 ,
		\core_c_psq_Iact_E_reg[8]/NET0131 ,
		_w20622_,
		_w20623_
	);
	LUT3 #(
		.INIT('ha2)
	) name16576 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w19945_,
		_w20623_,
		_w20624_
	);
	LUT2 #(
		.INIT('h4)
	) name16577 (
		_w19947_,
		_w20624_,
		_w20625_
	);
	LUT3 #(
		.INIT('hf8)
	) name16578 (
		_w19947_,
		_w20621_,
		_w20625_,
		_w20626_
	);
	LUT4 #(
		.INIT('h8a88)
	) name16579 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w6774_,
		_w6894_,
		_w6896_,
		_w20627_
	);
	LUT4 #(
		.INIT('h2000)
	) name16580 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001 ,
		_w20628_
	);
	LUT4 #(
		.INIT('h0800)
	) name16581 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001 ,
		_w20629_
	);
	LUT4 #(
		.INIT('h0100)
	) name16582 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001 ,
		_w20630_
	);
	LUT4 #(
		.INIT('h1000)
	) name16583 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001 ,
		_w20631_
	);
	LUT4 #(
		.INIT('h0001)
	) name16584 (
		_w20628_,
		_w20629_,
		_w20630_,
		_w20631_,
		_w20632_
	);
	LUT4 #(
		.INIT('h0200)
	) name16585 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001 ,
		_w20633_
	);
	LUT4 #(
		.INIT('h0400)
	) name16586 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001 ,
		_w20634_
	);
	LUT4 #(
		.INIT('h4000)
	) name16587 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001 ,
		_w20635_
	);
	LUT4 #(
		.INIT('h0001)
	) name16588 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w20633_,
		_w20634_,
		_w20635_,
		_w20636_
	);
	LUT2 #(
		.INIT('h8)
	) name16589 (
		_w20632_,
		_w20636_,
		_w20637_
	);
	LUT2 #(
		.INIT('h8)
	) name16590 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		_w20638_
	);
	LUT4 #(
		.INIT('h0045)
	) name16591 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4094_,
		_w4097_,
		_w20638_,
		_w20639_
	);
	LUT2 #(
		.INIT('h2)
	) name16592 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w20639_,
		_w20640_
	);
	LUT2 #(
		.INIT('h4)
	) name16593 (
		_w19947_,
		_w20640_,
		_w20641_
	);
	LUT4 #(
		.INIT('hff02)
	) name16594 (
		_w19947_,
		_w20627_,
		_w20637_,
		_w20641_,
		_w20642_
	);
	LUT4 #(
		.INIT('hb888)
	) name16595 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w4104_,
		_w19057_,
		_w19472_,
		_w20643_
	);
	LUT4 #(
		.INIT('hb888)
	) name16596 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w4104_,
		_w19049_,
		_w19472_,
		_w20644_
	);
	LUT4 #(
		.INIT('hb888)
	) name16597 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w4104_,
		_w19049_,
		_w19478_,
		_w20645_
	);
	LUT4 #(
		.INIT('hb888)
	) name16598 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w4104_,
		_w19057_,
		_w19478_,
		_w20646_
	);
	LUT4 #(
		.INIT('h2000)
	) name16599 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20647_
	);
	LUT4 #(
		.INIT('h4000)
	) name16600 (
		_w4104_,
		_w19058_,
		_w19050_,
		_w19057_,
		_w20648_
	);
	LUT2 #(
		.INIT('he)
	) name16601 (
		_w20647_,
		_w20648_,
		_w20649_
	);
	LUT4 #(
		.INIT('hb888)
	) name16602 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w4104_,
		_w19057_,
		_w19054_,
		_w20650_
	);
	LUT4 #(
		.INIT('hb888)
	) name16603 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w4104_,
		_w19049_,
		_w19054_,
		_w20651_
	);
	LUT4 #(
		.INIT('hb888)
	) name16604 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w4104_,
		_w19056_,
		_w19065_,
		_w20652_
	);
	LUT4 #(
		.INIT('h2000)
	) name16605 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20653_
	);
	LUT4 #(
		.INIT('h4000)
	) name16606 (
		_w4104_,
		_w19050_,
		_w19057_,
		_w19477_,
		_w20654_
	);
	LUT2 #(
		.INIT('he)
	) name16607 (
		_w20653_,
		_w20654_,
		_w20655_
	);
	LUT4 #(
		.INIT('hb888)
	) name16608 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w4104_,
		_w19065_,
		_w19048_,
		_w20656_
	);
	LUT3 #(
		.INIT('h40)
	) name16609 (
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		_w12828_,
		_w20082_,
		_w20657_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name16610 (
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[7]/NET0131 ,
		_w12828_,
		_w20082_,
		_w20658_
	);
	LUT4 #(
		.INIT('haba8)
	) name16611 (
		\sport1_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w19498_,
		_w20078_,
		_w20658_,
		_w20659_
	);
	LUT4 #(
		.INIT('h0100)
	) name16612 (
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[5]/NET0131 ,
		_w20082_,
		_w20660_
	);
	LUT3 #(
		.INIT('h31)
	) name16613 (
		\sport1_rxctl_Wcnt_reg[6]/NET0131 ,
		_w20657_,
		_w20660_,
		_w20661_
	);
	LUT3 #(
		.INIT('h2e)
	) name16614 (
		\sport1_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w20079_,
		_w20661_,
		_w20662_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name16615 (
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[5]/NET0131 ,
		_w20082_,
		_w20663_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16616 (
		\sport1_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w19498_,
		_w20078_,
		_w20663_,
		_w20664_
	);
	LUT2 #(
		.INIT('h9)
	) name16617 (
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		_w20082_,
		_w20665_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16618 (
		\sport1_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w19498_,
		_w20078_,
		_w20665_,
		_w20666_
	);
	LUT4 #(
		.INIT('h5595)
	) name16619 (
		\sport1_rxctl_Wcnt_reg[2]/NET0131 ,
		_w20074_,
		_w20075_,
		_w20077_,
		_w20667_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16620 (
		\sport1_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w19498_,
		_w20078_,
		_w20667_,
		_w20668_
	);
	LUT4 #(
		.INIT('h3363)
	) name16621 (
		\sport1_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[1]/NET0131 ,
		_w20074_,
		_w20077_,
		_w20669_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16622 (
		\sport1_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w19498_,
		_w20078_,
		_w20669_,
		_w20670_
	);
	LUT3 #(
		.INIT('h59)
	) name16623 (
		\sport1_rxctl_Wcnt_reg[0]/NET0131 ,
		_w20074_,
		_w20077_,
		_w20671_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16624 (
		\sport1_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w19498_,
		_w20078_,
		_w20671_,
		_w20672_
	);
	LUT3 #(
		.INIT('h40)
	) name16625 (
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		_w12840_,
		_w20112_,
		_w20673_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name16626 (
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[7]/NET0131 ,
		_w12840_,
		_w20112_,
		_w20674_
	);
	LUT4 #(
		.INIT('haba8)
	) name16627 (
		\sport0_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w19620_,
		_w20108_,
		_w20674_,
		_w20675_
	);
	LUT4 #(
		.INIT('h0100)
	) name16628 (
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[5]/NET0131 ,
		_w20112_,
		_w20676_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name16629 (
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[5]/NET0131 ,
		_w20112_,
		_w20677_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16630 (
		\sport0_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w19620_,
		_w20108_,
		_w20677_,
		_w20678_
	);
	LUT2 #(
		.INIT('h9)
	) name16631 (
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		_w20112_,
		_w20679_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16632 (
		\sport0_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w19620_,
		_w20108_,
		_w20679_,
		_w20680_
	);
	LUT4 #(
		.INIT('h3363)
	) name16633 (
		\sport0_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[1]/NET0131 ,
		_w20104_,
		_w20107_,
		_w20681_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16634 (
		\sport0_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w19620_,
		_w20108_,
		_w20681_,
		_w20682_
	);
	LUT3 #(
		.INIT('h59)
	) name16635 (
		\sport0_rxctl_Wcnt_reg[0]/NET0131 ,
		_w20104_,
		_w20107_,
		_w20683_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16636 (
		\sport0_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w19620_,
		_w20108_,
		_w20683_,
		_w20684_
	);
	LUT3 #(
		.INIT('h6c)
	) name16637 (
		\clkc_oscntr_reg_DO_reg[10]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[11]/NET0131 ,
		_w14700_,
		_w20685_
	);
	LUT4 #(
		.INIT('h5595)
	) name16638 (
		\sport0_rxctl_Wcnt_reg[2]/NET0131 ,
		_w20104_,
		_w20105_,
		_w20107_,
		_w20686_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name16639 (
		\sport0_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w19620_,
		_w20108_,
		_w20686_,
		_w20687_
	);
	LUT3 #(
		.INIT('h31)
	) name16640 (
		\sport0_rxctl_Wcnt_reg[6]/NET0131 ,
		_w20673_,
		_w20676_,
		_w20688_
	);
	LUT3 #(
		.INIT('h2e)
	) name16641 (
		\sport0_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w20109_,
		_w20688_,
		_w20689_
	);
	LUT2 #(
		.INIT('h6)
	) name16642 (
		\sice_IIRC_reg[16]/NET0131 ,
		_w14201_,
		_w20690_
	);
	LUT4 #(
		.INIT('h2000)
	) name16643 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20691_
	);
	LUT4 #(
		.INIT('h4000)
	) name16644 (
		_w4104_,
		_w19050_,
		_w19049_,
		_w19477_,
		_w20692_
	);
	LUT2 #(
		.INIT('he)
	) name16645 (
		_w20691_,
		_w20692_,
		_w20693_
	);
	LUT4 #(
		.INIT('h0020)
	) name16646 (
		\core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20694_
	);
	LUT3 #(
		.INIT('h0b)
	) name16647 (
		_w12398_,
		_w13536_,
		_w20694_,
		_w20695_
	);
	LUT4 #(
		.INIT('h0200)
	) name16648 (
		\core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20696_
	);
	LUT4 #(
		.INIT('h0002)
	) name16649 (
		\core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20697_
	);
	LUT4 #(
		.INIT('h2000)
	) name16650 (
		\core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20698_
	);
	LUT3 #(
		.INIT('h01)
	) name16651 (
		_w20697_,
		_w20698_,
		_w20696_,
		_w20699_
	);
	LUT2 #(
		.INIT('h8)
	) name16652 (
		_w20695_,
		_w20699_,
		_w20700_
	);
	LUT4 #(
		.INIT('hfe00)
	) name16653 (
		_w7140_,
		_w7240_,
		_w20281_,
		_w20700_,
		_w20701_
	);
	LUT3 #(
		.INIT('h10)
	) name16654 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20702_
	);
	LUT2 #(
		.INIT('h1)
	) name16655 (
		_w20701_,
		_w20702_,
		_w20703_
	);
	LUT4 #(
		.INIT('h0020)
	) name16656 (
		\core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20704_
	);
	LUT3 #(
		.INIT('h0b)
	) name16657 (
		_w12398_,
		_w13536_,
		_w20704_,
		_w20705_
	);
	LUT4 #(
		.INIT('h0200)
	) name16658 (
		\core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20706_
	);
	LUT4 #(
		.INIT('h0002)
	) name16659 (
		\core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20707_
	);
	LUT4 #(
		.INIT('h2000)
	) name16660 (
		\core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20708_
	);
	LUT3 #(
		.INIT('h01)
	) name16661 (
		_w20707_,
		_w20708_,
		_w20706_,
		_w20709_
	);
	LUT2 #(
		.INIT('h8)
	) name16662 (
		_w20705_,
		_w20709_,
		_w20710_
	);
	LUT4 #(
		.INIT('hfe00)
	) name16663 (
		_w7465_,
		_w7565_,
		_w20281_,
		_w20710_,
		_w20711_
	);
	LUT3 #(
		.INIT('h10)
	) name16664 (
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20712_
	);
	LUT2 #(
		.INIT('h1)
	) name16665 (
		_w20711_,
		_w20712_,
		_w20713_
	);
	LUT4 #(
		.INIT('h0020)
	) name16666 (
		\core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20714_
	);
	LUT3 #(
		.INIT('h0b)
	) name16667 (
		_w12398_,
		_w13536_,
		_w20714_,
		_w20715_
	);
	LUT4 #(
		.INIT('h0200)
	) name16668 (
		\core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20716_
	);
	LUT4 #(
		.INIT('h0002)
	) name16669 (
		\core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20717_
	);
	LUT4 #(
		.INIT('h2000)
	) name16670 (
		\core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20718_
	);
	LUT3 #(
		.INIT('h01)
	) name16671 (
		_w20717_,
		_w20718_,
		_w20716_,
		_w20719_
	);
	LUT2 #(
		.INIT('h8)
	) name16672 (
		_w20715_,
		_w20719_,
		_w20720_
	);
	LUT3 #(
		.INIT('h10)
	) name16673 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20721_
	);
	LUT4 #(
		.INIT('h002f)
	) name16674 (
		_w6758_,
		_w20281_,
		_w20720_,
		_w20721_,
		_w20722_
	);
	LUT4 #(
		.INIT('h0020)
	) name16675 (
		\core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w20723_
	);
	LUT3 #(
		.INIT('h0b)
	) name16676 (
		_w12398_,
		_w13536_,
		_w20723_,
		_w20724_
	);
	LUT4 #(
		.INIT('h0200)
	) name16677 (
		\core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w20725_
	);
	LUT4 #(
		.INIT('h0002)
	) name16678 (
		\core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w20726_
	);
	LUT4 #(
		.INIT('h2000)
	) name16679 (
		\core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w20727_
	);
	LUT3 #(
		.INIT('h01)
	) name16680 (
		_w20726_,
		_w20727_,
		_w20725_,
		_w20728_
	);
	LUT2 #(
		.INIT('h8)
	) name16681 (
		_w20724_,
		_w20728_,
		_w20729_
	);
	LUT4 #(
		.INIT('hfe00)
	) name16682 (
		_w6263_,
		_w6362_,
		_w20281_,
		_w20729_,
		_w20730_
	);
	LUT3 #(
		.INIT('h10)
	) name16683 (
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20731_
	);
	LUT2 #(
		.INIT('h1)
	) name16684 (
		_w20730_,
		_w20731_,
		_w20732_
	);
	LUT4 #(
		.INIT('h00e0)
	) name16685 (
		_w5013_,
		_w5014_,
		_w20274_,
		_w20278_,
		_w20733_
	);
	LUT4 #(
		.INIT('h000e)
	) name16686 (
		_w4976_,
		_w4978_,
		_w20274_,
		_w20278_,
		_w20734_
	);
	LUT4 #(
		.INIT('he000)
	) name16687 (
		_w5004_,
		_w5006_,
		_w20274_,
		_w20278_,
		_w20735_
	);
	LUT4 #(
		.INIT('h0e00)
	) name16688 (
		_w5020_,
		_w5021_,
		_w20274_,
		_w20278_,
		_w20736_
	);
	LUT4 #(
		.INIT('h0001)
	) name16689 (
		_w20733_,
		_w20734_,
		_w20735_,
		_w20736_,
		_w20737_
	);
	LUT4 #(
		.INIT('h0010)
	) name16690 (
		_w5013_,
		_w5014_,
		_w20274_,
		_w20278_,
		_w20738_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16691 (
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20739_
	);
	LUT4 #(
		.INIT('h0001)
	) name16692 (
		_w4976_,
		_w4978_,
		_w20274_,
		_w20278_,
		_w20740_
	);
	LUT2 #(
		.INIT('h8)
	) name16693 (
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		_w20740_,
		_w20741_
	);
	LUT4 #(
		.INIT('h1000)
	) name16694 (
		_w5004_,
		_w5006_,
		_w20274_,
		_w20278_,
		_w20742_
	);
	LUT4 #(
		.INIT('h0100)
	) name16695 (
		_w5020_,
		_w5021_,
		_w20274_,
		_w20278_,
		_w20743_
	);
	LUT4 #(
		.INIT('h153f)
	) name16696 (
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20744_
	);
	LUT3 #(
		.INIT('h40)
	) name16697 (
		_w20741_,
		_w20739_,
		_w20744_,
		_w20745_
	);
	LUT3 #(
		.INIT('h10)
	) name16698 (
		\core_dag_ilm2reg_I_reg[9]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20746_
	);
	LUT4 #(
		.INIT('h002f)
	) name16699 (
		_w13022_,
		_w20737_,
		_w20745_,
		_w20746_,
		_w20747_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16700 (
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20748_
	);
	LUT2 #(
		.INIT('h8)
	) name16701 (
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		_w20740_,
		_w20749_
	);
	LUT4 #(
		.INIT('h153f)
	) name16702 (
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20750_
	);
	LUT3 #(
		.INIT('h40)
	) name16703 (
		_w20749_,
		_w20748_,
		_w20750_,
		_w20751_
	);
	LUT3 #(
		.INIT('h10)
	) name16704 (
		\core_dag_ilm2reg_I_reg[6]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20752_
	);
	LUT4 #(
		.INIT('h002f)
	) name16705 (
		_w12931_,
		_w20737_,
		_w20751_,
		_w20752_,
		_w20753_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16706 (
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20754_
	);
	LUT2 #(
		.INIT('h8)
	) name16707 (
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		_w20740_,
		_w20755_
	);
	LUT4 #(
		.INIT('h153f)
	) name16708 (
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20756_
	);
	LUT3 #(
		.INIT('h40)
	) name16709 (
		_w20755_,
		_w20754_,
		_w20756_,
		_w20757_
	);
	LUT3 #(
		.INIT('h10)
	) name16710 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20758_
	);
	LUT4 #(
		.INIT('h002f)
	) name16711 (
		_w12939_,
		_w20737_,
		_w20757_,
		_w20758_,
		_w20759_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16712 (
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20760_
	);
	LUT2 #(
		.INIT('h8)
	) name16713 (
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		_w20740_,
		_w20761_
	);
	LUT4 #(
		.INIT('h153f)
	) name16714 (
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20762_
	);
	LUT3 #(
		.INIT('h40)
	) name16715 (
		_w20761_,
		_w20760_,
		_w20762_,
		_w20763_
	);
	LUT3 #(
		.INIT('h10)
	) name16716 (
		\core_dag_ilm2reg_I_reg[4]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20764_
	);
	LUT4 #(
		.INIT('h002f)
	) name16717 (
		_w12947_,
		_w20737_,
		_w20763_,
		_w20764_,
		_w20765_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16718 (
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20766_
	);
	LUT2 #(
		.INIT('h8)
	) name16719 (
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		_w20740_,
		_w20767_
	);
	LUT4 #(
		.INIT('h153f)
	) name16720 (
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20768_
	);
	LUT3 #(
		.INIT('h40)
	) name16721 (
		_w20767_,
		_w20766_,
		_w20768_,
		_w20769_
	);
	LUT3 #(
		.INIT('h10)
	) name16722 (
		\core_dag_ilm2reg_I_reg[3]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20770_
	);
	LUT4 #(
		.INIT('h002f)
	) name16723 (
		_w9156_,
		_w20737_,
		_w20769_,
		_w20770_,
		_w20771_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16724 (
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20772_
	);
	LUT2 #(
		.INIT('h8)
	) name16725 (
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		_w20740_,
		_w20773_
	);
	LUT4 #(
		.INIT('h153f)
	) name16726 (
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20774_
	);
	LUT3 #(
		.INIT('h40)
	) name16727 (
		_w20773_,
		_w20772_,
		_w20774_,
		_w20775_
	);
	LUT3 #(
		.INIT('h10)
	) name16728 (
		\core_dag_ilm2reg_I_reg[2]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20776_
	);
	LUT4 #(
		.INIT('h001f)
	) name16729 (
		_w12961_,
		_w20737_,
		_w20775_,
		_w20776_,
		_w20777_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16730 (
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20778_
	);
	LUT2 #(
		.INIT('h8)
	) name16731 (
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		_w20740_,
		_w20779_
	);
	LUT4 #(
		.INIT('h153f)
	) name16732 (
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20780_
	);
	LUT3 #(
		.INIT('h40)
	) name16733 (
		_w20779_,
		_w20778_,
		_w20780_,
		_w20781_
	);
	LUT3 #(
		.INIT('h10)
	) name16734 (
		\core_dag_ilm2reg_I_reg[1]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20782_
	);
	LUT4 #(
		.INIT('h001f)
	) name16735 (
		_w12969_,
		_w20737_,
		_w20781_,
		_w20782_,
		_w20783_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16736 (
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20784_
	);
	LUT2 #(
		.INIT('h8)
	) name16737 (
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		_w20740_,
		_w20785_
	);
	LUT4 #(
		.INIT('h153f)
	) name16738 (
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20786_
	);
	LUT3 #(
		.INIT('h40)
	) name16739 (
		_w20785_,
		_w20784_,
		_w20786_,
		_w20787_
	);
	LUT4 #(
		.INIT('hf100)
	) name16740 (
		_w12976_,
		_w12977_,
		_w20737_,
		_w20787_,
		_w20788_
	);
	LUT3 #(
		.INIT('h10)
	) name16741 (
		\core_dag_ilm2reg_I_reg[13]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20789_
	);
	LUT2 #(
		.INIT('h1)
	) name16742 (
		_w20788_,
		_w20789_,
		_w20790_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16743 (
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20791_
	);
	LUT2 #(
		.INIT('h8)
	) name16744 (
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		_w20740_,
		_w20792_
	);
	LUT4 #(
		.INIT('h153f)
	) name16745 (
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20793_
	);
	LUT3 #(
		.INIT('h40)
	) name16746 (
		_w20792_,
		_w20791_,
		_w20793_,
		_w20794_
	);
	LUT3 #(
		.INIT('h10)
	) name16747 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20795_
	);
	LUT4 #(
		.INIT('h001f)
	) name16748 (
		_w12984_,
		_w20737_,
		_w20794_,
		_w20795_,
		_w20796_
	);
	LUT4 #(
		.INIT('h45cf)
	) name16749 (
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w20797_
	);
	LUT2 #(
		.INIT('h8)
	) name16750 (
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		_w20740_,
		_w20798_
	);
	LUT4 #(
		.INIT('h153f)
	) name16751 (
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w20742_,
		_w20743_,
		_w20799_
	);
	LUT3 #(
		.INIT('h40)
	) name16752 (
		_w20798_,
		_w20797_,
		_w20799_,
		_w20800_
	);
	LUT3 #(
		.INIT('h10)
	) name16753 (
		\core_dag_ilm2reg_I_reg[0]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20801_
	);
	LUT4 #(
		.INIT('h001f)
	) name16754 (
		_w13008_,
		_w20737_,
		_w20800_,
		_w20801_,
		_w20802_
	);
	LUT3 #(
		.INIT('h20)
	) name16755 (
		\core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20803_
	);
	LUT3 #(
		.INIT('h20)
	) name16756 (
		\core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20804_
	);
	LUT3 #(
		.INIT('h20)
	) name16757 (
		\core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20805_
	);
	LUT3 #(
		.INIT('h20)
	) name16758 (
		\core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20806_
	);
	LUT4 #(
		.INIT('h0001)
	) name16759 (
		_w20803_,
		_w20804_,
		_w20805_,
		_w20806_,
		_w20807_
	);
	LUT2 #(
		.INIT('h4)
	) name16760 (
		_w13546_,
		_w20807_,
		_w20808_
	);
	LUT4 #(
		.INIT('hfe00)
	) name16761 (
		_w7140_,
		_w7240_,
		_w20366_,
		_w20808_,
		_w20809_
	);
	LUT2 #(
		.INIT('h4)
	) name16762 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w13546_,
		_w20810_
	);
	LUT2 #(
		.INIT('h1)
	) name16763 (
		_w20809_,
		_w20810_,
		_w20811_
	);
	LUT3 #(
		.INIT('h20)
	) name16764 (
		\core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20812_
	);
	LUT3 #(
		.INIT('h20)
	) name16765 (
		\core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20813_
	);
	LUT3 #(
		.INIT('h20)
	) name16766 (
		\core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20814_
	);
	LUT3 #(
		.INIT('h20)
	) name16767 (
		\core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20815_
	);
	LUT4 #(
		.INIT('h0001)
	) name16768 (
		_w20812_,
		_w20813_,
		_w20814_,
		_w20815_,
		_w20816_
	);
	LUT2 #(
		.INIT('h4)
	) name16769 (
		_w13546_,
		_w20816_,
		_w20817_
	);
	LUT4 #(
		.INIT('hfe00)
	) name16770 (
		_w7465_,
		_w7565_,
		_w20366_,
		_w20817_,
		_w20818_
	);
	LUT2 #(
		.INIT('h4)
	) name16771 (
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		_w13546_,
		_w20819_
	);
	LUT2 #(
		.INIT('h1)
	) name16772 (
		_w20818_,
		_w20819_,
		_w20820_
	);
	LUT3 #(
		.INIT('h20)
	) name16773 (
		\core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20821_
	);
	LUT3 #(
		.INIT('h20)
	) name16774 (
		\core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20822_
	);
	LUT3 #(
		.INIT('h20)
	) name16775 (
		\core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20823_
	);
	LUT3 #(
		.INIT('h20)
	) name16776 (
		\core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20824_
	);
	LUT4 #(
		.INIT('h0001)
	) name16777 (
		_w20821_,
		_w20822_,
		_w20823_,
		_w20824_,
		_w20825_
	);
	LUT2 #(
		.INIT('h4)
	) name16778 (
		_w13546_,
		_w20825_,
		_w20826_
	);
	LUT2 #(
		.INIT('h4)
	) name16779 (
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w13546_,
		_w20827_
	);
	LUT4 #(
		.INIT('h002f)
	) name16780 (
		_w5760_,
		_w20366_,
		_w20826_,
		_w20827_,
		_w20828_
	);
	LUT3 #(
		.INIT('h20)
	) name16781 (
		\core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20829_
	);
	LUT3 #(
		.INIT('h20)
	) name16782 (
		\core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20830_
	);
	LUT3 #(
		.INIT('h20)
	) name16783 (
		\core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20831_
	);
	LUT3 #(
		.INIT('h20)
	) name16784 (
		\core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20832_
	);
	LUT4 #(
		.INIT('h0001)
	) name16785 (
		_w20829_,
		_w20830_,
		_w20831_,
		_w20832_,
		_w20833_
	);
	LUT2 #(
		.INIT('h4)
	) name16786 (
		_w13546_,
		_w20833_,
		_w20834_
	);
	LUT2 #(
		.INIT('h4)
	) name16787 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		_w13546_,
		_w20835_
	);
	LUT4 #(
		.INIT('h002f)
	) name16788 (
		_w6758_,
		_w20366_,
		_w20834_,
		_w20835_,
		_w20836_
	);
	LUT3 #(
		.INIT('h20)
	) name16789 (
		\core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20837_
	);
	LUT3 #(
		.INIT('h20)
	) name16790 (
		\core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20838_
	);
	LUT3 #(
		.INIT('h20)
	) name16791 (
		\core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20839_
	);
	LUT3 #(
		.INIT('h20)
	) name16792 (
		\core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20840_
	);
	LUT4 #(
		.INIT('h0001)
	) name16793 (
		_w20837_,
		_w20838_,
		_w20839_,
		_w20840_,
		_w20841_
	);
	LUT2 #(
		.INIT('h4)
	) name16794 (
		_w13546_,
		_w20841_,
		_w20842_
	);
	LUT4 #(
		.INIT('hfe00)
	) name16795 (
		_w6263_,
		_w6362_,
		_w20366_,
		_w20842_,
		_w20843_
	);
	LUT2 #(
		.INIT('h4)
	) name16796 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		_w13546_,
		_w20844_
	);
	LUT2 #(
		.INIT('h1)
	) name16797 (
		_w20843_,
		_w20844_,
		_w20845_
	);
	LUT3 #(
		.INIT('h20)
	) name16798 (
		\core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131 ,
		_w16072_,
		_w20364_,
		_w20846_
	);
	LUT3 #(
		.INIT('h20)
	) name16799 (
		\core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131 ,
		_w16071_,
		_w20363_,
		_w20847_
	);
	LUT3 #(
		.INIT('h20)
	) name16800 (
		\core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131 ,
		_w16074_,
		_w20360_,
		_w20848_
	);
	LUT3 #(
		.INIT('h20)
	) name16801 (
		\core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131 ,
		_w16073_,
		_w20361_,
		_w20849_
	);
	LUT4 #(
		.INIT('h0001)
	) name16802 (
		_w20846_,
		_w20847_,
		_w20848_,
		_w20849_,
		_w20850_
	);
	LUT2 #(
		.INIT('h4)
	) name16803 (
		_w13546_,
		_w20850_,
		_w20851_
	);
	LUT4 #(
		.INIT('hfe00)
	) name16804 (
		_w5937_,
		_w6038_,
		_w20366_,
		_w20851_,
		_w20852_
	);
	LUT2 #(
		.INIT('h4)
	) name16805 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		_w13546_,
		_w20853_
	);
	LUT2 #(
		.INIT('h1)
	) name16806 (
		_w20852_,
		_w20853_,
		_w20854_
	);
	LUT3 #(
		.INIT('he0)
	) name16807 (
		_w5079_,
		_w5082_,
		_w20364_,
		_w20855_
	);
	LUT3 #(
		.INIT('he0)
	) name16808 (
		_w5087_,
		_w5090_,
		_w20360_,
		_w20856_
	);
	LUT3 #(
		.INIT('he0)
	) name16809 (
		_w5061_,
		_w5065_,
		_w20361_,
		_w20857_
	);
	LUT3 #(
		.INIT('he0)
	) name16810 (
		_w5070_,
		_w5073_,
		_w20363_,
		_w20858_
	);
	LUT4 #(
		.INIT('h0001)
	) name16811 (
		_w20855_,
		_w20856_,
		_w20857_,
		_w20858_,
		_w20859_
	);
	LUT4 #(
		.INIT('h00b1)
	) name16812 (
		_w5107_,
		_w7400_,
		_w7566_,
		_w20859_,
		_w20860_
	);
	LUT4 #(
		.INIT('h0200)
	) name16813 (
		\core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w20861_
	);
	LUT2 #(
		.INIT('h1)
	) name16814 (
		_w13546_,
		_w20861_,
		_w20862_
	);
	LUT4 #(
		.INIT('h0200)
	) name16815 (
		\core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w20863_
	);
	LUT4 #(
		.INIT('h0200)
	) name16816 (
		\core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w20864_
	);
	LUT4 #(
		.INIT('h0200)
	) name16817 (
		\core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w20865_
	);
	LUT3 #(
		.INIT('h01)
	) name16818 (
		_w20864_,
		_w20865_,
		_w20863_,
		_w20866_
	);
	LUT2 #(
		.INIT('h8)
	) name16819 (
		_w20862_,
		_w20866_,
		_w20867_
	);
	LUT2 #(
		.INIT('h4)
	) name16820 (
		\core_dag_ilm1reg_I_reg[8]/NET0131 ,
		_w13546_,
		_w20868_
	);
	LUT3 #(
		.INIT('h0b)
	) name16821 (
		_w20860_,
		_w20867_,
		_w20868_,
		_w20869_
	);
	LUT4 #(
		.INIT('h00b1)
	) name16822 (
		_w5107_,
		_w7579_,
		_w7710_,
		_w20859_,
		_w20870_
	);
	LUT4 #(
		.INIT('h0200)
	) name16823 (
		\core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w20871_
	);
	LUT2 #(
		.INIT('h1)
	) name16824 (
		_w13546_,
		_w20871_,
		_w20872_
	);
	LUT4 #(
		.INIT('h0200)
	) name16825 (
		\core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w20873_
	);
	LUT4 #(
		.INIT('h0200)
	) name16826 (
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w20874_
	);
	LUT4 #(
		.INIT('h0200)
	) name16827 (
		\core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w20875_
	);
	LUT3 #(
		.INIT('h01)
	) name16828 (
		_w20874_,
		_w20875_,
		_w20873_,
		_w20876_
	);
	LUT2 #(
		.INIT('h8)
	) name16829 (
		_w20872_,
		_w20876_,
		_w20877_
	);
	LUT2 #(
		.INIT('h4)
	) name16830 (
		\core_dag_ilm1reg_I_reg[5]/NET0131 ,
		_w13546_,
		_w20878_
	);
	LUT3 #(
		.INIT('h0b)
	) name16831 (
		_w20870_,
		_w20877_,
		_w20878_,
		_w20879_
	);
	LUT4 #(
		.INIT('h00b1)
	) name16832 (
		_w5107_,
		_w6591_,
		_w6897_,
		_w20859_,
		_w20880_
	);
	LUT4 #(
		.INIT('h0200)
	) name16833 (
		\core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w20881_
	);
	LUT2 #(
		.INIT('h1)
	) name16834 (
		_w13546_,
		_w20881_,
		_w20882_
	);
	LUT4 #(
		.INIT('h0200)
	) name16835 (
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w20883_
	);
	LUT4 #(
		.INIT('h0200)
	) name16836 (
		\core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w20884_
	);
	LUT4 #(
		.INIT('h0200)
	) name16837 (
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w20885_
	);
	LUT3 #(
		.INIT('h01)
	) name16838 (
		_w20884_,
		_w20885_,
		_w20883_,
		_w20886_
	);
	LUT2 #(
		.INIT('h8)
	) name16839 (
		_w20882_,
		_w20886_,
		_w20887_
	);
	LUT2 #(
		.INIT('h4)
	) name16840 (
		\core_dag_ilm1reg_I_reg[1]/NET0131 ,
		_w13546_,
		_w20888_
	);
	LUT3 #(
		.INIT('h0b)
	) name16841 (
		_w20880_,
		_w20887_,
		_w20888_,
		_w20889_
	);
	LUT4 #(
		.INIT('h0200)
	) name16842 (
		\core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w20890_
	);
	LUT2 #(
		.INIT('h1)
	) name16843 (
		_w13546_,
		_w20890_,
		_w20891_
	);
	LUT4 #(
		.INIT('h0200)
	) name16844 (
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w20892_
	);
	LUT4 #(
		.INIT('h0200)
	) name16845 (
		\core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w20893_
	);
	LUT4 #(
		.INIT('h0200)
	) name16846 (
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w20894_
	);
	LUT3 #(
		.INIT('h01)
	) name16847 (
		_w20893_,
		_w20894_,
		_w20892_,
		_w20895_
	);
	LUT2 #(
		.INIT('h8)
	) name16848 (
		_w20891_,
		_w20895_,
		_w20896_
	);
	LUT2 #(
		.INIT('h4)
	) name16849 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		_w13546_,
		_w20897_
	);
	LUT4 #(
		.INIT('h002f)
	) name16850 (
		_w15042_,
		_w20859_,
		_w20896_,
		_w20897_,
		_w20898_
	);
	LUT4 #(
		.INIT('h0200)
	) name16851 (
		\core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w20899_
	);
	LUT2 #(
		.INIT('h1)
	) name16852 (
		_w13546_,
		_w20899_,
		_w20900_
	);
	LUT4 #(
		.INIT('h0200)
	) name16853 (
		\core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w20901_
	);
	LUT4 #(
		.INIT('h0200)
	) name16854 (
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w20902_
	);
	LUT4 #(
		.INIT('h0200)
	) name16855 (
		\core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w20903_
	);
	LUT3 #(
		.INIT('h01)
	) name16856 (
		_w20902_,
		_w20903_,
		_w20901_,
		_w20904_
	);
	LUT2 #(
		.INIT('h8)
	) name16857 (
		_w20900_,
		_w20904_,
		_w20905_
	);
	LUT2 #(
		.INIT('h4)
	) name16858 (
		\core_dag_ilm1reg_I_reg[12]/NET0131 ,
		_w13546_,
		_w20906_
	);
	LUT4 #(
		.INIT('h001f)
	) name16859 (
		_w15045_,
		_w20859_,
		_w20905_,
		_w20906_,
		_w20907_
	);
	LUT4 #(
		.INIT('h0200)
	) name16860 (
		\core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w20908_
	);
	LUT2 #(
		.INIT('h1)
	) name16861 (
		_w13546_,
		_w20908_,
		_w20909_
	);
	LUT4 #(
		.INIT('h0200)
	) name16862 (
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w20910_
	);
	LUT4 #(
		.INIT('h0200)
	) name16863 (
		\core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w20911_
	);
	LUT4 #(
		.INIT('h0200)
	) name16864 (
		\core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w20912_
	);
	LUT3 #(
		.INIT('h01)
	) name16865 (
		_w20911_,
		_w20912_,
		_w20910_,
		_w20913_
	);
	LUT2 #(
		.INIT('h8)
	) name16866 (
		_w20909_,
		_w20913_,
		_w20914_
	);
	LUT2 #(
		.INIT('h4)
	) name16867 (
		\core_dag_ilm1reg_I_reg[11]/NET0131 ,
		_w13546_,
		_w20915_
	);
	LUT4 #(
		.INIT('h001f)
	) name16868 (
		_w15048_,
		_w20859_,
		_w20914_,
		_w20915_,
		_w20916_
	);
	LUT4 #(
		.INIT('h0200)
	) name16869 (
		\core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w20917_
	);
	LUT2 #(
		.INIT('h1)
	) name16870 (
		_w13546_,
		_w20917_,
		_w20918_
	);
	LUT4 #(
		.INIT('h0200)
	) name16871 (
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w20919_
	);
	LUT4 #(
		.INIT('h0200)
	) name16872 (
		\core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w20920_
	);
	LUT4 #(
		.INIT('h0200)
	) name16873 (
		\core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w20921_
	);
	LUT3 #(
		.INIT('h01)
	) name16874 (
		_w20920_,
		_w20921_,
		_w20919_,
		_w20922_
	);
	LUT2 #(
		.INIT('h8)
	) name16875 (
		_w20918_,
		_w20922_,
		_w20923_
	);
	LUT2 #(
		.INIT('h4)
	) name16876 (
		\core_dag_ilm1reg_I_reg[10]/NET0131 ,
		_w13546_,
		_w20924_
	);
	LUT4 #(
		.INIT('h002f)
	) name16877 (
		_w14869_,
		_w20859_,
		_w20923_,
		_w20924_,
		_w20925_
	);
	LUT2 #(
		.INIT('h6)
	) name16878 (
		\sice_ICYC_reg[16]/NET0131 ,
		_w13017_,
		_w20926_
	);
	LUT4 #(
		.INIT('h028a)
	) name16879 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		\core_c_dec_accPM_E_reg/P0001 ,
		_w6758_,
		_w8717_,
		_w20927_
	);
	LUT4 #(
		.INIT('h4000)
	) name16880 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w12695_,
		_w18495_,
		_w18481_,
		_w20928_
	);
	LUT4 #(
		.INIT('h222e)
	) name16881 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001 ,
		_w11830_,
		_w20927_,
		_w20928_,
		_w20929_
	);
	LUT4 #(
		.INIT('h222e)
	) name16882 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001 ,
		_w11329_,
		_w20927_,
		_w20928_,
		_w20930_
	);
	LUT3 #(
		.INIT('h13)
	) name16883 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001 ,
		_w9894_,
		_w20931_
	);
	LUT4 #(
		.INIT('h0002)
	) name16884 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w20931_,
		_w20932_
	);
	LUT4 #(
		.INIT('h313b)
	) name16885 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001 ,
		_w11631_,
		_w11635_,
		_w20933_
	);
	LUT4 #(
		.INIT('h2f00)
	) name16886 (
		_w11625_,
		_w12486_,
		_w20932_,
		_w20933_,
		_w20934_
	);
	LUT2 #(
		.INIT('h1)
	) name16887 (
		_w11624_,
		_w20934_,
		_w20935_
	);
	LUT4 #(
		.INIT('h80c4)
	) name16888 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w12343_,
		_w12345_,
		_w20936_
	);
	LUT2 #(
		.INIT('he)
	) name16889 (
		_w20935_,
		_w20936_,
		_w20937_
	);
	LUT3 #(
		.INIT('hca)
	) name16890 (
		\sport1_txctl_TXSHT_reg[10]/P0001 ,
		\sport1_txctl_TX_reg[11]/P0001 ,
		_w14269_,
		_w20938_
	);
	LUT4 #(
		.INIT('h4c08)
	) name16891 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w12343_,
		_w12345_,
		_w20939_
	);
	LUT2 #(
		.INIT('h2)
	) name16892 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001 ,
		_w11656_,
		_w20940_
	);
	LUT3 #(
		.INIT('h01)
	) name16893 (
		_w9946_,
		_w11659_,
		_w20940_,
		_w20941_
	);
	LUT3 #(
		.INIT('h70)
	) name16894 (
		_w11655_,
		_w12486_,
		_w20941_,
		_w20942_
	);
	LUT2 #(
		.INIT('h1)
	) name16895 (
		_w20939_,
		_w20942_,
		_w20943_
	);
	LUT3 #(
		.INIT('ha8)
	) name16896 (
		\sport1_rxctl_RCS_reg[1]/NET0131 ,
		_w19498_,
		_w19501_,
		_w20944_
	);
	LUT3 #(
		.INIT('ha8)
	) name16897 (
		\sport0_rxctl_RCS_reg[1]/NET0131 ,
		_w19620_,
		_w19623_,
		_w20945_
	);
	LUT3 #(
		.INIT('hca)
	) name16898 (
		\sport0_txctl_TXSHT_reg[10]/P0001 ,
		\sport0_txctl_TX_reg[11]/P0001 ,
		_w12552_,
		_w20946_
	);
	LUT4 #(
		.INIT('h78f0)
	) name16899 (
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		_w12301_,
		_w20947_
	);
	LUT3 #(
		.INIT('h20)
	) name16900 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w20947_,
		_w20948_
	);
	LUT2 #(
		.INIT('h6)
	) name16901 (
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		_w12301_,
		_w20949_
	);
	LUT3 #(
		.INIT('h20)
	) name16902 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w20949_,
		_w20950_
	);
	LUT4 #(
		.INIT('h1000)
	) name16903 (
		\core_c_dec_MFDAG2_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20951_
	);
	LUT3 #(
		.INIT('h01)
	) name16904 (
		_w19040_,
		_w19231_,
		_w19232_,
		_w20952_
	);
	LUT4 #(
		.INIT('h0002)
	) name16905 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w19040_,
		_w19231_,
		_w19232_,
		_w20953_
	);
	LUT2 #(
		.INIT('h4)
	) name16906 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w20953_,
		_w20954_
	);
	LUT2 #(
		.INIT('h4)
	) name16907 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w20955_
	);
	LUT4 #(
		.INIT('h0100)
	) name16908 (
		_w19040_,
		_w19231_,
		_w19232_,
		_w20955_,
		_w20956_
	);
	LUT4 #(
		.INIT('h6000)
	) name16909 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w19240_,
		_w20952_,
		_w20957_
	);
	LUT3 #(
		.INIT('ha8)
	) name16910 (
		_w5096_,
		_w19236_,
		_w19237_,
		_w20958_
	);
	LUT2 #(
		.INIT('h8)
	) name16911 (
		_w20953_,
		_w20958_,
		_w20959_
	);
	LUT4 #(
		.INIT('h0100)
	) name16912 (
		_w19040_,
		_w19231_,
		_w19232_,
		_w19234_,
		_w20960_
	);
	LUT2 #(
		.INIT('h8)
	) name16913 (
		_w19239_,
		_w20960_,
		_w20961_
	);
	LUT2 #(
		.INIT('h8)
	) name16914 (
		_w19720_,
		_w20960_,
		_w20962_
	);
	LUT3 #(
		.INIT('h1f)
	) name16915 (
		_w19239_,
		_w19720_,
		_w20960_,
		_w20963_
	);
	LUT3 #(
		.INIT('h10)
	) name16916 (
		_w20957_,
		_w20959_,
		_w20963_,
		_w20964_
	);
	LUT3 #(
		.INIT('h40)
	) name16917 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w19720_,
		_w20953_,
		_w20965_
	);
	LUT4 #(
		.INIT('h0400)
	) name16918 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w20966_
	);
	LUT3 #(
		.INIT('he0)
	) name16919 (
		_w19236_,
		_w19237_,
		_w20966_,
		_w20967_
	);
	LUT4 #(
		.INIT('hf040)
	) name16920 (
		_w19473_,
		_w19688_,
		_w20952_,
		_w20967_,
		_w20968_
	);
	LUT3 #(
		.INIT('h01)
	) name16921 (
		_w4104_,
		_w20965_,
		_w20968_,
		_w20969_
	);
	LUT3 #(
		.INIT('h15)
	) name16922 (
		_w20951_,
		_w20964_,
		_w20969_,
		_w20970_
	);
	LUT4 #(
		.INIT('h78f0)
	) name16923 (
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		_w12721_,
		_w20971_
	);
	LUT3 #(
		.INIT('h20)
	) name16924 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w20971_,
		_w20972_
	);
	LUT2 #(
		.INIT('h6)
	) name16925 (
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		_w12721_,
		_w20973_
	);
	LUT3 #(
		.INIT('h20)
	) name16926 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w20973_,
		_w20974_
	);
	LUT4 #(
		.INIT('h20aa)
	) name16927 (
		\core_c_psq_SSTAT_reg[2]/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w9438_,
		_w20975_
	);
	LUT4 #(
		.INIT('h00ba)
	) name16928 (
		_w4971_,
		_w17169_,
		_w17170_,
		_w20975_,
		_w20976_
	);
	LUT4 #(
		.INIT('h4500)
	) name16929 (
		_w4971_,
		_w17169_,
		_w17170_,
		_w20536_,
		_w20977_
	);
	LUT2 #(
		.INIT('h1)
	) name16930 (
		_w20976_,
		_w20977_,
		_w20978_
	);
	LUT3 #(
		.INIT('ha8)
	) name16931 (
		\bdma_BCTL_reg[0]/NET0131 ,
		\bdma_BCTL_reg[1]/NET0131 ,
		\bdma_DM_2nd_reg/NET0131 ,
		_w20979_
	);
	LUT4 #(
		.INIT('h00bf)
	) name16932 (
		_w4885_,
		_w4884_,
		_w4886_,
		_w20979_,
		_w20980_
	);
	LUT3 #(
		.INIT('h08)
	) name16933 (
		_w4761_,
		_w12533_,
		_w20980_,
		_w20981_
	);
	LUT2 #(
		.INIT('h4)
	) name16934 (
		\bdma_BCTL_reg[0]/NET0131 ,
		\bdma_BCTL_reg[1]/NET0131 ,
		_w20982_
	);
	LUT4 #(
		.INIT('h00f7)
	) name16935 (
		_w4761_,
		_w12533_,
		_w20980_,
		_w20982_,
		_w20983_
	);
	LUT3 #(
		.INIT('h46)
	) name16936 (
		\bdma_BCTL_reg[0]/NET0131 ,
		\bdma_BCTL_reg[1]/NET0131 ,
		\bdma_DM_2nd_reg/NET0131 ,
		_w20984_
	);
	LUT3 #(
		.INIT('h07)
	) name16937 (
		_w4884_,
		_w9075_,
		_w20984_,
		_w20985_
	);
	LUT3 #(
		.INIT('h08)
	) name16938 (
		_w4761_,
		_w12533_,
		_w20985_,
		_w20986_
	);
	LUT4 #(
		.INIT('h7f5f)
	) name16939 (
		_w4761_,
		_w9080_,
		_w12533_,
		_w20985_,
		_w20987_
	);
	LUT4 #(
		.INIT('h0080)
	) name16940 (
		\T_ED[0]_pad ,
		_w4761_,
		_w12533_,
		_w20980_,
		_w20988_
	);
	LUT4 #(
		.INIT('hfa8a)
	) name16941 (
		\bdma_BRdataBUF_reg[0]/P0001 ,
		_w20983_,
		_w20987_,
		_w20988_,
		_w20989_
	);
	LUT4 #(
		.INIT('h0603)
	) name16942 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		\bdma_BWCOUNT_reg[11]/NET0131 ,
		_w9432_,
		_w20504_,
		_w20990_
	);
	LUT3 #(
		.INIT('he0)
	) name16943 (
		_w6263_,
		_w6362_,
		_w9432_,
		_w20991_
	);
	LUT2 #(
		.INIT('h1)
	) name16944 (
		_w20990_,
		_w20991_,
		_w20992_
	);
	LUT3 #(
		.INIT('ha8)
	) name16945 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w9414_,
		_w9415_,
		_w20993_
	);
	LUT4 #(
		.INIT('h8880)
	) name16946 (
		\bdma_BIAD_reg[0]/NET0131 ,
		\bdma_BIAD_reg[1]/NET0131 ,
		_w9414_,
		_w9415_,
		_w20994_
	);
	LUT3 #(
		.INIT('h80)
	) name16947 (
		\bdma_BIAD_reg[2]/NET0131 ,
		\bdma_BIAD_reg[3]/NET0131 ,
		_w20994_,
		_w20995_
	);
	LUT4 #(
		.INIT('h8000)
	) name16948 (
		\bdma_BIAD_reg[2]/NET0131 ,
		\bdma_BIAD_reg[3]/NET0131 ,
		\bdma_BIAD_reg[4]/NET0131 ,
		_w20994_,
		_w20996_
	);
	LUT3 #(
		.INIT('h80)
	) name16949 (
		\bdma_BIAD_reg[5]/NET0131 ,
		\bdma_BIAD_reg[6]/NET0131 ,
		_w20996_,
		_w20997_
	);
	LUT4 #(
		.INIT('h8000)
	) name16950 (
		\bdma_BIAD_reg[5]/NET0131 ,
		\bdma_BIAD_reg[6]/NET0131 ,
		\bdma_BIAD_reg[7]/NET0131 ,
		_w20996_,
		_w20998_
	);
	LUT3 #(
		.INIT('h80)
	) name16951 (
		\bdma_BIAD_reg[8]/NET0131 ,
		\bdma_BIAD_reg[9]/NET0131 ,
		_w20998_,
		_w20999_
	);
	LUT4 #(
		.INIT('h8000)
	) name16952 (
		\bdma_BIAD_reg[10]/NET0131 ,
		\bdma_BIAD_reg[8]/NET0131 ,
		\bdma_BIAD_reg[9]/NET0131 ,
		_w20998_,
		_w21000_
	);
	LUT4 #(
		.INIT('h8000)
	) name16953 (
		_w5647_,
		_w5658_,
		_w9431_,
		_w12621_,
		_w21001_
	);
	LUT4 #(
		.INIT('h060c)
	) name16954 (
		\bdma_BIAD_reg[11]/NET0131 ,
		\bdma_BIAD_reg[12]/NET0131 ,
		_w21001_,
		_w21000_,
		_w21002_
	);
	LUT2 #(
		.INIT('h8)
	) name16955 (
		_w6758_,
		_w21001_,
		_w21003_
	);
	LUT2 #(
		.INIT('he)
	) name16956 (
		_w21002_,
		_w21003_,
		_w21004_
	);
	LUT3 #(
		.INIT('h10)
	) name16957 (
		_w6263_,
		_w6362_,
		_w21001_,
		_w21005_
	);
	LUT4 #(
		.INIT('hff12)
	) name16958 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w21001_,
		_w21000_,
		_w21005_,
		_w21006_
	);
	LUT4 #(
		.INIT('h870f)
	) name16959 (
		\bdma_BEAD_reg[11]/NET0131 ,
		\bdma_BEAD_reg[12]/NET0131 ,
		\bdma_BEAD_reg[13]/NET0131 ,
		_w20514_,
		_w21007_
	);
	LUT2 #(
		.INIT('h8)
	) name16960 (
		_w5760_,
		_w13032_,
		_w21008_
	);
	LUT3 #(
		.INIT('hf1)
	) name16961 (
		_w13032_,
		_w21007_,
		_w21008_,
		_w21009_
	);
	LUT3 #(
		.INIT('h10)
	) name16962 (
		_w6263_,
		_w6362_,
		_w13032_,
		_w21010_
	);
	LUT4 #(
		.INIT('hff12)
	) name16963 (
		\bdma_BEAD_reg[11]/NET0131 ,
		_w13032_,
		_w20514_,
		_w21010_,
		_w21011_
	);
	LUT4 #(
		.INIT('h4000)
	) name16964 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001 ,
		_w21012_
	);
	LUT4 #(
		.INIT('h0400)
	) name16965 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001 ,
		_w21013_
	);
	LUT4 #(
		.INIT('h0100)
	) name16966 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001 ,
		_w21014_
	);
	LUT4 #(
		.INIT('h0200)
	) name16967 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001 ,
		_w21015_
	);
	LUT4 #(
		.INIT('h0001)
	) name16968 (
		_w21012_,
		_w21013_,
		_w21014_,
		_w21015_,
		_w21016_
	);
	LUT4 #(
		.INIT('h0800)
	) name16969 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001 ,
		_w21017_
	);
	LUT4 #(
		.INIT('h2000)
	) name16970 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001 ,
		_w21018_
	);
	LUT4 #(
		.INIT('h1000)
	) name16971 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001 ,
		_w21019_
	);
	LUT4 #(
		.INIT('h0001)
	) name16972 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w21017_,
		_w21018_,
		_w21019_,
		_w21020_
	);
	LUT2 #(
		.INIT('h8)
	) name16973 (
		_w21016_,
		_w21020_,
		_w21021_
	);
	LUT4 #(
		.INIT('h0057)
	) name16974 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w7465_,
		_w7565_,
		_w21021_,
		_w21022_
	);
	LUT3 #(
		.INIT('h8a)
	) name16975 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[7]/NET0131 ,
		_w20622_,
		_w21023_
	);
	LUT3 #(
		.INIT('ha2)
	) name16976 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w19945_,
		_w21023_,
		_w21024_
	);
	LUT2 #(
		.INIT('h4)
	) name16977 (
		_w19947_,
		_w21024_,
		_w21025_
	);
	LUT3 #(
		.INIT('hf8)
	) name16978 (
		_w19947_,
		_w21022_,
		_w21025_,
		_w21026_
	);
	LUT3 #(
		.INIT('h8a)
	) name16979 (
		\bdma_BRdataBUF_reg[5]/P0001 ,
		_w20983_,
		_w20987_,
		_w21027_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name16980 (
		\T_ED[5]_pad ,
		_w4761_,
		_w9080_,
		_w12533_,
		_w21028_
	);
	LUT2 #(
		.INIT('h8)
	) name16981 (
		_w20981_,
		_w21028_,
		_w21029_
	);
	LUT2 #(
		.INIT('he)
	) name16982 (
		_w21027_,
		_w21029_,
		_w21030_
	);
	LUT3 #(
		.INIT('h8a)
	) name16983 (
		\bdma_BRdataBUF_reg[7]/P0001 ,
		_w20983_,
		_w20987_,
		_w21031_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name16984 (
		\T_ED[7]_pad ,
		_w4761_,
		_w9080_,
		_w12533_,
		_w21032_
	);
	LUT2 #(
		.INIT('h8)
	) name16985 (
		_w20981_,
		_w21032_,
		_w21033_
	);
	LUT2 #(
		.INIT('he)
	) name16986 (
		_w21031_,
		_w21033_,
		_w21034_
	);
	LUT3 #(
		.INIT('h8a)
	) name16987 (
		\bdma_BRdataBUF_reg[4]/P0001 ,
		_w20983_,
		_w20987_,
		_w21035_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name16988 (
		\T_ED[4]_pad ,
		_w4761_,
		_w9080_,
		_w12533_,
		_w21036_
	);
	LUT2 #(
		.INIT('h8)
	) name16989 (
		_w20981_,
		_w21036_,
		_w21037_
	);
	LUT2 #(
		.INIT('he)
	) name16990 (
		_w21035_,
		_w21037_,
		_w21038_
	);
	LUT3 #(
		.INIT('h8a)
	) name16991 (
		\bdma_BRdataBUF_reg[6]/P0001 ,
		_w20983_,
		_w20987_,
		_w21039_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name16992 (
		\T_ED[6]_pad ,
		_w4761_,
		_w9080_,
		_w12533_,
		_w21040_
	);
	LUT2 #(
		.INIT('h8)
	) name16993 (
		_w20981_,
		_w21040_,
		_w21041_
	);
	LUT2 #(
		.INIT('he)
	) name16994 (
		_w21039_,
		_w21041_,
		_w21042_
	);
	LUT3 #(
		.INIT('h8a)
	) name16995 (
		\bdma_BRdataBUF_reg[3]/P0001 ,
		_w20983_,
		_w20987_,
		_w21043_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name16996 (
		\T_ED[3]_pad ,
		_w4761_,
		_w9080_,
		_w12533_,
		_w21044_
	);
	LUT2 #(
		.INIT('h8)
	) name16997 (
		_w20981_,
		_w21044_,
		_w21045_
	);
	LUT2 #(
		.INIT('he)
	) name16998 (
		_w21043_,
		_w21045_,
		_w21046_
	);
	LUT3 #(
		.INIT('h8a)
	) name16999 (
		\bdma_BRdataBUF_reg[2]/P0001 ,
		_w20983_,
		_w20987_,
		_w21047_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name17000 (
		\T_ED[2]_pad ,
		_w4761_,
		_w9080_,
		_w12533_,
		_w21048_
	);
	LUT2 #(
		.INIT('h8)
	) name17001 (
		_w20981_,
		_w21048_,
		_w21049_
	);
	LUT2 #(
		.INIT('he)
	) name17002 (
		_w21047_,
		_w21049_,
		_w21050_
	);
	LUT3 #(
		.INIT('h8a)
	) name17003 (
		\bdma_BRdataBUF_reg[1]/P0001 ,
		_w20983_,
		_w20987_,
		_w21051_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name17004 (
		\T_ED[1]_pad ,
		_w4761_,
		_w9080_,
		_w12533_,
		_w21052_
	);
	LUT2 #(
		.INIT('h8)
	) name17005 (
		_w20981_,
		_w21052_,
		_w21053_
	);
	LUT2 #(
		.INIT('he)
	) name17006 (
		_w21051_,
		_w21053_,
		_w21054_
	);
	LUT3 #(
		.INIT('h6c)
	) name17007 (
		\sice_ICYC_reg[19]/NET0131 ,
		\sice_ICYC_reg[20]/NET0131 ,
		_w13018_,
		_w21055_
	);
	LUT4 #(
		.INIT('h8000)
	) name17008 (
		\sice_IIRC_reg[19]/NET0131 ,
		\sice_IIRC_reg[20]/NET0131 ,
		\sice_IIRC_reg[21]/NET0131 ,
		_w19741_,
		_w21056_
	);
	LUT3 #(
		.INIT('h6c)
	) name17009 (
		\sice_IIRC_reg[22]/NET0131 ,
		\sice_IIRC_reg[23]/NET0131 ,
		_w21056_,
		_w21057_
	);
	LUT2 #(
		.INIT('h6)
	) name17010 (
		\clkc_oscntr_reg_DO_reg[10]/NET0131 ,
		_w14700_,
		_w21058_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17011 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w7793_,
		_w7903_,
		_w7905_,
		_w21059_
	);
	LUT4 #(
		.INIT('h0400)
	) name17012 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001 ,
		_w21060_
	);
	LUT4 #(
		.INIT('h4000)
	) name17013 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001 ,
		_w21061_
	);
	LUT4 #(
		.INIT('h0200)
	) name17014 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001 ,
		_w21062_
	);
	LUT4 #(
		.INIT('h2000)
	) name17015 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001 ,
		_w21063_
	);
	LUT4 #(
		.INIT('h0001)
	) name17016 (
		_w21060_,
		_w21061_,
		_w21062_,
		_w21063_,
		_w21064_
	);
	LUT4 #(
		.INIT('h1000)
	) name17017 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001 ,
		_w21065_
	);
	LUT4 #(
		.INIT('h0800)
	) name17018 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001 ,
		_w21066_
	);
	LUT4 #(
		.INIT('h0100)
	) name17019 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001 ,
		_w21067_
	);
	LUT4 #(
		.INIT('h0001)
	) name17020 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w21065_,
		_w21066_,
		_w21067_,
		_w21068_
	);
	LUT2 #(
		.INIT('h8)
	) name17021 (
		_w21064_,
		_w21068_,
		_w21069_
	);
	LUT2 #(
		.INIT('h2)
	) name17022 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w20622_,
		_w21070_
	);
	LUT3 #(
		.INIT('ha2)
	) name17023 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w19945_,
		_w21070_,
		_w21071_
	);
	LUT2 #(
		.INIT('h4)
	) name17024 (
		_w19947_,
		_w21071_,
		_w21072_
	);
	LUT4 #(
		.INIT('hff02)
	) name17025 (
		_w19947_,
		_w21059_,
		_w21069_,
		_w21072_,
		_w21073_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17026 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w6378_,
		_w6498_,
		_w6500_,
		_w21074_
	);
	LUT4 #(
		.INIT('h0400)
	) name17027 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001 ,
		_w21075_
	);
	LUT4 #(
		.INIT('h4000)
	) name17028 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001 ,
		_w21076_
	);
	LUT4 #(
		.INIT('h0200)
	) name17029 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001 ,
		_w21077_
	);
	LUT4 #(
		.INIT('h2000)
	) name17030 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001 ,
		_w21078_
	);
	LUT4 #(
		.INIT('h0001)
	) name17031 (
		_w21075_,
		_w21076_,
		_w21077_,
		_w21078_,
		_w21079_
	);
	LUT4 #(
		.INIT('h1000)
	) name17032 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001 ,
		_w21080_
	);
	LUT4 #(
		.INIT('h0800)
	) name17033 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001 ,
		_w21081_
	);
	LUT4 #(
		.INIT('h0100)
	) name17034 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001 ,
		_w21082_
	);
	LUT4 #(
		.INIT('h0001)
	) name17035 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w21080_,
		_w21081_,
		_w21082_,
		_w21083_
	);
	LUT2 #(
		.INIT('h8)
	) name17036 (
		_w21079_,
		_w21083_,
		_w21084_
	);
	LUT3 #(
		.INIT('ha8)
	) name17037 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		_w21085_
	);
	LUT4 #(
		.INIT('h0045)
	) name17038 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4094_,
		_w4097_,
		_w21085_,
		_w21086_
	);
	LUT2 #(
		.INIT('h2)
	) name17039 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w21086_,
		_w21087_
	);
	LUT2 #(
		.INIT('h4)
	) name17040 (
		_w19947_,
		_w21087_,
		_w21088_
	);
	LUT4 #(
		.INIT('hff02)
	) name17041 (
		_w19947_,
		_w21074_,
		_w21084_,
		_w21088_,
		_w21089_
	);
	LUT3 #(
		.INIT('h6c)
	) name17042 (
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		_w14699_,
		_w21090_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17043 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w7257_,
		_w7375_,
		_w7377_,
		_w21091_
	);
	LUT4 #(
		.INIT('h0400)
	) name17044 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001 ,
		_w21092_
	);
	LUT4 #(
		.INIT('h4000)
	) name17045 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001 ,
		_w21093_
	);
	LUT4 #(
		.INIT('h0200)
	) name17046 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001 ,
		_w21094_
	);
	LUT4 #(
		.INIT('h2000)
	) name17047 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001 ,
		_w21095_
	);
	LUT4 #(
		.INIT('h0001)
	) name17048 (
		_w21092_,
		_w21093_,
		_w21094_,
		_w21095_,
		_w21096_
	);
	LUT4 #(
		.INIT('h1000)
	) name17049 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001 ,
		_w21097_
	);
	LUT4 #(
		.INIT('h0800)
	) name17050 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001 ,
		_w21098_
	);
	LUT4 #(
		.INIT('h0100)
	) name17051 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001 ,
		_w21099_
	);
	LUT4 #(
		.INIT('h0001)
	) name17052 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w21097_,
		_w21098_,
		_w21099_,
		_w21100_
	);
	LUT2 #(
		.INIT('h8)
	) name17053 (
		_w21096_,
		_w21100_,
		_w21101_
	);
	LUT2 #(
		.INIT('h2)
	) name17054 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w20466_,
		_w21102_
	);
	LUT4 #(
		.INIT('h0045)
	) name17055 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4094_,
		_w4097_,
		_w21102_,
		_w21103_
	);
	LUT2 #(
		.INIT('h2)
	) name17056 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w21103_,
		_w21104_
	);
	LUT2 #(
		.INIT('h4)
	) name17057 (
		_w19947_,
		_w21104_,
		_w21105_
	);
	LUT4 #(
		.INIT('hff02)
	) name17058 (
		_w19947_,
		_w21091_,
		_w21101_,
		_w21105_,
		_w21106_
	);
	LUT3 #(
		.INIT('h40)
	) name17059 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w21107_
	);
	LUT2 #(
		.INIT('h6)
	) name17060 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		_w17702_,
		_w21108_
	);
	LUT3 #(
		.INIT('hec)
	) name17061 (
		_w17734_,
		_w21107_,
		_w21108_,
		_w21109_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17062 (
		\sice_ICYC_reg[10]/NET0131 ,
		\sice_ICYC_reg[11]/NET0131 ,
		\sice_ICYC_reg[12]/NET0131 ,
		_w13015_,
		_w21110_
	);
	LUT3 #(
		.INIT('h40)
	) name17063 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w21111_
	);
	LUT2 #(
		.INIT('h6)
	) name17064 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		_w17666_,
		_w21112_
	);
	LUT3 #(
		.INIT('hec)
	) name17065 (
		_w17698_,
		_w21111_,
		_w21112_,
		_w21113_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17066 (
		\sice_IIRC_reg[10]/NET0131 ,
		\sice_IIRC_reg[11]/NET0131 ,
		\sice_IIRC_reg[12]/NET0131 ,
		_w13087_,
		_w21114_
	);
	LUT2 #(
		.INIT('h4)
	) name17067 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w21115_
	);
	LUT4 #(
		.INIT('h1055)
	) name17068 (
		_w6879_,
		_w16245_,
		_w16246_,
		_w16247_,
		_w21116_
	);
	LUT2 #(
		.INIT('h2)
	) name17069 (
		_w5882_,
		_w21116_,
		_w21117_
	);
	LUT4 #(
		.INIT('h8a00)
	) name17070 (
		_w6879_,
		_w16245_,
		_w16246_,
		_w16247_,
		_w21118_
	);
	LUT4 #(
		.INIT('h8088)
	) name17071 (
		_w6466_,
		_w16247_,
		_w16868_,
		_w16869_,
		_w21119_
	);
	LUT2 #(
		.INIT('h1)
	) name17072 (
		_w21118_,
		_w21119_,
		_w21120_
	);
	LUT3 #(
		.INIT('h51)
	) name17073 (
		_w6130_,
		_w16247_,
		_w18077_,
		_w21121_
	);
	LUT4 #(
		.INIT('h1511)
	) name17074 (
		_w6466_,
		_w16247_,
		_w16868_,
		_w16869_,
		_w21122_
	);
	LUT2 #(
		.INIT('h1)
	) name17075 (
		_w21121_,
		_w21122_,
		_w21123_
	);
	LUT4 #(
		.INIT('h4f00)
	) name17076 (
		_w14805_,
		_w21117_,
		_w21120_,
		_w21123_,
		_w21124_
	);
	LUT2 #(
		.INIT('h4)
	) name17077 (
		_w5742_,
		_w18071_,
		_w21125_
	);
	LUT3 #(
		.INIT('h08)
	) name17078 (
		_w6130_,
		_w16247_,
		_w18077_,
		_w21126_
	);
	LUT2 #(
		.INIT('h1)
	) name17079 (
		_w21125_,
		_w21126_,
		_w21127_
	);
	LUT2 #(
		.INIT('h2)
	) name17080 (
		_w5742_,
		_w18071_,
		_w21128_
	);
	LUT2 #(
		.INIT('h8)
	) name17081 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w21129_
	);
	LUT2 #(
		.INIT('h8)
	) name17082 (
		_w14774_,
		_w21129_,
		_w21130_
	);
	LUT3 #(
		.INIT('h10)
	) name17083 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w9453_,
		_w21130_,
		_w21131_
	);
	LUT2 #(
		.INIT('h4)
	) name17084 (
		_w21128_,
		_w21131_,
		_w21132_
	);
	LUT4 #(
		.INIT('h1055)
	) name17085 (
		_w21115_,
		_w21124_,
		_w21127_,
		_w21132_,
		_w21133_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17086 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w6774_,
		_w6894_,
		_w6896_,
		_w21134_
	);
	LUT4 #(
		.INIT('h1055)
	) name17087 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w16245_,
		_w16246_,
		_w16247_,
		_w21135_
	);
	LUT2 #(
		.INIT('h1)
	) name17088 (
		_w21134_,
		_w21135_,
		_w21136_
	);
	LUT4 #(
		.INIT('haea2)
	) name17089 (
		\core_eu_es_sht_es_reg_SBs_reg[1]/P0001 ,
		_w9893_,
		_w21133_,
		_w21136_,
		_w21137_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17090 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w5784_,
		_w5911_,
		_w5913_,
		_w21138_
	);
	LUT3 #(
		.INIT('h0b)
	) name17091 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w14805_,
		_w21138_,
		_w21139_
	);
	LUT4 #(
		.INIT('haea2)
	) name17092 (
		\core_eu_es_sht_es_reg_SBs_reg[0]/P0001 ,
		_w9893_,
		_w21133_,
		_w21139_,
		_w21140_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17093 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w6054_,
		_w6173_,
		_w6175_,
		_w21141_
	);
	LUT3 #(
		.INIT('h51)
	) name17094 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w16247_,
		_w18077_,
		_w21142_
	);
	LUT2 #(
		.INIT('h1)
	) name17095 (
		_w21141_,
		_w21142_,
		_w21143_
	);
	LUT4 #(
		.INIT('haea2)
	) name17096 (
		\core_eu_es_sht_es_reg_SBs_reg[3]/P0001 ,
		_w9893_,
		_w21133_,
		_w21143_,
		_w21144_
	);
	LUT4 #(
		.INIT('haea2)
	) name17097 (
		\core_eu_es_sht_es_reg_SBr_reg[3]/P0001 ,
		_w9452_,
		_w21133_,
		_w21143_,
		_w21145_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17098 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w6378_,
		_w6498_,
		_w6500_,
		_w21146_
	);
	LUT4 #(
		.INIT('h1511)
	) name17099 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w16247_,
		_w16868_,
		_w16869_,
		_w21147_
	);
	LUT2 #(
		.INIT('h1)
	) name17100 (
		_w21146_,
		_w21147_,
		_w21148_
	);
	LUT4 #(
		.INIT('haea2)
	) name17101 (
		\core_eu_es_sht_es_reg_SBs_reg[2]/P0001 ,
		_w9893_,
		_w21133_,
		_w21148_,
		_w21149_
	);
	LUT4 #(
		.INIT('haea2)
	) name17102 (
		\core_eu_es_sht_es_reg_SBr_reg[2]/P0001 ,
		_w9452_,
		_w21133_,
		_w21148_,
		_w21150_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17103 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w7257_,
		_w7375_,
		_w7377_,
		_w21151_
	);
	LUT2 #(
		.INIT('h4)
	) name17104 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w18071_,
		_w21152_
	);
	LUT2 #(
		.INIT('h1)
	) name17105 (
		_w21151_,
		_w21152_,
		_w21153_
	);
	LUT4 #(
		.INIT('haea2)
	) name17106 (
		\core_eu_es_sht_es_reg_SBr_reg[4]/P0001 ,
		_w9452_,
		_w21133_,
		_w21153_,
		_w21154_
	);
	LUT4 #(
		.INIT('haea2)
	) name17107 (
		\core_eu_es_sht_es_reg_SBr_reg[1]/P0001 ,
		_w9452_,
		_w21133_,
		_w21136_,
		_w21155_
	);
	LUT4 #(
		.INIT('haea2)
	) name17108 (
		\core_eu_es_sht_es_reg_SBs_reg[4]/P0001 ,
		_w9893_,
		_w21133_,
		_w21153_,
		_w21156_
	);
	LUT4 #(
		.INIT('haea2)
	) name17109 (
		\core_eu_es_sht_es_reg_SBr_reg[0]/P0001 ,
		_w9452_,
		_w21133_,
		_w21139_,
		_w21157_
	);
	LUT3 #(
		.INIT('h13)
	) name17110 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001 ,
		_w9894_,
		_w21158_
	);
	LUT4 #(
		.INIT('h0002)
	) name17111 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w21158_,
		_w21159_
	);
	LUT4 #(
		.INIT('h313b)
	) name17112 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001 ,
		_w11631_,
		_w11635_,
		_w21160_
	);
	LUT4 #(
		.INIT('h2f00)
	) name17113 (
		_w11625_,
		_w12284_,
		_w21159_,
		_w21160_,
		_w21161_
	);
	LUT2 #(
		.INIT('h1)
	) name17114 (
		_w11624_,
		_w21161_,
		_w21162_
	);
	LUT3 #(
		.INIT('hf2)
	) name17115 (
		_w11624_,
		_w12350_,
		_w21162_,
		_w21163_
	);
	LUT2 #(
		.INIT('h2)
	) name17116 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001 ,
		_w11656_,
		_w21164_
	);
	LUT3 #(
		.INIT('h01)
	) name17117 (
		_w9946_,
		_w11659_,
		_w21164_,
		_w21165_
	);
	LUT3 #(
		.INIT('h70)
	) name17118 (
		_w11655_,
		_w12284_,
		_w21165_,
		_w21166_
	);
	LUT3 #(
		.INIT('h07)
	) name17119 (
		_w9946_,
		_w12350_,
		_w21166_,
		_w21167_
	);
	LUT3 #(
		.INIT('h60)
	) name17120 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w21168_
	);
	LUT4 #(
		.INIT('h51a2)
	) name17121 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w21169_
	);
	LUT4 #(
		.INIT('h4544)
	) name17122 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13110_,
		_w21168_,
		_w21169_,
		_w21170_
	);
	LUT2 #(
		.INIT('h2)
	) name17123 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w21171_
	);
	LUT2 #(
		.INIT('h2)
	) name17124 (
		_w19097_,
		_w21171_,
		_w21172_
	);
	LUT3 #(
		.INIT('ha8)
	) name17125 (
		_w13098_,
		_w21170_,
		_w21172_,
		_w21173_
	);
	LUT3 #(
		.INIT('h10)
	) name17126 (
		_w13098_,
		_w19093_,
		_w19094_,
		_w21174_
	);
	LUT2 #(
		.INIT('h1)
	) name17127 (
		_w21173_,
		_w21174_,
		_w21175_
	);
	LUT4 #(
		.INIT('h8db1)
	) name17128 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w21176_
	);
	LUT4 #(
		.INIT('h1302)
	) name17129 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13122_,
		_w21176_,
		_w21177_
	);
	LUT4 #(
		.INIT('hfe54)
	) name17130 (
		_w13098_,
		_w21170_,
		_w21172_,
		_w21177_,
		_w21178_
	);
	LUT4 #(
		.INIT('h0040)
	) name17131 (
		_w13147_,
		_w13152_,
		_w21175_,
		_w21178_,
		_w21179_
	);
	LUT4 #(
		.INIT('h40bf)
	) name17132 (
		_w13147_,
		_w13152_,
		_w21175_,
		_w21178_,
		_w21180_
	);
	LUT4 #(
		.INIT('h1555)
	) name17133 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w19091_,
		_w19096_,
		_w21175_,
		_w21181_
	);
	LUT3 #(
		.INIT('h82)
	) name17134 (
		_w13155_,
		_w21180_,
		_w21181_,
		_w21182_
	);
	LUT3 #(
		.INIT('h40)
	) name17135 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[8]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w21183_
	);
	LUT2 #(
		.INIT('h1)
	) name17136 (
		_w13158_,
		_w21183_,
		_w21184_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17137 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w7465_,
		_w7565_,
		_w21184_,
		_w21185_
	);
	LUT4 #(
		.INIT('hafac)
	) name17138 (
		\sport0_rxctl_RXSHT_reg[8]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w21186_
	);
	LUT4 #(
		.INIT('h0002)
	) name17139 (
		\sport0_rxctl_RX_reg[8]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w21187_
	);
	LUT4 #(
		.INIT('hffb0)
	) name17140 (
		_w21182_,
		_w21185_,
		_w21186_,
		_w21187_,
		_w21188_
	);
	LUT4 #(
		.INIT('h7200)
	) name17141 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11294_,
		_w11296_,
		_w11624_,
		_w21189_
	);
	LUT2 #(
		.INIT('h1)
	) name17142 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001 ,
		_w17501_,
		_w21190_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17143 (
		_w11313_,
		_w11314_,
		_w12220_,
		_w17505_,
		_w21191_
	);
	LUT4 #(
		.INIT('h1311)
	) name17144 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001 ,
		_w11303_,
		_w11308_,
		_w21192_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17145 (
		_w12224_,
		_w21190_,
		_w21191_,
		_w21192_,
		_w21193_
	);
	LUT2 #(
		.INIT('h2)
	) name17146 (
		_w17500_,
		_w21193_,
		_w21194_
	);
	LUT2 #(
		.INIT('h1)
	) name17147 (
		_w21189_,
		_w21194_,
		_w21195_
	);
	LUT4 #(
		.INIT('h0804)
	) name17148 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w21196_
	);
	LUT4 #(
		.INIT('h0004)
	) name17149 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13098_,
		_w13143_,
		_w21196_,
		_w21197_
	);
	LUT3 #(
		.INIT('h0b)
	) name17150 (
		_w13098_,
		_w21177_,
		_w21197_,
		_w21198_
	);
	LUT2 #(
		.INIT('h8)
	) name17151 (
		_w21179_,
		_w21198_,
		_w21199_
	);
	LUT4 #(
		.INIT('h8000)
	) name17152 (
		_w19091_,
		_w19096_,
		_w21175_,
		_w21180_,
		_w21200_
	);
	LUT4 #(
		.INIT('h0001)
	) name17153 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w13098_,
		_w13143_,
		_w21196_,
		_w21201_
	);
	LUT3 #(
		.INIT('h20)
	) name17154 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w19092_,
		_w21202_
	);
	LUT2 #(
		.INIT('h1)
	) name17155 (
		_w21201_,
		_w21202_,
		_w21203_
	);
	LUT3 #(
		.INIT('h1e)
	) name17156 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w21200_,
		_w21203_,
		_w21204_
	);
	LUT3 #(
		.INIT('h40)
	) name17157 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[10]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w21205_
	);
	LUT2 #(
		.INIT('h1)
	) name17158 (
		_w13158_,
		_w21205_,
		_w21206_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17159 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w5937_,
		_w6038_,
		_w21206_,
		_w21207_
	);
	LUT4 #(
		.INIT('hd700)
	) name17160 (
		_w13155_,
		_w21199_,
		_w21204_,
		_w21207_,
		_w21208_
	);
	LUT4 #(
		.INIT('hafac)
	) name17161 (
		\sport0_rxctl_RXSHT_reg[10]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w21209_
	);
	LUT4 #(
		.INIT('h0002)
	) name17162 (
		\sport0_rxctl_RX_reg[10]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w21210_
	);
	LUT3 #(
		.INIT('hf4)
	) name17163 (
		_w21208_,
		_w21209_,
		_w21210_,
		_w21211_
	);
	LUT4 #(
		.INIT('h0001)
	) name17164 (
		\idma_DCTL_reg[11]/NET0131 ,
		\idma_DCTL_reg[12]/NET0131 ,
		\idma_DCTL_reg[13]/NET0131 ,
		\idma_DCTL_reg[1]/NET0131 ,
		_w21212_
	);
	LUT4 #(
		.INIT('h0001)
	) name17165 (
		\idma_DCTL_reg[0]/NET0131 ,
		\idma_DCTL_reg[10]/NET0131 ,
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		_w21213_
	);
	LUT4 #(
		.INIT('h0001)
	) name17166 (
		\idma_DCTL_reg[6]/NET0131 ,
		\idma_DCTL_reg[7]/NET0131 ,
		\idma_DCTL_reg[8]/NET0131 ,
		\idma_DCTL_reg[9]/NET0131 ,
		_w21214_
	);
	LUT4 #(
		.INIT('h0001)
	) name17167 (
		\idma_DCTL_reg[2]/NET0131 ,
		\idma_DCTL_reg[3]/NET0131 ,
		\idma_DCTL_reg[4]/NET0131 ,
		\idma_DCTL_reg[5]/NET0131 ,
		_w21215_
	);
	LUT4 #(
		.INIT('h8000)
	) name17168 (
		_w21214_,
		_w21215_,
		_w21212_,
		_w21213_,
		_w21216_
	);
	LUT3 #(
		.INIT('h15)
	) name17169 (
		_w4065_,
		_w19997_,
		_w21216_,
		_w21217_
	);
	LUT2 #(
		.INIT('h6)
	) name17170 (
		\clkc_OUTcnt_reg[4]/NET0131 ,
		_w12252_,
		_w21218_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17171 (
		_w12254_,
		_w12258_,
		_w12263_,
		_w21218_,
		_w21219_
	);
	LUT2 #(
		.INIT('h6)
	) name17172 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		_w19390_,
		_w21220_
	);
	LUT3 #(
		.INIT('h70)
	) name17173 (
		_w19400_,
		_w19405_,
		_w21220_,
		_w21221_
	);
	LUT4 #(
		.INIT('h3031)
	) name17174 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w4971_,
		_w9911_,
		_w21222_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17175 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w5784_,
		_w5911_,
		_w5913_,
		_w21223_
	);
	LUT4 #(
		.INIT('h4000)
	) name17176 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001 ,
		_w21224_
	);
	LUT4 #(
		.INIT('h0400)
	) name17177 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001 ,
		_w21225_
	);
	LUT4 #(
		.INIT('h0100)
	) name17178 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001 ,
		_w21226_
	);
	LUT4 #(
		.INIT('h0200)
	) name17179 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001 ,
		_w21227_
	);
	LUT4 #(
		.INIT('h0001)
	) name17180 (
		_w21224_,
		_w21225_,
		_w21226_,
		_w21227_,
		_w21228_
	);
	LUT4 #(
		.INIT('h0800)
	) name17181 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001 ,
		_w21229_
	);
	LUT4 #(
		.INIT('h2000)
	) name17182 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001 ,
		_w21230_
	);
	LUT4 #(
		.INIT('h1000)
	) name17183 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001 ,
		_w21231_
	);
	LUT4 #(
		.INIT('h0001)
	) name17184 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w21229_,
		_w21230_,
		_w21231_,
		_w21232_
	);
	LUT2 #(
		.INIT('h8)
	) name17185 (
		_w21228_,
		_w21232_,
		_w21233_
	);
	LUT4 #(
		.INIT('h1115)
	) name17186 (
		_w19945_,
		_w19946_,
		_w21223_,
		_w21233_,
		_w21234_
	);
	LUT2 #(
		.INIT('h4)
	) name17187 (
		_w21222_,
		_w21234_,
		_w21235_
	);
	LUT4 #(
		.INIT('h2000)
	) name17188 (
		\core_c_dec_MTTX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21236_
	);
	LUT4 #(
		.INIT('h1110)
	) name17189 (
		_w19710_,
		_w19711_,
		_w19713_,
		_w19714_,
		_w21237_
	);
	LUT4 #(
		.INIT('h00bf)
	) name17190 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19705_,
		_w21238_
	);
	LUT4 #(
		.INIT('h4000)
	) name17191 (
		_w19701_,
		_w19732_,
		_w21237_,
		_w21238_,
		_w21239_
	);
	LUT3 #(
		.INIT('ha8)
	) name17192 (
		_w4102_,
		_w21236_,
		_w21239_,
		_w21240_
	);
	LUT4 #(
		.INIT('h2000)
	) name17193 (
		\core_c_dec_MTTX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21241_
	);
	LUT4 #(
		.INIT('h4000)
	) name17194 (
		_w19701_,
		_w19729_,
		_w19732_,
		_w21238_,
		_w21242_
	);
	LUT3 #(
		.INIT('ha8)
	) name17195 (
		_w4102_,
		_w21241_,
		_w21242_,
		_w21243_
	);
	LUT4 #(
		.INIT('h2000)
	) name17196 (
		\core_c_dec_MTMreg_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21244_
	);
	LUT4 #(
		.INIT('h000e)
	) name17197 (
		_w19127_,
		_w19232_,
		_w19707_,
		_w19708_,
		_w21245_
	);
	LUT2 #(
		.INIT('h4)
	) name17198 (
		_w19712_,
		_w21245_,
		_w21246_
	);
	LUT4 #(
		.INIT('h1110)
	) name17199 (
		_w19713_,
		_w19714_,
		_w19703_,
		_w19704_,
		_w21247_
	);
	LUT4 #(
		.INIT('h5053)
	) name17200 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w19034_,
		_w19124_,
		_w21248_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17201 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21248_,
		_w21249_
	);
	LUT4 #(
		.INIT('h1555)
	) name17202 (
		_w21244_,
		_w21246_,
		_w21247_,
		_w21249_,
		_w21250_
	);
	LUT2 #(
		.INIT('h2)
	) name17203 (
		_w4102_,
		_w21250_,
		_w21251_
	);
	LUT2 #(
		.INIT('h9)
	) name17204 (
		\sport1_txctl_Bcnt_reg[4]/NET0131 ,
		_w14267_,
		_w21252_
	);
	LUT3 #(
		.INIT('h10)
	) name17205 (
		_w14590_,
		_w14591_,
		_w21252_,
		_w21253_
	);
	LUT4 #(
		.INIT('h2223)
	) name17206 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w14590_,
		_w14591_,
		_w21254_
	);
	LUT2 #(
		.INIT('h4)
	) name17207 (
		_w21253_,
		_w21254_,
		_w21255_
	);
	LUT2 #(
		.INIT('h9)
	) name17208 (
		\sport0_txctl_Bcnt_reg[4]/NET0131 ,
		_w12550_,
		_w21256_
	);
	LUT3 #(
		.INIT('h10)
	) name17209 (
		_w14596_,
		_w14597_,
		_w21256_,
		_w21257_
	);
	LUT4 #(
		.INIT('h2223)
	) name17210 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w14596_,
		_w14597_,
		_w21258_
	);
	LUT2 #(
		.INIT('h4)
	) name17211 (
		_w21257_,
		_w21258_,
		_w21259_
	);
	LUT3 #(
		.INIT('he0)
	) name17212 (
		_w7140_,
		_w7240_,
		_w9432_,
		_w21260_
	);
	LUT4 #(
		.INIT('h00de)
	) name17213 (
		\bdma_BWCOUNT_reg[9]/NET0131 ,
		_w9432_,
		_w20503_,
		_w21260_,
		_w21261_
	);
	LUT3 #(
		.INIT('he0)
	) name17214 (
		_w7465_,
		_w7565_,
		_w9432_,
		_w21262_
	);
	LUT4 #(
		.INIT('h0603)
	) name17215 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		\bdma_BWCOUNT_reg[8]/NET0131 ,
		_w9432_,
		_w20502_,
		_w21263_
	);
	LUT2 #(
		.INIT('h1)
	) name17216 (
		_w21262_,
		_w21263_,
		_w21264_
	);
	LUT2 #(
		.INIT('h4)
	) name17217 (
		_w6758_,
		_w9432_,
		_w21265_
	);
	LUT4 #(
		.INIT('h00de)
	) name17218 (
		\bdma_BWCOUNT_reg[12]/NET0131 ,
		_w9432_,
		_w20505_,
		_w21265_,
		_w21266_
	);
	LUT3 #(
		.INIT('he0)
	) name17219 (
		_w5937_,
		_w6038_,
		_w9432_,
		_w21267_
	);
	LUT4 #(
		.INIT('h00de)
	) name17220 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		_w9432_,
		_w20504_,
		_w21267_,
		_w21268_
	);
	LUT4 #(
		.INIT('h060c)
	) name17221 (
		\bdma_BIAD_reg[8]/NET0131 ,
		\bdma_BIAD_reg[9]/NET0131 ,
		_w21001_,
		_w20998_,
		_w21269_
	);
	LUT3 #(
		.INIT('h10)
	) name17222 (
		_w7140_,
		_w7240_,
		_w21001_,
		_w21270_
	);
	LUT2 #(
		.INIT('he)
	) name17223 (
		_w21269_,
		_w21270_,
		_w21271_
	);
	LUT3 #(
		.INIT('h10)
	) name17224 (
		_w7465_,
		_w7565_,
		_w21001_,
		_w21272_
	);
	LUT4 #(
		.INIT('hff12)
	) name17225 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w21001_,
		_w20998_,
		_w21272_,
		_w21273_
	);
	LUT4 #(
		.INIT('h870f)
	) name17226 (
		\bdma_BIAD_reg[11]/NET0131 ,
		\bdma_BIAD_reg[12]/NET0131 ,
		\bdma_BIAD_reg[13]/NET0131 ,
		_w21000_,
		_w21274_
	);
	LUT2 #(
		.INIT('h8)
	) name17227 (
		_w5760_,
		_w21001_,
		_w21275_
	);
	LUT3 #(
		.INIT('hf1)
	) name17228 (
		_w21001_,
		_w21274_,
		_w21275_,
		_w21276_
	);
	LUT3 #(
		.INIT('h10)
	) name17229 (
		_w5937_,
		_w6038_,
		_w21001_,
		_w21277_
	);
	LUT4 #(
		.INIT('hff12)
	) name17230 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w21001_,
		_w20999_,
		_w21277_,
		_w21278_
	);
	LUT4 #(
		.INIT('h060c)
	) name17231 (
		\bdma_BEAD_reg[8]/NET0131 ,
		\bdma_BEAD_reg[9]/NET0131 ,
		_w13032_,
		_w20512_,
		_w21279_
	);
	LUT3 #(
		.INIT('h10)
	) name17232 (
		_w7140_,
		_w7240_,
		_w13032_,
		_w21280_
	);
	LUT2 #(
		.INIT('he)
	) name17233 (
		_w21279_,
		_w21280_,
		_w21281_
	);
	LUT3 #(
		.INIT('h10)
	) name17234 (
		_w7465_,
		_w7565_,
		_w13032_,
		_w21282_
	);
	LUT4 #(
		.INIT('hff12)
	) name17235 (
		\bdma_BEAD_reg[8]/NET0131 ,
		_w13032_,
		_w20512_,
		_w21282_,
		_w21283_
	);
	LUT3 #(
		.INIT('h10)
	) name17236 (
		_w5937_,
		_w6038_,
		_w13032_,
		_w21284_
	);
	LUT4 #(
		.INIT('hff12)
	) name17237 (
		\bdma_BEAD_reg[10]/NET0131 ,
		_w13032_,
		_w20513_,
		_w21284_,
		_w21285_
	);
	LUT3 #(
		.INIT('hca)
	) name17238 (
		\sport1_txctl_TXSHT_reg[3]/P0001 ,
		\sport1_txctl_TX_reg[4]/P0001 ,
		_w14269_,
		_w21286_
	);
	LUT4 #(
		.INIT('h2000)
	) name17239 (
		\core_c_dec_MFSPT_Ei_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21287_
	);
	LUT4 #(
		.INIT('h1110)
	) name17240 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w19040_,
		_w19231_,
		_w19232_,
		_w21288_
	);
	LUT2 #(
		.INIT('h4)
	) name17241 (
		_w19238_,
		_w21288_,
		_w21289_
	);
	LUT3 #(
		.INIT('hec)
	) name17242 (
		_w16007_,
		_w21287_,
		_w21289_,
		_w21290_
	);
	LUT4 #(
		.INIT('hba00)
	) name17243 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w9432_,
		_w21291_
	);
	LUT4 #(
		.INIT('h00de)
	) name17244 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		_w9432_,
		_w20502_,
		_w21291_,
		_w21292_
	);
	LUT4 #(
		.INIT('hba00)
	) name17245 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w9432_,
		_w21293_
	);
	LUT2 #(
		.INIT('h1)
	) name17246 (
		_w9432_,
		_w20502_,
		_w21294_
	);
	LUT4 #(
		.INIT('h020f)
	) name17247 (
		\bdma_BWCOUNT_reg[6]/NET0131 ,
		_w9429_,
		_w21293_,
		_w21294_,
		_w21295_
	);
	LUT3 #(
		.INIT('hca)
	) name17248 (
		\sport0_txctl_TXSHT_reg[3]/P0001 ,
		\sport0_txctl_TX_reg[4]/P0001 ,
		_w12552_,
		_w21296_
	);
	LUT4 #(
		.INIT('he0f0)
	) name17249 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		\bdma_BWCOUNT_reg[3]/NET0131 ,
		\bdma_BWCOUNT_reg[4]/NET0131 ,
		_w9427_,
		_w21297_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name17250 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		_w9416_,
		_w9432_,
		_w9427_,
		_w21298_
	);
	LUT4 #(
		.INIT('hba00)
	) name17251 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w9432_,
		_w21299_
	);
	LUT3 #(
		.INIT('h0b)
	) name17252 (
		_w21297_,
		_w21298_,
		_w21299_,
		_w21300_
	);
	LUT4 #(
		.INIT('h0603)
	) name17253 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		\bdma_BWCOUNT_reg[3]/NET0131 ,
		_w9432_,
		_w9427_,
		_w21301_
	);
	LUT4 #(
		.INIT('hba00)
	) name17254 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w9432_,
		_w21302_
	);
	LUT2 #(
		.INIT('h1)
	) name17255 (
		_w21301_,
		_w21302_,
		_w21303_
	);
	LUT4 #(
		.INIT('hba00)
	) name17256 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w9432_,
		_w21304_
	);
	LUT4 #(
		.INIT('h00de)
	) name17257 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		_w9432_,
		_w9427_,
		_w21304_,
		_w21305_
	);
	LUT4 #(
		.INIT('h00a9)
	) name17258 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		_w9414_,
		_w9415_,
		_w9432_,
		_w21306_
	);
	LUT4 #(
		.INIT('hba00)
	) name17259 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w9432_,
		_w21307_
	);
	LUT2 #(
		.INIT('h1)
	) name17260 (
		_w21306_,
		_w21307_,
		_w21308_
	);
	LUT4 #(
		.INIT('h060c)
	) name17261 (
		\bdma_BIAD_reg[5]/NET0131 ,
		\bdma_BIAD_reg[6]/NET0131 ,
		_w21001_,
		_w20996_,
		_w21309_
	);
	LUT4 #(
		.INIT('h4500)
	) name17262 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w21001_,
		_w21310_
	);
	LUT2 #(
		.INIT('he)
	) name17263 (
		_w21309_,
		_w21310_,
		_w21311_
	);
	LUT4 #(
		.INIT('h4500)
	) name17264 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w21001_,
		_w21312_
	);
	LUT4 #(
		.INIT('hff12)
	) name17265 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w21001_,
		_w20997_,
		_w21312_,
		_w21313_
	);
	LUT4 #(
		.INIT('h4500)
	) name17266 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w21001_,
		_w21314_
	);
	LUT4 #(
		.INIT('hff12)
	) name17267 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w21001_,
		_w20996_,
		_w21314_,
		_w21315_
	);
	LUT4 #(
		.INIT('h4500)
	) name17268 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w21001_,
		_w21316_
	);
	LUT4 #(
		.INIT('hff12)
	) name17269 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w21001_,
		_w20995_,
		_w21316_,
		_w21317_
	);
	LUT4 #(
		.INIT('h060c)
	) name17270 (
		\bdma_BIAD_reg[2]/NET0131 ,
		\bdma_BIAD_reg[3]/NET0131 ,
		_w21001_,
		_w20994_,
		_w21318_
	);
	LUT4 #(
		.INIT('h4500)
	) name17271 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w21001_,
		_w21319_
	);
	LUT2 #(
		.INIT('he)
	) name17272 (
		_w21318_,
		_w21319_,
		_w21320_
	);
	LUT4 #(
		.INIT('h4500)
	) name17273 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w21001_,
		_w21321_
	);
	LUT4 #(
		.INIT('hff12)
	) name17274 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w21001_,
		_w20994_,
		_w21321_,
		_w21322_
	);
	LUT4 #(
		.INIT('h4500)
	) name17275 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w21001_,
		_w21323_
	);
	LUT4 #(
		.INIT('hff12)
	) name17276 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w21001_,
		_w20993_,
		_w21323_,
		_w21324_
	);
	LUT4 #(
		.INIT('h0056)
	) name17277 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w9414_,
		_w9415_,
		_w21001_,
		_w21325_
	);
	LUT4 #(
		.INIT('h4500)
	) name17278 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w21001_,
		_w21326_
	);
	LUT2 #(
		.INIT('he)
	) name17279 (
		_w21325_,
		_w21326_,
		_w21327_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name17280 (
		\sice_IIRC_reg[5]/NET0131 ,
		_w11935_,
		_w19738_,
		_w19739_,
		_w21328_
	);
	LUT3 #(
		.INIT('h6a)
	) name17281 (
		\sice_IIRC_reg[0]/NET0131 ,
		_w19738_,
		_w19739_,
		_w21329_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name17282 (
		\sice_IIRC_reg[18]/NET0131 ,
		_w14202_,
		_w19738_,
		_w19739_,
		_w21330_
	);
	LUT2 #(
		.INIT('h6)
	) name17283 (
		\sice_IIRC_reg[19]/NET0131 ,
		_w19741_,
		_w21331_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17284 (
		\sice_IIRC_reg[19]/NET0131 ,
		\sice_IIRC_reg[20]/NET0131 ,
		\sice_IIRC_reg[21]/NET0131 ,
		_w19741_,
		_w21332_
	);
	LUT2 #(
		.INIT('h6)
	) name17285 (
		\sice_IIRC_reg[22]/NET0131 ,
		_w21056_,
		_w21333_
	);
	LUT2 #(
		.INIT('h6)
	) name17286 (
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		_w14699_,
		_w21334_
	);
	LUT4 #(
		.INIT('h0200)
	) name17287 (
		\core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w21335_
	);
	LUT3 #(
		.INIT('h0b)
	) name17288 (
		_w12398_,
		_w13536_,
		_w21335_,
		_w21336_
	);
	LUT4 #(
		.INIT('h2000)
	) name17289 (
		\core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w21337_
	);
	LUT4 #(
		.INIT('h0020)
	) name17290 (
		\core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w21338_
	);
	LUT4 #(
		.INIT('h0002)
	) name17291 (
		\core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w21339_
	);
	LUT3 #(
		.INIT('h01)
	) name17292 (
		_w21338_,
		_w21339_,
		_w21337_,
		_w21340_
	);
	LUT2 #(
		.INIT('h8)
	) name17293 (
		_w21336_,
		_w21340_,
		_w21341_
	);
	LUT3 #(
		.INIT('h10)
	) name17294 (
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w12398_,
		_w13536_,
		_w21342_
	);
	LUT4 #(
		.INIT('h002f)
	) name17295 (
		_w5760_,
		_w20281_,
		_w21341_,
		_w21342_,
		_w21343_
	);
	LUT4 #(
		.INIT('h0200)
	) name17296 (
		\core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w21344_
	);
	LUT3 #(
		.INIT('h0b)
	) name17297 (
		_w12398_,
		_w13536_,
		_w21344_,
		_w21345_
	);
	LUT4 #(
		.INIT('h2000)
	) name17298 (
		\core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w21346_
	);
	LUT4 #(
		.INIT('h0020)
	) name17299 (
		\core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w21347_
	);
	LUT4 #(
		.INIT('h0002)
	) name17300 (
		\core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w21348_
	);
	LUT3 #(
		.INIT('h01)
	) name17301 (
		_w21347_,
		_w21348_,
		_w21346_,
		_w21349_
	);
	LUT2 #(
		.INIT('h8)
	) name17302 (
		_w21345_,
		_w21349_,
		_w21350_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17303 (
		_w5937_,
		_w6038_,
		_w20281_,
		_w21350_,
		_w21351_
	);
	LUT3 #(
		.INIT('h10)
	) name17304 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		_w12398_,
		_w13536_,
		_w21352_
	);
	LUT2 #(
		.INIT('h1)
	) name17305 (
		_w21351_,
		_w21352_,
		_w21353_
	);
	LUT4 #(
		.INIT('h45cf)
	) name17306 (
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w21354_
	);
	LUT2 #(
		.INIT('h8)
	) name17307 (
		\core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 ,
		_w20743_,
		_w21355_
	);
	LUT4 #(
		.INIT('h153f)
	) name17308 (
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 ,
		_w20742_,
		_w20740_,
		_w21356_
	);
	LUT3 #(
		.INIT('h40)
	) name17309 (
		_w21355_,
		_w21354_,
		_w21356_,
		_w21357_
	);
	LUT3 #(
		.INIT('h10)
	) name17310 (
		\core_dag_ilm2reg_I_reg[8]/NET0131 ,
		_w12398_,
		_w13536_,
		_w21358_
	);
	LUT4 #(
		.INIT('h002f)
	) name17311 (
		_w12913_,
		_w20737_,
		_w21357_,
		_w21358_,
		_w21359_
	);
	LUT4 #(
		.INIT('h45cf)
	) name17312 (
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w21360_
	);
	LUT2 #(
		.INIT('h8)
	) name17313 (
		\core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 ,
		_w20743_,
		_w21361_
	);
	LUT4 #(
		.INIT('h153f)
	) name17314 (
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 ,
		_w20742_,
		_w20740_,
		_w21362_
	);
	LUT3 #(
		.INIT('h40)
	) name17315 (
		_w21361_,
		_w21360_,
		_w21362_,
		_w21363_
	);
	LUT3 #(
		.INIT('h10)
	) name17316 (
		\core_dag_ilm2reg_I_reg[11]/NET0131 ,
		_w12398_,
		_w13536_,
		_w21364_
	);
	LUT4 #(
		.INIT('h001f)
	) name17317 (
		_w12991_,
		_w20737_,
		_w21363_,
		_w21364_,
		_w21365_
	);
	LUT4 #(
		.INIT('h45cf)
	) name17318 (
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w21366_
	);
	LUT2 #(
		.INIT('h8)
	) name17319 (
		\core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 ,
		_w20743_,
		_w21367_
	);
	LUT4 #(
		.INIT('h153f)
	) name17320 (
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 ,
		_w20742_,
		_w20740_,
		_w21368_
	);
	LUT3 #(
		.INIT('h40)
	) name17321 (
		_w21367_,
		_w21366_,
		_w21368_,
		_w21369_
	);
	LUT3 #(
		.INIT('h10)
	) name17322 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		_w12398_,
		_w13536_,
		_w21370_
	);
	LUT4 #(
		.INIT('h002f)
	) name17323 (
		_w13000_,
		_w20737_,
		_w21369_,
		_w21370_,
		_w21371_
	);
	LUT4 #(
		.INIT('h0200)
	) name17324 (
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w21372_
	);
	LUT2 #(
		.INIT('h1)
	) name17325 (
		_w13546_,
		_w21372_,
		_w21373_
	);
	LUT4 #(
		.INIT('h0200)
	) name17326 (
		\core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w21374_
	);
	LUT4 #(
		.INIT('h0200)
	) name17327 (
		\core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w21375_
	);
	LUT4 #(
		.INIT('h0200)
	) name17328 (
		\core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w21376_
	);
	LUT3 #(
		.INIT('h01)
	) name17329 (
		_w21375_,
		_w21376_,
		_w21374_,
		_w21377_
	);
	LUT2 #(
		.INIT('h8)
	) name17330 (
		_w21373_,
		_w21377_,
		_w21378_
	);
	LUT2 #(
		.INIT('h4)
	) name17331 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		_w13546_,
		_w21379_
	);
	LUT4 #(
		.INIT('h001f)
	) name17332 (
		_w15052_,
		_w20859_,
		_w21378_,
		_w21379_,
		_w21380_
	);
	LUT4 #(
		.INIT('h0045)
	) name17333 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w20281_,
		_w21381_
	);
	LUT4 #(
		.INIT('h2000)
	) name17334 (
		\core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131 ,
		_w16064_,
		_w20274_,
		_w20278_,
		_w21382_
	);
	LUT3 #(
		.INIT('h0b)
	) name17335 (
		_w12398_,
		_w13536_,
		_w21382_,
		_w21383_
	);
	LUT4 #(
		.INIT('h0200)
	) name17336 (
		\core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131 ,
		_w16061_,
		_w20274_,
		_w20278_,
		_w21384_
	);
	LUT4 #(
		.INIT('h0002)
	) name17337 (
		\core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131 ,
		_w16060_,
		_w20274_,
		_w20278_,
		_w21385_
	);
	LUT4 #(
		.INIT('h0020)
	) name17338 (
		\core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131 ,
		_w16068_,
		_w20274_,
		_w20278_,
		_w21386_
	);
	LUT3 #(
		.INIT('h01)
	) name17339 (
		_w21385_,
		_w21386_,
		_w21384_,
		_w21387_
	);
	LUT2 #(
		.INIT('h8)
	) name17340 (
		_w21383_,
		_w21387_,
		_w21388_
	);
	LUT3 #(
		.INIT('h10)
	) name17341 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		_w12398_,
		_w13536_,
		_w21389_
	);
	LUT3 #(
		.INIT('h0b)
	) name17342 (
		_w21381_,
		_w21388_,
		_w21389_,
		_w21390_
	);
	LUT4 #(
		.INIT('h45cf)
	) name17343 (
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		_w12398_,
		_w13536_,
		_w20738_,
		_w21391_
	);
	LUT2 #(
		.INIT('h8)
	) name17344 (
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		_w20740_,
		_w21392_
	);
	LUT4 #(
		.INIT('h153f)
	) name17345 (
		\core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 ,
		\core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 ,
		_w20742_,
		_w20743_,
		_w21393_
	);
	LUT3 #(
		.INIT('h40)
	) name17346 (
		_w21392_,
		_w21391_,
		_w21393_,
		_w21394_
	);
	LUT3 #(
		.INIT('h10)
	) name17347 (
		\core_dag_ilm2reg_I_reg[7]/NET0131 ,
		_w12398_,
		_w13536_,
		_w21395_
	);
	LUT4 #(
		.INIT('h002f)
	) name17348 (
		_w12923_,
		_w20737_,
		_w21394_,
		_w21395_,
		_w21396_
	);
	LUT4 #(
		.INIT('h00b1)
	) name17349 (
		_w5107_,
		_w7731_,
		_w7906_,
		_w20859_,
		_w21397_
	);
	LUT4 #(
		.INIT('h0200)
	) name17350 (
		\core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w21398_
	);
	LUT2 #(
		.INIT('h1)
	) name17351 (
		_w13546_,
		_w21398_,
		_w21399_
	);
	LUT4 #(
		.INIT('h0200)
	) name17352 (
		\core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w21400_
	);
	LUT4 #(
		.INIT('h0200)
	) name17353 (
		\core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w21401_
	);
	LUT4 #(
		.INIT('h0200)
	) name17354 (
		\core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w21402_
	);
	LUT3 #(
		.INIT('h01)
	) name17355 (
		_w21401_,
		_w21402_,
		_w21400_,
		_w21403_
	);
	LUT2 #(
		.INIT('h8)
	) name17356 (
		_w21399_,
		_w21403_,
		_w21404_
	);
	LUT2 #(
		.INIT('h4)
	) name17357 (
		\core_dag_ilm1reg_I_reg[7]/NET0131 ,
		_w13546_,
		_w21405_
	);
	LUT3 #(
		.INIT('h0b)
	) name17358 (
		_w21397_,
		_w21404_,
		_w21405_,
		_w21406_
	);
	LUT4 #(
		.INIT('h0200)
	) name17359 (
		\core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w21407_
	);
	LUT2 #(
		.INIT('h1)
	) name17360 (
		_w13546_,
		_w21407_,
		_w21408_
	);
	LUT4 #(
		.INIT('h0200)
	) name17361 (
		\core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w21409_
	);
	LUT4 #(
		.INIT('h0200)
	) name17362 (
		\core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w21410_
	);
	LUT4 #(
		.INIT('h0200)
	) name17363 (
		\core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w21411_
	);
	LUT3 #(
		.INIT('h01)
	) name17364 (
		_w21410_,
		_w21411_,
		_w21409_,
		_w21412_
	);
	LUT2 #(
		.INIT('h8)
	) name17365 (
		_w21408_,
		_w21412_,
		_w21413_
	);
	LUT2 #(
		.INIT('h4)
	) name17366 (
		\core_dag_ilm1reg_I_reg[6]/NET0131 ,
		_w13546_,
		_w21414_
	);
	LUT4 #(
		.INIT('h001f)
	) name17367 (
		_w15062_,
		_w20859_,
		_w21413_,
		_w21414_,
		_w21415_
	);
	LUT4 #(
		.INIT('h0200)
	) name17368 (
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w21416_
	);
	LUT2 #(
		.INIT('h1)
	) name17369 (
		_w13546_,
		_w21416_,
		_w21417_
	);
	LUT4 #(
		.INIT('h0200)
	) name17370 (
		\core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w21418_
	);
	LUT4 #(
		.INIT('h0200)
	) name17371 (
		\core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w21419_
	);
	LUT4 #(
		.INIT('h0200)
	) name17372 (
		\core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w21420_
	);
	LUT3 #(
		.INIT('h01)
	) name17373 (
		_w21419_,
		_w21420_,
		_w21418_,
		_w21421_
	);
	LUT2 #(
		.INIT('h8)
	) name17374 (
		_w21417_,
		_w21421_,
		_w21422_
	);
	LUT2 #(
		.INIT('h4)
	) name17375 (
		\core_dag_ilm1reg_I_reg[4]/NET0131 ,
		_w13546_,
		_w21423_
	);
	LUT4 #(
		.INIT('h001f)
	) name17376 (
		_w15068_,
		_w20859_,
		_w21422_,
		_w21423_,
		_w21424_
	);
	LUT4 #(
		.INIT('h0200)
	) name17377 (
		\core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w21425_
	);
	LUT2 #(
		.INIT('h1)
	) name17378 (
		_w13546_,
		_w21425_,
		_w21426_
	);
	LUT4 #(
		.INIT('h0200)
	) name17379 (
		\core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w21427_
	);
	LUT4 #(
		.INIT('h0200)
	) name17380 (
		\core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w21428_
	);
	LUT4 #(
		.INIT('h0200)
	) name17381 (
		\core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w21429_
	);
	LUT3 #(
		.INIT('h01)
	) name17382 (
		_w21428_,
		_w21429_,
		_w21427_,
		_w21430_
	);
	LUT2 #(
		.INIT('h8)
	) name17383 (
		_w21426_,
		_w21430_,
		_w21431_
	);
	LUT2 #(
		.INIT('h4)
	) name17384 (
		\core_dag_ilm1reg_I_reg[3]/NET0131 ,
		_w13546_,
		_w21432_
	);
	LUT4 #(
		.INIT('h002f)
	) name17385 (
		_w14929_,
		_w20859_,
		_w21431_,
		_w21432_,
		_w21433_
	);
	LUT4 #(
		.INIT('h008d)
	) name17386 (
		_w5107_,
		_w6501_,
		_w6555_,
		_w20859_,
		_w21434_
	);
	LUT4 #(
		.INIT('h0200)
	) name17387 (
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w21435_
	);
	LUT2 #(
		.INIT('h1)
	) name17388 (
		_w13546_,
		_w21435_,
		_w21436_
	);
	LUT4 #(
		.INIT('h0200)
	) name17389 (
		\core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w21437_
	);
	LUT4 #(
		.INIT('h0200)
	) name17390 (
		\core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w21438_
	);
	LUT4 #(
		.INIT('h0200)
	) name17391 (
		\core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w21439_
	);
	LUT3 #(
		.INIT('h01)
	) name17392 (
		_w21438_,
		_w21439_,
		_w21437_,
		_w21440_
	);
	LUT2 #(
		.INIT('h8)
	) name17393 (
		_w21436_,
		_w21440_,
		_w21441_
	);
	LUT2 #(
		.INIT('h4)
	) name17394 (
		\core_dag_ilm1reg_I_reg[2]/NET0131 ,
		_w13546_,
		_w21442_
	);
	LUT3 #(
		.INIT('h0b)
	) name17395 (
		_w21434_,
		_w21441_,
		_w21442_,
		_w21443_
	);
	LUT4 #(
		.INIT('h008d)
	) name17396 (
		_w5107_,
		_w5914_,
		_w5771_,
		_w20859_,
		_w21444_
	);
	LUT4 #(
		.INIT('h0200)
	) name17397 (
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w5070_,
		_w5073_,
		_w20363_,
		_w21445_
	);
	LUT2 #(
		.INIT('h1)
	) name17398 (
		_w13546_,
		_w21445_,
		_w21446_
	);
	LUT4 #(
		.INIT('h0200)
	) name17399 (
		\core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 ,
		_w5079_,
		_w5082_,
		_w20364_,
		_w21447_
	);
	LUT4 #(
		.INIT('h0200)
	) name17400 (
		\core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 ,
		_w5087_,
		_w5090_,
		_w20360_,
		_w21448_
	);
	LUT4 #(
		.INIT('h0200)
	) name17401 (
		\core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 ,
		_w5061_,
		_w5065_,
		_w20361_,
		_w21449_
	);
	LUT3 #(
		.INIT('h01)
	) name17402 (
		_w21448_,
		_w21449_,
		_w21447_,
		_w21450_
	);
	LUT2 #(
		.INIT('h8)
	) name17403 (
		_w21446_,
		_w21450_,
		_w21451_
	);
	LUT2 #(
		.INIT('h4)
	) name17404 (
		\core_dag_ilm1reg_I_reg[0]/NET0131 ,
		_w13546_,
		_w21452_
	);
	LUT3 #(
		.INIT('h0b)
	) name17405 (
		_w21444_,
		_w21451_,
		_w21452_,
		_w21453_
	);
	LUT3 #(
		.INIT('h0b)
	) name17406 (
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w17163_,
		_w21454_
	);
	LUT4 #(
		.INIT('h2022)
	) name17407 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w4971_,
		_w17169_,
		_w17170_,
		_w21455_
	);
	LUT3 #(
		.INIT('hce)
	) name17408 (
		\core_c_psq_CNTRval_reg/NET0131 ,
		_w21454_,
		_w21455_,
		_w21456_
	);
	LUT3 #(
		.INIT('h6c)
	) name17409 (
		\sice_IIRC_reg[7]/NET0131 ,
		\sice_IIRC_reg[8]/NET0131 ,
		_w11936_,
		_w21457_
	);
	LUT4 #(
		.INIT('h8200)
	) name17410 (
		T_IMS_pad,
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w21458_
	);
	LUT4 #(
		.INIT('h4000)
	) name17411 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[20]/P0001 ,
		_w21459_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17412 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[22]/P0001 ,
		_w21460_
	);
	LUT3 #(
		.INIT('h01)
	) name17413 (
		_w21459_,
		_w21458_,
		_w21460_,
		_w21461_
	);
	LUT4 #(
		.INIT('h153f)
	) name17414 (
		\sice_DMR2_reg[15]/NET0131 ,
		\sice_IIRC_reg[21]/NET0131 ,
		_w15161_,
		_w15519_,
		_w21462_
	);
	LUT4 #(
		.INIT('h135f)
	) name17415 (
		\sice_CLR_I_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[9]/P0001 ,
		_w14459_,
		_w16507_,
		_w21463_
	);
	LUT4 #(
		.INIT('h0100)
	) name17416 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w21464_
	);
	LUT3 #(
		.INIT('h13)
	) name17417 (
		\sice_IBR1_reg[15]/P0001 ,
		_w15568_,
		_w21464_,
		_w21465_
	);
	LUT4 #(
		.INIT('h153f)
	) name17418 (
		\sice_DBR1_reg[16]/P0001 ,
		\sice_IMR2_reg[15]/NET0131 ,
		_w15527_,
		_w15544_,
		_w21466_
	);
	LUT4 #(
		.INIT('h8000)
	) name17419 (
		_w21465_,
		_w21466_,
		_w21462_,
		_w21463_,
		_w21467_
	);
	LUT4 #(
		.INIT('h0400)
	) name17420 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w21468_
	);
	LUT2 #(
		.INIT('h8)
	) name17421 (
		\sice_IMR1_reg[15]/NET0131 ,
		_w21468_,
		_w21469_
	);
	LUT4 #(
		.INIT('h153f)
	) name17422 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\sice_IBR2_reg[15]/P0001 ,
		_w15559_,
		_w17323_,
		_w21470_
	);
	LUT4 #(
		.INIT('h153f)
	) name17423 (
		\sice_DMR1_reg[15]/NET0131 ,
		\sice_ICYC_reg[21]/NET0131 ,
		_w14695_,
		_w17158_,
		_w21471_
	);
	LUT4 #(
		.INIT('h0020)
	) name17424 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w21472_
	);
	LUT4 #(
		.INIT('h135f)
	) name17425 (
		\sice_DBR2_reg[16]/P0001 ,
		\sice_IRR_reg[11]/P0001 ,
		_w15508_,
		_w21472_,
		_w21473_
	);
	LUT4 #(
		.INIT('h4000)
	) name17426 (
		_w21469_,
		_w21471_,
		_w21473_,
		_w21470_,
		_w21474_
	);
	LUT4 #(
		.INIT('h1333)
	) name17427 (
		_w21458_,
		_w21461_,
		_w21467_,
		_w21474_,
		_w21475_
	);
	LUT2 #(
		.INIT('h1)
	) name17428 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001 ,
		_w17501_,
		_w21476_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17429 (
		_w12220_,
		_w12736_,
		_w12737_,
		_w17505_,
		_w21477_
	);
	LUT4 #(
		.INIT('h1311)
	) name17430 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001 ,
		_w11303_,
		_w11308_,
		_w21478_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17431 (
		_w12224_,
		_w21476_,
		_w21477_,
		_w21478_,
		_w21479_
	);
	LUT2 #(
		.INIT('h2)
	) name17432 (
		_w17500_,
		_w21479_,
		_w21480_
	);
	LUT4 #(
		.INIT('h0057)
	) name17433 (
		_w11624_,
		_w15367_,
		_w15372_,
		_w21480_,
		_w21481_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17434 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w7257_,
		_w7375_,
		_w7377_,
		_w21482_
	);
	LUT4 #(
		.INIT('h0200)
	) name17435 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001 ,
		_w21483_
	);
	LUT4 #(
		.INIT('h4000)
	) name17436 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001 ,
		_w21484_
	);
	LUT4 #(
		.INIT('h2000)
	) name17437 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001 ,
		_w21485_
	);
	LUT4 #(
		.INIT('h1000)
	) name17438 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001 ,
		_w21486_
	);
	LUT4 #(
		.INIT('h0001)
	) name17439 (
		_w21483_,
		_w21484_,
		_w21485_,
		_w21486_,
		_w21487_
	);
	LUT4 #(
		.INIT('h0100)
	) name17440 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001 ,
		_w21488_
	);
	LUT4 #(
		.INIT('h0400)
	) name17441 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001 ,
		_w21489_
	);
	LUT4 #(
		.INIT('h0800)
	) name17442 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001 ,
		_w21490_
	);
	LUT4 #(
		.INIT('h0001)
	) name17443 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w21488_,
		_w21489_,
		_w21490_,
		_w21491_
	);
	LUT4 #(
		.INIT('h2070)
	) name17444 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w21492_
	);
	LUT4 #(
		.INIT('h5540)
	) name17445 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w21487_,
		_w21491_,
		_w21492_,
		_w21493_
	);
	LUT2 #(
		.INIT('h1)
	) name17446 (
		_w21482_,
		_w21493_,
		_w21494_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17447 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w5784_,
		_w5911_,
		_w5913_,
		_w21495_
	);
	LUT4 #(
		.INIT('h4070)
	) name17448 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_dec_IRE_reg[7]/NET0131 ,
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w21496_
	);
	LUT4 #(
		.INIT('h0800)
	) name17449 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001 ,
		_w21497_
	);
	LUT4 #(
		.INIT('h1000)
	) name17450 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001 ,
		_w21498_
	);
	LUT4 #(
		.INIT('h2000)
	) name17451 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001 ,
		_w21499_
	);
	LUT4 #(
		.INIT('h0100)
	) name17452 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001 ,
		_w21500_
	);
	LUT4 #(
		.INIT('h0001)
	) name17453 (
		_w21497_,
		_w21498_,
		_w21499_,
		_w21500_,
		_w21501_
	);
	LUT4 #(
		.INIT('h4000)
	) name17454 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001 ,
		_w21502_
	);
	LUT4 #(
		.INIT('h0200)
	) name17455 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001 ,
		_w21503_
	);
	LUT4 #(
		.INIT('h0400)
	) name17456 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001 ,
		_w21504_
	);
	LUT4 #(
		.INIT('h0001)
	) name17457 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w21502_,
		_w21503_,
		_w21504_,
		_w21505_
	);
	LUT4 #(
		.INIT('h5444)
	) name17458 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w21496_,
		_w21501_,
		_w21505_,
		_w21506_
	);
	LUT2 #(
		.INIT('h1)
	) name17459 (
		_w21495_,
		_w21506_,
		_w21507_
	);
	LUT3 #(
		.INIT('h80)
	) name17460 (
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9079_,
		_w21508_
	);
	LUT4 #(
		.INIT('haa80)
	) name17461 (
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9075_,
		_w20984_,
		_w21509_
	);
	LUT4 #(
		.INIT('h3353)
	) name17462 (
		\bdma_BWdataBUF_h_reg[6]/P0001 ,
		\bdma_BWdataBUF_reg[6]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w20980_,
		_w21510_
	);
	LUT4 #(
		.INIT('h2023)
	) name17463 (
		\bdma_BWdataBUF_h_reg[14]/P0001 ,
		_w21508_,
		_w21509_,
		_w21510_,
		_w21511_
	);
	LUT4 #(
		.INIT('h8000)
	) name17464 (
		\bdma_BWdataBUF_h_reg[22]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9079_,
		_w21512_
	);
	LUT2 #(
		.INIT('he)
	) name17465 (
		_w21511_,
		_w21512_,
		_w21513_
	);
	LUT4 #(
		.INIT('h3353)
	) name17466 (
		\bdma_BWdataBUF_h_reg[5]/P0001 ,
		\bdma_BWdataBUF_reg[5]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w20980_,
		_w21514_
	);
	LUT4 #(
		.INIT('h2023)
	) name17467 (
		\bdma_BWdataBUF_h_reg[13]/P0001 ,
		_w21508_,
		_w21509_,
		_w21514_,
		_w21515_
	);
	LUT4 #(
		.INIT('h8000)
	) name17468 (
		\bdma_BWdataBUF_h_reg[21]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9079_,
		_w21516_
	);
	LUT2 #(
		.INIT('he)
	) name17469 (
		_w21515_,
		_w21516_,
		_w21517_
	);
	LUT4 #(
		.INIT('h3353)
	) name17470 (
		\bdma_BWdataBUF_h_reg[7]/P0001 ,
		\bdma_BWdataBUF_reg[7]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w20980_,
		_w21518_
	);
	LUT4 #(
		.INIT('h2023)
	) name17471 (
		\bdma_BWdataBUF_h_reg[15]/P0001 ,
		_w21508_,
		_w21509_,
		_w21518_,
		_w21519_
	);
	LUT4 #(
		.INIT('h8000)
	) name17472 (
		\bdma_BWdataBUF_h_reg[23]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9079_,
		_w21520_
	);
	LUT2 #(
		.INIT('he)
	) name17473 (
		_w21519_,
		_w21520_,
		_w21521_
	);
	LUT4 #(
		.INIT('h3353)
	) name17474 (
		\bdma_BWdataBUF_h_reg[4]/P0001 ,
		\bdma_BWdataBUF_reg[4]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w20980_,
		_w21522_
	);
	LUT4 #(
		.INIT('h2023)
	) name17475 (
		\bdma_BWdataBUF_h_reg[12]/P0001 ,
		_w21508_,
		_w21509_,
		_w21522_,
		_w21523_
	);
	LUT4 #(
		.INIT('h8000)
	) name17476 (
		\bdma_BWdataBUF_h_reg[20]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9079_,
		_w21524_
	);
	LUT2 #(
		.INIT('he)
	) name17477 (
		_w21523_,
		_w21524_,
		_w21525_
	);
	LUT4 #(
		.INIT('h3353)
	) name17478 (
		\bdma_BWdataBUF_h_reg[3]/P0001 ,
		\bdma_BWdataBUF_reg[3]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w20980_,
		_w21526_
	);
	LUT4 #(
		.INIT('h2023)
	) name17479 (
		\bdma_BWdataBUF_h_reg[11]/P0001 ,
		_w21508_,
		_w21509_,
		_w21526_,
		_w21527_
	);
	LUT4 #(
		.INIT('h8000)
	) name17480 (
		\bdma_BWdataBUF_h_reg[19]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9079_,
		_w21528_
	);
	LUT2 #(
		.INIT('he)
	) name17481 (
		_w21527_,
		_w21528_,
		_w21529_
	);
	LUT4 #(
		.INIT('h3353)
	) name17482 (
		\bdma_BWdataBUF_h_reg[2]/P0001 ,
		\bdma_BWdataBUF_reg[2]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w20980_,
		_w21530_
	);
	LUT4 #(
		.INIT('h2023)
	) name17483 (
		\bdma_BWdataBUF_h_reg[10]/P0001 ,
		_w21508_,
		_w21509_,
		_w21530_,
		_w21531_
	);
	LUT4 #(
		.INIT('h8000)
	) name17484 (
		\bdma_BWdataBUF_h_reg[18]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9079_,
		_w21532_
	);
	LUT2 #(
		.INIT('he)
	) name17485 (
		_w21531_,
		_w21532_,
		_w21533_
	);
	LUT4 #(
		.INIT('h3353)
	) name17486 (
		\bdma_BWdataBUF_h_reg[1]/P0001 ,
		\bdma_BWdataBUF_reg[1]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w20980_,
		_w21534_
	);
	LUT4 #(
		.INIT('h2023)
	) name17487 (
		\bdma_BWdataBUF_h_reg[9]/P0001 ,
		_w21508_,
		_w21509_,
		_w21534_,
		_w21535_
	);
	LUT4 #(
		.INIT('h8000)
	) name17488 (
		\bdma_BWdataBUF_h_reg[17]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9079_,
		_w21536_
	);
	LUT2 #(
		.INIT('he)
	) name17489 (
		_w21535_,
		_w21536_,
		_w21537_
	);
	LUT4 #(
		.INIT('h3353)
	) name17490 (
		\bdma_BWdataBUF_h_reg[0]/P0001 ,
		\bdma_BWdataBUF_reg[0]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w20980_,
		_w21538_
	);
	LUT4 #(
		.INIT('h2023)
	) name17491 (
		\bdma_BWdataBUF_h_reg[8]/P0001 ,
		_w21508_,
		_w21509_,
		_w21538_,
		_w21539_
	);
	LUT4 #(
		.INIT('h8000)
	) name17492 (
		\bdma_BWdataBUF_h_reg[16]/P0001 ,
		\bdma_WRlat_reg/P0001 ,
		_w4884_,
		_w9079_,
		_w21540_
	);
	LUT2 #(
		.INIT('he)
	) name17493 (
		_w21539_,
		_w21540_,
		_w21541_
	);
	LUT4 #(
		.INIT('h4000)
	) name17494 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[11]/P0001 ,
		_w21542_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17495 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[13]/P0001 ,
		_w21543_
	);
	LUT3 #(
		.INIT('h01)
	) name17496 (
		_w21458_,
		_w21542_,
		_w21543_,
		_w21544_
	);
	LUT4 #(
		.INIT('h153f)
	) name17497 (
		\sice_IMR1_reg[6]/NET0131 ,
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w16507_,
		_w21468_,
		_w21545_
	);
	LUT4 #(
		.INIT('h153f)
	) name17498 (
		\sice_DMR1_reg[6]/NET0131 ,
		\sice_IIRC_reg[12]/NET0131 ,
		_w15161_,
		_w17158_,
		_w21546_
	);
	LUT2 #(
		.INIT('h8)
	) name17499 (
		\sice_ITR_reg[2]/NET0131 ,
		_w15568_,
		_w21547_
	);
	LUT4 #(
		.INIT('h153f)
	) name17500 (
		\sice_DBR1_reg[7]/P0001 ,
		\sice_DMR2_reg[6]/NET0131 ,
		_w15519_,
		_w15544_,
		_w21548_
	);
	LUT4 #(
		.INIT('h4000)
	) name17501 (
		_w21547_,
		_w21548_,
		_w21545_,
		_w21546_,
		_w21549_
	);
	LUT4 #(
		.INIT('h0001)
	) name17502 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w21550_
	);
	LUT3 #(
		.INIT('h07)
	) name17503 (
		\sice_ICYC_reg[12]/NET0131 ,
		_w14695_,
		_w21550_,
		_w21551_
	);
	LUT4 #(
		.INIT('h153f)
	) name17504 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		\sice_IBR2_reg[6]/P0001 ,
		_w15559_,
		_w17323_,
		_w21552_
	);
	LUT4 #(
		.INIT('h153f)
	) name17505 (
		\sice_IBR1_reg[6]/P0001 ,
		\sice_IMR2_reg[6]/NET0131 ,
		_w15527_,
		_w21464_,
		_w21553_
	);
	LUT4 #(
		.INIT('h135f)
	) name17506 (
		\sice_DBR2_reg[7]/P0001 ,
		\sice_IRR_reg[2]/P0001 ,
		_w15508_,
		_w21472_,
		_w21554_
	);
	LUT4 #(
		.INIT('h8000)
	) name17507 (
		_w21553_,
		_w21554_,
		_w21551_,
		_w21552_,
		_w21555_
	);
	LUT4 #(
		.INIT('h1333)
	) name17508 (
		_w21458_,
		_w21544_,
		_w21549_,
		_w21555_,
		_w21556_
	);
	LUT4 #(
		.INIT('h4000)
	) name17509 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[10]/P0001 ,
		_w21557_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17510 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[12]/P0001 ,
		_w21558_
	);
	LUT3 #(
		.INIT('h01)
	) name17511 (
		_w21458_,
		_w21557_,
		_w21558_,
		_w21559_
	);
	LUT4 #(
		.INIT('h135f)
	) name17512 (
		\sice_ICYC_reg[11]/NET0131 ,
		\sice_IMR2_reg[5]/NET0131 ,
		_w14695_,
		_w15527_,
		_w21560_
	);
	LUT4 #(
		.INIT('h153f)
	) name17513 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\sice_DBR1_reg[6]/P0001 ,
		_w15544_,
		_w17323_,
		_w21561_
	);
	LUT2 #(
		.INIT('h8)
	) name17514 (
		\sice_ITR_reg[1]/NET0131 ,
		_w15568_,
		_w21562_
	);
	LUT3 #(
		.INIT('h07)
	) name17515 (
		\sice_IBR2_reg[5]/P0001 ,
		_w15559_,
		_w21550_,
		_w21563_
	);
	LUT4 #(
		.INIT('h4000)
	) name17516 (
		_w21562_,
		_w21563_,
		_w21560_,
		_w21561_,
		_w21564_
	);
	LUT4 #(
		.INIT('h153f)
	) name17517 (
		\sice_DBR2_reg[6]/P0001 ,
		\sice_IIRC_reg[11]/NET0131 ,
		_w15161_,
		_w15508_,
		_w21565_
	);
	LUT4 #(
		.INIT('h135f)
	) name17518 (
		\sice_DMR1_reg[5]/NET0131 ,
		\sice_IRR_reg[1]/P0001 ,
		_w17158_,
		_w21472_,
		_w21566_
	);
	LUT4 #(
		.INIT('h135f)
	) name17519 (
		\sice_DMR2_reg[5]/NET0131 ,
		\sice_IMR1_reg[5]/NET0131 ,
		_w15519_,
		_w21468_,
		_w21567_
	);
	LUT4 #(
		.INIT('h153f)
	) name17520 (
		\sice_IBR1_reg[5]/P0001 ,
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w16507_,
		_w21464_,
		_w21568_
	);
	LUT4 #(
		.INIT('h8000)
	) name17521 (
		_w21567_,
		_w21568_,
		_w21565_,
		_w21566_,
		_w21569_
	);
	LUT4 #(
		.INIT('h1333)
	) name17522 (
		_w21458_,
		_w21559_,
		_w21564_,
		_w21569_,
		_w21570_
	);
	LUT4 #(
		.INIT('h4000)
	) name17523 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[9]/P0001 ,
		_w21571_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17524 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[11]/P0001 ,
		_w21572_
	);
	LUT3 #(
		.INIT('h01)
	) name17525 (
		_w21458_,
		_w21571_,
		_w21572_,
		_w21573_
	);
	LUT4 #(
		.INIT('h135f)
	) name17526 (
		\sice_IIRC_reg[10]/NET0131 ,
		\sice_IMR2_reg[4]/NET0131 ,
		_w15161_,
		_w15527_,
		_w21574_
	);
	LUT4 #(
		.INIT('h153f)
	) name17527 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\sice_DBR1_reg[5]/P0001 ,
		_w15544_,
		_w17323_,
		_w21575_
	);
	LUT2 #(
		.INIT('h8)
	) name17528 (
		\sice_ITR_reg[0]/NET0131 ,
		_w15568_,
		_w21576_
	);
	LUT3 #(
		.INIT('h07)
	) name17529 (
		\sice_IBR2_reg[4]/P0001 ,
		_w15559_,
		_w21550_,
		_w21577_
	);
	LUT4 #(
		.INIT('h4000)
	) name17530 (
		_w21576_,
		_w21577_,
		_w21574_,
		_w21575_,
		_w21578_
	);
	LUT4 #(
		.INIT('h135f)
	) name17531 (
		\sice_DBR2_reg[5]/P0001 ,
		\sice_DMR2_reg[4]/NET0131 ,
		_w15508_,
		_w15519_,
		_w21579_
	);
	LUT4 #(
		.INIT('h135f)
	) name17532 (
		\sice_DMR1_reg[4]/NET0131 ,
		\sice_IRR_reg[0]/P0001 ,
		_w17158_,
		_w21472_,
		_w21580_
	);
	LUT4 #(
		.INIT('h135f)
	) name17533 (
		\sice_ICYC_reg[10]/NET0131 ,
		\sice_IMR1_reg[4]/NET0131 ,
		_w14695_,
		_w21468_,
		_w21581_
	);
	LUT4 #(
		.INIT('h153f)
	) name17534 (
		\sice_IBR1_reg[4]/P0001 ,
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w16507_,
		_w21464_,
		_w21582_
	);
	LUT4 #(
		.INIT('h8000)
	) name17535 (
		_w21581_,
		_w21582_,
		_w21579_,
		_w21580_,
		_w21583_
	);
	LUT4 #(
		.INIT('h1333)
	) name17536 (
		_w21458_,
		_w21573_,
		_w21578_,
		_w21583_,
		_w21584_
	);
	LUT3 #(
		.INIT('h6c)
	) name17537 (
		\sice_ICYC_reg[7]/NET0131 ,
		\sice_ICYC_reg[8]/NET0131 ,
		_w11932_,
		_w21585_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17538 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		_w14698_,
		_w21586_
	);
	LUT2 #(
		.INIT('h1)
	) name17539 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001 ,
		_w17501_,
		_w21587_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17540 (
		_w12220_,
		_w12626_,
		_w12627_,
		_w17505_,
		_w21588_
	);
	LUT4 #(
		.INIT('h1311)
	) name17541 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001 ,
		_w11303_,
		_w11308_,
		_w21589_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17542 (
		_w12224_,
		_w21587_,
		_w21588_,
		_w21589_,
		_w21590_
	);
	LUT2 #(
		.INIT('h2)
	) name17543 (
		_w17500_,
		_w21590_,
		_w21591_
	);
	LUT3 #(
		.INIT('h07)
	) name17544 (
		_w11624_,
		_w15554_,
		_w21591_,
		_w21592_
	);
	LUT2 #(
		.INIT('h1)
	) name17545 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 ,
		_w17501_,
		_w21593_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17546 (
		_w12220_,
		_w12315_,
		_w12316_,
		_w17505_,
		_w21594_
	);
	LUT4 #(
		.INIT('h1311)
	) name17547 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 ,
		_w11303_,
		_w11308_,
		_w21595_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17548 (
		_w12224_,
		_w21593_,
		_w21594_,
		_w21595_,
		_w21596_
	);
	LUT2 #(
		.INIT('h2)
	) name17549 (
		_w17500_,
		_w21596_,
		_w21597_
	);
	LUT4 #(
		.INIT('h0057)
	) name17550 (
		_w11624_,
		_w15570_,
		_w15571_,
		_w21597_,
		_w21598_
	);
	LUT4 #(
		.INIT('h8000)
	) name17551 (
		_w5344_,
		_w5346_,
		_w5348_,
		_w5374_,
		_w21599_
	);
	LUT4 #(
		.INIT('haaa8)
	) name17552 (
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w5434_,
		_w6210_,
		_w21599_,
		_w21600_
	);
	LUT3 #(
		.INIT('h40)
	) name17553 (
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w5127_,
		_w5148_,
		_w21601_
	);
	LUT4 #(
		.INIT('h5501)
	) name17554 (
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w5767_,
		_w5918_,
		_w21601_,
		_w21602_
	);
	LUT3 #(
		.INIT('h02)
	) name17555 (
		\auctl_T0Sack_reg/NET0131 ,
		_w21600_,
		_w21602_,
		_w21603_
	);
	LUT3 #(
		.INIT('h02)
	) name17556 (
		\auctl_R0Sack_reg/NET0131 ,
		_w21600_,
		_w21602_,
		_w21604_
	);
	LUT3 #(
		.INIT('h02)
	) name17557 (
		\auctl_T1Sack_reg/NET0131 ,
		_w21600_,
		_w21602_,
		_w21605_
	);
	LUT3 #(
		.INIT('h02)
	) name17558 (
		\auctl_R1Sack_reg/NET0131 ,
		_w21600_,
		_w21602_,
		_w21606_
	);
	LUT4 #(
		.INIT('h2000)
	) name17559 (
		\core_c_dec_MTIreg_E_reg[4]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21607_
	);
	LUT4 #(
		.INIT('h5053)
	) name17560 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[18]/NET0131 ,
		_w19034_,
		_w19124_,
		_w21608_
	);
	LUT2 #(
		.INIT('h8)
	) name17561 (
		_w19709_,
		_w21608_,
		_w21609_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17562 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19705_,
		_w21610_
	);
	LUT4 #(
		.INIT('h4000)
	) name17563 (
		_w19701_,
		_w19729_,
		_w21609_,
		_w21610_,
		_w21611_
	);
	LUT3 #(
		.INIT('ha8)
	) name17564 (
		_w4102_,
		_w21607_,
		_w21611_,
		_w21612_
	);
	LUT3 #(
		.INIT('h01)
	) name17565 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		\core_c_dec_IRE_reg[1]/NET0131 ,
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w21613_
	);
	LUT2 #(
		.INIT('h2)
	) name17566 (
		\clkc_SIDLE_s1_reg/NET0131 ,
		\clkc_SIDLE_s2_reg/NET0131 ,
		_w21614_
	);
	LUT3 #(
		.INIT('h45)
	) name17567 (
		\clkc_SlowDn_reg/NET0131 ,
		_w21613_,
		_w21614_,
		_w21615_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name17568 (
		\clkc_STBY_reg/NET0131 ,
		_w14453_,
		_w21613_,
		_w21614_,
		_w21616_
	);
	LUT2 #(
		.INIT('h4)
	) name17569 (
		_w21615_,
		_w21616_,
		_w21617_
	);
	LUT3 #(
		.INIT('h80)
	) name17570 (
		_w20441_,
		_w20450_,
		_w21617_,
		_w21618_
	);
	LUT4 #(
		.INIT('h152a)
	) name17571 (
		\clkc_STDcnt_reg[7]/NET0131 ,
		_w19400_,
		_w19405_,
		_w19393_,
		_w21619_
	);
	LUT4 #(
		.INIT('h2000)
	) name17572 (
		\core_c_dec_MTIreg_E_reg[7]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21620_
	);
	LUT4 #(
		.INIT('h4000)
	) name17573 (
		_w19701_,
		_w21237_,
		_w21238_,
		_w21609_,
		_w21621_
	);
	LUT3 #(
		.INIT('ha8)
	) name17574 (
		_w4102_,
		_w21620_,
		_w21621_,
		_w21622_
	);
	LUT4 #(
		.INIT('h2000)
	) name17575 (
		\core_c_dec_MTDMOVL_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21623_
	);
	LUT4 #(
		.INIT('haa80)
	) name17576 (
		_w4102_,
		_w19734_,
		_w21238_,
		_w21623_,
		_w21624_
	);
	LUT3 #(
		.INIT('h15)
	) name17577 (
		_w4104_,
		_w19730_,
		_w19731_,
		_w21625_
	);
	LUT4 #(
		.INIT('h1000)
	) name17578 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21626_
	);
	LUT2 #(
		.INIT('h2)
	) name17579 (
		_w4102_,
		_w21626_,
		_w21627_
	);
	LUT2 #(
		.INIT('h4)
	) name17580 (
		_w21625_,
		_w21627_,
		_w21628_
	);
	LUT4 #(
		.INIT('h2000)
	) name17581 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21629_
	);
	LUT2 #(
		.INIT('h8)
	) name17582 (
		_w19702_,
		_w21610_,
		_w21630_
	);
	LUT2 #(
		.INIT('h8)
	) name17583 (
		_w19709_,
		_w19716_,
		_w21631_
	);
	LUT4 #(
		.INIT('h070f)
	) name17584 (
		_w19702_,
		_w21610_,
		_w21629_,
		_w21631_,
		_w21632_
	);
	LUT2 #(
		.INIT('h2)
	) name17585 (
		_w4102_,
		_w21632_,
		_w21633_
	);
	LUT4 #(
		.INIT('h2000)
	) name17586 (
		\core_c_dec_MTRX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21634_
	);
	LUT4 #(
		.INIT('h4000)
	) name17587 (
		_w19701_,
		_w19732_,
		_w21237_,
		_w21610_,
		_w21635_
	);
	LUT3 #(
		.INIT('ha8)
	) name17588 (
		_w4102_,
		_w21634_,
		_w21635_,
		_w21636_
	);
	LUT4 #(
		.INIT('h2000)
	) name17589 (
		\core_c_dec_MTRX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21637_
	);
	LUT4 #(
		.INIT('h4000)
	) name17590 (
		_w19701_,
		_w19729_,
		_w19732_,
		_w21610_,
		_w21638_
	);
	LUT3 #(
		.INIT('ha8)
	) name17591 (
		_w4102_,
		_w21637_,
		_w21638_,
		_w21639_
	);
	LUT4 #(
		.INIT('h2000)
	) name17592 (
		\core_c_dec_MTPMOVL_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21640_
	);
	LUT4 #(
		.INIT('haa80)
	) name17593 (
		_w4102_,
		_w19734_,
		_w21610_,
		_w21640_,
		_w21641_
	);
	LUT4 #(
		.INIT('h2000)
	) name17594 (
		\core_c_dec_MTOWRCNTR_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21642_
	);
	LUT4 #(
		.INIT('h000e)
	) name17595 (
		_w19710_,
		_w19711_,
		_w19713_,
		_w19714_,
		_w21643_
	);
	LUT4 #(
		.INIT('h1000)
	) name17596 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4428_,
		_w8172_,
		_w21643_,
		_w21644_
	);
	LUT2 #(
		.INIT('h8)
	) name17597 (
		_w19702_,
		_w21238_,
		_w21645_
	);
	LUT4 #(
		.INIT('h2333)
	) name17598 (
		_w19709_,
		_w21642_,
		_w21644_,
		_w21645_,
		_w21646_
	);
	LUT2 #(
		.INIT('h2)
	) name17599 (
		_w4102_,
		_w21646_,
		_w21647_
	);
	LUT4 #(
		.INIT('h2000)
	) name17600 (
		\core_c_dec_MTMreg_E_reg[7]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21648_
	);
	LUT4 #(
		.INIT('h2000)
	) name17601 (
		_w19716_,
		_w19701_,
		_w21238_,
		_w21609_,
		_w21649_
	);
	LUT3 #(
		.INIT('ha8)
	) name17602 (
		_w4102_,
		_w21648_,
		_w21649_,
		_w21650_
	);
	LUT4 #(
		.INIT('h2000)
	) name17603 (
		\core_c_dec_MTMreg_E_reg[6]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21651_
	);
	LUT4 #(
		.INIT('h2000)
	) name17604 (
		_w19716_,
		_w19701_,
		_w21609_,
		_w21610_,
		_w21652_
	);
	LUT3 #(
		.INIT('ha8)
	) name17605 (
		_w4102_,
		_w21651_,
		_w21652_,
		_w21653_
	);
	LUT4 #(
		.INIT('h2000)
	) name17606 (
		\core_c_dec_MTMreg_E_reg[5]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21654_
	);
	LUT4 #(
		.INIT('h4000)
	) name17607 (
		_w19701_,
		_w21238_,
		_w21609_,
		_w21643_,
		_w21655_
	);
	LUT3 #(
		.INIT('ha8)
	) name17608 (
		_w4102_,
		_w21654_,
		_w21655_,
		_w21656_
	);
	LUT4 #(
		.INIT('h2000)
	) name17609 (
		\core_c_dec_MTMreg_E_reg[4]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21657_
	);
	LUT4 #(
		.INIT('h4000)
	) name17610 (
		_w19701_,
		_w21609_,
		_w21610_,
		_w21643_,
		_w21658_
	);
	LUT3 #(
		.INIT('ha8)
	) name17611 (
		_w4102_,
		_w21657_,
		_w21658_,
		_w21659_
	);
	LUT4 #(
		.INIT('heee0)
	) name17612 (
		_w19713_,
		_w19714_,
		_w19703_,
		_w19704_,
		_w21660_
	);
	LUT4 #(
		.INIT('h2000)
	) name17613 (
		\core_c_dec_MTMreg_E_reg[3]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21661_
	);
	LUT4 #(
		.INIT('h007f)
	) name17614 (
		_w21246_,
		_w21249_,
		_w21660_,
		_w21661_,
		_w21662_
	);
	LUT2 #(
		.INIT('h2)
	) name17615 (
		_w4102_,
		_w21662_,
		_w21663_
	);
	LUT4 #(
		.INIT('h000e)
	) name17616 (
		_w19713_,
		_w19714_,
		_w19703_,
		_w19704_,
		_w21664_
	);
	LUT4 #(
		.INIT('h2000)
	) name17617 (
		\core_c_dec_MTMreg_E_reg[2]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21665_
	);
	LUT4 #(
		.INIT('h007f)
	) name17618 (
		_w21246_,
		_w21249_,
		_w21664_,
		_w21665_,
		_w21666_
	);
	LUT2 #(
		.INIT('h2)
	) name17619 (
		_w4102_,
		_w21666_,
		_w21667_
	);
	LUT4 #(
		.INIT('h2000)
	) name17620 (
		\core_c_dec_MTMreg_E_reg[0]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21668_
	);
	LUT2 #(
		.INIT('h8)
	) name17621 (
		_w19705_,
		_w21643_,
		_w21669_
	);
	LUT4 #(
		.INIT('h070f)
	) name17622 (
		_w21245_,
		_w21249_,
		_w21668_,
		_w21669_,
		_w21670_
	);
	LUT2 #(
		.INIT('h2)
	) name17623 (
		_w4102_,
		_w21670_,
		_w21671_
	);
	LUT2 #(
		.INIT('h4)
	) name17624 (
		_w19709_,
		_w21608_,
		_w21672_
	);
	LUT4 #(
		.INIT('h4000)
	) name17625 (
		_w19701_,
		_w21237_,
		_w21238_,
		_w21672_,
		_w21673_
	);
	LUT4 #(
		.INIT('h2000)
	) name17626 (
		\core_c_dec_MTLreg_E_reg[7]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21674_
	);
	LUT3 #(
		.INIT('ha8)
	) name17627 (
		_w4102_,
		_w21673_,
		_w21674_,
		_w21675_
	);
	LUT4 #(
		.INIT('h4000)
	) name17628 (
		_w19701_,
		_w21237_,
		_w21610_,
		_w21672_,
		_w21676_
	);
	LUT4 #(
		.INIT('h2000)
	) name17629 (
		\core_c_dec_MTLreg_E_reg[6]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21677_
	);
	LUT3 #(
		.INIT('ha8)
	) name17630 (
		_w4102_,
		_w21676_,
		_w21677_,
		_w21678_
	);
	LUT4 #(
		.INIT('h4000)
	) name17631 (
		_w19701_,
		_w19729_,
		_w21238_,
		_w21672_,
		_w21679_
	);
	LUT4 #(
		.INIT('h2000)
	) name17632 (
		\core_c_dec_MTLreg_E_reg[5]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21680_
	);
	LUT3 #(
		.INIT('ha8)
	) name17633 (
		_w4102_,
		_w21679_,
		_w21680_,
		_w21681_
	);
	LUT4 #(
		.INIT('h2000)
	) name17634 (
		\core_c_dec_MTLreg_E_reg[4]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21682_
	);
	LUT4 #(
		.INIT('h4000)
	) name17635 (
		_w19701_,
		_w19729_,
		_w21610_,
		_w21672_,
		_w21683_
	);
	LUT3 #(
		.INIT('ha8)
	) name17636 (
		_w4102_,
		_w21682_,
		_w21683_,
		_w21684_
	);
	LUT4 #(
		.INIT('h2000)
	) name17637 (
		\core_c_dec_MTLreg_E_reg[3]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21685_
	);
	LUT4 #(
		.INIT('h4000)
	) name17638 (
		_w4104_,
		_w19712_,
		_w19733_,
		_w21660_,
		_w21686_
	);
	LUT3 #(
		.INIT('ha8)
	) name17639 (
		_w4102_,
		_w21685_,
		_w21686_,
		_w21687_
	);
	LUT4 #(
		.INIT('h2000)
	) name17640 (
		\core_c_dec_MTLreg_E_reg[2]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21688_
	);
	LUT4 #(
		.INIT('h4000)
	) name17641 (
		_w4104_,
		_w19712_,
		_w19733_,
		_w21664_,
		_w21689_
	);
	LUT3 #(
		.INIT('ha8)
	) name17642 (
		_w4102_,
		_w21688_,
		_w21689_,
		_w21690_
	);
	LUT4 #(
		.INIT('h2000)
	) name17643 (
		\core_c_dec_MTLreg_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21691_
	);
	LUT4 #(
		.INIT('h4000)
	) name17644 (
		_w4104_,
		_w19712_,
		_w19733_,
		_w21247_,
		_w21692_
	);
	LUT3 #(
		.INIT('ha8)
	) name17645 (
		_w4102_,
		_w21691_,
		_w21692_,
		_w21693_
	);
	LUT4 #(
		.INIT('h4777)
	) name17646 (
		\core_c_dec_MTLreg_E_reg[0]/P0001 ,
		_w4104_,
		_w19730_,
		_w19733_,
		_w21694_
	);
	LUT2 #(
		.INIT('h2)
	) name17647 (
		_w4102_,
		_w21694_,
		_w21695_
	);
	LUT4 #(
		.INIT('h2000)
	) name17648 (
		\core_c_dec_MTIreg_E_reg[6]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21696_
	);
	LUT4 #(
		.INIT('h4000)
	) name17649 (
		_w19701_,
		_w21237_,
		_w21609_,
		_w21610_,
		_w21697_
	);
	LUT3 #(
		.INIT('ha8)
	) name17650 (
		_w4102_,
		_w21696_,
		_w21697_,
		_w21698_
	);
	LUT4 #(
		.INIT('h2000)
	) name17651 (
		\core_c_dec_MTIreg_E_reg[5]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21699_
	);
	LUT4 #(
		.INIT('h4000)
	) name17652 (
		_w19701_,
		_w19729_,
		_w21238_,
		_w21609_,
		_w21700_
	);
	LUT3 #(
		.INIT('ha8)
	) name17653 (
		_w4102_,
		_w21699_,
		_w21700_,
		_w21701_
	);
	LUT2 #(
		.INIT('h8)
	) name17654 (
		_w19712_,
		_w21245_,
		_w21702_
	);
	LUT4 #(
		.INIT('h2000)
	) name17655 (
		\core_c_dec_MTIreg_E_reg[3]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21703_
	);
	LUT4 #(
		.INIT('h007f)
	) name17656 (
		_w21249_,
		_w21660_,
		_w21702_,
		_w21703_,
		_w21704_
	);
	LUT2 #(
		.INIT('h2)
	) name17657 (
		_w4102_,
		_w21704_,
		_w21705_
	);
	LUT4 #(
		.INIT('h2000)
	) name17658 (
		\core_c_dec_MTIreg_E_reg[2]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21706_
	);
	LUT4 #(
		.INIT('h007f)
	) name17659 (
		_w21249_,
		_w21664_,
		_w21702_,
		_w21706_,
		_w21707_
	);
	LUT2 #(
		.INIT('h2)
	) name17660 (
		_w4102_,
		_w21707_,
		_w21708_
	);
	LUT4 #(
		.INIT('h2000)
	) name17661 (
		\core_c_dec_MTIreg_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21709_
	);
	LUT4 #(
		.INIT('h007f)
	) name17662 (
		_w21247_,
		_w21249_,
		_w21702_,
		_w21709_,
		_w21710_
	);
	LUT2 #(
		.INIT('h2)
	) name17663 (
		_w4102_,
		_w21710_,
		_w21711_
	);
	LUT3 #(
		.INIT('h13)
	) name17664 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001 ,
		_w11300_,
		_w21712_
	);
	LUT4 #(
		.INIT('hccc8)
	) name17665 (
		_w11310_,
		_w11312_,
		_w12626_,
		_w12627_,
		_w21713_
	);
	LUT4 #(
		.INIT('h2322)
	) name17666 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001 ,
		_w11303_,
		_w11308_,
		_w21714_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17667 (
		_w11320_,
		_w21712_,
		_w21713_,
		_w21714_,
		_w21715_
	);
	LUT2 #(
		.INIT('h2)
	) name17668 (
		_w11325_,
		_w21715_,
		_w21716_
	);
	LUT3 #(
		.INIT('h07)
	) name17669 (
		_w9946_,
		_w15554_,
		_w21716_,
		_w21717_
	);
	LUT4 #(
		.INIT('h2000)
	) name17670 (
		\core_c_dec_MTIreg_E_reg[0]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21718_
	);
	LUT4 #(
		.INIT('h007f)
	) name17671 (
		_w19730_,
		_w21245_,
		_w21249_,
		_w21718_,
		_w21719_
	);
	LUT2 #(
		.INIT('h2)
	) name17672 (
		_w4102_,
		_w21719_,
		_w21720_
	);
	LUT4 #(
		.INIT('h2000)
	) name17673 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21721_
	);
	LUT4 #(
		.INIT('h00bf)
	) name17674 (
		_w19709_,
		_w21630_,
		_w21644_,
		_w21721_,
		_w21722_
	);
	LUT2 #(
		.INIT('h2)
	) name17675 (
		_w4102_,
		_w21722_,
		_w21723_
	);
	LUT4 #(
		.INIT('h4777)
	) name17676 (
		\core_c_dec_MTIDR_E_reg/P0001 ,
		_w4104_,
		_w19733_,
		_w21669_,
		_w21724_
	);
	LUT2 #(
		.INIT('h2)
	) name17677 (
		_w4102_,
		_w21724_,
		_w21725_
	);
	LUT4 #(
		.INIT('h2000)
	) name17678 (
		\core_c_dec_MTICNTL_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21726_
	);
	LUT4 #(
		.INIT('h007f)
	) name17679 (
		_w19709_,
		_w21630_,
		_w21644_,
		_w21726_,
		_w21727_
	);
	LUT2 #(
		.INIT('h2)
	) name17680 (
		_w4102_,
		_w21727_,
		_w21728_
	);
	LUT4 #(
		.INIT('h2000)
	) name17681 (
		\core_c_dec_MTCNTR_Eg_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21729_
	);
	LUT4 #(
		.INIT('h007f)
	) name17682 (
		_w19709_,
		_w21644_,
		_w21645_,
		_w21729_,
		_w21730_
	);
	LUT2 #(
		.INIT('h2)
	) name17683 (
		_w4102_,
		_w21730_,
		_w21731_
	);
	LUT4 #(
		.INIT('hba00)
	) name17684 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w9432_,
		_w21732_
	);
	LUT4 #(
		.INIT('h00de)
	) name17685 (
		\bdma_BWCOUNT_reg[1]/NET0131 ,
		_w9432_,
		_w9426_,
		_w21732_,
		_w21733_
	);
	LUT4 #(
		.INIT('h333b)
	) name17686 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		_w9422_,
		_w9414_,
		_w9415_,
		_w21734_
	);
	LUT3 #(
		.INIT('h8c)
	) name17687 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w4142_,
		_w12114_,
		_w21735_
	);
	LUT4 #(
		.INIT('hef00)
	) name17688 (
		_w12114_,
		_w12164_,
		_w12177_,
		_w21735_,
		_w21736_
	);
	LUT2 #(
		.INIT('h2)
	) name17689 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w12486_,
		_w21737_
	);
	LUT4 #(
		.INIT('h4000)
	) name17690 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11837_,
		_w18362_,
		_w18368_,
		_w21738_
	);
	LUT4 #(
		.INIT('h222e)
	) name17691 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001 ,
		_w11830_,
		_w21737_,
		_w21738_,
		_w21739_
	);
	LUT4 #(
		.INIT('h222e)
	) name17692 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001 ,
		_w11329_,
		_w21737_,
		_w21738_,
		_w21740_
	);
	LUT2 #(
		.INIT('h2)
	) name17693 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w14918_,
		_w21741_
	);
	LUT4 #(
		.INIT('h4000)
	) name17694 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w18113_,
		_w18684_,
		_w18692_,
		_w21742_
	);
	LUT4 #(
		.INIT('h222e)
	) name17695 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001 ,
		_w11946_,
		_w21741_,
		_w21742_,
		_w21743_
	);
	LUT4 #(
		.INIT('h222e)
	) name17696 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001 ,
		_w12048_,
		_w21741_,
		_w21742_,
		_w21744_
	);
	LUT3 #(
		.INIT('h13)
	) name17697 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001 ,
		_w11300_,
		_w21745_
	);
	LUT4 #(
		.INIT('hccc8)
	) name17698 (
		_w11310_,
		_w11312_,
		_w12736_,
		_w12737_,
		_w21746_
	);
	LUT4 #(
		.INIT('h2322)
	) name17699 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001 ,
		_w11303_,
		_w11308_,
		_w21747_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17700 (
		_w11320_,
		_w21745_,
		_w21746_,
		_w21747_,
		_w21748_
	);
	LUT2 #(
		.INIT('h2)
	) name17701 (
		_w11325_,
		_w21748_,
		_w21749_
	);
	LUT4 #(
		.INIT('h0057)
	) name17702 (
		_w9946_,
		_w15367_,
		_w15372_,
		_w21749_,
		_w21750_
	);
	LUT3 #(
		.INIT('h13)
	) name17703 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001 ,
		_w9894_,
		_w21751_
	);
	LUT4 #(
		.INIT('h0002)
	) name17704 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w21751_,
		_w21752_
	);
	LUT4 #(
		.INIT('h313b)
	) name17705 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001 ,
		_w11631_,
		_w11635_,
		_w21753_
	);
	LUT4 #(
		.INIT('h2f00)
	) name17706 (
		_w11625_,
		_w14918_,
		_w21752_,
		_w21753_,
		_w21754_
	);
	LUT2 #(
		.INIT('h1)
	) name17707 (
		_w11624_,
		_w21754_,
		_w21755_
	);
	LUT4 #(
		.INIT('hc840)
	) name17708 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11624_,
		_w12351_,
		_w12349_,
		_w21756_
	);
	LUT2 #(
		.INIT('he)
	) name17709 (
		_w21755_,
		_w21756_,
		_w21757_
	);
	LUT4 #(
		.INIT('h048c)
	) name17710 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w12351_,
		_w12349_,
		_w21758_
	);
	LUT2 #(
		.INIT('h2)
	) name17711 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001 ,
		_w11656_,
		_w21759_
	);
	LUT3 #(
		.INIT('h01)
	) name17712 (
		_w9946_,
		_w11659_,
		_w21759_,
		_w21760_
	);
	LUT3 #(
		.INIT('h70)
	) name17713 (
		_w11655_,
		_w14918_,
		_w21760_,
		_w21761_
	);
	LUT2 #(
		.INIT('h1)
	) name17714 (
		_w21758_,
		_w21761_,
		_w21762_
	);
	LUT2 #(
		.INIT('h2)
	) name17715 (
		\bdma_BWRn_reg/NET0131 ,
		\bdma_WRlat_reg/P0001 ,
		_w21763_
	);
	LUT4 #(
		.INIT('he000)
	) name17716 (
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		\bdma_BCTL_reg[6]/NET0131 ,
		\bdma_BCTL_reg[7]/NET0131 ,
		_w21764_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name17717 (
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		\bdma_BCTL_reg[6]/NET0131 ,
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w21765_
	);
	LUT3 #(
		.INIT('h90)
	) name17718 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w21764_,
		_w21765_,
		_w21766_
	);
	LUT4 #(
		.INIT('h001f)
	) name17719 (
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		\bdma_BCTL_reg[6]/NET0131 ,
		\bdma_BCTL_reg[7]/NET0131 ,
		_w21767_
	);
	LUT2 #(
		.INIT('h1)
	) name17720 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w21767_,
		_w21768_
	);
	LUT2 #(
		.INIT('h6)
	) name17721 (
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		_w21769_
	);
	LUT3 #(
		.INIT('h28)
	) name17722 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BWcnt_reg[0]/NET0131 ,
		_w21770_
	);
	LUT3 #(
		.INIT('h60)
	) name17723 (
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w21769_,
		_w21770_,
		_w21771_
	);
	LUT4 #(
		.INIT('h9000)
	) name17724 (
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w21768_,
		_w21771_,
		_w21766_,
		_w21772_
	);
	LUT2 #(
		.INIT('he)
	) name17725 (
		_w21763_,
		_w21772_,
		_w21773_
	);
	LUT4 #(
		.INIT('haa8a)
	) name17726 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w21774_
	);
	LUT4 #(
		.INIT('h00ba)
	) name17727 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w19092_,
		_w21774_,
		_w21775_
	);
	LUT4 #(
		.INIT('h00ea)
	) name17728 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w19091_,
		_w19096_,
		_w21775_,
		_w21776_
	);
	LUT4 #(
		.INIT('h1500)
	) name17729 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w19091_,
		_w19096_,
		_w21775_,
		_w21777_
	);
	LUT3 #(
		.INIT('h02)
	) name17730 (
		_w13155_,
		_w21777_,
		_w21776_,
		_w21778_
	);
	LUT3 #(
		.INIT('h40)
	) name17731 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[11]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w21779_
	);
	LUT2 #(
		.INIT('h1)
	) name17732 (
		_w13158_,
		_w21779_,
		_w21780_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17733 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w6263_,
		_w6362_,
		_w21780_,
		_w21781_
	);
	LUT4 #(
		.INIT('hafac)
	) name17734 (
		\sport0_rxctl_RXSHT_reg[11]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w21782_
	);
	LUT4 #(
		.INIT('h0002)
	) name17735 (
		\sport0_rxctl_RX_reg[11]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w21783_
	);
	LUT4 #(
		.INIT('hffb0)
	) name17736 (
		_w21778_,
		_w21781_,
		_w21782_,
		_w21783_,
		_w21784_
	);
	LUT3 #(
		.INIT('h45)
	) name17737 (
		IACKn_pad,
		\idma_WRCMD_d1_reg/P0001 ,
		\idma_WRCMD_reg/P0001 ,
		_w21785_
	);
	LUT2 #(
		.INIT('h4)
	) name17738 (
		_w13074_,
		_w21785_,
		_w21786_
	);
	LUT3 #(
		.INIT('h01)
	) name17739 (
		_w12821_,
		_w19997_,
		_w21786_,
		_w21787_
	);
	LUT4 #(
		.INIT('h00bf)
	) name17740 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w15506_,
		_w21788_
	);
	LUT3 #(
		.INIT('hca)
	) name17741 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		_w20243_,
		_w21788_,
		_w21789_
	);
	LUT4 #(
		.INIT('h03aa)
	) name17742 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		_w20167_,
		_w20174_,
		_w21788_,
		_w21790_
	);
	LUT4 #(
		.INIT('h03aa)
	) name17743 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		_w20222_,
		_w20229_,
		_w21788_,
		_w21791_
	);
	LUT4 #(
		.INIT('h03aa)
	) name17744 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		_w20155_,
		_w20162_,
		_w21788_,
		_w21792_
	);
	LUT4 #(
		.INIT('h03aa)
	) name17745 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		_w20209_,
		_w20216_,
		_w21788_,
		_w21793_
	);
	LUT3 #(
		.INIT('h0e)
	) name17746 (
		_w7062_,
		_w7067_,
		_w19745_,
		_w21794_
	);
	LUT4 #(
		.INIT('h4f00)
	) name17747 (
		_w7122_,
		_w7126_,
		_w19745_,
		_w19748_,
		_w21795_
	);
	LUT2 #(
		.INIT('h4)
	) name17748 (
		_w21794_,
		_w21795_,
		_w21796_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name17749 (
		_w5041_,
		_w5049_,
		_w7110_,
		_w7096_,
		_w21797_
	);
	LUT3 #(
		.INIT('he0)
	) name17750 (
		_w19746_,
		_w19747_,
		_w21797_,
		_w21798_
	);
	LUT4 #(
		.INIT('hf400)
	) name17751 (
		_w7083_,
		_w7086_,
		_w19745_,
		_w21798_,
		_w21799_
	);
	LUT4 #(
		.INIT('h0203)
	) name17752 (
		_w5041_,
		_w5108_,
		_w7108_,
		_w19744_,
		_w21800_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name17753 (
		_w5041_,
		_w5108_,
		_w7077_,
		_w19744_,
		_w21801_
	);
	LUT4 #(
		.INIT('h000e)
	) name17754 (
		_w19746_,
		_w19747_,
		_w21801_,
		_w21800_,
		_w21802_
	);
	LUT4 #(
		.INIT('h4500)
	) name17755 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w19745_,
		_w21803_
	);
	LUT3 #(
		.INIT('h01)
	) name17756 (
		_w7140_,
		_w7240_,
		_w19745_,
		_w21804_
	);
	LUT4 #(
		.INIT('h3331)
	) name17757 (
		_w19748_,
		_w21802_,
		_w21804_,
		_w21803_,
		_w21805_
	);
	LUT2 #(
		.INIT('h2)
	) name17758 (
		_w19757_,
		_w21805_,
		_w21806_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17759 (
		_w19757_,
		_w21796_,
		_w21799_,
		_w21806_,
		_w21807_
	);
	LUT3 #(
		.INIT('he2)
	) name17760 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w21788_,
		_w21807_,
		_w21808_
	);
	LUT3 #(
		.INIT('hb0)
	) name17761 (
		_w6204_,
		_w6207_,
		_w19745_,
		_w21809_
	);
	LUT4 #(
		.INIT('hf400)
	) name17762 (
		_w5920_,
		_w5924_,
		_w19745_,
		_w19748_,
		_w21810_
	);
	LUT2 #(
		.INIT('h4)
	) name17763 (
		_w21809_,
		_w21810_,
		_w21811_
	);
	LUT4 #(
		.INIT('h00fd)
	) name17764 (
		_w5041_,
		_w5049_,
		_w7034_,
		_w7050_,
		_w21812_
	);
	LUT3 #(
		.INIT('he0)
	) name17765 (
		_w19746_,
		_w19747_,
		_w21812_,
		_w21813_
	);
	LUT4 #(
		.INIT('hf400)
	) name17766 (
		_w7044_,
		_w7048_,
		_w19745_,
		_w21813_,
		_w21814_
	);
	LUT4 #(
		.INIT('h0203)
	) name17767 (
		_w5041_,
		_w5108_,
		_w6237_,
		_w19744_,
		_w21815_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name17768 (
		_w5041_,
		_w5108_,
		_w6197_,
		_w19744_,
		_w21816_
	);
	LUT4 #(
		.INIT('h000e)
	) name17769 (
		_w19746_,
		_w19747_,
		_w21816_,
		_w21815_,
		_w21817_
	);
	LUT4 #(
		.INIT('h4500)
	) name17770 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w19745_,
		_w21818_
	);
	LUT3 #(
		.INIT('h01)
	) name17771 (
		_w5937_,
		_w6038_,
		_w19745_,
		_w21819_
	);
	LUT4 #(
		.INIT('h3331)
	) name17772 (
		_w19748_,
		_w21817_,
		_w21819_,
		_w21818_,
		_w21820_
	);
	LUT2 #(
		.INIT('h2)
	) name17773 (
		_w19757_,
		_w21820_,
		_w21821_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17774 (
		_w19757_,
		_w21811_,
		_w21814_,
		_w21821_,
		_w21822_
	);
	LUT3 #(
		.INIT('he2)
	) name17775 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w21788_,
		_w21822_,
		_w21823_
	);
	LUT3 #(
		.INIT('h0b)
	) name17776 (
		_w6245_,
		_w6250_,
		_w19745_,
		_w21824_
	);
	LUT4 #(
		.INIT('h00b0)
	) name17777 (
		_w6555_,
		_w19745_,
		_w19748_,
		_w21824_,
		_w21825_
	);
	LUT4 #(
		.INIT('h00fd)
	) name17778 (
		_w5041_,
		_w5049_,
		_w6996_,
		_w7010_,
		_w21826_
	);
	LUT3 #(
		.INIT('he0)
	) name17779 (
		_w19746_,
		_w19747_,
		_w21826_,
		_w21827_
	);
	LUT4 #(
		.INIT('hf400)
	) name17780 (
		_w7004_,
		_w7008_,
		_w19745_,
		_w21827_,
		_w21828_
	);
	LUT4 #(
		.INIT('h0203)
	) name17781 (
		_w5041_,
		_w5108_,
		_w6566_,
		_w19744_,
		_w21829_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name17782 (
		_w5041_,
		_w5108_,
		_w6522_,
		_w19744_,
		_w21830_
	);
	LUT4 #(
		.INIT('h000e)
	) name17783 (
		_w19746_,
		_w19747_,
		_w21830_,
		_w21829_,
		_w21831_
	);
	LUT4 #(
		.INIT('h4500)
	) name17784 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w19745_,
		_w21832_
	);
	LUT3 #(
		.INIT('h01)
	) name17785 (
		_w6263_,
		_w6362_,
		_w19745_,
		_w21833_
	);
	LUT4 #(
		.INIT('h3331)
	) name17786 (
		_w19748_,
		_w21831_,
		_w21833_,
		_w21832_,
		_w21834_
	);
	LUT2 #(
		.INIT('h2)
	) name17787 (
		_w19757_,
		_w21834_,
		_w21835_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17788 (
		_w19757_,
		_w21825_,
		_w21828_,
		_w21835_,
		_w21836_
	);
	LUT3 #(
		.INIT('he2)
	) name17789 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		_w21788_,
		_w21836_,
		_w21837_
	);
	LUT3 #(
		.INIT('h0b)
	) name17790 (
		_w6643_,
		_w6646_,
		_w19745_,
		_w21838_
	);
	LUT4 #(
		.INIT('h00b0)
	) name17791 (
		_w6591_,
		_w19745_,
		_w19748_,
		_w21838_,
		_w21839_
	);
	LUT4 #(
		.INIT('h00fd)
	) name17792 (
		_w5041_,
		_w5049_,
		_w6955_,
		_w6972_,
		_w21840_
	);
	LUT3 #(
		.INIT('he0)
	) name17793 (
		_w19746_,
		_w19747_,
		_w21840_,
		_w21841_
	);
	LUT4 #(
		.INIT('hf400)
	) name17794 (
		_w6965_,
		_w6970_,
		_w19745_,
		_w21841_,
		_w21842_
	);
	LUT4 #(
		.INIT('h0203)
	) name17795 (
		_w5041_,
		_w5108_,
		_w6637_,
		_w19744_,
		_w21843_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name17796 (
		_w5041_,
		_w5108_,
		_w6602_,
		_w19744_,
		_w21844_
	);
	LUT4 #(
		.INIT('h000e)
	) name17797 (
		_w19746_,
		_w19747_,
		_w21844_,
		_w21843_,
		_w21845_
	);
	LUT4 #(
		.INIT('h4500)
	) name17798 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w19745_,
		_w21846_
	);
	LUT4 #(
		.INIT('h000d)
	) name17799 (
		_w6758_,
		_w19745_,
		_w19746_,
		_w19747_,
		_w21847_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17800 (
		_w19757_,
		_w21845_,
		_w21846_,
		_w21847_,
		_w21848_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17801 (
		_w19757_,
		_w21839_,
		_w21842_,
		_w21848_,
		_w21849_
	);
	LUT3 #(
		.INIT('he2)
	) name17802 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w21788_,
		_w21849_,
		_w21850_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name17803 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		_w19758_,
		_w19765_,
		_w21788_,
		_w21851_
	);
	LUT4 #(
		.INIT('h03aa)
	) name17804 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		_w20181_,
		_w20188_,
		_w21788_,
		_w21852_
	);
	LUT4 #(
		.INIT('h03aa)
	) name17805 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w20194_,
		_w20201_,
		_w21788_,
		_w21853_
	);
	LUT3 #(
		.INIT('hca)
	) name17806 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w20256_,
		_w21788_,
		_w21854_
	);
	LUT4 #(
		.INIT('hf400)
	) name17807 (
		_w5312_,
		_w5315_,
		_w19745_,
		_w19748_,
		_w21855_
	);
	LUT3 #(
		.INIT('hb0)
	) name17808 (
		_w5771_,
		_w19745_,
		_w21855_,
		_w21856_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name17809 (
		_w5041_,
		_w5049_,
		_w5565_,
		_w5549_,
		_w21857_
	);
	LUT3 #(
		.INIT('he0)
	) name17810 (
		_w19746_,
		_w19747_,
		_w21857_,
		_w21858_
	);
	LUT4 #(
		.INIT('hf400)
	) name17811 (
		_w5439_,
		_w5529_,
		_w19745_,
		_w21858_,
		_w21859_
	);
	LUT4 #(
		.INIT('h0203)
	) name17812 (
		_w5041_,
		_w5108_,
		_w5562_,
		_w19744_,
		_w21860_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name17813 (
		_w5041_,
		_w5108_,
		_w5325_,
		_w19744_,
		_w21861_
	);
	LUT4 #(
		.INIT('h000e)
	) name17814 (
		_w19746_,
		_w19747_,
		_w21861_,
		_w21860_,
		_w21862_
	);
	LUT4 #(
		.INIT('h4500)
	) name17815 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w19745_,
		_w21863_
	);
	LUT4 #(
		.INIT('h000d)
	) name17816 (
		_w5760_,
		_w19745_,
		_w19746_,
		_w19747_,
		_w21864_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17817 (
		_w19757_,
		_w21862_,
		_w21863_,
		_w21864_,
		_w21865_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17818 (
		_w19757_,
		_w21856_,
		_w21859_,
		_w21865_,
		_w21866_
	);
	LUT3 #(
		.INIT('he2)
	) name17819 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		_w21788_,
		_w21866_,
		_w21867_
	);
	LUT2 #(
		.INIT('h8)
	) name17820 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w4106_,
		_w21868_
	);
	LUT4 #(
		.INIT('hff80)
	) name17821 (
		_w14570_,
		_w19715_,
		_w19728_,
		_w21868_,
		_w21869_
	);
	LUT4 #(
		.INIT('h4500)
	) name17822 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w13032_,
		_w21870_
	);
	LUT4 #(
		.INIT('hff12)
	) name17823 (
		\bdma_BEAD_reg[7]/NET0131 ,
		_w13032_,
		_w20511_,
		_w21870_,
		_w21871_
	);
	LUT4 #(
		.INIT('h060c)
	) name17824 (
		\bdma_BEAD_reg[5]/NET0131 ,
		\bdma_BEAD_reg[6]/NET0131 ,
		_w13032_,
		_w20510_,
		_w21872_
	);
	LUT4 #(
		.INIT('h4500)
	) name17825 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w13032_,
		_w21873_
	);
	LUT2 #(
		.INIT('he)
	) name17826 (
		_w21872_,
		_w21873_,
		_w21874_
	);
	LUT4 #(
		.INIT('h4500)
	) name17827 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w13032_,
		_w21875_
	);
	LUT4 #(
		.INIT('hff12)
	) name17828 (
		\bdma_BEAD_reg[5]/NET0131 ,
		_w13032_,
		_w20510_,
		_w21875_,
		_w21876_
	);
	LUT3 #(
		.INIT('h40)
	) name17829 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w21877_
	);
	LUT2 #(
		.INIT('h6)
	) name17830 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w21878_
	);
	LUT3 #(
		.INIT('hec)
	) name17831 (
		_w17698_,
		_w21877_,
		_w21878_,
		_w21879_
	);
	LUT3 #(
		.INIT('h40)
	) name17832 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w21880_
	);
	LUT2 #(
		.INIT('h6)
	) name17833 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w21881_
	);
	LUT3 #(
		.INIT('hec)
	) name17834 (
		_w17734_,
		_w21880_,
		_w21881_,
		_w21882_
	);
	LUT3 #(
		.INIT('h13)
	) name17835 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 ,
		_w11300_,
		_w21883_
	);
	LUT4 #(
		.INIT('hccc8)
	) name17836 (
		_w11310_,
		_w11312_,
		_w12315_,
		_w12316_,
		_w21884_
	);
	LUT4 #(
		.INIT('h2322)
	) name17837 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 ,
		_w11303_,
		_w11308_,
		_w21885_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17838 (
		_w11320_,
		_w21883_,
		_w21884_,
		_w21885_,
		_w21886_
	);
	LUT2 #(
		.INIT('h2)
	) name17839 (
		_w11325_,
		_w21886_,
		_w21887_
	);
	LUT4 #(
		.INIT('h0057)
	) name17840 (
		_w9946_,
		_w15570_,
		_w15571_,
		_w21887_,
		_w21888_
	);
	LUT3 #(
		.INIT('h6c)
	) name17841 (
		\sice_ICYC_reg[22]/NET0131 ,
		\sice_ICYC_reg[23]/NET0131 ,
		_w13019_,
		_w21889_
	);
	LUT2 #(
		.INIT('h8)
	) name17842 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w4106_,
		_w21890_
	);
	LUT3 #(
		.INIT('hf8)
	) name17843 (
		_w14570_,
		_w19718_,
		_w21890_,
		_w21891_
	);
	LUT3 #(
		.INIT('h40)
	) name17844 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w21892_
	);
	LUT3 #(
		.INIT('h6c)
	) name17845 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w21893_
	);
	LUT3 #(
		.INIT('hec)
	) name17846 (
		_w17734_,
		_w21892_,
		_w21893_,
		_w21894_
	);
	LUT3 #(
		.INIT('h40)
	) name17847 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w21895_
	);
	LUT3 #(
		.INIT('h6c)
	) name17848 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w21896_
	);
	LUT3 #(
		.INIT('hec)
	) name17849 (
		_w17698_,
		_w21895_,
		_w21896_,
		_w21897_
	);
	LUT3 #(
		.INIT('h40)
	) name17850 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w21898_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17851 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w21899_
	);
	LUT3 #(
		.INIT('hec)
	) name17852 (
		_w17698_,
		_w21898_,
		_w21899_,
		_w21900_
	);
	LUT3 #(
		.INIT('h40)
	) name17853 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w21901_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17854 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[5]/NET0131 ,
		_w17666_,
		_w21902_
	);
	LUT3 #(
		.INIT('hec)
	) name17855 (
		_w17698_,
		_w21901_,
		_w21902_,
		_w21903_
	);
	LUT3 #(
		.INIT('h40)
	) name17856 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w21904_
	);
	LUT4 #(
		.INIT('hff48)
	) name17857 (
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w17698_,
		_w17669_,
		_w21904_,
		_w21905_
	);
	LUT3 #(
		.INIT('h40)
	) name17858 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w21906_
	);
	LUT4 #(
		.INIT('h60c0)
	) name17859 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[13]/NET0131 ,
		_w17734_,
		_w17708_,
		_w21907_
	);
	LUT2 #(
		.INIT('he)
	) name17860 (
		_w21906_,
		_w21907_,
		_w21908_
	);
	LUT3 #(
		.INIT('h40)
	) name17861 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w21909_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17862 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w21910_
	);
	LUT3 #(
		.INIT('hec)
	) name17863 (
		_w17734_,
		_w21909_,
		_w21910_,
		_w21911_
	);
	LUT3 #(
		.INIT('h40)
	) name17864 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w21912_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17865 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[5]/NET0131 ,
		_w17702_,
		_w21913_
	);
	LUT3 #(
		.INIT('hec)
	) name17866 (
		_w17734_,
		_w21912_,
		_w21913_,
		_w21914_
	);
	LUT2 #(
		.INIT('h6)
	) name17867 (
		\sice_ICYC_reg[4]/NET0131 ,
		_w11931_,
		_w21915_
	);
	LUT3 #(
		.INIT('h40)
	) name17868 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w21916_
	);
	LUT4 #(
		.INIT('hff48)
	) name17869 (
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w17734_,
		_w17705_,
		_w21916_,
		_w21917_
	);
	LUT2 #(
		.INIT('h6)
	) name17870 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		_w14698_,
		_w21918_
	);
	LUT2 #(
		.INIT('h6)
	) name17871 (
		\sice_IIRC_reg[4]/NET0131 ,
		_w11934_,
		_w21919_
	);
	LUT3 #(
		.INIT('h40)
	) name17872 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w21920_
	);
	LUT4 #(
		.INIT('h60c0)
	) name17873 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[13]/NET0131 ,
		_w17698_,
		_w17672_,
		_w21921_
	);
	LUT2 #(
		.INIT('he)
	) name17874 (
		_w21920_,
		_w21921_,
		_w21922_
	);
	LUT4 #(
		.INIT('h3555)
	) name17875 (
		\sice_IRR_reg[4]/P0001 ,
		\sice_SPC_reg[14]/P0001 ,
		_w16506_,
		_w21472_,
		_w21923_
	);
	LUT3 #(
		.INIT('h2e)
	) name17876 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		_w4084_,
		_w21923_,
		_w21924_
	);
	LUT4 #(
		.INIT('h3555)
	) name17877 (
		\sice_IRR_reg[9]/P0001 ,
		\sice_SPC_reg[19]/P0001 ,
		_w16506_,
		_w21472_,
		_w21925_
	);
	LUT3 #(
		.INIT('h2e)
	) name17878 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		_w4084_,
		_w21925_,
		_w21926_
	);
	LUT4 #(
		.INIT('h3555)
	) name17879 (
		\sice_IRR_reg[8]/P0001 ,
		\sice_SPC_reg[18]/P0001 ,
		_w16506_,
		_w21472_,
		_w21927_
	);
	LUT3 #(
		.INIT('h2e)
	) name17880 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		_w4084_,
		_w21927_,
		_w21928_
	);
	LUT4 #(
		.INIT('h3555)
	) name17881 (
		\sice_IRR_reg[7]/P0001 ,
		\sice_SPC_reg[17]/P0001 ,
		_w16506_,
		_w21472_,
		_w21929_
	);
	LUT3 #(
		.INIT('h2e)
	) name17882 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		_w4084_,
		_w21929_,
		_w21930_
	);
	LUT4 #(
		.INIT('h3555)
	) name17883 (
		\sice_IRR_reg[6]/P0001 ,
		\sice_SPC_reg[16]/P0001 ,
		_w16506_,
		_w21472_,
		_w21931_
	);
	LUT3 #(
		.INIT('h2e)
	) name17884 (
		\core_c_psq_EXA_reg[6]/P0001 ,
		_w4084_,
		_w21931_,
		_w21932_
	);
	LUT4 #(
		.INIT('h3555)
	) name17885 (
		\sice_IRR_reg[5]/P0001 ,
		\sice_SPC_reg[15]/P0001 ,
		_w16506_,
		_w21472_,
		_w21933_
	);
	LUT3 #(
		.INIT('h2e)
	) name17886 (
		\core_c_psq_EXA_reg[5]/P0001 ,
		_w4084_,
		_w21933_,
		_w21934_
	);
	LUT4 #(
		.INIT('h3555)
	) name17887 (
		\sice_IRR_reg[3]/P0001 ,
		\sice_SPC_reg[13]/P0001 ,
		_w16506_,
		_w21472_,
		_w21935_
	);
	LUT3 #(
		.INIT('h2e)
	) name17888 (
		\core_c_psq_EXA_reg[3]/P0001 ,
		_w4084_,
		_w21935_,
		_w21936_
	);
	LUT4 #(
		.INIT('h3555)
	) name17889 (
		\sice_IRR_reg[2]/P0001 ,
		\sice_SPC_reg[12]/P0001 ,
		_w16506_,
		_w21472_,
		_w21937_
	);
	LUT3 #(
		.INIT('h2e)
	) name17890 (
		\core_c_psq_EXA_reg[2]/P0001 ,
		_w4084_,
		_w21937_,
		_w21938_
	);
	LUT4 #(
		.INIT('h3555)
	) name17891 (
		\sice_IRR_reg[13]/P0001 ,
		\sice_SPC_reg[23]/P0001 ,
		_w16506_,
		_w21472_,
		_w21939_
	);
	LUT3 #(
		.INIT('h2e)
	) name17892 (
		\core_c_psq_EXA_reg[13]/P0001 ,
		_w4084_,
		_w21939_,
		_w21940_
	);
	LUT4 #(
		.INIT('h3555)
	) name17893 (
		\sice_IRR_reg[1]/P0001 ,
		\sice_SPC_reg[11]/P0001 ,
		_w16506_,
		_w21472_,
		_w21941_
	);
	LUT3 #(
		.INIT('h2e)
	) name17894 (
		\core_c_psq_EXA_reg[1]/P0001 ,
		_w4084_,
		_w21941_,
		_w21942_
	);
	LUT4 #(
		.INIT('h3555)
	) name17895 (
		\sice_IRR_reg[12]/P0001 ,
		\sice_SPC_reg[22]/P0001 ,
		_w16506_,
		_w21472_,
		_w21943_
	);
	LUT3 #(
		.INIT('h2e)
	) name17896 (
		\core_c_psq_EXA_reg[12]/P0001 ,
		_w4084_,
		_w21943_,
		_w21944_
	);
	LUT4 #(
		.INIT('h3555)
	) name17897 (
		\sice_IRR_reg[11]/P0001 ,
		\sice_SPC_reg[21]/P0001 ,
		_w16506_,
		_w21472_,
		_w21945_
	);
	LUT3 #(
		.INIT('h2e)
	) name17898 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		_w4084_,
		_w21945_,
		_w21946_
	);
	LUT4 #(
		.INIT('h3555)
	) name17899 (
		\sice_IRR_reg[10]/P0001 ,
		\sice_SPC_reg[20]/P0001 ,
		_w16506_,
		_w21472_,
		_w21947_
	);
	LUT3 #(
		.INIT('h2e)
	) name17900 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		_w4084_,
		_w21947_,
		_w21948_
	);
	LUT4 #(
		.INIT('h3555)
	) name17901 (
		\sice_IRR_reg[0]/P0001 ,
		\sice_SPC_reg[10]/P0001 ,
		_w16506_,
		_w21472_,
		_w21949_
	);
	LUT3 #(
		.INIT('h2e)
	) name17902 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		_w4084_,
		_w21949_,
		_w21950_
	);
	LUT4 #(
		.INIT('h5400)
	) name17903 (
		_w19040_,
		_w19231_,
		_w19232_,
		_w20955_,
		_w21951_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17904 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w19240_,
		_w21952_
	);
	LUT4 #(
		.INIT('h2000)
	) name17905 (
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w21953_
	);
	LUT3 #(
		.INIT('hf8)
	) name17906 (
		_w21951_,
		_w21952_,
		_w21953_,
		_w21954_
	);
	LUT3 #(
		.INIT('hca)
	) name17907 (
		\sport0_txctl_TXSHT_reg[13]/P0001 ,
		\sport0_txctl_TX_reg[14]/P0001 ,
		_w12552_,
		_w21955_
	);
	LUT3 #(
		.INIT('hca)
	) name17908 (
		\sport0_txctl_TXSHT_reg[9]/P0001 ,
		\sport0_txctl_TX_reg[10]/P0001 ,
		_w12552_,
		_w21956_
	);
	LUT3 #(
		.INIT('hca)
	) name17909 (
		\sport0_txctl_TXSHT_reg[8]/P0001 ,
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w12552_,
		_w21957_
	);
	LUT3 #(
		.INIT('hca)
	) name17910 (
		\sport0_txctl_TXSHT_reg[7]/P0001 ,
		\sport0_txctl_TX_reg[8]/P0001 ,
		_w12552_,
		_w21958_
	);
	LUT3 #(
		.INIT('hca)
	) name17911 (
		\sport1_txctl_TXSHT_reg[8]/P0001 ,
		\sport1_txctl_TX_reg[9]/P0001 ,
		_w14269_,
		_w21959_
	);
	LUT3 #(
		.INIT('hca)
	) name17912 (
		\sport0_txctl_TXSHT_reg[5]/P0001 ,
		\sport0_txctl_TX_reg[6]/P0001 ,
		_w12552_,
		_w21960_
	);
	LUT3 #(
		.INIT('hca)
	) name17913 (
		\sport1_txctl_TXSHT_reg[7]/P0001 ,
		\sport1_txctl_TX_reg[8]/P0001 ,
		_w14269_,
		_w21961_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17914 (
		\sice_ICYC_reg[13]/NET0131 ,
		\sice_ICYC_reg[14]/NET0131 ,
		\sice_ICYC_reg[15]/NET0131 ,
		_w13016_,
		_w21962_
	);
	LUT3 #(
		.INIT('hca)
	) name17915 (
		\sport0_txctl_TXSHT_reg[4]/P0001 ,
		\sport0_txctl_TX_reg[5]/P0001 ,
		_w12552_,
		_w21963_
	);
	LUT4 #(
		.INIT('h78f0)
	) name17916 (
		\sice_IIRC_reg[13]/NET0131 ,
		\sice_IIRC_reg[14]/NET0131 ,
		\sice_IIRC_reg[15]/NET0131 ,
		_w13088_,
		_w21964_
	);
	LUT3 #(
		.INIT('hca)
	) name17917 (
		\sport1_txctl_TXSHT_reg[5]/P0001 ,
		\sport1_txctl_TX_reg[6]/P0001 ,
		_w14269_,
		_w21965_
	);
	LUT3 #(
		.INIT('hca)
	) name17918 (
		\sport1_txctl_TXSHT_reg[4]/P0001 ,
		\sport1_txctl_TX_reg[5]/P0001 ,
		_w14269_,
		_w21966_
	);
	LUT3 #(
		.INIT('hca)
	) name17919 (
		\sport0_txctl_TXSHT_reg[2]/P0001 ,
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w12552_,
		_w21967_
	);
	LUT2 #(
		.INIT('h6)
	) name17920 (
		\sice_ICYC_reg[0]/NET0131 ,
		_w19738_,
		_w21968_
	);
	LUT2 #(
		.INIT('h2)
	) name17921 (
		\sice_SPC_reg[5]/P0001 ,
		_w16259_,
		_w21969_
	);
	LUT4 #(
		.INIT('h153f)
	) name17922 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\sice_DBR2_reg[0]/P0001 ,
		_w15508_,
		_w17323_,
		_w21970_
	);
	LUT4 #(
		.INIT('h135f)
	) name17923 (
		\sice_ICYC_reg[5]/NET0131 ,
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w14695_,
		_w16507_,
		_w21971_
	);
	LUT4 #(
		.INIT('h153f)
	) name17924 (
		\sice_DBR1_reg[0]/P0001 ,
		\sice_IIRC_reg[5]/NET0131 ,
		_w15161_,
		_w15544_,
		_w21972_
	);
	LUT4 #(
		.INIT('h8000)
	) name17925 (
		_w21458_,
		_w21970_,
		_w21971_,
		_w21972_,
		_w21973_
	);
	LUT4 #(
		.INIT('h4000)
	) name17926 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[4]/P0001 ,
		_w21974_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17927 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[6]/P0001 ,
		_w21975_
	);
	LUT4 #(
		.INIT('haaa8)
	) name17928 (
		_w16259_,
		_w21458_,
		_w21974_,
		_w21975_,
		_w21976_
	);
	LUT3 #(
		.INIT('hba)
	) name17929 (
		_w21969_,
		_w21973_,
		_w21976_,
		_w21977_
	);
	LUT4 #(
		.INIT('h4000)
	) name17930 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[8]/P0001 ,
		_w21978_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17931 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[10]/P0001 ,
		_w21979_
	);
	LUT3 #(
		.INIT('h01)
	) name17932 (
		_w21458_,
		_w21978_,
		_w21979_,
		_w21980_
	);
	LUT4 #(
		.INIT('h135f)
	) name17933 (
		\sice_DBR1_reg[4]/P0001 ,
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w15544_,
		_w16507_,
		_w21981_
	);
	LUT4 #(
		.INIT('h153f)
	) name17934 (
		\sice_DMR1_reg[3]/NET0131 ,
		\sice_ICYC_reg[9]/NET0131 ,
		_w14695_,
		_w17158_,
		_w21982_
	);
	LUT2 #(
		.INIT('h8)
	) name17935 (
		_w21981_,
		_w21982_,
		_w21983_
	);
	LUT4 #(
		.INIT('h135f)
	) name17936 (
		\sice_DMR2_reg[3]/NET0131 ,
		\sice_IBR1_reg[3]/P0001 ,
		_w15519_,
		_w21464_,
		_w21984_
	);
	LUT4 #(
		.INIT('h135f)
	) name17937 (
		\sice_IIRC_reg[9]/NET0131 ,
		\sice_IMR2_reg[3]/NET0131 ,
		_w15161_,
		_w15527_,
		_w21985_
	);
	LUT4 #(
		.INIT('h153f)
	) name17938 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		\sice_DBR2_reg[4]/P0001 ,
		_w15508_,
		_w17323_,
		_w21986_
	);
	LUT4 #(
		.INIT('h135f)
	) name17939 (
		\sice_IBR2_reg[3]/P0001 ,
		\sice_IMR1_reg[3]/NET0131 ,
		_w15559_,
		_w21468_,
		_w21987_
	);
	LUT4 #(
		.INIT('h8000)
	) name17940 (
		_w21986_,
		_w21987_,
		_w21984_,
		_w21985_,
		_w21988_
	);
	LUT4 #(
		.INIT('h1333)
	) name17941 (
		_w21458_,
		_w21980_,
		_w21983_,
		_w21988_,
		_w21989_
	);
	LUT3 #(
		.INIT('hca)
	) name17942 (
		\sport0_txctl_TXSHT_reg[1]/P0001 ,
		\sport0_txctl_TX_reg[2]/P0001 ,
		_w12552_,
		_w21990_
	);
	LUT4 #(
		.INIT('h4000)
	) name17943 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[5]/P0001 ,
		_w21991_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17944 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[7]/P0001 ,
		_w21992_
	);
	LUT3 #(
		.INIT('h01)
	) name17945 (
		_w21458_,
		_w21991_,
		_w21992_,
		_w21993_
	);
	LUT4 #(
		.INIT('h135f)
	) name17946 (
		\sice_IBR2_reg[0]/P0001 ,
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w15559_,
		_w16507_,
		_w21994_
	);
	LUT4 #(
		.INIT('h153f)
	) name17947 (
		\sice_DBR2_reg[1]/P0001 ,
		\sice_ICYC_reg[6]/NET0131 ,
		_w14695_,
		_w15508_,
		_w21995_
	);
	LUT2 #(
		.INIT('h8)
	) name17948 (
		_w21994_,
		_w21995_,
		_w21996_
	);
	LUT4 #(
		.INIT('h153f)
	) name17949 (
		\sice_IBR1_reg[0]/P0001 ,
		\sice_IMR2_reg[0]/NET0131 ,
		_w15527_,
		_w21464_,
		_w21997_
	);
	LUT4 #(
		.INIT('h135f)
	) name17950 (
		\sice_IIRC_reg[6]/NET0131 ,
		\sice_IMR1_reg[0]/NET0131 ,
		_w15161_,
		_w21468_,
		_w21998_
	);
	LUT4 #(
		.INIT('h153f)
	) name17951 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		\sice_DMR1_reg[0]/NET0131 ,
		_w17158_,
		_w17323_,
		_w21999_
	);
	LUT4 #(
		.INIT('h153f)
	) name17952 (
		\sice_DBR1_reg[1]/P0001 ,
		\sice_DMR2_reg[0]/NET0131 ,
		_w15519_,
		_w15544_,
		_w22000_
	);
	LUT4 #(
		.INIT('h8000)
	) name17953 (
		_w21999_,
		_w22000_,
		_w21997_,
		_w21998_,
		_w22001_
	);
	LUT4 #(
		.INIT('h1333)
	) name17954 (
		_w21458_,
		_w21993_,
		_w21996_,
		_w22001_,
		_w22002_
	);
	LUT3 #(
		.INIT('hca)
	) name17955 (
		\sport0_txctl_TXSHT_reg[0]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w12552_,
		_w22003_
	);
	LUT3 #(
		.INIT('hca)
	) name17956 (
		\sport1_txctl_TXSHT_reg[2]/P0001 ,
		\sport1_txctl_TX_reg[3]/P0001 ,
		_w14269_,
		_w22004_
	);
	LUT3 #(
		.INIT('hca)
	) name17957 (
		\sport1_txctl_TXSHT_reg[1]/P0001 ,
		\sport1_txctl_TX_reg[2]/P0001 ,
		_w14269_,
		_w22005_
	);
	LUT4 #(
		.INIT('h10b0)
	) name17958 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w11294_,
		_w11624_,
		_w15552_,
		_w22006_
	);
	LUT2 #(
		.INIT('h1)
	) name17959 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001 ,
		_w17501_,
		_w22007_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17960 (
		_w12220_,
		_w13610_,
		_w13611_,
		_w17505_,
		_w22008_
	);
	LUT4 #(
		.INIT('h1311)
	) name17961 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001 ,
		_w11303_,
		_w11308_,
		_w22009_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17962 (
		_w12224_,
		_w22007_,
		_w22008_,
		_w22009_,
		_w22010_
	);
	LUT2 #(
		.INIT('h2)
	) name17963 (
		_w17500_,
		_w22010_,
		_w22011_
	);
	LUT2 #(
		.INIT('h1)
	) name17964 (
		_w22006_,
		_w22011_,
		_w22012_
	);
	LUT2 #(
		.INIT('h8)
	) name17965 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		_w12552_,
		_w22013_
	);
	LUT3 #(
		.INIT('hca)
	) name17966 (
		\sport1_txctl_TXSHT_reg[0]/P0001 ,
		\sport1_txctl_TX_reg[1]/P0001 ,
		_w14269_,
		_w22014_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name17967 (
		_w4785_,
		_w4787_,
		_w8596_,
		_w12703_,
		_w22015_
	);
	LUT3 #(
		.INIT('ha8)
	) name17968 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w4721_,
		_w4805_,
		_w22016_
	);
	LUT2 #(
		.INIT('h2)
	) name17969 (
		\memc_Dwrite_E_reg/NET0131 ,
		_w4799_,
		_w22017_
	);
	LUT3 #(
		.INIT('hfe)
	) name17970 (
		_w22016_,
		_w22015_,
		_w22017_,
		_w22018_
	);
	LUT2 #(
		.INIT('h1)
	) name17971 (
		_w4781_,
		_w4796_,
		_w22019_
	);
	LUT4 #(
		.INIT('h4000)
	) name17972 (
		_w4747_,
		_w4768_,
		_w4787_,
		_w22019_,
		_w22020_
	);
	LUT2 #(
		.INIT('h8)
	) name17973 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w22020_,
		_w22021_
	);
	LUT3 #(
		.INIT('h10)
	) name17974 (
		_w4787_,
		_w8596_,
		_w12703_,
		_w22022_
	);
	LUT4 #(
		.INIT('h00b0)
	) name17975 (
		_w4747_,
		_w4768_,
		_w4798_,
		_w9938_,
		_w22023_
	);
	LUT4 #(
		.INIT('h0007)
	) name17976 (
		\memc_Pread_E_reg/NET0131 ,
		_w4805_,
		_w22020_,
		_w22023_,
		_w22024_
	);
	LUT3 #(
		.INIT('hba)
	) name17977 (
		_w22021_,
		_w22022_,
		_w22024_,
		_w22025_
	);
	LUT3 #(
		.INIT('h40)
	) name17978 (
		_w4787_,
		_w8596_,
		_w12703_,
		_w22026_
	);
	LUT4 #(
		.INIT('h8a00)
	) name17979 (
		\memc_Dwrite_E_reg/NET0131 ,
		_w4747_,
		_w4768_,
		_w4798_,
		_w22027_
	);
	LUT3 #(
		.INIT('h07)
	) name17980 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w4805_,
		_w22027_,
		_w22028_
	);
	LUT2 #(
		.INIT('h4)
	) name17981 (
		_w22026_,
		_w22028_,
		_w22029_
	);
	LUT2 #(
		.INIT('h8)
	) name17982 (
		\sport1_txctl_TX_reg[0]/P0001 ,
		_w14269_,
		_w22030_
	);
	LUT4 #(
		.INIT('hdccc)
	) name17983 (
		_w4747_,
		_w4766_,
		_w4768_,
		_w22019_,
		_w22031_
	);
	LUT2 #(
		.INIT('h2)
	) name17984 (
		\core_c_psq_PCS_reg[12]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w22032_
	);
	LUT4 #(
		.INIT('ha820)
	) name17985 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		_w22033_
	);
	LUT2 #(
		.INIT('h1)
	) name17986 (
		_w22032_,
		_w22033_,
		_w22034_
	);
	LUT2 #(
		.INIT('he)
	) name17987 (
		_w22032_,
		_w22033_,
		_w22035_
	);
	LUT4 #(
		.INIT('h5455)
	) name17988 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4862_,
		_w4864_,
		_w22034_,
		_w22036_
	);
	LUT4 #(
		.INIT('h00d8)
	) name17989 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4069_,
		_w12054_,
		_w22036_,
		_w22037_
	);
	LUT2 #(
		.INIT('h2)
	) name17990 (
		_w4106_,
		_w22037_,
		_w22038_
	);
	LUT2 #(
		.INIT('h2)
	) name17991 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12284_,
		_w22039_
	);
	LUT4 #(
		.INIT('h0400)
	) name17992 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w18113_,
		_w18118_,
		_w18135_,
		_w22040_
	);
	LUT4 #(
		.INIT('h222e)
	) name17993 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001 ,
		_w11946_,
		_w22039_,
		_w22040_,
		_w22041_
	);
	LUT4 #(
		.INIT('h222e)
	) name17994 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001 ,
		_w12048_,
		_w22039_,
		_w22040_,
		_w22042_
	);
	LUT4 #(
		.INIT('h8808)
	) name17995 (
		_w11710_,
		_w11713_,
		_w11735_,
		_w14466_,
		_w22043_
	);
	LUT3 #(
		.INIT('h48)
	) name17996 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w22043_,
		_w22044_
	);
	LUT4 #(
		.INIT('h00ba)
	) name17997 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w11739_,
		_w22045_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name17998 (
		\auctl_T0Sack_reg/NET0131 ,
		\sport0_txctl_TX_reg[5]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w11738_,
		_w22046_
	);
	LUT2 #(
		.INIT('h4)
	) name17999 (
		_w22045_,
		_w22046_,
		_w22047_
	);
	LUT2 #(
		.INIT('he)
	) name18000 (
		_w22044_,
		_w22047_,
		_w22048_
	);
	LUT4 #(
		.INIT('hb1e4)
	) name18001 (
		\ISCLK0_pad ,
		\T_SCLK0_pad ,
		\sport0_cfg_SCLKi_h_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w22049_
	);
	LUT4 #(
		.INIT('hb1e4)
	) name18002 (
		\ISCLK1_pad ,
		\T_SCLK1_pad ,
		\sport1_cfg_SCLKi_h_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w22050_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18003 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11830_,
		_w14918_,
		_w18663_,
		_w22051_
	);
	LUT4 #(
		.INIT('h5545)
	) name18004 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w22052_
	);
	LUT2 #(
		.INIT('h1)
	) name18005 (
		_w22051_,
		_w22052_,
		_w22053_
	);
	LUT4 #(
		.INIT('h5401)
	) name18006 (
		_w9455_,
		_w9456_,
		_w12116_,
		_w12119_,
		_w22054_
	);
	LUT2 #(
		.INIT('h8)
	) name18007 (
		_w9455_,
		_w9828_,
		_w22055_
	);
	LUT4 #(
		.INIT('heee2)
	) name18008 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001 ,
		_w9895_,
		_w22054_,
		_w22055_,
		_w22056_
	);
	LUT4 #(
		.INIT('heee2)
	) name18009 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001 ,
		_w9454_,
		_w22054_,
		_w22055_,
		_w22057_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18010 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11830_,
		_w14866_,
		_w18311_,
		_w22058_
	);
	LUT4 #(
		.INIT('h5545)
	) name18011 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w22059_
	);
	LUT2 #(
		.INIT('h1)
	) name18012 (
		_w22058_,
		_w22059_,
		_w22060_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18013 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11329_,
		_w14918_,
		_w18663_,
		_w22061_
	);
	LUT2 #(
		.INIT('h1)
	) name18014 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001 ,
		_w11329_,
		_w22062_
	);
	LUT2 #(
		.INIT('h1)
	) name18015 (
		_w22061_,
		_w22062_,
		_w22063_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18016 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11329_,
		_w14866_,
		_w18311_,
		_w22064_
	);
	LUT2 #(
		.INIT('h1)
	) name18017 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001 ,
		_w11329_,
		_w22065_
	);
	LUT2 #(
		.INIT('h1)
	) name18018 (
		_w22064_,
		_w22065_,
		_w22066_
	);
	LUT2 #(
		.INIT('h2)
	) name18019 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w11318_,
		_w22067_
	);
	LUT4 #(
		.INIT('h4000)
	) name18020 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12451_,
		_w17953_,
		_w17977_,
		_w22068_
	);
	LUT4 #(
		.INIT('h222e)
	) name18021 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001 ,
		_w11946_,
		_w22067_,
		_w22068_,
		_w22069_
	);
	LUT4 #(
		.INIT('h01fe)
	) name18022 (
		\sport0_txctl_Bcnt_reg[0]/NET0131 ,
		\sport0_txctl_Bcnt_reg[1]/NET0131 ,
		\sport0_txctl_Bcnt_reg[2]/NET0131 ,
		\sport0_txctl_Bcnt_reg[3]/NET0131 ,
		_w22070_
	);
	LUT3 #(
		.INIT('h01)
	) name18023 (
		_w14596_,
		_w14597_,
		_w22070_,
		_w22071_
	);
	LUT4 #(
		.INIT('h1113)
	) name18024 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w14596_,
		_w14597_,
		_w22072_
	);
	LUT2 #(
		.INIT('hb)
	) name18025 (
		_w22071_,
		_w22072_,
		_w22073_
	);
	LUT4 #(
		.INIT('h01fe)
	) name18026 (
		\sport1_txctl_Bcnt_reg[0]/NET0131 ,
		\sport1_txctl_Bcnt_reg[1]/NET0131 ,
		\sport1_txctl_Bcnt_reg[2]/NET0131 ,
		\sport1_txctl_Bcnt_reg[3]/NET0131 ,
		_w22074_
	);
	LUT3 #(
		.INIT('h01)
	) name18027 (
		_w14590_,
		_w14591_,
		_w22074_,
		_w22075_
	);
	LUT4 #(
		.INIT('h1113)
	) name18028 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w14590_,
		_w14591_,
		_w22076_
	);
	LUT2 #(
		.INIT('hb)
	) name18029 (
		_w22075_,
		_w22076_,
		_w22077_
	);
	LUT3 #(
		.INIT('h1e)
	) name18030 (
		\sport1_txctl_Bcnt_reg[0]/NET0131 ,
		\sport1_txctl_Bcnt_reg[1]/NET0131 ,
		\sport1_txctl_Bcnt_reg[2]/NET0131 ,
		_w22078_
	);
	LUT3 #(
		.INIT('h01)
	) name18031 (
		_w14590_,
		_w14591_,
		_w22078_,
		_w22079_
	);
	LUT4 #(
		.INIT('h1113)
	) name18032 (
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w14590_,
		_w14591_,
		_w22080_
	);
	LUT2 #(
		.INIT('hb)
	) name18033 (
		_w22079_,
		_w22080_,
		_w22081_
	);
	LUT4 #(
		.INIT('h222e)
	) name18034 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001 ,
		_w12048_,
		_w22067_,
		_w22068_,
		_w22082_
	);
	LUT2 #(
		.INIT('h6)
	) name18035 (
		\sport1_txctl_Bcnt_reg[0]/NET0131 ,
		\sport1_txctl_Bcnt_reg[1]/NET0131 ,
		_w22083_
	);
	LUT3 #(
		.INIT('h01)
	) name18036 (
		_w14590_,
		_w14591_,
		_w22083_,
		_w22084_
	);
	LUT4 #(
		.INIT('h1113)
	) name18037 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w14590_,
		_w14591_,
		_w22085_
	);
	LUT2 #(
		.INIT('hb)
	) name18038 (
		_w22084_,
		_w22085_,
		_w22086_
	);
	LUT2 #(
		.INIT('h1)
	) name18039 (
		T_IRDn_pad,
		T_ISn_pad,
		_w22087_
	);
	LUT3 #(
		.INIT('ha8)
	) name18040 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w14590_,
		_w14591_,
		_w22088_
	);
	LUT4 #(
		.INIT('h5554)
	) name18041 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		\sport1_txctl_Bcnt_reg[0]/NET0131 ,
		_w14590_,
		_w14591_,
		_w22089_
	);
	LUT2 #(
		.INIT('hb)
	) name18042 (
		_w22088_,
		_w22089_,
		_w22090_
	);
	LUT2 #(
		.INIT('h6)
	) name18043 (
		\sport0_txctl_Bcnt_reg[0]/NET0131 ,
		\sport0_txctl_Bcnt_reg[1]/NET0131 ,
		_w22091_
	);
	LUT3 #(
		.INIT('h01)
	) name18044 (
		_w14596_,
		_w14597_,
		_w22091_,
		_w22092_
	);
	LUT4 #(
		.INIT('h1113)
	) name18045 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w14596_,
		_w14597_,
		_w22093_
	);
	LUT2 #(
		.INIT('hb)
	) name18046 (
		_w22092_,
		_w22093_,
		_w22094_
	);
	LUT3 #(
		.INIT('ha8)
	) name18047 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w14596_,
		_w14597_,
		_w22095_
	);
	LUT4 #(
		.INIT('h5554)
	) name18048 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		\sport0_txctl_Bcnt_reg[0]/NET0131 ,
		_w14596_,
		_w14597_,
		_w22096_
	);
	LUT2 #(
		.INIT('hb)
	) name18049 (
		_w22095_,
		_w22096_,
		_w22097_
	);
	LUT3 #(
		.INIT('h1e)
	) name18050 (
		\sport0_txctl_Bcnt_reg[0]/NET0131 ,
		\sport0_txctl_Bcnt_reg[1]/NET0131 ,
		\sport0_txctl_Bcnt_reg[2]/NET0131 ,
		_w22098_
	);
	LUT3 #(
		.INIT('h01)
	) name18051 (
		_w14596_,
		_w14597_,
		_w22098_,
		_w22099_
	);
	LUT4 #(
		.INIT('h1113)
	) name18052 (
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w14596_,
		_w14597_,
		_w22100_
	);
	LUT2 #(
		.INIT('hb)
	) name18053 (
		_w22099_,
		_w22100_,
		_w22101_
	);
	LUT3 #(
		.INIT('h2a)
	) name18054 (
		_w14835_,
		_w20441_,
		_w20450_,
		_w22102_
	);
	LUT4 #(
		.INIT('h7f80)
	) name18055 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_OUTcnt_reg[1]/NET0131 ,
		\clkc_OUTcnt_reg[2]/NET0131 ,
		\clkc_OUTcnt_reg[3]/NET0131 ,
		_w22103_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18056 (
		_w12254_,
		_w12258_,
		_w12263_,
		_w22103_,
		_w22104_
	);
	LUT4 #(
		.INIT('h7f80)
	) name18057 (
		\clkc_STDcnt_reg[0]/NET0131 ,
		\clkc_STDcnt_reg[1]/NET0131 ,
		\clkc_STDcnt_reg[2]/NET0131 ,
		\clkc_STDcnt_reg[3]/NET0131 ,
		_w22105_
	);
	LUT3 #(
		.INIT('h70)
	) name18058 (
		_w19400_,
		_w19405_,
		_w22105_,
		_w22106_
	);
	LUT3 #(
		.INIT('h80)
	) name18059 (
		_w5028_,
		_w5044_,
		_w5045_,
		_w22107_
	);
	LUT3 #(
		.INIT('h01)
	) name18060 (
		_w5029_,
		_w12917_,
		_w22107_,
		_w22108_
	);
	LUT4 #(
		.INIT('h2000)
	) name18061 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w5027_,
		_w5028_,
		_w22109_
	);
	LUT2 #(
		.INIT('h1)
	) name18062 (
		_w13450_,
		_w22109_,
		_w22110_
	);
	LUT2 #(
		.INIT('h8)
	) name18063 (
		_w22108_,
		_w22110_,
		_w22111_
	);
	LUT4 #(
		.INIT('h1000)
	) name18064 (
		\core_c_dec_Usecond_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22112_
	);
	LUT4 #(
		.INIT('h020a)
	) name18065 (
		_w4102_,
		_w9933_,
		_w22112_,
		_w22111_,
		_w22113_
	);
	LUT4 #(
		.INIT('h7f80)
	) name18066 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		_w22114_
	);
	LUT3 #(
		.INIT('h20)
	) name18067 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w12108_,
		_w22114_,
		_w22115_
	);
	LUT3 #(
		.INIT('hb0)
	) name18068 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		\idma_WRcyc_reg/NET0131 ,
		_w22116_
	);
	LUT4 #(
		.INIT('h0e00)
	) name18069 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		\idma_RDCMD_d1_reg/P0001 ,
		\idma_RDCMD_reg/P0001 ,
		_w22117_
	);
	LUT4 #(
		.INIT('hffea)
	) name18070 (
		\idma_DSreq_reg/NET0131 ,
		_w12812_,
		_w22116_,
		_w22117_,
		_w22118_
	);
	LUT2 #(
		.INIT('h8)
	) name18071 (
		_w12621_,
		_w14140_,
		_w22119_
	);
	LUT3 #(
		.INIT('h10)
	) name18072 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22120_
	);
	LUT3 #(
		.INIT('h2a)
	) name18073 (
		\IRFS1_pad ,
		_w12621_,
		_w14140_,
		_w22121_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18074 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22121_,
		_w22122_
	);
	LUT4 #(
		.INIT('h10ff)
	) name18075 (
		_w7465_,
		_w7565_,
		_w22119_,
		_w22122_,
		_w22123_
	);
	LUT3 #(
		.INIT('h2a)
	) name18076 (
		\ITFS1_pad ,
		_w12621_,
		_w14140_,
		_w22124_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18077 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22124_,
		_w22125_
	);
	LUT4 #(
		.INIT('h10ff)
	) name18078 (
		_w7140_,
		_w7240_,
		_w22119_,
		_w22125_,
		_w22126_
	);
	LUT4 #(
		.INIT('h4500)
	) name18079 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w22119_,
		_w22127_
	);
	LUT3 #(
		.INIT('h2a)
	) name18080 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w12621_,
		_w14140_,
		_w22128_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18081 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22128_,
		_w22129_
	);
	LUT2 #(
		.INIT('hb)
	) name18082 (
		_w22127_,
		_w22129_,
		_w22130_
	);
	LUT3 #(
		.INIT('h2a)
	) name18083 (
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w12621_,
		_w14140_,
		_w22131_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18084 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22131_,
		_w22132_
	);
	LUT4 #(
		.INIT('h10ff)
	) name18085 (
		_w6263_,
		_w6362_,
		_w22119_,
		_w22132_,
		_w22133_
	);
	LUT3 #(
		.INIT('h2a)
	) name18086 (
		\sport1_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w12621_,
		_w14140_,
		_w22134_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18087 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22134_,
		_w22135_
	);
	LUT4 #(
		.INIT('h10ff)
	) name18088 (
		_w5937_,
		_w6038_,
		_w22119_,
		_w22135_,
		_w22136_
	);
	LUT4 #(
		.INIT('h4500)
	) name18089 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w22119_,
		_w22137_
	);
	LUT3 #(
		.INIT('h2a)
	) name18090 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w12621_,
		_w14140_,
		_w22138_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18091 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22138_,
		_w22139_
	);
	LUT2 #(
		.INIT('hb)
	) name18092 (
		_w22137_,
		_w22139_,
		_w22140_
	);
	LUT2 #(
		.INIT('h1)
	) name18093 (
		\sport1_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w11984_,
		_w22141_
	);
	LUT4 #(
		.INIT('hba00)
	) name18094 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w11986_,
		_w22142_
	);
	LUT2 #(
		.INIT('h1)
	) name18095 (
		_w22141_,
		_w22142_,
		_w22143_
	);
	LUT2 #(
		.INIT('h1)
	) name18096 (
		\sport1_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w11984_,
		_w22144_
	);
	LUT4 #(
		.INIT('hba00)
	) name18097 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w11986_,
		_w22145_
	);
	LUT2 #(
		.INIT('h1)
	) name18098 (
		_w22144_,
		_w22145_,
		_w22146_
	);
	LUT2 #(
		.INIT('h1)
	) name18099 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w11984_,
		_w22147_
	);
	LUT3 #(
		.INIT('h0b)
	) name18100 (
		_w8802_,
		_w11986_,
		_w22147_,
		_w22148_
	);
	LUT4 #(
		.INIT('h4000)
	) name18101 (
		\memc_MMR_web_reg/NET0131 ,
		_w9431_,
		_w11604_,
		_w12622_,
		_w22149_
	);
	LUT4 #(
		.INIT('h4500)
	) name18102 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w22149_,
		_w22150_
	);
	LUT2 #(
		.INIT('h2)
	) name18103 (
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w22149_,
		_w22151_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18104 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22151_,
		_w22152_
	);
	LUT2 #(
		.INIT('hb)
	) name18105 (
		_w22150_,
		_w22152_,
		_w22153_
	);
	LUT4 #(
		.INIT('h4500)
	) name18106 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w22149_,
		_w22154_
	);
	LUT2 #(
		.INIT('h2)
	) name18107 (
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w22149_,
		_w22155_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18108 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22155_,
		_w22156_
	);
	LUT2 #(
		.INIT('hb)
	) name18109 (
		_w22154_,
		_w22156_,
		_w22157_
	);
	LUT4 #(
		.INIT('h4500)
	) name18110 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w22149_,
		_w22158_
	);
	LUT2 #(
		.INIT('h2)
	) name18111 (
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w22149_,
		_w22159_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18112 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22159_,
		_w22160_
	);
	LUT2 #(
		.INIT('hb)
	) name18113 (
		_w22158_,
		_w22160_,
		_w22161_
	);
	LUT4 #(
		.INIT('h4500)
	) name18114 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w22149_,
		_w22162_
	);
	LUT2 #(
		.INIT('h2)
	) name18115 (
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w22149_,
		_w22163_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18116 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22163_,
		_w22164_
	);
	LUT2 #(
		.INIT('hb)
	) name18117 (
		_w22162_,
		_w22164_,
		_w22165_
	);
	LUT4 #(
		.INIT('h4500)
	) name18118 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w22149_,
		_w22166_
	);
	LUT2 #(
		.INIT('h2)
	) name18119 (
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w22149_,
		_w22167_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18120 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22167_,
		_w22168_
	);
	LUT2 #(
		.INIT('hb)
	) name18121 (
		_w22166_,
		_w22168_,
		_w22169_
	);
	LUT4 #(
		.INIT('h4500)
	) name18122 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w22149_,
		_w22170_
	);
	LUT2 #(
		.INIT('h2)
	) name18123 (
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w22149_,
		_w22171_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18124 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22171_,
		_w22172_
	);
	LUT2 #(
		.INIT('hb)
	) name18125 (
		_w22170_,
		_w22172_,
		_w22173_
	);
	LUT4 #(
		.INIT('h4500)
	) name18126 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w22149_,
		_w22174_
	);
	LUT2 #(
		.INIT('h2)
	) name18127 (
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w22149_,
		_w22175_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18128 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22175_,
		_w22176_
	);
	LUT2 #(
		.INIT('hb)
	) name18129 (
		_w22174_,
		_w22176_,
		_w22177_
	);
	LUT4 #(
		.INIT('h4500)
	) name18130 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w22149_,
		_w22178_
	);
	LUT2 #(
		.INIT('h2)
	) name18131 (
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w22149_,
		_w22179_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18132 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22179_,
		_w22180_
	);
	LUT2 #(
		.INIT('hb)
	) name18133 (
		_w22178_,
		_w22180_,
		_w22181_
	);
	LUT4 #(
		.INIT('h7f80)
	) name18134 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		_w22182_
	);
	LUT3 #(
		.INIT('h20)
	) name18135 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w12086_,
		_w22182_,
		_w22183_
	);
	LUT2 #(
		.INIT('h2)
	) name18136 (
		\ITFS0_pad ,
		_w11607_,
		_w22184_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18137 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22184_,
		_w22185_
	);
	LUT4 #(
		.INIT('h10ff)
	) name18138 (
		_w7140_,
		_w7240_,
		_w11607_,
		_w22185_,
		_w22186_
	);
	LUT2 #(
		.INIT('h2)
	) name18139 (
		\IRFS0_pad ,
		_w11607_,
		_w22187_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18140 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22187_,
		_w22188_
	);
	LUT4 #(
		.INIT('h10ff)
	) name18141 (
		_w7465_,
		_w7565_,
		_w11607_,
		_w22188_,
		_w22189_
	);
	LUT4 #(
		.INIT('h4500)
	) name18142 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w11607_,
		_w22190_
	);
	LUT2 #(
		.INIT('h2)
	) name18143 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w11607_,
		_w22191_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18144 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22191_,
		_w22192_
	);
	LUT2 #(
		.INIT('hb)
	) name18145 (
		_w22190_,
		_w22192_,
		_w22193_
	);
	LUT2 #(
		.INIT('h2)
	) name18146 (
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w11607_,
		_w22194_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18147 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22194_,
		_w22195_
	);
	LUT4 #(
		.INIT('h10ff)
	) name18148 (
		_w6263_,
		_w6362_,
		_w11607_,
		_w22195_,
		_w22196_
	);
	LUT2 #(
		.INIT('h2)
	) name18149 (
		\sport0_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w11607_,
		_w22197_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18150 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22197_,
		_w22198_
	);
	LUT4 #(
		.INIT('h10ff)
	) name18151 (
		_w5937_,
		_w6038_,
		_w11607_,
		_w22198_,
		_w22199_
	);
	LUT4 #(
		.INIT('h4500)
	) name18152 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w11607_,
		_w22200_
	);
	LUT2 #(
		.INIT('h2)
	) name18153 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w11607_,
		_w22201_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18154 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22201_,
		_w22202_
	);
	LUT2 #(
		.INIT('hb)
	) name18155 (
		_w22200_,
		_w22202_,
		_w22203_
	);
	LUT2 #(
		.INIT('h1)
	) name18156 (
		\sport0_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w11609_,
		_w22204_
	);
	LUT4 #(
		.INIT('hba00)
	) name18157 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w12031_,
		_w22205_
	);
	LUT2 #(
		.INIT('h1)
	) name18158 (
		_w22204_,
		_w22205_,
		_w22206_
	);
	LUT2 #(
		.INIT('h1)
	) name18159 (
		\sport0_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w11609_,
		_w22207_
	);
	LUT4 #(
		.INIT('hba00)
	) name18160 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w12031_,
		_w22208_
	);
	LUT2 #(
		.INIT('h1)
	) name18161 (
		_w22207_,
		_w22208_,
		_w22209_
	);
	LUT2 #(
		.INIT('h1)
	) name18162 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w11609_,
		_w22210_
	);
	LUT3 #(
		.INIT('h0b)
	) name18163 (
		_w8802_,
		_w12031_,
		_w22210_,
		_w22211_
	);
	LUT4 #(
		.INIT('h4500)
	) name18164 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w11787_,
		_w22212_
	);
	LUT2 #(
		.INIT('h2)
	) name18165 (
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w11787_,
		_w22213_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18166 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22213_,
		_w22214_
	);
	LUT2 #(
		.INIT('hb)
	) name18167 (
		_w22212_,
		_w22214_,
		_w22215_
	);
	LUT4 #(
		.INIT('h4500)
	) name18168 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w11787_,
		_w22216_
	);
	LUT2 #(
		.INIT('h2)
	) name18169 (
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w11787_,
		_w22217_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18170 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22217_,
		_w22218_
	);
	LUT2 #(
		.INIT('hb)
	) name18171 (
		_w22216_,
		_w22218_,
		_w22219_
	);
	LUT4 #(
		.INIT('h4500)
	) name18172 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w11787_,
		_w22220_
	);
	LUT2 #(
		.INIT('h2)
	) name18173 (
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w11787_,
		_w22221_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18174 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22221_,
		_w22222_
	);
	LUT2 #(
		.INIT('hb)
	) name18175 (
		_w22220_,
		_w22222_,
		_w22223_
	);
	LUT4 #(
		.INIT('h4500)
	) name18176 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w11787_,
		_w22224_
	);
	LUT2 #(
		.INIT('h2)
	) name18177 (
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w11787_,
		_w22225_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18178 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22225_,
		_w22226_
	);
	LUT2 #(
		.INIT('hb)
	) name18179 (
		_w22224_,
		_w22226_,
		_w22227_
	);
	LUT4 #(
		.INIT('h4500)
	) name18180 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w11787_,
		_w22228_
	);
	LUT2 #(
		.INIT('h2)
	) name18181 (
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w11787_,
		_w22229_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18182 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22229_,
		_w22230_
	);
	LUT2 #(
		.INIT('hb)
	) name18183 (
		_w22228_,
		_w22230_,
		_w22231_
	);
	LUT4 #(
		.INIT('h4500)
	) name18184 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w11787_,
		_w22232_
	);
	LUT2 #(
		.INIT('h2)
	) name18185 (
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w11787_,
		_w22233_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18186 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22233_,
		_w22234_
	);
	LUT2 #(
		.INIT('hb)
	) name18187 (
		_w22232_,
		_w22234_,
		_w22235_
	);
	LUT4 #(
		.INIT('h4500)
	) name18188 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w11787_,
		_w22236_
	);
	LUT2 #(
		.INIT('h2)
	) name18189 (
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w11787_,
		_w22237_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18190 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22237_,
		_w22238_
	);
	LUT2 #(
		.INIT('hb)
	) name18191 (
		_w22236_,
		_w22238_,
		_w22239_
	);
	LUT4 #(
		.INIT('h4500)
	) name18192 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w11787_,
		_w22240_
	);
	LUT2 #(
		.INIT('h2)
	) name18193 (
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w11787_,
		_w22241_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18194 (
		_w8757_,
		_w8760_,
		_w11609_,
		_w22241_,
		_w22242_
	);
	LUT2 #(
		.INIT('hb)
	) name18195 (
		_w22240_,
		_w22242_,
		_w22243_
	);
	LUT4 #(
		.INIT('h0020)
	) name18196 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w22244_
	);
	LUT4 #(
		.INIT('h0800)
	) name18197 (
		_w5658_,
		_w9431_,
		_w15880_,
		_w22244_,
		_w22245_
	);
	LUT2 #(
		.INIT('h2)
	) name18198 (
		\PIO_out[6]_pad ,
		_w22245_,
		_w22246_
	);
	LUT4 #(
		.INIT('h4500)
	) name18199 (
		_w7927_,
		_w8040_,
		_w8042_,
		_w22245_,
		_w22247_
	);
	LUT4 #(
		.INIT('heee4)
	) name18200 (
		\PIO_oe[6]_pad ,
		\pio_PIO_RES_reg[6]/NET0131 ,
		_w22246_,
		_w22247_,
		_w22248_
	);
	LUT4 #(
		.INIT('h0800)
	) name18201 (
		_w5658_,
		_w9431_,
		_w15888_,
		_w22244_,
		_w22249_
	);
	LUT2 #(
		.INIT('h2)
	) name18202 (
		\PIO_out[4]_pad ,
		_w22249_,
		_w22250_
	);
	LUT4 #(
		.INIT('h4500)
	) name18203 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w22249_,
		_w22251_
	);
	LUT4 #(
		.INIT('heee4)
	) name18204 (
		\PIO_oe[4]_pad ,
		\pio_PIO_RES_reg[4]/NET0131 ,
		_w22250_,
		_w22251_,
		_w22252_
	);
	LUT4 #(
		.INIT('h0800)
	) name18205 (
		_w5658_,
		_w9431_,
		_w15875_,
		_w22244_,
		_w22253_
	);
	LUT2 #(
		.INIT('h2)
	) name18206 (
		\PIO_out[2]_pad ,
		_w22253_,
		_w22254_
	);
	LUT4 #(
		.INIT('h4500)
	) name18207 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w22253_,
		_w22255_
	);
	LUT4 #(
		.INIT('heee4)
	) name18208 (
		\PIO_oe[2]_pad ,
		\pio_PIO_RES_reg[2]/NET0131 ,
		_w22254_,
		_w22255_,
		_w22256_
	);
	LUT4 #(
		.INIT('h0800)
	) name18209 (
		_w5658_,
		_w9431_,
		_w15870_,
		_w22244_,
		_w22257_
	);
	LUT4 #(
		.INIT('hfc55)
	) name18210 (
		\PIO_out[10]_pad ,
		_w8757_,
		_w8760_,
		_w22257_,
		_w22258_
	);
	LUT3 #(
		.INIT('h4e)
	) name18211 (
		\PIO_oe[10]_pad ,
		\pio_PIO_RES_reg[10]/NET0131 ,
		_w22258_,
		_w22259_
	);
	LUT4 #(
		.INIT('h0800)
	) name18212 (
		_w5658_,
		_w9431_,
		_w15865_,
		_w22244_,
		_w22260_
	);
	LUT2 #(
		.INIT('h2)
	) name18213 (
		\PIO_out[0]_pad ,
		_w22260_,
		_w22261_
	);
	LUT4 #(
		.INIT('h4500)
	) name18214 (
		_w5784_,
		_w5911_,
		_w5913_,
		_w22260_,
		_w22262_
	);
	LUT4 #(
		.INIT('heee4)
	) name18215 (
		\PIO_oe[0]_pad ,
		\pio_PIO_RES_reg[0]/NET0131 ,
		_w22261_,
		_w22262_,
		_w22263_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name18216 (
		\sice_DMR1_reg[8]/NET0131 ,
		\sice_SPC_reg[14]/P0001 ,
		_w14460_,
		_w17158_,
		_w22264_
	);
	LUT3 #(
		.INIT('he8)
	) name18217 (
		\core_c_psq_T_IRQL0p_reg/P0001 ,
		\core_c_psq_irql0_de_IN_syn_reg/P0001 ,
		\core_c_psq_irql0_de_OUT_reg/P0001 ,
		_w22265_
	);
	LUT4 #(
		.INIT('h0800)
	) name18218 (
		_w5658_,
		_w9431_,
		_w15860_,
		_w22244_,
		_w22266_
	);
	LUT4 #(
		.INIT('ha088)
	) name18219 (
		\PIO_oe[9]_pad ,
		\PIO_out[9]_pad ,
		_w5760_,
		_w22266_,
		_w22267_
	);
	LUT2 #(
		.INIT('h4)
	) name18220 (
		\PIO_oe[9]_pad ,
		\pio_PIO_RES_reg[9]/NET0131 ,
		_w22268_
	);
	LUT2 #(
		.INIT('he)
	) name18221 (
		_w22267_,
		_w22268_,
		_w22269_
	);
	LUT4 #(
		.INIT('ha088)
	) name18222 (
		\PIO_oe[8]_pad ,
		\PIO_out[8]_pad ,
		_w6758_,
		_w22266_,
		_w22270_
	);
	LUT2 #(
		.INIT('h4)
	) name18223 (
		\PIO_oe[8]_pad ,
		\pio_PIO_RES_reg[8]/NET0131 ,
		_w22271_
	);
	LUT2 #(
		.INIT('he)
	) name18224 (
		_w22270_,
		_w22271_,
		_w22272_
	);
	LUT2 #(
		.INIT('h2)
	) name18225 (
		\PIO_out[5]_pad ,
		_w22249_,
		_w22273_
	);
	LUT4 #(
		.INIT('h4500)
	) name18226 (
		_w7592_,
		_w7707_,
		_w7709_,
		_w22249_,
		_w22274_
	);
	LUT4 #(
		.INIT('heee4)
	) name18227 (
		\PIO_oe[5]_pad ,
		\pio_PIO_RES_reg[5]/NET0131 ,
		_w22273_,
		_w22274_,
		_w22275_
	);
	LUT2 #(
		.INIT('h2)
	) name18228 (
		\PIO_out[7]_pad ,
		_w22245_,
		_w22276_
	);
	LUT4 #(
		.INIT('h4500)
	) name18229 (
		_w7793_,
		_w7903_,
		_w7905_,
		_w22245_,
		_w22277_
	);
	LUT4 #(
		.INIT('heee4)
	) name18230 (
		\PIO_oe[7]_pad ,
		\pio_PIO_RES_reg[7]/NET0131 ,
		_w22276_,
		_w22277_,
		_w22278_
	);
	LUT2 #(
		.INIT('h2)
	) name18231 (
		\PIO_out[3]_pad ,
		_w22253_,
		_w22279_
	);
	LUT4 #(
		.INIT('h4500)
	) name18232 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w22253_,
		_w22280_
	);
	LUT4 #(
		.INIT('heee4)
	) name18233 (
		\PIO_oe[3]_pad ,
		\pio_PIO_RES_reg[3]/NET0131 ,
		_w22279_,
		_w22280_,
		_w22281_
	);
	LUT2 #(
		.INIT('h2)
	) name18234 (
		\PIO_out[1]_pad ,
		_w22260_,
		_w22282_
	);
	LUT4 #(
		.INIT('h4500)
	) name18235 (
		_w6774_,
		_w6894_,
		_w6896_,
		_w22260_,
		_w22283_
	);
	LUT4 #(
		.INIT('heee4)
	) name18236 (
		\PIO_oe[1]_pad ,
		\pio_PIO_RES_reg[1]/NET0131 ,
		_w22282_,
		_w22283_,
		_w22284_
	);
	LUT2 #(
		.INIT('h2)
	) name18237 (
		\sice_SPC_reg[7]/P0001 ,
		_w16259_,
		_w22285_
	);
	LUT4 #(
		.INIT('h135f)
	) name18238 (
		\sice_DBR1_reg[2]/P0001 ,
		\sice_IMR1_reg[1]/NET0131 ,
		_w15544_,
		_w21468_,
		_w22286_
	);
	LUT4 #(
		.INIT('h135f)
	) name18239 (
		\sice_ICYC_reg[7]/NET0131 ,
		\sice_IIRC_reg[7]/NET0131 ,
		_w14695_,
		_w15161_,
		_w22287_
	);
	LUT2 #(
		.INIT('h8)
	) name18240 (
		_w22286_,
		_w22287_,
		_w22288_
	);
	LUT4 #(
		.INIT('h135f)
	) name18241 (
		\sice_DBR2_reg[2]/P0001 ,
		\sice_DMR2_reg[1]/NET0131 ,
		_w15508_,
		_w15519_,
		_w22289_
	);
	LUT4 #(
		.INIT('h135f)
	) name18242 (
		\sice_IBR2_reg[1]/P0001 ,
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w15559_,
		_w16507_,
		_w22290_
	);
	LUT4 #(
		.INIT('h153f)
	) name18243 (
		\sice_DMR1_reg[1]/NET0131 ,
		\sice_IMR2_reg[1]/NET0131 ,
		_w15527_,
		_w17158_,
		_w22291_
	);
	LUT4 #(
		.INIT('h135f)
	) name18244 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		\sice_IBR1_reg[1]/P0001 ,
		_w17323_,
		_w21464_,
		_w22292_
	);
	LUT4 #(
		.INIT('h8000)
	) name18245 (
		_w22291_,
		_w22292_,
		_w22289_,
		_w22290_,
		_w22293_
	);
	LUT4 #(
		.INIT('h4000)
	) name18246 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[6]/P0001 ,
		_w22294_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18247 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[8]/P0001 ,
		_w22295_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18248 (
		_w16259_,
		_w21458_,
		_w22294_,
		_w22295_,
		_w22296_
	);
	LUT4 #(
		.INIT('h7f00)
	) name18249 (
		_w21458_,
		_w22288_,
		_w22293_,
		_w22296_,
		_w22297_
	);
	LUT2 #(
		.INIT('he)
	) name18250 (
		_w22285_,
		_w22297_,
		_w22298_
	);
	LUT2 #(
		.INIT('h2)
	) name18251 (
		\sice_SPC_reg[8]/P0001 ,
		_w16259_,
		_w22299_
	);
	LUT4 #(
		.INIT('h135f)
	) name18252 (
		\sice_DBR1_reg[3]/P0001 ,
		\sice_IMR1_reg[2]/NET0131 ,
		_w15544_,
		_w21468_,
		_w22300_
	);
	LUT4 #(
		.INIT('h135f)
	) name18253 (
		\sice_ICYC_reg[8]/NET0131 ,
		\sice_IIRC_reg[8]/NET0131 ,
		_w14695_,
		_w15161_,
		_w22301_
	);
	LUT2 #(
		.INIT('h8)
	) name18254 (
		_w22300_,
		_w22301_,
		_w22302_
	);
	LUT4 #(
		.INIT('h135f)
	) name18255 (
		\sice_DBR2_reg[3]/P0001 ,
		\sice_DMR2_reg[2]/NET0131 ,
		_w15508_,
		_w15519_,
		_w22303_
	);
	LUT4 #(
		.INIT('h135f)
	) name18256 (
		\sice_IBR2_reg[2]/P0001 ,
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w15559_,
		_w16507_,
		_w22304_
	);
	LUT4 #(
		.INIT('h153f)
	) name18257 (
		\sice_DMR1_reg[2]/NET0131 ,
		\sice_IMR2_reg[2]/NET0131 ,
		_w15527_,
		_w17158_,
		_w22305_
	);
	LUT4 #(
		.INIT('h135f)
	) name18258 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\sice_IBR1_reg[2]/P0001 ,
		_w17323_,
		_w21464_,
		_w22306_
	);
	LUT4 #(
		.INIT('h8000)
	) name18259 (
		_w22305_,
		_w22306_,
		_w22303_,
		_w22304_,
		_w22307_
	);
	LUT4 #(
		.INIT('h4000)
	) name18260 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[7]/P0001 ,
		_w22308_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18261 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[9]/P0001 ,
		_w22309_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18262 (
		_w16259_,
		_w21458_,
		_w22308_,
		_w22309_,
		_w22310_
	);
	LUT4 #(
		.INIT('h7f00)
	) name18263 (
		_w21458_,
		_w22302_,
		_w22307_,
		_w22310_,
		_w22311_
	);
	LUT2 #(
		.INIT('he)
	) name18264 (
		_w22299_,
		_w22311_,
		_w22312_
	);
	LUT4 #(
		.INIT('h0c44)
	) name18265 (
		\auctl_DSack_reg/NET0131 ,
		\idma_WRcyc_reg/NET0131 ,
		_w12812_,
		_w19996_,
		_w22313_
	);
	LUT2 #(
		.INIT('he)
	) name18266 (
		_w12814_,
		_w22313_,
		_w22314_
	);
	LUT4 #(
		.INIT('hfc55)
	) name18267 (
		\PIO_out[11]_pad ,
		_w8798_,
		_w8801_,
		_w22257_,
		_w22315_
	);
	LUT3 #(
		.INIT('h4e)
	) name18268 (
		\PIO_oe[11]_pad ,
		\pio_PIO_RES_reg[11]/NET0131 ,
		_w22315_,
		_w22316_
	);
	LUT3 #(
		.INIT('h80)
	) name18269 (
		_w11922_,
		_w11926_,
		_w13447_,
		_w22317_
	);
	LUT4 #(
		.INIT('h2a00)
	) name18270 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w11917_,
		_w11920_,
		_w11924_,
		_w22318_
	);
	LUT4 #(
		.INIT('h31f5)
	) name18271 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w4554_,
		_w11926_,
		_w22318_,
		_w22319_
	);
	LUT2 #(
		.INIT('hb)
	) name18272 (
		_w22317_,
		_w22319_,
		_w22320_
	);
	LUT4 #(
		.INIT('h00ba)
	) name18273 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4084_,
		_w5575_,
		_w22321_
	);
	LUT4 #(
		.INIT('h00b8)
	) name18274 (
		\memc_Dwrite_C_reg/NET0131 ,
		_w4971_,
		_w5571_,
		_w22321_,
		_w22322_
	);
	LUT3 #(
		.INIT('h04)
	) name18275 (
		_w8190_,
		_w8192_,
		_w22322_,
		_w22323_
	);
	LUT4 #(
		.INIT('hff4e)
	) name18276 (
		_w6944_,
		_w8170_,
		_w8465_,
		_w22323_,
		_w22324_
	);
	LUT2 #(
		.INIT('h8)
	) name18277 (
		_w14460_,
		_w21468_,
		_w22325_
	);
	LUT3 #(
		.INIT('h0d)
	) name18278 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w22326_
	);
	LUT3 #(
		.INIT('he2)
	) name18279 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w11926_,
		_w22326_,
		_w22327_
	);
	LUT4 #(
		.INIT('hc444)
	) name18280 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		_w4073_,
		_w4084_,
		_w22328_
	);
	LUT4 #(
		.INIT('h002a)
	) name18281 (
		\core_c_psq_INT_en_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20447_,
		_w22329_
	);
	LUT4 #(
		.INIT('h4000)
	) name18282 (
		_w12270_,
		_w12279_,
		_w20443_,
		_w20440_,
		_w22330_
	);
	LUT3 #(
		.INIT('hea)
	) name18283 (
		_w22328_,
		_w22329_,
		_w22330_,
		_w22331_
	);
	LUT3 #(
		.INIT('h6a)
	) name18284 (
		\clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131 ,
		_w19400_,
		_w19405_,
		_w22332_
	);
	LUT2 #(
		.INIT('h8)
	) name18285 (
		_w14460_,
		_w21464_,
		_w22333_
	);
	LUT4 #(
		.INIT('h0010)
	) name18286 (
		\sport1_txctl_Wcnt_reg[0]/NET0131 ,
		\sport1_txctl_Wcnt_reg[1]/NET0131 ,
		_w14591_,
		_w14594_,
		_w22334_
	);
	LUT4 #(
		.INIT('h0100)
	) name18287 (
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		\sport1_txctl_Wcnt_reg[3]/NET0131 ,
		\sport1_txctl_Wcnt_reg[4]/NET0131 ,
		_w22334_,
		_w22335_
	);
	LUT2 #(
		.INIT('h4)
	) name18288 (
		\sport1_txctl_Wcnt_reg[5]/NET0131 ,
		_w22335_,
		_w22336_
	);
	LUT3 #(
		.INIT('h10)
	) name18289 (
		\sport1_txctl_Wcnt_reg[5]/NET0131 ,
		\sport1_txctl_Wcnt_reg[6]/NET0131 ,
		_w22335_,
		_w22337_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18290 (
		\sport1_regs_MWORDreg_DO_reg[7]/NET0131 ,
		\sport1_txctl_Wcnt_reg[7]/NET0131 ,
		_w14595_,
		_w22337_,
		_w22338_
	);
	LUT2 #(
		.INIT('h9)
	) name18291 (
		\sport1_txctl_Wcnt_reg[5]/NET0131 ,
		_w22335_,
		_w22339_
	);
	LUT3 #(
		.INIT('h8b)
	) name18292 (
		\sport1_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w14595_,
		_w22339_,
		_w22340_
	);
	LUT4 #(
		.INIT('h0010)
	) name18293 (
		\sport0_txctl_Wcnt_reg[0]/NET0131 ,
		\sport0_txctl_Wcnt_reg[1]/NET0131 ,
		_w14597_,
		_w14600_,
		_w22341_
	);
	LUT4 #(
		.INIT('h0100)
	) name18294 (
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		\sport0_txctl_Wcnt_reg[3]/NET0131 ,
		\sport0_txctl_Wcnt_reg[4]/NET0131 ,
		_w22341_,
		_w22342_
	);
	LUT2 #(
		.INIT('h4)
	) name18295 (
		\sport0_txctl_Wcnt_reg[5]/NET0131 ,
		_w22342_,
		_w22343_
	);
	LUT3 #(
		.INIT('h10)
	) name18296 (
		\sport0_txctl_Wcnt_reg[5]/NET0131 ,
		\sport0_txctl_Wcnt_reg[6]/NET0131 ,
		_w22342_,
		_w22344_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18297 (
		\sport0_regs_MWORDreg_DO_reg[7]/NET0131 ,
		\sport0_txctl_Wcnt_reg[7]/NET0131 ,
		_w14601_,
		_w22344_,
		_w22345_
	);
	LUT2 #(
		.INIT('h9)
	) name18298 (
		\sport0_txctl_Wcnt_reg[5]/NET0131 ,
		_w22342_,
		_w22346_
	);
	LUT3 #(
		.INIT('h8b)
	) name18299 (
		\sport0_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w14601_,
		_w22346_,
		_w22347_
	);
	LUT3 #(
		.INIT('h6a)
	) name18300 (
		\idma_WRcnt_reg[2]/NET0131 ,
		_w12811_,
		_w12854_,
		_w22348_
	);
	LUT3 #(
		.INIT('hb8)
	) name18301 (
		\memc_usysr_DO_reg[9]/NET0131 ,
		_w12856_,
		_w22348_,
		_w22349_
	);
	LUT2 #(
		.INIT('h1)
	) name18302 (
		_w13258_,
		_w13259_,
		_w22350_
	);
	LUT3 #(
		.INIT('h13)
	) name18303 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w22351_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name18304 (
		\core_c_dec_RET_Ed_reg/P0001 ,
		_w4160_,
		_w4158_,
		_w4167_,
		_w22352_
	);
	LUT2 #(
		.INIT('h2)
	) name18305 (
		_w22351_,
		_w22352_,
		_w22353_
	);
	LUT3 #(
		.INIT('h23)
	) name18306 (
		_w4507_,
		_w4971_,
		_w22353_,
		_w22354_
	);
	LUT4 #(
		.INIT('h0405)
	) name18307 (
		\core_c_psq_pcstk_ptr_reg[4]/NET0131 ,
		_w4507_,
		_w4971_,
		_w22353_,
		_w22355_
	);
	LUT4 #(
		.INIT('h0001)
	) name18308 (
		\core_c_dec_Call_Ed_reg/P0001 ,
		\core_c_dec_RET_Ed_reg/P0001 ,
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22356_
	);
	LUT3 #(
		.INIT('h80)
	) name18309 (
		_w13257_,
		_w22351_,
		_w22356_,
		_w22357_
	);
	LUT4 #(
		.INIT('hc8ca)
	) name18310 (
		_w4111_,
		_w4109_,
		_w13258_,
		_w13259_,
		_w22358_
	);
	LUT4 #(
		.INIT('hae00)
	) name18311 (
		_w22350_,
		_w22355_,
		_w22357_,
		_w22358_,
		_w22359_
	);
	LUT2 #(
		.INIT('h6)
	) name18312 (
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w22359_,
		_w22360_
	);
	LUT4 #(
		.INIT('h4454)
	) name18313 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		_w22350_,
		_w22355_,
		_w22357_,
		_w22361_
	);
	LUT3 #(
		.INIT('h02)
	) name18314 (
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		_w13258_,
		_w13259_,
		_w22362_
	);
	LUT4 #(
		.INIT('h4445)
	) name18315 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		_w13258_,
		_w13259_,
		_w22363_
	);
	LUT4 #(
		.INIT('haa56)
	) name18316 (
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		_w22361_,
		_w22362_,
		_w22363_,
		_w22364_
	);
	LUT3 #(
		.INIT('ha9)
	) name18317 (
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		_w13258_,
		_w13259_,
		_w22365_
	);
	LUT2 #(
		.INIT('h6)
	) name18318 (
		_w22361_,
		_w22365_,
		_w22366_
	);
	LUT4 #(
		.INIT('h6656)
	) name18319 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		_w22350_,
		_w22355_,
		_w22357_,
		_w22367_
	);
	LUT4 #(
		.INIT('hc444)
	) name18320 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		_w4073_,
		_w4084_,
		_w22368_
	);
	LUT3 #(
		.INIT('h10)
	) name18321 (
		_w20442_,
		_w20444_,
		_w20445_,
		_w22369_
	);
	LUT4 #(
		.INIT('h4000)
	) name18322 (
		_w12270_,
		_w12279_,
		_w20440_,
		_w22369_,
		_w22370_
	);
	LUT3 #(
		.INIT('hec)
	) name18323 (
		_w22329_,
		_w22368_,
		_w22370_,
		_w22371_
	);
	LUT4 #(
		.INIT('hc444)
	) name18324 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		_w4073_,
		_w4084_,
		_w22372_
	);
	LUT4 #(
		.INIT('h135f)
	) name18325 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_Iflag_reg[0]/NET0131 ,
		\core_c_psq_Iflag_reg[6]/NET0131 ,
		_w22373_
	);
	LUT3 #(
		.INIT('h40)
	) name18326 (
		_w12273_,
		_w20448_,
		_w22373_,
		_w22374_
	);
	LUT3 #(
		.INIT('h80)
	) name18327 (
		_w12278_,
		_w20446_,
		_w22374_,
		_w22375_
	);
	LUT4 #(
		.INIT('hf2f0)
	) name18328 (
		_w12271_,
		_w12272_,
		_w22372_,
		_w22375_,
		_w22376_
	);
	LUT2 #(
		.INIT('h8)
	) name18329 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w4106_,
		_w22377_
	);
	LUT4 #(
		.INIT('hff20)
	) name18330 (
		_w14570_,
		_w19715_,
		_w19728_,
		_w22377_,
		_w22378_
	);
	LUT4 #(
		.INIT('h2000)
	) name18331 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22379_
	);
	LUT4 #(
		.INIT('hff80)
	) name18332 (
		_w15936_,
		_w19720_,
		_w21288_,
		_w22379_,
		_w22380_
	);
	LUT4 #(
		.INIT('h2000)
	) name18333 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22381_
	);
	LUT2 #(
		.INIT('h8)
	) name18334 (
		_w19235_,
		_w19719_,
		_w22382_
	);
	LUT3 #(
		.INIT('hec)
	) name18335 (
		_w16161_,
		_w22381_,
		_w22382_,
		_w22383_
	);
	LUT4 #(
		.INIT('h2000)
	) name18336 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22384_
	);
	LUT4 #(
		.INIT('hff80)
	) name18337 (
		_w15936_,
		_w19240_,
		_w21288_,
		_w22384_,
		_w22385_
	);
	LUT4 #(
		.INIT('h2000)
	) name18338 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22386_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18339 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w20967_,
		_w22387_
	);
	LUT3 #(
		.INIT('hec)
	) name18340 (
		_w19233_,
		_w22386_,
		_w22387_,
		_w22388_
	);
	LUT4 #(
		.INIT('h2000)
	) name18341 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22389_
	);
	LUT3 #(
		.INIT('hf8)
	) name18342 (
		_w15933_,
		_w22382_,
		_w22389_,
		_w22390_
	);
	LUT3 #(
		.INIT('hb8)
	) name18343 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		_w4104_,
		_w20493_,
		_w22391_
	);
	LUT4 #(
		.INIT('h2000)
	) name18344 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22392_
	);
	LUT3 #(
		.INIT('hf8)
	) name18345 (
		_w16161_,
		_w20959_,
		_w22392_,
		_w22393_
	);
	LUT4 #(
		.INIT('h2000)
	) name18346 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22394_
	);
	LUT3 #(
		.INIT('hf8)
	) name18347 (
		_w15933_,
		_w20959_,
		_w22394_,
		_w22395_
	);
	LUT4 #(
		.INIT('h2000)
	) name18348 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22396_
	);
	LUT4 #(
		.INIT('hff80)
	) name18349 (
		_w16161_,
		_w19687_,
		_w20956_,
		_w22396_,
		_w22397_
	);
	LUT4 #(
		.INIT('h2000)
	) name18350 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22398_
	);
	LUT3 #(
		.INIT('hf8)
	) name18351 (
		_w20956_,
		_w21952_,
		_w22398_,
		_w22399_
	);
	LUT4 #(
		.INIT('h2000)
	) name18352 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22400_
	);
	LUT3 #(
		.INIT('ha8)
	) name18353 (
		_w5096_,
		_w19231_,
		_w19232_,
		_w22401_
	);
	LUT4 #(
		.INIT('h0002)
	) name18354 (
		_w12156_,
		_w19040_,
		_w19236_,
		_w19237_,
		_w22402_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18355 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22402_,
		_w22403_
	);
	LUT3 #(
		.INIT('hea)
	) name18356 (
		_w22400_,
		_w22401_,
		_w22403_,
		_w22404_
	);
	LUT4 #(
		.INIT('h2000)
	) name18357 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22405_
	);
	LUT4 #(
		.INIT('h0002)
	) name18358 (
		_w12158_,
		_w19040_,
		_w19236_,
		_w19237_,
		_w22406_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18359 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22406_,
		_w22407_
	);
	LUT3 #(
		.INIT('hec)
	) name18360 (
		_w22401_,
		_w22405_,
		_w22407_,
		_w22408_
	);
	LUT4 #(
		.INIT('h2000)
	) name18361 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22409_
	);
	LUT4 #(
		.INIT('h0002)
	) name18362 (
		_w12153_,
		_w19040_,
		_w19236_,
		_w19237_,
		_w22410_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18363 (
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22410_,
		_w22411_
	);
	LUT3 #(
		.INIT('hec)
	) name18364 (
		_w22401_,
		_w22409_,
		_w22411_,
		_w22412_
	);
	LUT4 #(
		.INIT('h2000)
	) name18365 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22413_
	);
	LUT3 #(
		.INIT('h80)
	) name18366 (
		_w12150_,
		_w19681_,
		_w19693_,
		_w22414_
	);
	LUT3 #(
		.INIT('hec)
	) name18367 (
		_w16002_,
		_w22413_,
		_w22414_,
		_w22415_
	);
	LUT4 #(
		.INIT('h2000)
	) name18368 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22416_
	);
	LUT4 #(
		.INIT('hff80)
	) name18369 (
		_w16161_,
		_w19235_,
		_w19687_,
		_w22416_,
		_w22417_
	);
	LUT3 #(
		.INIT('hb8)
	) name18370 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		_w4104_,
		_w20965_,
		_w22418_
	);
	LUT4 #(
		.INIT('h2000)
	) name18371 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22419_
	);
	LUT3 #(
		.INIT('hf8)
	) name18372 (
		_w20952_,
		_w22387_,
		_w22419_,
		_w22420_
	);
	LUT3 #(
		.INIT('hb8)
	) name18373 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		_w4104_,
		_w20962_,
		_w22421_
	);
	LUT4 #(
		.INIT('h2000)
	) name18374 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22422_
	);
	LUT3 #(
		.INIT('hf8)
	) name18375 (
		_w16007_,
		_w20961_,
		_w22422_,
		_w22423_
	);
	LUT3 #(
		.INIT('hb8)
	) name18376 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		_w4104_,
		_w19684_,
		_w22424_
	);
	LUT3 #(
		.INIT('hb8)
	) name18377 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		_w4104_,
		_w19695_,
		_w22425_
	);
	LUT3 #(
		.INIT('hb8)
	) name18378 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		_w4104_,
		_w19692_,
		_w22426_
	);
	LUT4 #(
		.INIT('h2000)
	) name18379 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22427_
	);
	LUT4 #(
		.INIT('hff80)
	) name18380 (
		_w16161_,
		_w19687_,
		_w20954_,
		_w22427_,
		_w22428_
	);
	LUT4 #(
		.INIT('h2000)
	) name18381 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22429_
	);
	LUT3 #(
		.INIT('hf8)
	) name18382 (
		_w20954_,
		_w21952_,
		_w22429_,
		_w22430_
	);
	LUT4 #(
		.INIT('h2000)
	) name18383 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22431_
	);
	LUT4 #(
		.INIT('hff80)
	) name18384 (
		_w16161_,
		_w19687_,
		_w20960_,
		_w22431_,
		_w22432_
	);
	LUT4 #(
		.INIT('h2000)
	) name18385 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22433_
	);
	LUT3 #(
		.INIT('hf8)
	) name18386 (
		_w20960_,
		_w21952_,
		_w22433_,
		_w22434_
	);
	LUT4 #(
		.INIT('h2000)
	) name18387 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22435_
	);
	LUT3 #(
		.INIT('ha8)
	) name18388 (
		_w5098_,
		_w19231_,
		_w19232_,
		_w22436_
	);
	LUT3 #(
		.INIT('hec)
	) name18389 (
		_w22403_,
		_w22435_,
		_w22436_,
		_w22437_
	);
	LUT4 #(
		.INIT('h2000)
	) name18390 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22438_
	);
	LUT3 #(
		.INIT('hf8)
	) name18391 (
		_w22411_,
		_w22436_,
		_w22438_,
		_w22439_
	);
	LUT4 #(
		.INIT('h2000)
	) name18392 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22440_
	);
	LUT3 #(
		.INIT('h80)
	) name18393 (
		_w19234_,
		_w19681_,
		_w19693_,
		_w22441_
	);
	LUT3 #(
		.INIT('hec)
	) name18394 (
		_w15933_,
		_w22440_,
		_w22441_,
		_w22442_
	);
	LUT4 #(
		.INIT('h2000)
	) name18395 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22443_
	);
	LUT4 #(
		.INIT('hff80)
	) name18396 (
		_w15936_,
		_w19688_,
		_w21288_,
		_w22443_,
		_w22444_
	);
	LUT3 #(
		.INIT('hb8)
	) name18397 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		_w4104_,
		_w20494_,
		_w22445_
	);
	LUT3 #(
		.INIT('hb8)
	) name18398 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		_w4104_,
		_w20497_,
		_w22446_
	);
	LUT4 #(
		.INIT('h2000)
	) name18399 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22447_
	);
	LUT3 #(
		.INIT('hf8)
	) name18400 (
		_w19235_,
		_w21952_,
		_w22447_,
		_w22448_
	);
	LUT4 #(
		.INIT('h4500)
	) name18401 (
		_w7257_,
		_w7375_,
		_w7377_,
		_w13032_,
		_w22449_
	);
	LUT4 #(
		.INIT('hff12)
	) name18402 (
		\bdma_BEAD_reg[4]/NET0131 ,
		_w13032_,
		_w20509_,
		_w22449_,
		_w22450_
	);
	LUT4 #(
		.INIT('h060c)
	) name18403 (
		\bdma_BEAD_reg[2]/NET0131 ,
		\bdma_BEAD_reg[3]/NET0131 ,
		_w13032_,
		_w13031_,
		_w22451_
	);
	LUT4 #(
		.INIT('h4500)
	) name18404 (
		_w6054_,
		_w6173_,
		_w6175_,
		_w13032_,
		_w22452_
	);
	LUT2 #(
		.INIT('he)
	) name18405 (
		_w22451_,
		_w22452_,
		_w22453_
	);
	LUT4 #(
		.INIT('h2000)
	) name18406 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22454_
	);
	LUT3 #(
		.INIT('hf8)
	) name18407 (
		_w22407_,
		_w22436_,
		_w22454_,
		_w22455_
	);
	LUT3 #(
		.INIT('h08)
	) name18408 (
		\core_c_psq_pcstk_ptr_reg[4]/NET0131 ,
		_w4114_,
		_w13258_,
		_w22456_
	);
	LUT3 #(
		.INIT('ha8)
	) name18409 (
		_w4115_,
		_w13258_,
		_w13259_,
		_w22457_
	);
	LUT4 #(
		.INIT('h5155)
	) name18410 (
		\core_c_psq_pcstk_ptr_reg[4]/NET0131 ,
		_w22354_,
		_w22357_,
		_w22457_,
		_w22458_
	);
	LUT2 #(
		.INIT('h1)
	) name18411 (
		_w22456_,
		_w22458_,
		_w22459_
	);
	LUT2 #(
		.INIT('h6)
	) name18412 (
		\sice_ICYC_reg[19]/NET0131 ,
		_w13018_,
		_w22460_
	);
	LUT2 #(
		.INIT('h8)
	) name18413 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4106_,
		_w22461_
	);
	LUT3 #(
		.INIT('hf8)
	) name18414 (
		_w14570_,
		_w19721_,
		_w22461_,
		_w22462_
	);
	LUT4 #(
		.INIT('h4000)
	) name18415 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[22]/P0001 ,
		_w22463_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name18416 (
		T_ID_pad,
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w22464_
	);
	LUT3 #(
		.INIT('h01)
	) name18417 (
		_w21458_,
		_w22463_,
		_w22464_,
		_w22465_
	);
	LUT2 #(
		.INIT('h8)
	) name18418 (
		\emc_eRDY_reg/NET0131 ,
		_w21550_,
		_w22466_
	);
	LUT3 #(
		.INIT('h13)
	) name18419 (
		\sice_IMR1_reg[17]/NET0131 ,
		_w15568_,
		_w21468_,
		_w22467_
	);
	LUT4 #(
		.INIT('h135f)
	) name18420 (
		\sice_CMRW_reg/NET0131 ,
		\sice_DMR1_reg[17]/NET0131 ,
		_w14459_,
		_w17158_,
		_w22468_
	);
	LUT3 #(
		.INIT('h40)
	) name18421 (
		_w22466_,
		_w22467_,
		_w22468_,
		_w22469_
	);
	LUT2 #(
		.INIT('h8)
	) name18422 (
		\sice_DMR2_reg[17]/NET0131 ,
		_w15519_,
		_w22470_
	);
	LUT4 #(
		.INIT('h153f)
	) name18423 (
		\sice_IBR1_reg[17]/P0001 ,
		\sice_ICYC_reg[23]/NET0131 ,
		_w14695_,
		_w21464_,
		_w22471_
	);
	LUT2 #(
		.INIT('h4)
	) name18424 (
		_w22470_,
		_w22471_,
		_w22472_
	);
	LUT4 #(
		.INIT('h135f)
	) name18425 (
		\core_c_dec_IR_reg[23]/NET0131 ,
		\sice_IRR_reg[13]/P0001 ,
		_w17323_,
		_w21472_,
		_w22473_
	);
	LUT4 #(
		.INIT('h135f)
	) name18426 (
		\sice_IIRC_reg[23]/NET0131 ,
		\sice_IMR2_reg[17]/NET0131 ,
		_w15161_,
		_w15527_,
		_w22474_
	);
	LUT4 #(
		.INIT('h153f)
	) name18427 (
		\sice_DBR1_reg[18]/P0001 ,
		\sice_DBR2_reg[18]/P0001 ,
		_w15508_,
		_w15544_,
		_w22475_
	);
	LUT4 #(
		.INIT('h135f)
	) name18428 (
		\sice_IBR2_reg[17]/P0001 ,
		\sice_idr1_reg_DO_reg[11]/P0001 ,
		_w15559_,
		_w16507_,
		_w22476_
	);
	LUT4 #(
		.INIT('h8000)
	) name18429 (
		_w22475_,
		_w22476_,
		_w22473_,
		_w22474_,
		_w22477_
	);
	LUT4 #(
		.INIT('h8000)
	) name18430 (
		_w21458_,
		_w22472_,
		_w22469_,
		_w22477_,
		_w22478_
	);
	LUT2 #(
		.INIT('h1)
	) name18431 (
		_w22465_,
		_w22478_,
		_w22479_
	);
	LUT4 #(
		.INIT('h4000)
	) name18432 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[21]/P0001 ,
		_w22480_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18433 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[23]/P0001 ,
		_w22481_
	);
	LUT3 #(
		.INIT('h01)
	) name18434 (
		_w21458_,
		_w22480_,
		_w22481_,
		_w22482_
	);
	LUT2 #(
		.INIT('h8)
	) name18435 (
		\sice_IDONE_reg/NET0131 ,
		_w21550_,
		_w22483_
	);
	LUT3 #(
		.INIT('h13)
	) name18436 (
		\sice_IMR1_reg[16]/NET0131 ,
		_w15568_,
		_w21468_,
		_w22484_
	);
	LUT4 #(
		.INIT('h153f)
	) name18437 (
		\sice_DMR1_reg[16]/NET0131 ,
		\sice_IIRC_reg[22]/NET0131 ,
		_w15161_,
		_w17158_,
		_w22485_
	);
	LUT3 #(
		.INIT('h40)
	) name18438 (
		_w22483_,
		_w22484_,
		_w22485_,
		_w22486_
	);
	LUT2 #(
		.INIT('h8)
	) name18439 (
		\sice_DMR2_reg[16]/NET0131 ,
		_w15519_,
		_w22487_
	);
	LUT4 #(
		.INIT('h153f)
	) name18440 (
		\sice_IBR1_reg[16]/P0001 ,
		\sice_IBR2_reg[16]/P0001 ,
		_w15559_,
		_w21464_,
		_w22488_
	);
	LUT2 #(
		.INIT('h4)
	) name18441 (
		_w22487_,
		_w22488_,
		_w22489_
	);
	LUT4 #(
		.INIT('h135f)
	) name18442 (
		\core_c_dec_IR_reg[22]/NET0131 ,
		\sice_IRR_reg[12]/P0001 ,
		_w17323_,
		_w21472_,
		_w22490_
	);
	LUT4 #(
		.INIT('h135f)
	) name18443 (
		\sice_ICYC_reg[22]/NET0131 ,
		\sice_IMR2_reg[16]/NET0131 ,
		_w14695_,
		_w15527_,
		_w22491_
	);
	LUT4 #(
		.INIT('h153f)
	) name18444 (
		\sice_DBR1_reg[17]/P0001 ,
		\sice_DBR2_reg[17]/P0001 ,
		_w15508_,
		_w15544_,
		_w22492_
	);
	LUT4 #(
		.INIT('h135f)
	) name18445 (
		\sice_CLR_M_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[10]/P0001 ,
		_w14459_,
		_w16507_,
		_w22493_
	);
	LUT4 #(
		.INIT('h8000)
	) name18446 (
		_w22492_,
		_w22493_,
		_w22490_,
		_w22491_,
		_w22494_
	);
	LUT4 #(
		.INIT('h8000)
	) name18447 (
		_w21458_,
		_w22489_,
		_w22486_,
		_w22494_,
		_w22495_
	);
	LUT2 #(
		.INIT('h1)
	) name18448 (
		_w22482_,
		_w22495_,
		_w22496_
	);
	LUT4 #(
		.INIT('h4000)
	) name18449 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[19]/P0001 ,
		_w22497_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18450 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[21]/P0001 ,
		_w22498_
	);
	LUT3 #(
		.INIT('h01)
	) name18451 (
		_w21458_,
		_w22497_,
		_w22498_,
		_w22499_
	);
	LUT2 #(
		.INIT('h4)
	) name18452 (
		_w4069_,
		_w21550_,
		_w22500_
	);
	LUT3 #(
		.INIT('h13)
	) name18453 (
		\sice_IMR1_reg[14]/NET0131 ,
		_w15568_,
		_w21468_,
		_w22501_
	);
	LUT4 #(
		.INIT('h153f)
	) name18454 (
		\sice_DMR1_reg[14]/NET0131 ,
		\sice_IIRC_reg[20]/NET0131 ,
		_w15161_,
		_w17158_,
		_w22502_
	);
	LUT3 #(
		.INIT('h40)
	) name18455 (
		_w22500_,
		_w22501_,
		_w22502_,
		_w22503_
	);
	LUT2 #(
		.INIT('h8)
	) name18456 (
		\sice_DMR2_reg[14]/NET0131 ,
		_w15519_,
		_w22504_
	);
	LUT4 #(
		.INIT('h153f)
	) name18457 (
		\sice_IBR1_reg[14]/P0001 ,
		\sice_IBR2_reg[14]/P0001 ,
		_w15559_,
		_w21464_,
		_w22505_
	);
	LUT2 #(
		.INIT('h4)
	) name18458 (
		_w22504_,
		_w22505_,
		_w22506_
	);
	LUT4 #(
		.INIT('h135f)
	) name18459 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\sice_IRR_reg[10]/P0001 ,
		_w17323_,
		_w21472_,
		_w22507_
	);
	LUT4 #(
		.INIT('h135f)
	) name18460 (
		\sice_ICYC_reg[20]/NET0131 ,
		\sice_IMR2_reg[14]/NET0131 ,
		_w14695_,
		_w15527_,
		_w22508_
	);
	LUT4 #(
		.INIT('h153f)
	) name18461 (
		\sice_DBR1_reg[15]/P0001 ,
		\sice_DBR2_reg[15]/P0001 ,
		_w15508_,
		_w15544_,
		_w22509_
	);
	LUT4 #(
		.INIT('h135f)
	) name18462 (
		\sice_GO_NX_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[8]/P0001 ,
		_w14459_,
		_w16507_,
		_w22510_
	);
	LUT4 #(
		.INIT('h8000)
	) name18463 (
		_w22509_,
		_w22510_,
		_w22507_,
		_w22508_,
		_w22511_
	);
	LUT4 #(
		.INIT('h8000)
	) name18464 (
		_w21458_,
		_w22506_,
		_w22503_,
		_w22511_,
		_w22512_
	);
	LUT2 #(
		.INIT('h1)
	) name18465 (
		_w22499_,
		_w22512_,
		_w22513_
	);
	LUT4 #(
		.INIT('h4000)
	) name18466 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[18]/P0001 ,
		_w22514_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18467 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[20]/P0001 ,
		_w22515_
	);
	LUT3 #(
		.INIT('h01)
	) name18468 (
		_w21458_,
		_w22514_,
		_w22515_,
		_w22516_
	);
	LUT2 #(
		.INIT('h8)
	) name18469 (
		\core_c_psq_MGNT_reg/NET0131 ,
		_w21550_,
		_w22517_
	);
	LUT3 #(
		.INIT('h13)
	) name18470 (
		\sice_IMR1_reg[13]/NET0131 ,
		_w15568_,
		_w21468_,
		_w22518_
	);
	LUT4 #(
		.INIT('h153f)
	) name18471 (
		\sice_DMR1_reg[13]/NET0131 ,
		\sice_IIRC_reg[19]/NET0131 ,
		_w15161_,
		_w17158_,
		_w22519_
	);
	LUT3 #(
		.INIT('h40)
	) name18472 (
		_w22517_,
		_w22518_,
		_w22519_,
		_w22520_
	);
	LUT2 #(
		.INIT('h8)
	) name18473 (
		\sice_DMR2_reg[13]/NET0131 ,
		_w15519_,
		_w22521_
	);
	LUT4 #(
		.INIT('h153f)
	) name18474 (
		\sice_IBR1_reg[13]/P0001 ,
		\sice_IBR2_reg[13]/P0001 ,
		_w15559_,
		_w21464_,
		_w22522_
	);
	LUT2 #(
		.INIT('h4)
	) name18475 (
		_w22521_,
		_w22522_,
		_w22523_
	);
	LUT4 #(
		.INIT('h135f)
	) name18476 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		\sice_IRR_reg[9]/P0001 ,
		_w17323_,
		_w21472_,
		_w22524_
	);
	LUT4 #(
		.INIT('h135f)
	) name18477 (
		\sice_ICYC_reg[19]/NET0131 ,
		\sice_IMR2_reg[13]/NET0131 ,
		_w14695_,
		_w15527_,
		_w22525_
	);
	LUT4 #(
		.INIT('h153f)
	) name18478 (
		\sice_DBR1_reg[14]/P0001 ,
		\sice_DBR2_reg[14]/P0001 ,
		_w15508_,
		_w15544_,
		_w22526_
	);
	LUT4 #(
		.INIT('h45cf)
	) name18479 (
		\sice_idr1_reg_DO_reg[7]/P0001 ,
		_w14453_,
		_w14459_,
		_w16507_,
		_w22527_
	);
	LUT4 #(
		.INIT('h8000)
	) name18480 (
		_w22526_,
		_w22527_,
		_w22524_,
		_w22525_,
		_w22528_
	);
	LUT4 #(
		.INIT('h8000)
	) name18481 (
		_w21458_,
		_w22523_,
		_w22520_,
		_w22528_,
		_w22529_
	);
	LUT2 #(
		.INIT('h1)
	) name18482 (
		_w22516_,
		_w22529_,
		_w22530_
	);
	LUT4 #(
		.INIT('h4000)
	) name18483 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[17]/P0001 ,
		_w22531_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18484 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[19]/P0001 ,
		_w22532_
	);
	LUT3 #(
		.INIT('h01)
	) name18485 (
		_w21458_,
		_w22531_,
		_w22532_,
		_w22533_
	);
	LUT2 #(
		.INIT('h8)
	) name18486 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w21550_,
		_w22534_
	);
	LUT3 #(
		.INIT('h13)
	) name18487 (
		\sice_IMR1_reg[12]/NET0131 ,
		_w15568_,
		_w21468_,
		_w22535_
	);
	LUT4 #(
		.INIT('h153f)
	) name18488 (
		\sice_DMR1_reg[12]/NET0131 ,
		\sice_IIRC_reg[18]/NET0131 ,
		_w15161_,
		_w17158_,
		_w22536_
	);
	LUT3 #(
		.INIT('h40)
	) name18489 (
		_w22534_,
		_w22535_,
		_w22536_,
		_w22537_
	);
	LUT2 #(
		.INIT('h8)
	) name18490 (
		\sice_DMR2_reg[12]/NET0131 ,
		_w15519_,
		_w22538_
	);
	LUT4 #(
		.INIT('h153f)
	) name18491 (
		\sice_IBR1_reg[12]/P0001 ,
		\sice_IBR2_reg[12]/P0001 ,
		_w15559_,
		_w21464_,
		_w22539_
	);
	LUT2 #(
		.INIT('h4)
	) name18492 (
		_w22538_,
		_w22539_,
		_w22540_
	);
	LUT4 #(
		.INIT('h135f)
	) name18493 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\sice_IRR_reg[8]/P0001 ,
		_w17323_,
		_w21472_,
		_w22541_
	);
	LUT4 #(
		.INIT('h135f)
	) name18494 (
		\sice_ICYC_reg[18]/NET0131 ,
		\sice_IMR2_reg[12]/NET0131 ,
		_w14695_,
		_w15527_,
		_w22542_
	);
	LUT4 #(
		.INIT('h153f)
	) name18495 (
		\sice_DBR1_reg[13]/P0001 ,
		\sice_DBR2_reg[13]/P0001 ,
		_w15508_,
		_w15544_,
		_w22543_
	);
	LUT4 #(
		.INIT('h135f)
	) name18496 (
		\sice_IRST_reg/NET0131 ,
		\sice_idr1_reg_DO_reg[6]/P0001 ,
		_w14459_,
		_w16507_,
		_w22544_
	);
	LUT4 #(
		.INIT('h8000)
	) name18497 (
		_w22543_,
		_w22544_,
		_w22541_,
		_w22542_,
		_w22545_
	);
	LUT4 #(
		.INIT('h8000)
	) name18498 (
		_w21458_,
		_w22540_,
		_w22537_,
		_w22545_,
		_w22546_
	);
	LUT2 #(
		.INIT('h1)
	) name18499 (
		_w22533_,
		_w22546_,
		_w22547_
	);
	LUT4 #(
		.INIT('h2000)
	) name18500 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22548_
	);
	LUT3 #(
		.INIT('hf8)
	) name18501 (
		_w19474_,
		_w21952_,
		_w22548_,
		_w22549_
	);
	LUT3 #(
		.INIT('hb8)
	) name18502 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		_w4104_,
		_w19686_,
		_w22550_
	);
	LUT4 #(
		.INIT('h2000)
	) name18503 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\sice_GO_NX_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w22551_
	);
	LUT4 #(
		.INIT('hff80)
	) name18504 (
		_w16161_,
		_w19687_,
		_w21951_,
		_w22551_,
		_w22552_
	);
	LUT4 #(
		.INIT('h4000)
	) name18505 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[12]/P0001 ,
		_w22553_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18506 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[14]/P0001 ,
		_w22554_
	);
	LUT3 #(
		.INIT('h01)
	) name18507 (
		_w21458_,
		_w22553_,
		_w22554_,
		_w22555_
	);
	LUT3 #(
		.INIT('h07)
	) name18508 (
		\sice_IMR2_reg[7]/NET0131 ,
		_w15527_,
		_w15567_,
		_w22556_
	);
	LUT4 #(
		.INIT('h135f)
	) name18509 (
		\sice_IBR1_reg[7]/P0001 ,
		\sice_IRR_reg[3]/P0001 ,
		_w21464_,
		_w21472_,
		_w22557_
	);
	LUT4 #(
		.INIT('h153f)
	) name18510 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\sice_IBR2_reg[7]/P0001 ,
		_w15559_,
		_w17323_,
		_w22558_
	);
	LUT3 #(
		.INIT('h80)
	) name18511 (
		_w22556_,
		_w22557_,
		_w22558_,
		_w22559_
	);
	LUT4 #(
		.INIT('h153f)
	) name18512 (
		\sice_DBR1_reg[8]/P0001 ,
		\sice_DBR2_reg[8]/P0001 ,
		_w15508_,
		_w15544_,
		_w22560_
	);
	LUT4 #(
		.INIT('h135f)
	) name18513 (
		\sice_IIRC_reg[13]/NET0131 ,
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w15161_,
		_w16507_,
		_w22561_
	);
	LUT4 #(
		.INIT('h153f)
	) name18514 (
		\sice_DMR2_reg[7]/NET0131 ,
		\sice_ICYC_reg[13]/NET0131 ,
		_w14695_,
		_w15519_,
		_w22562_
	);
	LUT4 #(
		.INIT('h135f)
	) name18515 (
		\sice_DMR1_reg[7]/NET0131 ,
		\sice_IMR1_reg[7]/NET0131 ,
		_w17158_,
		_w21468_,
		_w22563_
	);
	LUT4 #(
		.INIT('h8000)
	) name18516 (
		_w22562_,
		_w22563_,
		_w22560_,
		_w22561_,
		_w22564_
	);
	LUT4 #(
		.INIT('h1333)
	) name18517 (
		_w21458_,
		_w22555_,
		_w22559_,
		_w22564_,
		_w22565_
	);
	LUT4 #(
		.INIT('h4000)
	) name18518 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[13]/P0001 ,
		_w22566_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18519 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[15]/P0001 ,
		_w22567_
	);
	LUT3 #(
		.INIT('h01)
	) name18520 (
		_w21458_,
		_w22566_,
		_w22567_,
		_w22568_
	);
	LUT3 #(
		.INIT('h07)
	) name18521 (
		\sice_DBR1_reg[9]/P0001 ,
		_w15544_,
		_w15567_,
		_w22569_
	);
	LUT4 #(
		.INIT('h135f)
	) name18522 (
		\sice_IMR2_reg[8]/NET0131 ,
		\sice_IRR_reg[4]/P0001 ,
		_w15527_,
		_w21472_,
		_w22570_
	);
	LUT4 #(
		.INIT('h153f)
	) name18523 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		\sice_IBR2_reg[8]/P0001 ,
		_w15559_,
		_w17323_,
		_w22571_
	);
	LUT3 #(
		.INIT('h80)
	) name18524 (
		_w22569_,
		_w22570_,
		_w22571_,
		_w22572_
	);
	LUT4 #(
		.INIT('h153f)
	) name18525 (
		\sice_DBR2_reg[9]/P0001 ,
		\sice_IIRC_reg[14]/NET0131 ,
		_w15161_,
		_w15508_,
		_w22573_
	);
	LUT4 #(
		.INIT('h153f)
	) name18526 (
		\sice_DMR1_reg[8]/NET0131 ,
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w16507_,
		_w17158_,
		_w22574_
	);
	LUT4 #(
		.INIT('h153f)
	) name18527 (
		\sice_DMR2_reg[8]/NET0131 ,
		\sice_ICYC_reg[14]/NET0131 ,
		_w14695_,
		_w15519_,
		_w22575_
	);
	LUT4 #(
		.INIT('h135f)
	) name18528 (
		\sice_IBR1_reg[8]/P0001 ,
		\sice_IMR1_reg[8]/NET0131 ,
		_w21464_,
		_w21468_,
		_w22576_
	);
	LUT4 #(
		.INIT('h8000)
	) name18529 (
		_w22575_,
		_w22576_,
		_w22573_,
		_w22574_,
		_w22577_
	);
	LUT4 #(
		.INIT('h1333)
	) name18530 (
		_w21458_,
		_w22568_,
		_w22572_,
		_w22577_,
		_w22578_
	);
	LUT4 #(
		.INIT('h4000)
	) name18531 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[14]/P0001 ,
		_w22579_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18532 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[16]/P0001 ,
		_w22580_
	);
	LUT3 #(
		.INIT('h01)
	) name18533 (
		_w21458_,
		_w22579_,
		_w22580_,
		_w22581_
	);
	LUT3 #(
		.INIT('h07)
	) name18534 (
		\sice_DBR1_reg[10]/P0001 ,
		_w15544_,
		_w15567_,
		_w22582_
	);
	LUT4 #(
		.INIT('h135f)
	) name18535 (
		\sice_IMR2_reg[9]/NET0131 ,
		\sice_IRR_reg[5]/P0001 ,
		_w15527_,
		_w21472_,
		_w22583_
	);
	LUT4 #(
		.INIT('h153f)
	) name18536 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\sice_IBR2_reg[9]/P0001 ,
		_w15559_,
		_w17323_,
		_w22584_
	);
	LUT3 #(
		.INIT('h80)
	) name18537 (
		_w22582_,
		_w22583_,
		_w22584_,
		_w22585_
	);
	LUT4 #(
		.INIT('h153f)
	) name18538 (
		\sice_DBR2_reg[10]/P0001 ,
		\sice_IIRC_reg[15]/NET0131 ,
		_w15161_,
		_w15508_,
		_w22586_
	);
	LUT4 #(
		.INIT('h153f)
	) name18539 (
		\sice_DMR1_reg[9]/NET0131 ,
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w16507_,
		_w17158_,
		_w22587_
	);
	LUT4 #(
		.INIT('h153f)
	) name18540 (
		\sice_DMR2_reg[9]/NET0131 ,
		\sice_ICYC_reg[15]/NET0131 ,
		_w14695_,
		_w15519_,
		_w22588_
	);
	LUT4 #(
		.INIT('h135f)
	) name18541 (
		\sice_IBR1_reg[9]/P0001 ,
		\sice_IMR1_reg[9]/NET0131 ,
		_w21464_,
		_w21468_,
		_w22589_
	);
	LUT4 #(
		.INIT('h8000)
	) name18542 (
		_w22588_,
		_w22589_,
		_w22586_,
		_w22587_,
		_w22590_
	);
	LUT4 #(
		.INIT('h1333)
	) name18543 (
		_w21458_,
		_w22581_,
		_w22585_,
		_w22590_,
		_w22591_
	);
	LUT3 #(
		.INIT('h6c)
	) name18544 (
		\sice_ICYC_reg[10]/NET0131 ,
		\sice_ICYC_reg[11]/NET0131 ,
		_w13015_,
		_w22592_
	);
	LUT3 #(
		.INIT('h6c)
	) name18545 (
		\sice_IIRC_reg[10]/NET0131 ,
		\sice_IIRC_reg[11]/NET0131 ,
		_w13087_,
		_w22593_
	);
	LUT4 #(
		.INIT('h4000)
	) name18546 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[16]/P0001 ,
		_w22594_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18547 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[18]/P0001 ,
		_w22595_
	);
	LUT3 #(
		.INIT('h01)
	) name18548 (
		_w21458_,
		_w22594_,
		_w22595_,
		_w22596_
	);
	LUT3 #(
		.INIT('h07)
	) name18549 (
		\sice_DBR1_reg[12]/P0001 ,
		_w15544_,
		_w15567_,
		_w22597_
	);
	LUT4 #(
		.INIT('h135f)
	) name18550 (
		\sice_IMR2_reg[11]/NET0131 ,
		\sice_IRR_reg[7]/P0001 ,
		_w15527_,
		_w21472_,
		_w22598_
	);
	LUT4 #(
		.INIT('h135f)
	) name18551 (
		\sice_IBR2_reg[11]/P0001 ,
		\sice_idr1_reg_DO_reg[5]/P0001 ,
		_w15559_,
		_w16507_,
		_w22599_
	);
	LUT3 #(
		.INIT('h80)
	) name18552 (
		_w22597_,
		_w22598_,
		_w22599_,
		_w22600_
	);
	LUT4 #(
		.INIT('h153f)
	) name18553 (
		\sice_DBR2_reg[12]/P0001 ,
		\sice_IIRC_reg[17]/NET0131 ,
		_w15161_,
		_w15508_,
		_w22601_
	);
	LUT4 #(
		.INIT('h153f)
	) name18554 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		\sice_DMR1_reg[11]/NET0131 ,
		_w17158_,
		_w17323_,
		_w22602_
	);
	LUT4 #(
		.INIT('h153f)
	) name18555 (
		\sice_DMR2_reg[11]/NET0131 ,
		\sice_ICYC_reg[17]/NET0131 ,
		_w14695_,
		_w15519_,
		_w22603_
	);
	LUT4 #(
		.INIT('h135f)
	) name18556 (
		\sice_IBR1_reg[11]/P0001 ,
		\sice_IMR1_reg[11]/NET0131 ,
		_w21464_,
		_w21468_,
		_w22604_
	);
	LUT4 #(
		.INIT('h8000)
	) name18557 (
		_w22603_,
		_w22604_,
		_w22601_,
		_w22602_,
		_w22605_
	);
	LUT4 #(
		.INIT('h1333)
	) name18558 (
		_w21458_,
		_w22596_,
		_w22600_,
		_w22605_,
		_w22606_
	);
	LUT4 #(
		.INIT('h2220)
	) name18559 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\memc_Dread_E_reg/NET0131 ,
		\memc_Dwrite_E_reg/NET0131 ,
		_w22607_
	);
	LUT2 #(
		.INIT('h4)
	) name18560 (
		_w4069_,
		_w22607_,
		_w22608_
	);
	LUT3 #(
		.INIT('ha2)
	) name18561 (
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w9936_,
		_w22609_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name18562 (
		_w12058_,
		_w12060_,
		_w22608_,
		_w22609_,
		_w22610_
	);
	LUT4 #(
		.INIT('h4000)
	) name18563 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[15]/P0001 ,
		_w22611_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18564 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[17]/P0001 ,
		_w22612_
	);
	LUT3 #(
		.INIT('h01)
	) name18565 (
		_w21458_,
		_w22611_,
		_w22612_,
		_w22613_
	);
	LUT3 #(
		.INIT('h07)
	) name18566 (
		\sice_DBR1_reg[11]/P0001 ,
		_w15544_,
		_w15567_,
		_w22614_
	);
	LUT4 #(
		.INIT('h135f)
	) name18567 (
		\sice_IMR2_reg[10]/NET0131 ,
		\sice_IRR_reg[6]/P0001 ,
		_w15527_,
		_w21472_,
		_w22615_
	);
	LUT4 #(
		.INIT('h135f)
	) name18568 (
		\sice_IBR2_reg[10]/P0001 ,
		\sice_idr1_reg_DO_reg[4]/P0001 ,
		_w15559_,
		_w16507_,
		_w22616_
	);
	LUT3 #(
		.INIT('h80)
	) name18569 (
		_w22614_,
		_w22615_,
		_w22616_,
		_w22617_
	);
	LUT4 #(
		.INIT('h153f)
	) name18570 (
		\sice_DBR2_reg[11]/P0001 ,
		\sice_IIRC_reg[16]/NET0131 ,
		_w15161_,
		_w15508_,
		_w22618_
	);
	LUT4 #(
		.INIT('h153f)
	) name18571 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\sice_DMR1_reg[10]/NET0131 ,
		_w17158_,
		_w17323_,
		_w22619_
	);
	LUT4 #(
		.INIT('h153f)
	) name18572 (
		\sice_DMR2_reg[10]/NET0131 ,
		\sice_ICYC_reg[16]/NET0131 ,
		_w14695_,
		_w15519_,
		_w22620_
	);
	LUT4 #(
		.INIT('h135f)
	) name18573 (
		\sice_IBR1_reg[10]/P0001 ,
		\sice_IMR1_reg[10]/NET0131 ,
		_w21464_,
		_w21468_,
		_w22621_
	);
	LUT4 #(
		.INIT('h8000)
	) name18574 (
		_w22620_,
		_w22621_,
		_w22618_,
		_w22619_,
		_w22622_
	);
	LUT4 #(
		.INIT('h1333)
	) name18575 (
		_w21458_,
		_w22613_,
		_w22617_,
		_w22622_,
		_w22623_
	);
	LUT2 #(
		.INIT('h2)
	) name18576 (
		\sice_SPC_reg[4]/P0001 ,
		_w16259_,
		_w22624_
	);
	LUT4 #(
		.INIT('h153f)
	) name18577 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w16507_,
		_w17323_,
		_w22625_
	);
	LUT4 #(
		.INIT('h135f)
	) name18578 (
		\sice_ICYC_reg[4]/NET0131 ,
		\sice_IIRC_reg[4]/NET0131 ,
		_w14695_,
		_w15161_,
		_w22626_
	);
	LUT4 #(
		.INIT('h4000)
	) name18579 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[3]/P0001 ,
		_w22627_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18580 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[5]/P0001 ,
		_w22628_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18581 (
		_w16259_,
		_w21458_,
		_w22627_,
		_w22628_,
		_w22629_
	);
	LUT4 #(
		.INIT('h7f00)
	) name18582 (
		_w21458_,
		_w22625_,
		_w22626_,
		_w22629_,
		_w22630_
	);
	LUT2 #(
		.INIT('he)
	) name18583 (
		_w22624_,
		_w22630_,
		_w22631_
	);
	LUT2 #(
		.INIT('h2)
	) name18584 (
		\sice_SPC_reg[3]/P0001 ,
		_w16259_,
		_w22632_
	);
	LUT4 #(
		.INIT('h153f)
	) name18585 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w16507_,
		_w17323_,
		_w22633_
	);
	LUT4 #(
		.INIT('h135f)
	) name18586 (
		\sice_ICYC_reg[3]/NET0131 ,
		\sice_IIRC_reg[3]/NET0131 ,
		_w14695_,
		_w15161_,
		_w22634_
	);
	LUT4 #(
		.INIT('h4000)
	) name18587 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[2]/P0001 ,
		_w22635_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18588 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[4]/P0001 ,
		_w22636_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18589 (
		_w16259_,
		_w21458_,
		_w22635_,
		_w22636_,
		_w22637_
	);
	LUT4 #(
		.INIT('h7f00)
	) name18590 (
		_w21458_,
		_w22633_,
		_w22634_,
		_w22637_,
		_w22638_
	);
	LUT2 #(
		.INIT('he)
	) name18591 (
		_w22632_,
		_w22638_,
		_w22639_
	);
	LUT2 #(
		.INIT('h2)
	) name18592 (
		\sice_SPC_reg[2]/P0001 ,
		_w16259_,
		_w22640_
	);
	LUT4 #(
		.INIT('h153f)
	) name18593 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w16507_,
		_w17323_,
		_w22641_
	);
	LUT4 #(
		.INIT('h135f)
	) name18594 (
		\sice_ICYC_reg[2]/NET0131 ,
		\sice_IIRC_reg[2]/NET0131 ,
		_w14695_,
		_w15161_,
		_w22642_
	);
	LUT4 #(
		.INIT('h4000)
	) name18595 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[1]/P0001 ,
		_w22643_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18596 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[3]/P0001 ,
		_w22644_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18597 (
		_w16259_,
		_w21458_,
		_w22643_,
		_w22644_,
		_w22645_
	);
	LUT4 #(
		.INIT('h7f00)
	) name18598 (
		_w21458_,
		_w22641_,
		_w22642_,
		_w22645_,
		_w22646_
	);
	LUT2 #(
		.INIT('he)
	) name18599 (
		_w22640_,
		_w22646_,
		_w22647_
	);
	LUT2 #(
		.INIT('h2)
	) name18600 (
		\sice_SPC_reg[1]/P0001 ,
		_w16259_,
		_w22648_
	);
	LUT4 #(
		.INIT('h153f)
	) name18601 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w16507_,
		_w17323_,
		_w22649_
	);
	LUT4 #(
		.INIT('h135f)
	) name18602 (
		\sice_ICYC_reg[1]/NET0131 ,
		\sice_IIRC_reg[1]/NET0131 ,
		_w14695_,
		_w15161_,
		_w22650_
	);
	LUT4 #(
		.INIT('h4000)
	) name18603 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[0]/P0001 ,
		_w22651_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18604 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		\sice_SPC_reg[2]/P0001 ,
		_w22652_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18605 (
		_w16259_,
		_w21458_,
		_w22651_,
		_w22652_,
		_w22653_
	);
	LUT4 #(
		.INIT('h7f00)
	) name18606 (
		_w21458_,
		_w22649_,
		_w22650_,
		_w22653_,
		_w22654_
	);
	LUT2 #(
		.INIT('he)
	) name18607 (
		_w22648_,
		_w22654_,
		_w22655_
	);
	LUT4 #(
		.INIT('h048c)
	) name18608 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w9946_,
		_w11294_,
		_w15552_,
		_w22656_
	);
	LUT3 #(
		.INIT('h13)
	) name18609 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001 ,
		_w11300_,
		_w22657_
	);
	LUT4 #(
		.INIT('hccc8)
	) name18610 (
		_w11310_,
		_w11312_,
		_w13610_,
		_w13611_,
		_w22658_
	);
	LUT4 #(
		.INIT('h2322)
	) name18611 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001 ,
		_w11303_,
		_w11308_,
		_w22659_
	);
	LUT4 #(
		.INIT('h00ab)
	) name18612 (
		_w11320_,
		_w22657_,
		_w22658_,
		_w22659_,
		_w22660_
	);
	LUT2 #(
		.INIT('h2)
	) name18613 (
		_w11325_,
		_w22660_,
		_w22661_
	);
	LUT2 #(
		.INIT('h1)
	) name18614 (
		_w22656_,
		_w22661_,
		_w22662_
	);
	LUT3 #(
		.INIT('h15)
	) name18615 (
		\clkc_STDcnt_reg[0]/NET0131 ,
		_w19400_,
		_w19405_,
		_w22663_
	);
	LUT3 #(
		.INIT('h12)
	) name18616 (
		\clkc_STDcnt_reg[9]/NET0131 ,
		_w19406_,
		_w19395_,
		_w22664_
	);
	LUT3 #(
		.INIT('hb4)
	) name18617 (
		_w13147_,
		_w13152_,
		_w21175_,
		_w22665_
	);
	LUT4 #(
		.INIT('hea00)
	) name18618 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w19091_,
		_w19096_,
		_w22665_,
		_w22666_
	);
	LUT4 #(
		.INIT('h0015)
	) name18619 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w19091_,
		_w19096_,
		_w22665_,
		_w22667_
	);
	LUT3 #(
		.INIT('h02)
	) name18620 (
		_w13155_,
		_w22667_,
		_w22666_,
		_w22668_
	);
	LUT4 #(
		.INIT('h1011)
	) name18621 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w7793_,
		_w7903_,
		_w7905_,
		_w22669_
	);
	LUT3 #(
		.INIT('h40)
	) name18622 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[7]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w22670_
	);
	LUT2 #(
		.INIT('h1)
	) name18623 (
		_w13158_,
		_w22670_,
		_w22671_
	);
	LUT4 #(
		.INIT('hafac)
	) name18624 (
		\sport0_rxctl_RXSHT_reg[7]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w22672_
	);
	LUT4 #(
		.INIT('hef00)
	) name18625 (
		_w22668_,
		_w22669_,
		_w22671_,
		_w22672_,
		_w22673_
	);
	LUT4 #(
		.INIT('h0002)
	) name18626 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w22674_
	);
	LUT2 #(
		.INIT('he)
	) name18627 (
		_w22673_,
		_w22674_,
		_w22675_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18628 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11830_,
		_w12738_,
		_w17826_,
		_w22676_
	);
	LUT4 #(
		.INIT('h5545)
	) name18629 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w22677_
	);
	LUT2 #(
		.INIT('h1)
	) name18630 (
		_w22676_,
		_w22677_,
		_w22678_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18631 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11830_,
		_w12317_,
		_w18799_,
		_w22679_
	);
	LUT4 #(
		.INIT('h5545)
	) name18632 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001 ,
		_w9453_,
		_w9894_,
		_w11328_,
		_w22680_
	);
	LUT2 #(
		.INIT('h1)
	) name18633 (
		_w22679_,
		_w22680_,
		_w22681_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18634 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11329_,
		_w12317_,
		_w18799_,
		_w22682_
	);
	LUT2 #(
		.INIT('h1)
	) name18635 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001 ,
		_w11329_,
		_w22683_
	);
	LUT2 #(
		.INIT('h1)
	) name18636 (
		_w22682_,
		_w22683_,
		_w22684_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18637 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w11946_,
		_w14949_,
		_w18477_,
		_w22685_
	);
	LUT4 #(
		.INIT('h5545)
	) name18638 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001 ,
		_w9453_,
		_w9894_,
		_w11945_,
		_w22686_
	);
	LUT2 #(
		.INIT('h1)
	) name18639 (
		_w22685_,
		_w22686_,
		_w22687_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18640 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12048_,
		_w14949_,
		_w18477_,
		_w22688_
	);
	LUT2 #(
		.INIT('h1)
	) name18641 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001 ,
		_w12048_,
		_w22689_
	);
	LUT2 #(
		.INIT('h1)
	) name18642 (
		_w22688_,
		_w22689_,
		_w22690_
	);
	LUT3 #(
		.INIT('h13)
	) name18643 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001 ,
		_w9894_,
		_w22691_
	);
	LUT4 #(
		.INIT('h0002)
	) name18644 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w11631_,
		_w11632_,
		_w22691_,
		_w22692_
	);
	LUT4 #(
		.INIT('h5700)
	) name18645 (
		_w11625_,
		_w12560_,
		_w12561_,
		_w22692_,
		_w22693_
	);
	LUT4 #(
		.INIT('h313b)
	) name18646 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001 ,
		_w11631_,
		_w11635_,
		_w22694_
	);
	LUT4 #(
		.INIT('h7277)
	) name18647 (
		_w11624_,
		_w12355_,
		_w22693_,
		_w22694_,
		_w22695_
	);
	LUT2 #(
		.INIT('h2)
	) name18648 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001 ,
		_w11656_,
		_w22696_
	);
	LUT3 #(
		.INIT('h01)
	) name18649 (
		_w9946_,
		_w11659_,
		_w22696_,
		_w22697_
	);
	LUT4 #(
		.INIT('hfd00)
	) name18650 (
		_w11655_,
		_w12560_,
		_w12561_,
		_w22697_,
		_w22698_
	);
	LUT3 #(
		.INIT('h07)
	) name18651 (
		_w9946_,
		_w12355_,
		_w22698_,
		_w22699_
	);
	LUT2 #(
		.INIT('h6)
	) name18652 (
		_w21179_,
		_w21198_,
		_w22700_
	);
	LUT4 #(
		.INIT('h04c8)
	) name18653 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w13155_,
		_w21200_,
		_w22700_,
		_w22701_
	);
	LUT3 #(
		.INIT('h40)
	) name18654 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[9]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w22702_
	);
	LUT2 #(
		.INIT('h1)
	) name18655 (
		_w13158_,
		_w22702_,
		_w22703_
	);
	LUT4 #(
		.INIT('hfe00)
	) name18656 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w7140_,
		_w7240_,
		_w22703_,
		_w22704_
	);
	LUT4 #(
		.INIT('hafac)
	) name18657 (
		\sport0_rxctl_RXSHT_reg[9]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w22705_
	);
	LUT4 #(
		.INIT('h0002)
	) name18658 (
		\sport0_rxctl_RX_reg[9]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w22706_
	);
	LUT4 #(
		.INIT('hffb0)
	) name18659 (
		_w22701_,
		_w22704_,
		_w22705_,
		_w22706_,
		_w22707_
	);
	LUT4 #(
		.INIT('h4c08)
	) name18660 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w11329_,
		_w12738_,
		_w17826_,
		_w22708_
	);
	LUT2 #(
		.INIT('h1)
	) name18661 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001 ,
		_w11329_,
		_w22709_
	);
	LUT2 #(
		.INIT('h1)
	) name18662 (
		_w22708_,
		_w22709_,
		_w22710_
	);
	LUT3 #(
		.INIT('ha8)
	) name18663 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w12560_,
		_w12561_,
		_w22711_
	);
	LUT4 #(
		.INIT('h00bf)
	) name18664 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w18555_,
		_w18560_,
		_w22711_,
		_w22712_
	);
	LUT3 #(
		.INIT('he2)
	) name18665 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001 ,
		_w11946_,
		_w22712_,
		_w22713_
	);
	LUT2 #(
		.INIT('h2)
	) name18666 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w14866_,
		_w22714_
	);
	LUT4 #(
		.INIT('h4000)
	) name18667 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w18250_,
		_w18259_,
		_w18270_,
		_w22715_
	);
	LUT4 #(
		.INIT('h222e)
	) name18668 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001 ,
		_w11946_,
		_w22714_,
		_w22715_,
		_w22716_
	);
	LUT3 #(
		.INIT('he2)
	) name18669 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001 ,
		_w12048_,
		_w22712_,
		_w22717_
	);
	LUT4 #(
		.INIT('h222e)
	) name18670 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001 ,
		_w12048_,
		_w22714_,
		_w22715_,
		_w22718_
	);
	LUT4 #(
		.INIT('h152a)
	) name18671 (
		\clkc_STDcnt_reg[5]/NET0131 ,
		_w19400_,
		_w19405_,
		_w19391_,
		_w22719_
	);
	LUT3 #(
		.INIT('h78)
	) name18672 (
		\clkc_STDcnt_reg[0]/NET0131 ,
		\clkc_STDcnt_reg[1]/NET0131 ,
		\clkc_STDcnt_reg[2]/NET0131 ,
		_w22720_
	);
	LUT3 #(
		.INIT('h70)
	) name18673 (
		_w19400_,
		_w19405_,
		_w22720_,
		_w22721_
	);
	LUT4 #(
		.INIT('h5995)
	) name18674 (
		\tm_TCR_TMP_reg[11]/NET0131 ,
		_w14108_,
		_w14112_,
		_w14115_,
		_w22722_
	);
	LUT4 #(
		.INIT('h2023)
	) name18675 (
		\tm_tpr_reg_DO_reg[11]/NET0131 ,
		_w12803_,
		_w14103_,
		_w22722_,
		_w22723_
	);
	LUT4 #(
		.INIT('h0400)
	) name18676 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		\tm_tcr_reg_DO_reg[11]/NET0131 ,
		_w22724_
	);
	LUT2 #(
		.INIT('he)
	) name18677 (
		_w22723_,
		_w22724_,
		_w22725_
	);
	LUT2 #(
		.INIT('h8)
	) name18678 (
		\bdma_BCTL_reg[0]/NET0131 ,
		\bdma_BCTL_reg[1]/NET0131 ,
		_w22726_
	);
	LUT4 #(
		.INIT('hf700)
	) name18679 (
		_w4761_,
		_w12533_,
		_w20980_,
		_w22726_,
		_w22727_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18680 (
		\T_ED[1]_pad ,
		\bdma_BRdataBUF_reg[9]/P0001 ,
		_w20986_,
		_w22727_,
		_w22728_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18681 (
		\T_ED[0]_pad ,
		\bdma_BRdataBUF_reg[8]/P0001 ,
		_w20986_,
		_w22727_,
		_w22729_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18682 (
		\T_ED[7]_pad ,
		\bdma_BRdataBUF_reg[15]/P0001 ,
		_w20986_,
		_w22727_,
		_w22730_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18683 (
		\T_ED[6]_pad ,
		\bdma_BRdataBUF_reg[14]/P0001 ,
		_w20986_,
		_w22727_,
		_w22731_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18684 (
		\T_ED[5]_pad ,
		\bdma_BRdataBUF_reg[13]/P0001 ,
		_w20986_,
		_w22727_,
		_w22732_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18685 (
		\T_ED[4]_pad ,
		\bdma_BRdataBUF_reg[12]/P0001 ,
		_w20986_,
		_w22727_,
		_w22733_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18686 (
		\T_ED[3]_pad ,
		\bdma_BRdataBUF_reg[11]/P0001 ,
		_w20986_,
		_w22727_,
		_w22734_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name18687 (
		\T_ED[2]_pad ,
		\bdma_BRdataBUF_reg[10]/P0001 ,
		_w20986_,
		_w22727_,
		_w22735_
	);
	LUT4 #(
		.INIT('h135f)
	) name18688 (
		\sice_ICYC_reg[0]/NET0131 ,
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w14695_,
		_w16507_,
		_w22736_
	);
	LUT4 #(
		.INIT('h153f)
	) name18689 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\sice_IIRC_reg[0]/NET0131 ,
		_w15161_,
		_w17323_,
		_w22737_
	);
	LUT2 #(
		.INIT('h2)
	) name18690 (
		\sice_SPC_reg[1]/P0001 ,
		_w17747_,
		_w22738_
	);
	LUT4 #(
		.INIT('h00d5)
	) name18691 (
		_w21458_,
		_w22736_,
		_w22737_,
		_w22738_,
		_w22739_
	);
	LUT3 #(
		.INIT('h2e)
	) name18692 (
		\sice_SPC_reg[0]/P0001 ,
		_w16259_,
		_w22739_,
		_w22740_
	);
	LUT2 #(
		.INIT('h6)
	) name18693 (
		\clkc_STDcnt_reg[0]/NET0131 ,
		\clkc_STDcnt_reg[1]/NET0131 ,
		_w22741_
	);
	LUT3 #(
		.INIT('h70)
	) name18694 (
		_w19400_,
		_w19405_,
		_w22741_,
		_w22742_
	);
	LUT4 #(
		.INIT('ha800)
	) name18695 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w17711_,
		_w17732_,
		_w17733_,
		_w22743_
	);
	LUT4 #(
		.INIT('ha800)
	) name18696 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w17675_,
		_w17696_,
		_w17697_,
		_w22744_
	);
	LUT4 #(
		.INIT('hf888)
	) name18697 (
		\core_c_dec_updMF_E_reg/P0001 ,
		_w4106_,
		_w11926_,
		_w12808_,
		_w22745_
	);
	LUT2 #(
		.INIT('h8)
	) name18698 (
		\core_c_psq_SSTAT_reg[0]/NET0131 ,
		_w13258_,
		_w22746_
	);
	LUT4 #(
		.INIT('hefe0)
	) name18699 (
		\core_c_psq_pcstk_ptr_reg[4]/NET0131 ,
		_w4115_,
		_w22354_,
		_w22746_,
		_w22747_
	);
	LUT4 #(
		.INIT('h00ef)
	) name18700 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22119_,
		_w22748_
	);
	LUT2 #(
		.INIT('h8)
	) name18701 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w22748_,
		_w22749_
	);
	LUT4 #(
		.INIT('h0200)
	) name18702 (
		_w5672_,
		_w8757_,
		_w8760_,
		_w11605_,
		_w22750_
	);
	LUT2 #(
		.INIT('h2)
	) name18703 (
		_w22119_,
		_w22750_,
		_w22751_
	);
	LUT3 #(
		.INIT('hec)
	) name18704 (
		_w6176_,
		_w22749_,
		_w22751_,
		_w22752_
	);
	LUT2 #(
		.INIT('h8)
	) name18705 (
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w22748_,
		_w22753_
	);
	LUT3 #(
		.INIT('hf8)
	) name18706 (
		_w6501_,
		_w22751_,
		_w22753_,
		_w22754_
	);
	LUT2 #(
		.INIT('h8)
	) name18707 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w11610_,
		_w22755_
	);
	LUT3 #(
		.INIT('hf8)
	) name18708 (
		_w6176_,
		_w11614_,
		_w22755_,
		_w22756_
	);
	LUT2 #(
		.INIT('h8)
	) name18709 (
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w11610_,
		_w22757_
	);
	LUT3 #(
		.INIT('hf8)
	) name18710 (
		_w6501_,
		_w11614_,
		_w22757_,
		_w22758_
	);
	LUT4 #(
		.INIT('h7774)
	) name18711 (
		\idma_IADi_reg[14]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w8757_,
		_w8760_,
		_w22759_
	);
	LUT3 #(
		.INIT('h2e)
	) name18712 (
		\idma_DCTL_reg[14]/NET0131 ,
		_w19994_,
		_w22759_,
		_w22760_
	);
	LUT4 #(
		.INIT('hc444)
	) name18713 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		_w4073_,
		_w4084_,
		_w22761_
	);
	LUT2 #(
		.INIT('h4)
	) name18714 (
		_w12274_,
		_w12277_,
		_w22762_
	);
	LUT4 #(
		.INIT('hf2f0)
	) name18715 (
		_w12271_,
		_w12272_,
		_w22761_,
		_w22762_,
		_w22763_
	);
	LUT2 #(
		.INIT('h8)
	) name18716 (
		\bdma_BEAD_reg[11]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w22764_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18717 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		_w4721_,
		_w4804_,
		_w4805_,
		_w22765_
	);
	LUT4 #(
		.INIT('h8088)
	) name18718 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		\emc_DMcst_reg/NET0131 ,
		_w4718_,
		_w4799_,
		_w22766_
	);
	LUT2 #(
		.INIT('h8)
	) name18719 (
		\emc_ECMA_reg[11]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w22767_
	);
	LUT4 #(
		.INIT('h5554)
	) name18720 (
		\bdma_BM_cyc_reg/P0001 ,
		_w22766_,
		_w22767_,
		_w22765_,
		_w22768_
	);
	LUT2 #(
		.INIT('he)
	) name18721 (
		_w22764_,
		_w22768_,
		_w22769_
	);
	LUT4 #(
		.INIT('h0002)
	) name18722 (
		_w4128_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w22770_
	);
	LUT3 #(
		.INIT('h14)
	) name18723 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[7]/P0001 ,
		_w4528_,
		_w22771_
	);
	LUT4 #(
		.INIT('h2022)
	) name18724 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w7793_,
		_w7903_,
		_w7905_,
		_w22772_
	);
	LUT4 #(
		.INIT('h4447)
	) name18725 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22771_,
		_w22772_,
		_w22773_
	);
	LUT3 #(
		.INIT('h2e)
	) name18726 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001 ,
		_w22770_,
		_w22773_,
		_w22774_
	);
	LUT4 #(
		.INIT('h1450)
	) name18727 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[4]/P0001 ,
		\core_c_psq_EXA_reg[5]/P0001 ,
		_w4527_,
		_w22775_
	);
	LUT4 #(
		.INIT('h2022)
	) name18728 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w7592_,
		_w7707_,
		_w7709_,
		_w22776_
	);
	LUT4 #(
		.INIT('h4447)
	) name18729 (
		\core_c_psq_EXA_reg[5]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22775_,
		_w22776_,
		_w22777_
	);
	LUT3 #(
		.INIT('h2e)
	) name18730 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001 ,
		_w22770_,
		_w22777_,
		_w22778_
	);
	LUT3 #(
		.INIT('h14)
	) name18731 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[4]/P0001 ,
		_w4527_,
		_w22779_
	);
	LUT4 #(
		.INIT('h2022)
	) name18732 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w7257_,
		_w7375_,
		_w7377_,
		_w22780_
	);
	LUT4 #(
		.INIT('h4447)
	) name18733 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22779_,
		_w22780_,
		_w22781_
	);
	LUT3 #(
		.INIT('h2e)
	) name18734 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001 ,
		_w22770_,
		_w22781_,
		_w22782_
	);
	LUT2 #(
		.INIT('h4)
	) name18735 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w4601_,
		_w22783_
	);
	LUT4 #(
		.INIT('h2022)
	) name18736 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w6054_,
		_w6173_,
		_w6175_,
		_w22784_
	);
	LUT4 #(
		.INIT('h4447)
	) name18737 (
		\core_c_psq_EXA_reg[3]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22783_,
		_w22784_,
		_w22785_
	);
	LUT3 #(
		.INIT('h2e)
	) name18738 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001 ,
		_w22770_,
		_w22785_,
		_w22786_
	);
	LUT3 #(
		.INIT('h14)
	) name18739 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_EXA_reg[1]/P0001 ,
		_w22787_
	);
	LUT4 #(
		.INIT('h2022)
	) name18740 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w6774_,
		_w6894_,
		_w6896_,
		_w22788_
	);
	LUT4 #(
		.INIT('h4447)
	) name18741 (
		\core_c_psq_EXA_reg[1]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22787_,
		_w22788_,
		_w22789_
	);
	LUT3 #(
		.INIT('h2e)
	) name18742 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001 ,
		_w22770_,
		_w22789_,
		_w22790_
	);
	LUT2 #(
		.INIT('h2)
	) name18743 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001 ,
		_w22770_,
		_w22791_
	);
	LUT4 #(
		.INIT('h1450)
	) name18744 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_EXA_reg[11]/P0001 ,
		_w4529_,
		_w22792_
	);
	LUT4 #(
		.INIT('h00fd)
	) name18745 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w6263_,
		_w6362_,
		_w22792_,
		_w22793_
	);
	LUT4 #(
		.INIT('h80b0)
	) name18746 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22770_,
		_w22793_,
		_w22794_
	);
	LUT2 #(
		.INIT('he)
	) name18747 (
		_w22791_,
		_w22794_,
		_w22795_
	);
	LUT2 #(
		.INIT('h2)
	) name18748 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001 ,
		_w22770_,
		_w22796_
	);
	LUT3 #(
		.INIT('h14)
	) name18749 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[10]/P0001 ,
		_w4529_,
		_w22797_
	);
	LUT4 #(
		.INIT('h00fd)
	) name18750 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5937_,
		_w6038_,
		_w22797_,
		_w22798_
	);
	LUT4 #(
		.INIT('h80b0)
	) name18751 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22770_,
		_w22798_,
		_w22799_
	);
	LUT2 #(
		.INIT('he)
	) name18752 (
		_w22796_,
		_w22799_,
		_w22800_
	);
	LUT4 #(
		.INIT('h2022)
	) name18753 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5784_,
		_w5911_,
		_w5913_,
		_w22801_
	);
	LUT4 #(
		.INIT('h303e)
	) name18754 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22801_,
		_w22802_
	);
	LUT3 #(
		.INIT('h2e)
	) name18755 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001 ,
		_w22770_,
		_w22802_,
		_w22803_
	);
	LUT4 #(
		.INIT('h0002)
	) name18756 (
		_w4115_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w22804_
	);
	LUT2 #(
		.INIT('h2)
	) name18757 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001 ,
		_w22804_,
		_w22805_
	);
	LUT2 #(
		.INIT('h4)
	) name18758 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w4704_,
		_w22806_
	);
	LUT4 #(
		.INIT('h00fd)
	) name18759 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w7140_,
		_w7240_,
		_w22806_,
		_w22807_
	);
	LUT4 #(
		.INIT('h80b0)
	) name18760 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22804_,
		_w22807_,
		_w22808_
	);
	LUT2 #(
		.INIT('he)
	) name18761 (
		_w22805_,
		_w22808_,
		_w22809_
	);
	LUT2 #(
		.INIT('h2)
	) name18762 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001 ,
		_w22804_,
		_w22810_
	);
	LUT4 #(
		.INIT('h1450)
	) name18763 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[7]/P0001 ,
		\core_c_psq_EXA_reg[8]/P0001 ,
		_w4528_,
		_w22811_
	);
	LUT4 #(
		.INIT('h00fd)
	) name18764 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w7465_,
		_w7565_,
		_w22811_,
		_w22812_
	);
	LUT4 #(
		.INIT('h80b0)
	) name18765 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22804_,
		_w22812_,
		_w22813_
	);
	LUT2 #(
		.INIT('he)
	) name18766 (
		_w22810_,
		_w22813_,
		_w22814_
	);
	LUT3 #(
		.INIT('h3a)
	) name18767 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001 ,
		_w22773_,
		_w22804_,
		_w22815_
	);
	LUT2 #(
		.INIT('h4)
	) name18768 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w4659_,
		_w22816_
	);
	LUT4 #(
		.INIT('h2022)
	) name18769 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w7927_,
		_w8040_,
		_w8042_,
		_w22817_
	);
	LUT4 #(
		.INIT('h4447)
	) name18770 (
		\core_c_psq_EXA_reg[6]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22816_,
		_w22817_,
		_w22818_
	);
	LUT3 #(
		.INIT('h2e)
	) name18771 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001 ,
		_w22804_,
		_w22818_,
		_w22819_
	);
	LUT3 #(
		.INIT('h3a)
	) name18772 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001 ,
		_w22785_,
		_w22804_,
		_w22820_
	);
	LUT4 #(
		.INIT('h1540)
	) name18773 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_EXA_reg[1]/P0001 ,
		\core_c_psq_EXA_reg[2]/P0001 ,
		_w22821_
	);
	LUT4 #(
		.INIT('h2022)
	) name18774 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w6378_,
		_w6498_,
		_w6500_,
		_w22822_
	);
	LUT4 #(
		.INIT('h4447)
	) name18775 (
		\core_c_psq_EXA_reg[2]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22821_,
		_w22822_,
		_w22823_
	);
	LUT3 #(
		.INIT('h2e)
	) name18776 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001 ,
		_w22804_,
		_w22823_,
		_w22824_
	);
	LUT3 #(
		.INIT('h3a)
	) name18777 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001 ,
		_w22789_,
		_w22804_,
		_w22825_
	);
	LUT4 #(
		.INIT('h3210)
	) name18778 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4828_,
		_w5760_,
		_w22826_
	);
	LUT2 #(
		.INIT('h8)
	) name18779 (
		\core_c_psq_EXA_reg[13]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22827_
	);
	LUT4 #(
		.INIT('heee2)
	) name18780 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001 ,
		_w22804_,
		_w22826_,
		_w22827_,
		_w22828_
	);
	LUT4 #(
		.INIT('h3210)
	) name18781 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4811_,
		_w6758_,
		_w22829_
	);
	LUT2 #(
		.INIT('h8)
	) name18782 (
		\core_c_psq_EXA_reg[12]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22830_
	);
	LUT4 #(
		.INIT('heee2)
	) name18783 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001 ,
		_w22804_,
		_w22829_,
		_w22830_,
		_w22831_
	);
	LUT2 #(
		.INIT('h2)
	) name18784 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001 ,
		_w22804_,
		_w22832_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18785 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w22804_,
		_w22833_
	);
	LUT2 #(
		.INIT('he)
	) name18786 (
		_w22832_,
		_w22833_,
		_w22834_
	);
	LUT2 #(
		.INIT('h2)
	) name18787 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001 ,
		_w22804_,
		_w22835_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18788 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w22804_,
		_w22836_
	);
	LUT2 #(
		.INIT('he)
	) name18789 (
		_w22835_,
		_w22836_,
		_w22837_
	);
	LUT3 #(
		.INIT('h3a)
	) name18790 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001 ,
		_w22802_,
		_w22804_,
		_w22838_
	);
	LUT4 #(
		.INIT('h0002)
	) name18791 (
		_w4125_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w22839_
	);
	LUT2 #(
		.INIT('h2)
	) name18792 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001 ,
		_w22839_,
		_w22840_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18793 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w22839_,
		_w22841_
	);
	LUT2 #(
		.INIT('he)
	) name18794 (
		_w22840_,
		_w22841_,
		_w22842_
	);
	LUT2 #(
		.INIT('h2)
	) name18795 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001 ,
		_w22839_,
		_w22843_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18796 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w22839_,
		_w22844_
	);
	LUT2 #(
		.INIT('he)
	) name18797 (
		_w22843_,
		_w22844_,
		_w22845_
	);
	LUT3 #(
		.INIT('h3a)
	) name18798 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001 ,
		_w22773_,
		_w22839_,
		_w22846_
	);
	LUT3 #(
		.INIT('h3a)
	) name18799 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001 ,
		_w22818_,
		_w22839_,
		_w22847_
	);
	LUT3 #(
		.INIT('h3a)
	) name18800 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001 ,
		_w22777_,
		_w22839_,
		_w22848_
	);
	LUT3 #(
		.INIT('h3a)
	) name18801 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001 ,
		_w22781_,
		_w22839_,
		_w22849_
	);
	LUT3 #(
		.INIT('h3a)
	) name18802 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001 ,
		_w22785_,
		_w22839_,
		_w22850_
	);
	LUT3 #(
		.INIT('h3a)
	) name18803 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001 ,
		_w22823_,
		_w22839_,
		_w22851_
	);
	LUT3 #(
		.INIT('h3a)
	) name18804 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001 ,
		_w22789_,
		_w22839_,
		_w22852_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18805 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w22839_,
		_w22853_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18806 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w22839_,
		_w22854_
	);
	LUT2 #(
		.INIT('h2)
	) name18807 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001 ,
		_w22839_,
		_w22855_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18808 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w22839_,
		_w22856_
	);
	LUT2 #(
		.INIT('he)
	) name18809 (
		_w22855_,
		_w22856_,
		_w22857_
	);
	LUT2 #(
		.INIT('h2)
	) name18810 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001 ,
		_w22839_,
		_w22858_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18811 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w22839_,
		_w22859_
	);
	LUT2 #(
		.INIT('he)
	) name18812 (
		_w22858_,
		_w22859_,
		_w22860_
	);
	LUT3 #(
		.INIT('h3a)
	) name18813 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001 ,
		_w22802_,
		_w22839_,
		_w22861_
	);
	LUT4 #(
		.INIT('h0002)
	) name18814 (
		_w4118_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w22862_
	);
	LUT2 #(
		.INIT('h2)
	) name18815 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001 ,
		_w22862_,
		_w22863_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18816 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w22862_,
		_w22864_
	);
	LUT2 #(
		.INIT('he)
	) name18817 (
		_w22863_,
		_w22864_,
		_w22865_
	);
	LUT2 #(
		.INIT('h2)
	) name18818 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001 ,
		_w22862_,
		_w22866_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18819 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w22862_,
		_w22867_
	);
	LUT2 #(
		.INIT('he)
	) name18820 (
		_w22866_,
		_w22867_,
		_w22868_
	);
	LUT3 #(
		.INIT('h3a)
	) name18821 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001 ,
		_w22773_,
		_w22862_,
		_w22869_
	);
	LUT3 #(
		.INIT('h3a)
	) name18822 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001 ,
		_w22818_,
		_w22862_,
		_w22870_
	);
	LUT3 #(
		.INIT('h3a)
	) name18823 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001 ,
		_w22777_,
		_w22862_,
		_w22871_
	);
	LUT3 #(
		.INIT('h3a)
	) name18824 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001 ,
		_w22781_,
		_w22862_,
		_w22872_
	);
	LUT3 #(
		.INIT('h3a)
	) name18825 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001 ,
		_w22785_,
		_w22862_,
		_w22873_
	);
	LUT3 #(
		.INIT('h3a)
	) name18826 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001 ,
		_w22823_,
		_w22862_,
		_w22874_
	);
	LUT3 #(
		.INIT('h3a)
	) name18827 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001 ,
		_w22789_,
		_w22862_,
		_w22875_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18828 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w22862_,
		_w22876_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18829 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w22862_,
		_w22877_
	);
	LUT2 #(
		.INIT('h2)
	) name18830 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001 ,
		_w22862_,
		_w22878_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18831 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w22862_,
		_w22879_
	);
	LUT2 #(
		.INIT('he)
	) name18832 (
		_w22878_,
		_w22879_,
		_w22880_
	);
	LUT2 #(
		.INIT('h2)
	) name18833 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001 ,
		_w22862_,
		_w22881_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18834 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w22862_,
		_w22882_
	);
	LUT2 #(
		.INIT('he)
	) name18835 (
		_w22881_,
		_w22882_,
		_w22883_
	);
	LUT3 #(
		.INIT('h3a)
	) name18836 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001 ,
		_w22802_,
		_w22862_,
		_w22884_
	);
	LUT4 #(
		.INIT('h0002)
	) name18837 (
		_w4135_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w22885_
	);
	LUT2 #(
		.INIT('h2)
	) name18838 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001 ,
		_w22885_,
		_w22886_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18839 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w22885_,
		_w22887_
	);
	LUT2 #(
		.INIT('he)
	) name18840 (
		_w22886_,
		_w22887_,
		_w22888_
	);
	LUT2 #(
		.INIT('h2)
	) name18841 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001 ,
		_w22885_,
		_w22889_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18842 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w22885_,
		_w22890_
	);
	LUT2 #(
		.INIT('he)
	) name18843 (
		_w22889_,
		_w22890_,
		_w22891_
	);
	LUT3 #(
		.INIT('h3a)
	) name18844 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001 ,
		_w22773_,
		_w22885_,
		_w22892_
	);
	LUT3 #(
		.INIT('h3a)
	) name18845 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001 ,
		_w22818_,
		_w22885_,
		_w22893_
	);
	LUT3 #(
		.INIT('h3a)
	) name18846 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001 ,
		_w22777_,
		_w22885_,
		_w22894_
	);
	LUT3 #(
		.INIT('h3a)
	) name18847 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001 ,
		_w22781_,
		_w22885_,
		_w22895_
	);
	LUT3 #(
		.INIT('h3a)
	) name18848 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001 ,
		_w22785_,
		_w22885_,
		_w22896_
	);
	LUT3 #(
		.INIT('h3a)
	) name18849 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001 ,
		_w22823_,
		_w22885_,
		_w22897_
	);
	LUT3 #(
		.INIT('h3a)
	) name18850 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001 ,
		_w22789_,
		_w22885_,
		_w22898_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18851 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w22885_,
		_w22899_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18852 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w22885_,
		_w22900_
	);
	LUT2 #(
		.INIT('h2)
	) name18853 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001 ,
		_w22885_,
		_w22901_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18854 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w22885_,
		_w22902_
	);
	LUT2 #(
		.INIT('he)
	) name18855 (
		_w22901_,
		_w22902_,
		_w22903_
	);
	LUT2 #(
		.INIT('h2)
	) name18856 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001 ,
		_w22885_,
		_w22904_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18857 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w22885_,
		_w22905_
	);
	LUT2 #(
		.INIT('he)
	) name18858 (
		_w22904_,
		_w22905_,
		_w22906_
	);
	LUT3 #(
		.INIT('h3a)
	) name18859 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001 ,
		_w22802_,
		_w22885_,
		_w22907_
	);
	LUT4 #(
		.INIT('h0002)
	) name18860 (
		_w4121_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w22908_
	);
	LUT2 #(
		.INIT('h2)
	) name18861 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001 ,
		_w22908_,
		_w22909_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18862 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w22908_,
		_w22910_
	);
	LUT2 #(
		.INIT('he)
	) name18863 (
		_w22909_,
		_w22910_,
		_w22911_
	);
	LUT2 #(
		.INIT('h2)
	) name18864 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001 ,
		_w22908_,
		_w22912_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18865 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w22908_,
		_w22913_
	);
	LUT2 #(
		.INIT('he)
	) name18866 (
		_w22912_,
		_w22913_,
		_w22914_
	);
	LUT3 #(
		.INIT('h3a)
	) name18867 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001 ,
		_w22773_,
		_w22908_,
		_w22915_
	);
	LUT3 #(
		.INIT('h3a)
	) name18868 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001 ,
		_w22818_,
		_w22908_,
		_w22916_
	);
	LUT3 #(
		.INIT('h3a)
	) name18869 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001 ,
		_w22777_,
		_w22908_,
		_w22917_
	);
	LUT3 #(
		.INIT('h3a)
	) name18870 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001 ,
		_w22781_,
		_w22908_,
		_w22918_
	);
	LUT3 #(
		.INIT('h3a)
	) name18871 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001 ,
		_w22785_,
		_w22908_,
		_w22919_
	);
	LUT3 #(
		.INIT('h3a)
	) name18872 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001 ,
		_w22823_,
		_w22908_,
		_w22920_
	);
	LUT3 #(
		.INIT('h3a)
	) name18873 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001 ,
		_w22789_,
		_w22908_,
		_w22921_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18874 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w22908_,
		_w22922_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18875 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w22908_,
		_w22923_
	);
	LUT2 #(
		.INIT('h2)
	) name18876 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001 ,
		_w22908_,
		_w22924_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18877 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w22908_,
		_w22925_
	);
	LUT2 #(
		.INIT('he)
	) name18878 (
		_w22924_,
		_w22925_,
		_w22926_
	);
	LUT2 #(
		.INIT('h2)
	) name18879 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001 ,
		_w22908_,
		_w22927_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18880 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w22908_,
		_w22928_
	);
	LUT2 #(
		.INIT('he)
	) name18881 (
		_w22927_,
		_w22928_,
		_w22929_
	);
	LUT3 #(
		.INIT('h3a)
	) name18882 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001 ,
		_w22802_,
		_w22908_,
		_w22930_
	);
	LUT4 #(
		.INIT('h0002)
	) name18883 (
		_w4119_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w22931_
	);
	LUT2 #(
		.INIT('h2)
	) name18884 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001 ,
		_w22931_,
		_w22932_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18885 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w22931_,
		_w22933_
	);
	LUT2 #(
		.INIT('he)
	) name18886 (
		_w22932_,
		_w22933_,
		_w22934_
	);
	LUT2 #(
		.INIT('h2)
	) name18887 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001 ,
		_w22931_,
		_w22935_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18888 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w22931_,
		_w22936_
	);
	LUT2 #(
		.INIT('he)
	) name18889 (
		_w22935_,
		_w22936_,
		_w22937_
	);
	LUT3 #(
		.INIT('h3a)
	) name18890 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001 ,
		_w22773_,
		_w22931_,
		_w22938_
	);
	LUT3 #(
		.INIT('h3a)
	) name18891 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001 ,
		_w22818_,
		_w22931_,
		_w22939_
	);
	LUT3 #(
		.INIT('h3a)
	) name18892 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001 ,
		_w22777_,
		_w22931_,
		_w22940_
	);
	LUT3 #(
		.INIT('h3a)
	) name18893 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001 ,
		_w22781_,
		_w22931_,
		_w22941_
	);
	LUT3 #(
		.INIT('h3a)
	) name18894 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001 ,
		_w22785_,
		_w22931_,
		_w22942_
	);
	LUT3 #(
		.INIT('h3a)
	) name18895 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001 ,
		_w22823_,
		_w22931_,
		_w22943_
	);
	LUT3 #(
		.INIT('h3a)
	) name18896 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001 ,
		_w22789_,
		_w22931_,
		_w22944_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18897 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w22931_,
		_w22945_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18898 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w22931_,
		_w22946_
	);
	LUT2 #(
		.INIT('h2)
	) name18899 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001 ,
		_w22931_,
		_w22947_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18900 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w22931_,
		_w22948_
	);
	LUT2 #(
		.INIT('he)
	) name18901 (
		_w22947_,
		_w22948_,
		_w22949_
	);
	LUT2 #(
		.INIT('h2)
	) name18902 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001 ,
		_w22931_,
		_w22950_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18903 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w22931_,
		_w22951_
	);
	LUT2 #(
		.INIT('he)
	) name18904 (
		_w22950_,
		_w22951_,
		_w22952_
	);
	LUT3 #(
		.INIT('h3a)
	) name18905 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001 ,
		_w22802_,
		_w22931_,
		_w22953_
	);
	LUT4 #(
		.INIT('h0002)
	) name18906 (
		_w4131_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w22954_
	);
	LUT2 #(
		.INIT('h2)
	) name18907 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001 ,
		_w22954_,
		_w22955_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18908 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w22954_,
		_w22956_
	);
	LUT2 #(
		.INIT('he)
	) name18909 (
		_w22955_,
		_w22956_,
		_w22957_
	);
	LUT2 #(
		.INIT('h2)
	) name18910 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001 ,
		_w22954_,
		_w22958_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18911 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w22954_,
		_w22959_
	);
	LUT2 #(
		.INIT('he)
	) name18912 (
		_w22958_,
		_w22959_,
		_w22960_
	);
	LUT3 #(
		.INIT('h3a)
	) name18913 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001 ,
		_w22773_,
		_w22954_,
		_w22961_
	);
	LUT3 #(
		.INIT('h3a)
	) name18914 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001 ,
		_w22818_,
		_w22954_,
		_w22962_
	);
	LUT3 #(
		.INIT('h3a)
	) name18915 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001 ,
		_w22777_,
		_w22954_,
		_w22963_
	);
	LUT3 #(
		.INIT('h3a)
	) name18916 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001 ,
		_w22781_,
		_w22954_,
		_w22964_
	);
	LUT3 #(
		.INIT('h3a)
	) name18917 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001 ,
		_w22785_,
		_w22954_,
		_w22965_
	);
	LUT3 #(
		.INIT('h3a)
	) name18918 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001 ,
		_w22823_,
		_w22954_,
		_w22966_
	);
	LUT3 #(
		.INIT('h3a)
	) name18919 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001 ,
		_w22789_,
		_w22954_,
		_w22967_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18920 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w22954_,
		_w22968_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18921 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w22954_,
		_w22969_
	);
	LUT2 #(
		.INIT('h2)
	) name18922 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001 ,
		_w22954_,
		_w22970_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18923 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w22954_,
		_w22971_
	);
	LUT2 #(
		.INIT('he)
	) name18924 (
		_w22970_,
		_w22971_,
		_w22972_
	);
	LUT2 #(
		.INIT('h2)
	) name18925 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001 ,
		_w22954_,
		_w22973_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18926 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w22954_,
		_w22974_
	);
	LUT2 #(
		.INIT('he)
	) name18927 (
		_w22973_,
		_w22974_,
		_w22975_
	);
	LUT3 #(
		.INIT('h3a)
	) name18928 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001 ,
		_w22802_,
		_w22954_,
		_w22976_
	);
	LUT4 #(
		.INIT('h0008)
	) name18929 (
		\core_c_psq_pcstk_ptr_reg[4]/NET0131 ,
		_w4114_,
		_w13258_,
		_w22357_,
		_w22977_
	);
	LUT2 #(
		.INIT('h2)
	) name18930 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001 ,
		_w22977_,
		_w22978_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18931 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w22977_,
		_w22979_
	);
	LUT2 #(
		.INIT('he)
	) name18932 (
		_w22978_,
		_w22979_,
		_w22980_
	);
	LUT2 #(
		.INIT('h2)
	) name18933 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001 ,
		_w22977_,
		_w22981_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18934 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w22977_,
		_w22982_
	);
	LUT2 #(
		.INIT('he)
	) name18935 (
		_w22981_,
		_w22982_,
		_w22983_
	);
	LUT3 #(
		.INIT('h3a)
	) name18936 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001 ,
		_w22773_,
		_w22977_,
		_w22984_
	);
	LUT3 #(
		.INIT('h3a)
	) name18937 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001 ,
		_w22818_,
		_w22977_,
		_w22985_
	);
	LUT3 #(
		.INIT('h3a)
	) name18938 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001 ,
		_w22777_,
		_w22977_,
		_w22986_
	);
	LUT3 #(
		.INIT('h3a)
	) name18939 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001 ,
		_w22781_,
		_w22977_,
		_w22987_
	);
	LUT3 #(
		.INIT('h3a)
	) name18940 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001 ,
		_w22785_,
		_w22977_,
		_w22988_
	);
	LUT3 #(
		.INIT('h3a)
	) name18941 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001 ,
		_w22823_,
		_w22977_,
		_w22989_
	);
	LUT3 #(
		.INIT('h3a)
	) name18942 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001 ,
		_w22789_,
		_w22977_,
		_w22990_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18943 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w22977_,
		_w22991_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name18944 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w22977_,
		_w22992_
	);
	LUT2 #(
		.INIT('h2)
	) name18945 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001 ,
		_w22977_,
		_w22993_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18946 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w22977_,
		_w22994_
	);
	LUT2 #(
		.INIT('he)
	) name18947 (
		_w22993_,
		_w22994_,
		_w22995_
	);
	LUT2 #(
		.INIT('h2)
	) name18948 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001 ,
		_w22977_,
		_w22996_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18949 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w22977_,
		_w22997_
	);
	LUT2 #(
		.INIT('he)
	) name18950 (
		_w22996_,
		_w22997_,
		_w22998_
	);
	LUT3 #(
		.INIT('h3a)
	) name18951 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001 ,
		_w22802_,
		_w22977_,
		_w22999_
	);
	LUT4 #(
		.INIT('hc444)
	) name18952 (
		\core_c_psq_INT_en_reg/NET0131 ,
		\core_c_psq_Iact_E_reg[3]/NET0131 ,
		_w4073_,
		_w4084_,
		_w23000_
	);
	LUT2 #(
		.INIT('h8)
	) name18953 (
		_w12269_,
		_w20447_,
		_w23001_
	);
	LUT3 #(
		.INIT('h80)
	) name18954 (
		_w12279_,
		_w20440_,
		_w23001_,
		_w23002_
	);
	LUT4 #(
		.INIT('h2a00)
	) name18955 (
		\core_c_psq_INT_en_reg/NET0131 ,
		_w4073_,
		_w4084_,
		_w23002_,
		_w23003_
	);
	LUT2 #(
		.INIT('he)
	) name18956 (
		_w23000_,
		_w23003_,
		_w23004_
	);
	LUT3 #(
		.INIT('h2e)
	) name18957 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001 ,
		_w22770_,
		_w22818_,
		_w23005_
	);
	LUT4 #(
		.INIT('h5444)
	) name18958 (
		\sport1_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w14590_,
		_w14591_,
		_w14594_,
		_w23006_
	);
	LUT4 #(
		.INIT('h0121)
	) name18959 (
		\sport1_txctl_Wcnt_reg[0]/NET0131 ,
		_w14590_,
		_w14591_,
		_w14594_,
		_w23007_
	);
	LUT2 #(
		.INIT('h1)
	) name18960 (
		_w23006_,
		_w23007_,
		_w23008_
	);
	LUT4 #(
		.INIT('ha3ac)
	) name18961 (
		\sport1_regs_MWORDreg_DO_reg[6]/NET0131 ,
		\sport1_txctl_Wcnt_reg[6]/NET0131 ,
		_w14595_,
		_w22336_,
		_w23009_
	);
	LUT3 #(
		.INIT('h63)
	) name18962 (
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		\sport1_txctl_Wcnt_reg[3]/NET0131 ,
		_w22334_,
		_w23010_
	);
	LUT4 #(
		.INIT('h1500)
	) name18963 (
		_w14590_,
		_w14591_,
		_w14594_,
		_w23010_,
		_w23011_
	);
	LUT4 #(
		.INIT('h5444)
	) name18964 (
		\sport1_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w14590_,
		_w14591_,
		_w14594_,
		_w23012_
	);
	LUT2 #(
		.INIT('h1)
	) name18965 (
		_w23011_,
		_w23012_,
		_w23013_
	);
	LUT2 #(
		.INIT('h9)
	) name18966 (
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		_w22334_,
		_w23014_
	);
	LUT4 #(
		.INIT('h1500)
	) name18967 (
		_w14590_,
		_w14591_,
		_w14594_,
		_w23014_,
		_w23015_
	);
	LUT4 #(
		.INIT('h5444)
	) name18968 (
		\sport1_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w14590_,
		_w14591_,
		_w14594_,
		_w23016_
	);
	LUT2 #(
		.INIT('h1)
	) name18969 (
		_w23015_,
		_w23016_,
		_w23017_
	);
	LUT4 #(
		.INIT('ha3ac)
	) name18970 (
		\sport0_regs_MWORDreg_DO_reg[6]/NET0131 ,
		\sport0_txctl_Wcnt_reg[6]/NET0131 ,
		_w14601_,
		_w22343_,
		_w23018_
	);
	LUT3 #(
		.INIT('h63)
	) name18971 (
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		\sport0_txctl_Wcnt_reg[3]/NET0131 ,
		_w22341_,
		_w23019_
	);
	LUT4 #(
		.INIT('h1500)
	) name18972 (
		_w14596_,
		_w14597_,
		_w14600_,
		_w23019_,
		_w23020_
	);
	LUT4 #(
		.INIT('h5444)
	) name18973 (
		\sport0_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w14596_,
		_w14597_,
		_w14600_,
		_w23021_
	);
	LUT2 #(
		.INIT('h1)
	) name18974 (
		_w23020_,
		_w23021_,
		_w23022_
	);
	LUT2 #(
		.INIT('h9)
	) name18975 (
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		_w22341_,
		_w23023_
	);
	LUT4 #(
		.INIT('h1500)
	) name18976 (
		_w14596_,
		_w14597_,
		_w14600_,
		_w23023_,
		_w23024_
	);
	LUT4 #(
		.INIT('h5444)
	) name18977 (
		\sport0_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w14596_,
		_w14597_,
		_w14600_,
		_w23025_
	);
	LUT2 #(
		.INIT('h1)
	) name18978 (
		_w23024_,
		_w23025_,
		_w23026_
	);
	LUT4 #(
		.INIT('h5444)
	) name18979 (
		\sport0_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w14596_,
		_w14597_,
		_w14600_,
		_w23027_
	);
	LUT4 #(
		.INIT('h0121)
	) name18980 (
		\sport0_txctl_Wcnt_reg[0]/NET0131 ,
		_w14596_,
		_w14597_,
		_w14600_,
		_w23028_
	);
	LUT2 #(
		.INIT('h1)
	) name18981 (
		_w23027_,
		_w23028_,
		_w23029_
	);
	LUT2 #(
		.INIT('h1)
	) name18982 (
		_w12619_,
		_w19993_,
		_w23030_
	);
	LUT3 #(
		.INIT('hca)
	) name18983 (
		\idma_DOVL_reg[9]/NET0131 ,
		_w20007_,
		_w23030_,
		_w23031_
	);
	LUT3 #(
		.INIT('hca)
	) name18984 (
		\idma_DOVL_reg[8]/NET0131 ,
		_w19995_,
		_w23030_,
		_w23032_
	);
	LUT3 #(
		.INIT('hca)
	) name18985 (
		\idma_DOVL_reg[10]/NET0131 ,
		_w20026_,
		_w23030_,
		_w23033_
	);
	LUT3 #(
		.INIT('hca)
	) name18986 (
		\idma_DOVL_reg[11]/NET0131 ,
		_w20023_,
		_w23030_,
		_w23034_
	);
	LUT4 #(
		.INIT('heee2)
	) name18987 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001 ,
		_w22770_,
		_w22829_,
		_w22830_,
		_w23035_
	);
	LUT4 #(
		.INIT('heee2)
	) name18988 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001 ,
		_w22770_,
		_w22826_,
		_w22827_,
		_w23036_
	);
	LUT3 #(
		.INIT('h3a)
	) name18989 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001 ,
		_w22777_,
		_w22804_,
		_w23037_
	);
	LUT3 #(
		.INIT('h2e)
	) name18990 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001 ,
		_w22770_,
		_w22823_,
		_w23038_
	);
	LUT4 #(
		.INIT('h0002)
	) name18991 (
		_w4110_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w23039_
	);
	LUT2 #(
		.INIT('h2)
	) name18992 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001 ,
		_w23039_,
		_w23040_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18993 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w23039_,
		_w23041_
	);
	LUT2 #(
		.INIT('he)
	) name18994 (
		_w23040_,
		_w23041_,
		_w23042_
	);
	LUT2 #(
		.INIT('h2)
	) name18995 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001 ,
		_w23039_,
		_w23043_
	);
	LUT4 #(
		.INIT('h8b00)
	) name18996 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w23039_,
		_w23044_
	);
	LUT2 #(
		.INIT('he)
	) name18997 (
		_w23043_,
		_w23044_,
		_w23045_
	);
	LUT3 #(
		.INIT('h3a)
	) name18998 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001 ,
		_w22773_,
		_w23039_,
		_w23046_
	);
	LUT3 #(
		.INIT('h3a)
	) name18999 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001 ,
		_w22818_,
		_w23039_,
		_w23047_
	);
	LUT3 #(
		.INIT('h3a)
	) name19000 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001 ,
		_w22777_,
		_w23039_,
		_w23048_
	);
	LUT3 #(
		.INIT('h3a)
	) name19001 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001 ,
		_w22781_,
		_w23039_,
		_w23049_
	);
	LUT3 #(
		.INIT('h3a)
	) name19002 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001 ,
		_w22785_,
		_w23039_,
		_w23050_
	);
	LUT3 #(
		.INIT('h3a)
	) name19003 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001 ,
		_w22823_,
		_w23039_,
		_w23051_
	);
	LUT3 #(
		.INIT('h3a)
	) name19004 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001 ,
		_w22789_,
		_w23039_,
		_w23052_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19005 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w23039_,
		_w23053_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19006 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w23039_,
		_w23054_
	);
	LUT2 #(
		.INIT('h2)
	) name19007 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001 ,
		_w23039_,
		_w23055_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19008 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w23039_,
		_w23056_
	);
	LUT2 #(
		.INIT('he)
	) name19009 (
		_w23055_,
		_w23056_,
		_w23057_
	);
	LUT2 #(
		.INIT('h2)
	) name19010 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001 ,
		_w23039_,
		_w23058_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19011 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w23039_,
		_w23059_
	);
	LUT2 #(
		.INIT('he)
	) name19012 (
		_w23058_,
		_w23059_,
		_w23060_
	);
	LUT3 #(
		.INIT('h3a)
	) name19013 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001 ,
		_w22802_,
		_w23039_,
		_w23061_
	);
	LUT4 #(
		.INIT('h0002)
	) name19014 (
		_w4112_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w23062_
	);
	LUT2 #(
		.INIT('h2)
	) name19015 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001 ,
		_w23062_,
		_w23063_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19016 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w23062_,
		_w23064_
	);
	LUT2 #(
		.INIT('he)
	) name19017 (
		_w23063_,
		_w23064_,
		_w23065_
	);
	LUT2 #(
		.INIT('h2)
	) name19018 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001 ,
		_w23062_,
		_w23066_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19019 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w23062_,
		_w23067_
	);
	LUT2 #(
		.INIT('he)
	) name19020 (
		_w23066_,
		_w23067_,
		_w23068_
	);
	LUT3 #(
		.INIT('h3a)
	) name19021 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001 ,
		_w22773_,
		_w23062_,
		_w23069_
	);
	LUT3 #(
		.INIT('h3a)
	) name19022 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001 ,
		_w22818_,
		_w23062_,
		_w23070_
	);
	LUT3 #(
		.INIT('h3a)
	) name19023 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001 ,
		_w22777_,
		_w23062_,
		_w23071_
	);
	LUT3 #(
		.INIT('h3a)
	) name19024 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001 ,
		_w22781_,
		_w23062_,
		_w23072_
	);
	LUT3 #(
		.INIT('h3a)
	) name19025 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001 ,
		_w22785_,
		_w23062_,
		_w23073_
	);
	LUT3 #(
		.INIT('h3a)
	) name19026 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001 ,
		_w22823_,
		_w23062_,
		_w23074_
	);
	LUT3 #(
		.INIT('h3a)
	) name19027 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001 ,
		_w22789_,
		_w23062_,
		_w23075_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19028 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w23062_,
		_w23076_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19029 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w23062_,
		_w23077_
	);
	LUT2 #(
		.INIT('h2)
	) name19030 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001 ,
		_w23062_,
		_w23078_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19031 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w23062_,
		_w23079_
	);
	LUT2 #(
		.INIT('he)
	) name19032 (
		_w23078_,
		_w23079_,
		_w23080_
	);
	LUT2 #(
		.INIT('h2)
	) name19033 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001 ,
		_w23062_,
		_w23081_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19034 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w23062_,
		_w23082_
	);
	LUT2 #(
		.INIT('he)
	) name19035 (
		_w23081_,
		_w23082_,
		_w23083_
	);
	LUT3 #(
		.INIT('h3a)
	) name19036 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001 ,
		_w22802_,
		_w23062_,
		_w23084_
	);
	LUT4 #(
		.INIT('h0002)
	) name19037 (
		_w4129_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w23085_
	);
	LUT2 #(
		.INIT('h2)
	) name19038 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001 ,
		_w23085_,
		_w23086_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19039 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w23085_,
		_w23087_
	);
	LUT2 #(
		.INIT('he)
	) name19040 (
		_w23086_,
		_w23087_,
		_w23088_
	);
	LUT2 #(
		.INIT('h2)
	) name19041 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001 ,
		_w23085_,
		_w23089_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19042 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w23085_,
		_w23090_
	);
	LUT2 #(
		.INIT('he)
	) name19043 (
		_w23089_,
		_w23090_,
		_w23091_
	);
	LUT3 #(
		.INIT('h3a)
	) name19044 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001 ,
		_w22773_,
		_w23085_,
		_w23092_
	);
	LUT3 #(
		.INIT('h3a)
	) name19045 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001 ,
		_w22818_,
		_w23085_,
		_w23093_
	);
	LUT3 #(
		.INIT('h3a)
	) name19046 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001 ,
		_w22777_,
		_w23085_,
		_w23094_
	);
	LUT3 #(
		.INIT('h3a)
	) name19047 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001 ,
		_w22781_,
		_w23085_,
		_w23095_
	);
	LUT3 #(
		.INIT('h3a)
	) name19048 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001 ,
		_w22785_,
		_w23085_,
		_w23096_
	);
	LUT3 #(
		.INIT('h3a)
	) name19049 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001 ,
		_w22823_,
		_w23085_,
		_w23097_
	);
	LUT3 #(
		.INIT('h3a)
	) name19050 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001 ,
		_w22789_,
		_w23085_,
		_w23098_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19051 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w23085_,
		_w23099_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19052 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w23085_,
		_w23100_
	);
	LUT2 #(
		.INIT('h2)
	) name19053 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001 ,
		_w23085_,
		_w23101_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19054 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w23085_,
		_w23102_
	);
	LUT2 #(
		.INIT('he)
	) name19055 (
		_w23101_,
		_w23102_,
		_w23103_
	);
	LUT2 #(
		.INIT('h2)
	) name19056 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001 ,
		_w23085_,
		_w23104_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19057 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w23085_,
		_w23105_
	);
	LUT2 #(
		.INIT('he)
	) name19058 (
		_w23104_,
		_w23105_,
		_w23106_
	);
	LUT3 #(
		.INIT('h3a)
	) name19059 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001 ,
		_w22802_,
		_w23085_,
		_w23107_
	);
	LUT4 #(
		.INIT('h0002)
	) name19060 (
		_w4132_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w23108_
	);
	LUT2 #(
		.INIT('h2)
	) name19061 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001 ,
		_w23108_,
		_w23109_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19062 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w23108_,
		_w23110_
	);
	LUT2 #(
		.INIT('he)
	) name19063 (
		_w23109_,
		_w23110_,
		_w23111_
	);
	LUT2 #(
		.INIT('h2)
	) name19064 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001 ,
		_w23108_,
		_w23112_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19065 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w23108_,
		_w23113_
	);
	LUT2 #(
		.INIT('he)
	) name19066 (
		_w23112_,
		_w23113_,
		_w23114_
	);
	LUT3 #(
		.INIT('h3a)
	) name19067 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001 ,
		_w22773_,
		_w23108_,
		_w23115_
	);
	LUT3 #(
		.INIT('h3a)
	) name19068 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001 ,
		_w22818_,
		_w23108_,
		_w23116_
	);
	LUT3 #(
		.INIT('h3a)
	) name19069 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001 ,
		_w22781_,
		_w23108_,
		_w23117_
	);
	LUT3 #(
		.INIT('h3a)
	) name19070 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001 ,
		_w22785_,
		_w23108_,
		_w23118_
	);
	LUT3 #(
		.INIT('h3a)
	) name19071 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001 ,
		_w22777_,
		_w23108_,
		_w23119_
	);
	LUT3 #(
		.INIT('h3a)
	) name19072 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001 ,
		_w22823_,
		_w23108_,
		_w23120_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19073 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w23108_,
		_w23121_
	);
	LUT3 #(
		.INIT('h3a)
	) name19074 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001 ,
		_w22789_,
		_w23108_,
		_w23122_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19075 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w23108_,
		_w23123_
	);
	LUT2 #(
		.INIT('h2)
	) name19076 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001 ,
		_w23108_,
		_w23124_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19077 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w23108_,
		_w23125_
	);
	LUT2 #(
		.INIT('he)
	) name19078 (
		_w23124_,
		_w23125_,
		_w23126_
	);
	LUT2 #(
		.INIT('h2)
	) name19079 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001 ,
		_w23108_,
		_w23127_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19080 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w23108_,
		_w23128_
	);
	LUT2 #(
		.INIT('he)
	) name19081 (
		_w23127_,
		_w23128_,
		_w23129_
	);
	LUT3 #(
		.INIT('h3a)
	) name19082 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001 ,
		_w22802_,
		_w23108_,
		_w23130_
	);
	LUT4 #(
		.INIT('h0002)
	) name19083 (
		_w4126_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w23131_
	);
	LUT2 #(
		.INIT('h2)
	) name19084 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001 ,
		_w23131_,
		_w23132_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19085 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w23131_,
		_w23133_
	);
	LUT2 #(
		.INIT('he)
	) name19086 (
		_w23132_,
		_w23133_,
		_w23134_
	);
	LUT2 #(
		.INIT('h2)
	) name19087 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001 ,
		_w23131_,
		_w23135_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19088 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w23131_,
		_w23136_
	);
	LUT2 #(
		.INIT('he)
	) name19089 (
		_w23135_,
		_w23136_,
		_w23137_
	);
	LUT3 #(
		.INIT('h3a)
	) name19090 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001 ,
		_w22773_,
		_w23131_,
		_w23138_
	);
	LUT3 #(
		.INIT('h3a)
	) name19091 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001 ,
		_w22818_,
		_w23131_,
		_w23139_
	);
	LUT3 #(
		.INIT('h3a)
	) name19092 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001 ,
		_w22777_,
		_w23131_,
		_w23140_
	);
	LUT3 #(
		.INIT('h3a)
	) name19093 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001 ,
		_w22781_,
		_w23131_,
		_w23141_
	);
	LUT3 #(
		.INIT('h3a)
	) name19094 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001 ,
		_w22785_,
		_w23131_,
		_w23142_
	);
	LUT3 #(
		.INIT('h3a)
	) name19095 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001 ,
		_w22823_,
		_w23131_,
		_w23143_
	);
	LUT3 #(
		.INIT('h3a)
	) name19096 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001 ,
		_w22789_,
		_w23131_,
		_w23144_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19097 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w23131_,
		_w23145_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19098 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w23131_,
		_w23146_
	);
	LUT2 #(
		.INIT('h2)
	) name19099 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001 ,
		_w23131_,
		_w23147_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19100 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w23131_,
		_w23148_
	);
	LUT2 #(
		.INIT('he)
	) name19101 (
		_w23147_,
		_w23148_,
		_w23149_
	);
	LUT3 #(
		.INIT('h3a)
	) name19102 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001 ,
		_w22802_,
		_w23131_,
		_w23150_
	);
	LUT2 #(
		.INIT('h2)
	) name19103 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001 ,
		_w23131_,
		_w23151_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19104 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w23131_,
		_w23152_
	);
	LUT2 #(
		.INIT('he)
	) name19105 (
		_w23151_,
		_w23152_,
		_w23153_
	);
	LUT4 #(
		.INIT('h0002)
	) name19106 (
		_w4134_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w23154_
	);
	LUT2 #(
		.INIT('h2)
	) name19107 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001 ,
		_w23154_,
		_w23155_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19108 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w23154_,
		_w23156_
	);
	LUT2 #(
		.INIT('he)
	) name19109 (
		_w23155_,
		_w23156_,
		_w23157_
	);
	LUT2 #(
		.INIT('h2)
	) name19110 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001 ,
		_w23154_,
		_w23158_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19111 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w23154_,
		_w23159_
	);
	LUT2 #(
		.INIT('he)
	) name19112 (
		_w23158_,
		_w23159_,
		_w23160_
	);
	LUT3 #(
		.INIT('h3a)
	) name19113 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001 ,
		_w22773_,
		_w23154_,
		_w23161_
	);
	LUT3 #(
		.INIT('h3a)
	) name19114 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001 ,
		_w22818_,
		_w23154_,
		_w23162_
	);
	LUT3 #(
		.INIT('h3a)
	) name19115 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001 ,
		_w22777_,
		_w23154_,
		_w23163_
	);
	LUT3 #(
		.INIT('h3a)
	) name19116 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001 ,
		_w22781_,
		_w23154_,
		_w23164_
	);
	LUT3 #(
		.INIT('h3a)
	) name19117 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001 ,
		_w22785_,
		_w23154_,
		_w23165_
	);
	LUT3 #(
		.INIT('h3a)
	) name19118 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001 ,
		_w22823_,
		_w23154_,
		_w23166_
	);
	LUT3 #(
		.INIT('h3a)
	) name19119 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001 ,
		_w22789_,
		_w23154_,
		_w23167_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19120 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w23154_,
		_w23168_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19121 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w23154_,
		_w23169_
	);
	LUT2 #(
		.INIT('h2)
	) name19122 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001 ,
		_w23154_,
		_w23170_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19123 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w23154_,
		_w23171_
	);
	LUT2 #(
		.INIT('he)
	) name19124 (
		_w23170_,
		_w23171_,
		_w23172_
	);
	LUT2 #(
		.INIT('h2)
	) name19125 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001 ,
		_w23154_,
		_w23173_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19126 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w23154_,
		_w23174_
	);
	LUT2 #(
		.INIT('he)
	) name19127 (
		_w23173_,
		_w23174_,
		_w23175_
	);
	LUT3 #(
		.INIT('h3a)
	) name19128 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001 ,
		_w22802_,
		_w23154_,
		_w23176_
	);
	LUT4 #(
		.INIT('h0002)
	) name19129 (
		_w4122_,
		_w13258_,
		_w13259_,
		_w22357_,
		_w23177_
	);
	LUT2 #(
		.INIT('h2)
	) name19130 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001 ,
		_w23177_,
		_w23178_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19131 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22807_,
		_w23177_,
		_w23179_
	);
	LUT2 #(
		.INIT('he)
	) name19132 (
		_w23178_,
		_w23179_,
		_w23180_
	);
	LUT2 #(
		.INIT('h2)
	) name19133 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001 ,
		_w23177_,
		_w23181_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19134 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22812_,
		_w23177_,
		_w23182_
	);
	LUT2 #(
		.INIT('he)
	) name19135 (
		_w23181_,
		_w23182_,
		_w23183_
	);
	LUT3 #(
		.INIT('h3a)
	) name19136 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001 ,
		_w22773_,
		_w23177_,
		_w23184_
	);
	LUT3 #(
		.INIT('h3a)
	) name19137 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001 ,
		_w22781_,
		_w22804_,
		_w23185_
	);
	LUT3 #(
		.INIT('h3a)
	) name19138 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001 ,
		_w22818_,
		_w23177_,
		_w23186_
	);
	LUT3 #(
		.INIT('h3a)
	) name19139 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001 ,
		_w22777_,
		_w23177_,
		_w23187_
	);
	LUT3 #(
		.INIT('h3a)
	) name19140 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001 ,
		_w22781_,
		_w23177_,
		_w23188_
	);
	LUT3 #(
		.INIT('h3a)
	) name19141 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001 ,
		_w22785_,
		_w23177_,
		_w23189_
	);
	LUT3 #(
		.INIT('h3a)
	) name19142 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001 ,
		_w22823_,
		_w23177_,
		_w23190_
	);
	LUT3 #(
		.INIT('h3a)
	) name19143 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001 ,
		_w22789_,
		_w23177_,
		_w23191_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19144 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001 ,
		_w22826_,
		_w22827_,
		_w23177_,
		_w23192_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name19145 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001 ,
		_w22829_,
		_w22830_,
		_w23177_,
		_w23193_
	);
	LUT2 #(
		.INIT('h2)
	) name19146 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001 ,
		_w23177_,
		_w23194_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19147 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22793_,
		_w23177_,
		_w23195_
	);
	LUT2 #(
		.INIT('he)
	) name19148 (
		_w23194_,
		_w23195_,
		_w23196_
	);
	LUT2 #(
		.INIT('h2)
	) name19149 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001 ,
		_w23177_,
		_w23197_
	);
	LUT4 #(
		.INIT('h8b00)
	) name19150 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22798_,
		_w23177_,
		_w23198_
	);
	LUT2 #(
		.INIT('he)
	) name19151 (
		_w23197_,
		_w23198_,
		_w23199_
	);
	LUT3 #(
		.INIT('h3a)
	) name19152 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001 ,
		_w22802_,
		_w23177_,
		_w23200_
	);
	LUT2 #(
		.INIT('h2)
	) name19153 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001 ,
		_w22770_,
		_w23201_
	);
	LUT4 #(
		.INIT('h80b0)
	) name19154 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22770_,
		_w22807_,
		_w23202_
	);
	LUT2 #(
		.INIT('he)
	) name19155 (
		_w23201_,
		_w23202_,
		_w23203_
	);
	LUT2 #(
		.INIT('h2)
	) name19156 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001 ,
		_w22770_,
		_w23204_
	);
	LUT4 #(
		.INIT('h80b0)
	) name19157 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w22770_,
		_w22812_,
		_w23205_
	);
	LUT2 #(
		.INIT('he)
	) name19158 (
		_w23204_,
		_w23205_,
		_w23206_
	);
	LUT4 #(
		.INIT('h03aa)
	) name19159 (
		\idma_DOVL_reg[7]/NET0131 ,
		_w20037_,
		_w20038_,
		_w23030_,
		_w23207_
	);
	LUT4 #(
		.INIT('h03aa)
	) name19160 (
		\idma_DOVL_reg[6]/NET0131 ,
		_w20046_,
		_w20047_,
		_w23030_,
		_w23208_
	);
	LUT4 #(
		.INIT('h03aa)
	) name19161 (
		\idma_DOVL_reg[5]/NET0131 ,
		_w20041_,
		_w20042_,
		_w23030_,
		_w23209_
	);
	LUT4 #(
		.INIT('h03aa)
	) name19162 (
		\idma_DOVL_reg[3]/NET0131 ,
		_w20055_,
		_w20056_,
		_w23030_,
		_w23210_
	);
	LUT4 #(
		.INIT('h03aa)
	) name19163 (
		\idma_DOVL_reg[4]/NET0131 ,
		_w20050_,
		_w20051_,
		_w23030_,
		_w23211_
	);
	LUT4 #(
		.INIT('h03aa)
	) name19164 (
		\idma_DOVL_reg[2]/NET0131 ,
		_w20060_,
		_w20061_,
		_w23030_,
		_w23212_
	);
	LUT4 #(
		.INIT('h03aa)
	) name19165 (
		\idma_DOVL_reg[1]/NET0131 ,
		_w20117_,
		_w20118_,
		_w23030_,
		_w23213_
	);
	LUT4 #(
		.INIT('h03aa)
	) name19166 (
		\idma_DOVL_reg[0]/NET0131 ,
		_w20065_,
		_w20066_,
		_w23030_,
		_w23214_
	);
	LUT2 #(
		.INIT('h8)
	) name19167 (
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w11610_,
		_w23215_
	);
	LUT3 #(
		.INIT('hf8)
	) name19168 (
		_w7906_,
		_w11614_,
		_w23215_,
		_w23216_
	);
	LUT2 #(
		.INIT('h8)
	) name19169 (
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w11610_,
		_w23217_
	);
	LUT3 #(
		.INIT('hf8)
	) name19170 (
		_w8043_,
		_w11614_,
		_w23217_,
		_w23218_
	);
	LUT2 #(
		.INIT('h8)
	) name19171 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w11610_,
		_w23219_
	);
	LUT3 #(
		.INIT('hf8)
	) name19172 (
		_w7710_,
		_w11614_,
		_w23219_,
		_w23220_
	);
	LUT2 #(
		.INIT('h8)
	) name19173 (
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w11610_,
		_w23221_
	);
	LUT3 #(
		.INIT('h08)
	) name19174 (
		_w8802_,
		_w11607_,
		_w11613_,
		_w23222_
	);
	LUT2 #(
		.INIT('he)
	) name19175 (
		_w23221_,
		_w23222_,
		_w23223_
	);
	LUT2 #(
		.INIT('h8)
	) name19176 (
		\ISCLK0_pad ,
		_w11610_,
		_w23224_
	);
	LUT3 #(
		.INIT('h08)
	) name19177 (
		_w8761_,
		_w11607_,
		_w11613_,
		_w23225_
	);
	LUT2 #(
		.INIT('he)
	) name19178 (
		_w23224_,
		_w23225_,
		_w23226_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name19179 (
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		\sport0_txctl_Wcnt_reg[3]/NET0131 ,
		\sport0_txctl_Wcnt_reg[4]/NET0131 ,
		_w22341_,
		_w23227_
	);
	LUT4 #(
		.INIT('h1500)
	) name19180 (
		_w14596_,
		_w14597_,
		_w14600_,
		_w23227_,
		_w23228_
	);
	LUT4 #(
		.INIT('h5444)
	) name19181 (
		\sport0_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w14596_,
		_w14597_,
		_w14600_,
		_w23229_
	);
	LUT2 #(
		.INIT('h1)
	) name19182 (
		_w23228_,
		_w23229_,
		_w23230_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name19183 (
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		\sport1_txctl_Wcnt_reg[3]/NET0131 ,
		\sport1_txctl_Wcnt_reg[4]/NET0131 ,
		_w22334_,
		_w23231_
	);
	LUT4 #(
		.INIT('h1500)
	) name19184 (
		_w14590_,
		_w14591_,
		_w14594_,
		_w23231_,
		_w23232_
	);
	LUT4 #(
		.INIT('h5444)
	) name19185 (
		\sport1_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w14590_,
		_w14591_,
		_w14594_,
		_w23233_
	);
	LUT2 #(
		.INIT('h1)
	) name19186 (
		_w23232_,
		_w23233_,
		_w23234_
	);
	LUT3 #(
		.INIT('h12)
	) name19187 (
		\bdma_BEAD_reg[2]/NET0131 ,
		_w13032_,
		_w13031_,
		_w23235_
	);
	LUT4 #(
		.INIT('h4500)
	) name19188 (
		_w6378_,
		_w6498_,
		_w6500_,
		_w13032_,
		_w23236_
	);
	LUT2 #(
		.INIT('he)
	) name19189 (
		_w23235_,
		_w23236_,
		_w23237_
	);
	LUT4 #(
		.INIT('h3363)
	) name19190 (
		\sport1_txctl_Wcnt_reg[0]/NET0131 ,
		\sport1_txctl_Wcnt_reg[1]/NET0131 ,
		_w14591_,
		_w14594_,
		_w23238_
	);
	LUT4 #(
		.INIT('h1500)
	) name19191 (
		_w14590_,
		_w14591_,
		_w14594_,
		_w23238_,
		_w23239_
	);
	LUT4 #(
		.INIT('h5444)
	) name19192 (
		\sport1_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w14590_,
		_w14591_,
		_w14594_,
		_w23240_
	);
	LUT2 #(
		.INIT('h1)
	) name19193 (
		_w23239_,
		_w23240_,
		_w23241_
	);
	LUT4 #(
		.INIT('h3363)
	) name19194 (
		\sport0_txctl_Wcnt_reg[0]/NET0131 ,
		\sport0_txctl_Wcnt_reg[1]/NET0131 ,
		_w14597_,
		_w14600_,
		_w23242_
	);
	LUT4 #(
		.INIT('h1500)
	) name19195 (
		_w14596_,
		_w14597_,
		_w14600_,
		_w23242_,
		_w23243_
	);
	LUT4 #(
		.INIT('h5444)
	) name19196 (
		\sport0_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w14596_,
		_w14597_,
		_w14600_,
		_w23244_
	);
	LUT2 #(
		.INIT('h1)
	) name19197 (
		_w23243_,
		_w23244_,
		_w23245_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name19198 (
		\idma_RDcnt_reg[2]/NET0131 ,
		\memc_usysr_DO_reg[6]/NET0131 ,
		_w13075_,
		_w13076_,
		_w23246_
	);
	LUT2 #(
		.INIT('h8)
	) name19199 (
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w22748_,
		_w23247_
	);
	LUT3 #(
		.INIT('hf8)
	) name19200 (
		_w7906_,
		_w22751_,
		_w23247_,
		_w23248_
	);
	LUT2 #(
		.INIT('h8)
	) name19201 (
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w22748_,
		_w23249_
	);
	LUT3 #(
		.INIT('hf8)
	) name19202 (
		_w8043_,
		_w22751_,
		_w23249_,
		_w23250_
	);
	LUT2 #(
		.INIT('h8)
	) name19203 (
		\sport1_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w22748_,
		_w23251_
	);
	LUT3 #(
		.INIT('hf8)
	) name19204 (
		_w7710_,
		_w22751_,
		_w23251_,
		_w23252_
	);
	LUT2 #(
		.INIT('h8)
	) name19205 (
		\sport1_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w22748_,
		_w23253_
	);
	LUT3 #(
		.INIT('hf8)
	) name19206 (
		_w7378_,
		_w22751_,
		_w23253_,
		_w23254_
	);
	LUT2 #(
		.INIT('h8)
	) name19207 (
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w22748_,
		_w23255_
	);
	LUT3 #(
		.INIT('h08)
	) name19208 (
		_w8802_,
		_w22119_,
		_w22750_,
		_w23256_
	);
	LUT2 #(
		.INIT('he)
	) name19209 (
		_w23255_,
		_w23256_,
		_w23257_
	);
	LUT4 #(
		.INIT('h0103)
	) name19210 (
		_w5672_,
		_w8757_,
		_w8760_,
		_w11605_,
		_w23258_
	);
	LUT4 #(
		.INIT('hce02)
	) name19211 (
		\ISCLK1_pad ,
		_w22119_,
		_w22120_,
		_w23258_,
		_w23259_
	);
	LUT2 #(
		.INIT('h8)
	) name19212 (
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w22748_,
		_w23260_
	);
	LUT3 #(
		.INIT('h08)
	) name19213 (
		_w5760_,
		_w22119_,
		_w22750_,
		_w23261_
	);
	LUT2 #(
		.INIT('he)
	) name19214 (
		_w23260_,
		_w23261_,
		_w23262_
	);
	LUT2 #(
		.INIT('h8)
	) name19215 (
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w22748_,
		_w23263_
	);
	LUT3 #(
		.INIT('h08)
	) name19216 (
		_w6758_,
		_w22119_,
		_w22750_,
		_w23264_
	);
	LUT2 #(
		.INIT('he)
	) name19217 (
		_w23263_,
		_w23264_,
		_w23265_
	);
	LUT4 #(
		.INIT('h00ef)
	) name19218 (
		_w8757_,
		_w8760_,
		_w11984_,
		_w22149_,
		_w23266_
	);
	LUT2 #(
		.INIT('h8)
	) name19219 (
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w23266_,
		_w23267_
	);
	LUT4 #(
		.INIT('h0010)
	) name19220 (
		_w7140_,
		_w7240_,
		_w22149_,
		_w22750_,
		_w23268_
	);
	LUT2 #(
		.INIT('he)
	) name19221 (
		_w23267_,
		_w23268_,
		_w23269_
	);
	LUT2 #(
		.INIT('h8)
	) name19222 (
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w23266_,
		_w23270_
	);
	LUT4 #(
		.INIT('h0010)
	) name19223 (
		_w7465_,
		_w7565_,
		_w22149_,
		_w22750_,
		_w23271_
	);
	LUT2 #(
		.INIT('he)
	) name19224 (
		_w23270_,
		_w23271_,
		_w23272_
	);
	LUT2 #(
		.INIT('h8)
	) name19225 (
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w23266_,
		_w23273_
	);
	LUT3 #(
		.INIT('h08)
	) name19226 (
		_w8802_,
		_w22149_,
		_w22750_,
		_w23274_
	);
	LUT2 #(
		.INIT('he)
	) name19227 (
		_w23273_,
		_w23274_,
		_w23275_
	);
	LUT4 #(
		.INIT('hf202)
	) name19228 (
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w22120_,
		_w22149_,
		_w23258_,
		_w23276_
	);
	LUT2 #(
		.INIT('h8)
	) name19229 (
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w23266_,
		_w23277_
	);
	LUT3 #(
		.INIT('h08)
	) name19230 (
		_w5760_,
		_w22149_,
		_w22750_,
		_w23278_
	);
	LUT2 #(
		.INIT('he)
	) name19231 (
		_w23277_,
		_w23278_,
		_w23279_
	);
	LUT2 #(
		.INIT('h8)
	) name19232 (
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w23266_,
		_w23280_
	);
	LUT3 #(
		.INIT('h08)
	) name19233 (
		_w6758_,
		_w22149_,
		_w22750_,
		_w23281_
	);
	LUT2 #(
		.INIT('he)
	) name19234 (
		_w23280_,
		_w23281_,
		_w23282_
	);
	LUT2 #(
		.INIT('h8)
	) name19235 (
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w23266_,
		_w23283_
	);
	LUT4 #(
		.INIT('h0010)
	) name19236 (
		_w5937_,
		_w6038_,
		_w22149_,
		_w22750_,
		_w23284_
	);
	LUT2 #(
		.INIT('he)
	) name19237 (
		_w23283_,
		_w23284_,
		_w23285_
	);
	LUT2 #(
		.INIT('h8)
	) name19238 (
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w23266_,
		_w23286_
	);
	LUT4 #(
		.INIT('h0010)
	) name19239 (
		_w6263_,
		_w6362_,
		_w22149_,
		_w22750_,
		_w23287_
	);
	LUT2 #(
		.INIT('he)
	) name19240 (
		_w23286_,
		_w23287_,
		_w23288_
	);
	LUT4 #(
		.INIT('hccac)
	) name19241 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001 ,
		_w9919_,
		_w11602_,
		_w23289_
	);
	LUT4 #(
		.INIT('hccac)
	) name19242 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001 ,
		_w9919_,
		_w11602_,
		_w23290_
	);
	LUT4 #(
		.INIT('haaca)
	) name19243 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001 ,
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w9919_,
		_w11602_,
		_w23291_
	);
	LUT4 #(
		.INIT('haa3a)
	) name19244 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001 ,
		_w4155_,
		_w9919_,
		_w11602_,
		_w23292_
	);
	LUT4 #(
		.INIT('haaca)
	) name19245 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w9919_,
		_w11602_,
		_w23293_
	);
	LUT4 #(
		.INIT('haaca)
	) name19246 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w9919_,
		_w11602_,
		_w23294_
	);
	LUT4 #(
		.INIT('haaca)
	) name19247 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w9919_,
		_w11602_,
		_w23295_
	);
	LUT4 #(
		.INIT('haaca)
	) name19248 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w9919_,
		_w11602_,
		_w23296_
	);
	LUT4 #(
		.INIT('hccac)
	) name19249 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001 ,
		_w9919_,
		_w11602_,
		_w23297_
	);
	LUT4 #(
		.INIT('hccac)
	) name19250 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001 ,
		_w9919_,
		_w11602_,
		_w23298_
	);
	LUT4 #(
		.INIT('hccac)
	) name19251 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001 ,
		_w9919_,
		_w11602_,
		_w23299_
	);
	LUT4 #(
		.INIT('hccac)
	) name19252 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001 ,
		_w9919_,
		_w11602_,
		_w23300_
	);
	LUT4 #(
		.INIT('hccac)
	) name19253 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001 ,
		_w9919_,
		_w11602_,
		_w23301_
	);
	LUT4 #(
		.INIT('haaca)
	) name19254 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001 ,
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w9919_,
		_w11602_,
		_w23302_
	);
	LUT4 #(
		.INIT('hccac)
	) name19255 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001 ,
		_w9919_,
		_w11602_,
		_w23303_
	);
	LUT4 #(
		.INIT('hccac)
	) name19256 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001 ,
		_w9919_,
		_w11602_,
		_w23304_
	);
	LUT4 #(
		.INIT('hccac)
	) name19257 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001 ,
		_w9919_,
		_w11602_,
		_w23305_
	);
	LUT4 #(
		.INIT('hccac)
	) name19258 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001 ,
		_w9919_,
		_w11602_,
		_w23306_
	);
	LUT4 #(
		.INIT('hccac)
	) name19259 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001 ,
		_w9919_,
		_w11602_,
		_w23307_
	);
	LUT4 #(
		.INIT('hccac)
	) name19260 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001 ,
		_w9919_,
		_w11602_,
		_w23308_
	);
	LUT4 #(
		.INIT('hccac)
	) name19261 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001 ,
		_w9919_,
		_w11602_,
		_w23309_
	);
	LUT4 #(
		.INIT('h04c8)
	) name19262 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w13155_,
		_w19091_,
		_w19096_,
		_w23310_
	);
	LUT4 #(
		.INIT('h1011)
	) name19263 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w7927_,
		_w8040_,
		_w8042_,
		_w23311_
	);
	LUT3 #(
		.INIT('h40)
	) name19264 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w23312_
	);
	LUT2 #(
		.INIT('h1)
	) name19265 (
		_w13158_,
		_w23312_,
		_w23313_
	);
	LUT4 #(
		.INIT('hafac)
	) name19266 (
		\sport0_rxctl_RXSHT_reg[6]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w23314_
	);
	LUT4 #(
		.INIT('hef00)
	) name19267 (
		_w23310_,
		_w23311_,
		_w23313_,
		_w23314_,
		_w23315_
	);
	LUT4 #(
		.INIT('h0002)
	) name19268 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w13158_,
		_w13161_,
		_w23316_
	);
	LUT2 #(
		.INIT('he)
	) name19269 (
		_w23315_,
		_w23316_,
		_w23317_
	);
	LUT4 #(
		.INIT('hccac)
	) name19270 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001 ,
		_w9919_,
		_w11602_,
		_w23318_
	);
	LUT4 #(
		.INIT('hccac)
	) name19271 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001 ,
		_w9919_,
		_w11602_,
		_w23319_
	);
	LUT4 #(
		.INIT('hccac)
	) name19272 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001 ,
		_w9919_,
		_w11602_,
		_w23320_
	);
	LUT4 #(
		.INIT('haaca)
	) name19273 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w9919_,
		_w11602_,
		_w23321_
	);
	LUT4 #(
		.INIT('hccac)
	) name19274 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001 ,
		_w9925_,
		_w11602_,
		_w23322_
	);
	LUT4 #(
		.INIT('hccac)
	) name19275 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001 ,
		_w9925_,
		_w11602_,
		_w23323_
	);
	LUT4 #(
		.INIT('haaca)
	) name19276 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001 ,
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w9925_,
		_w11602_,
		_w23324_
	);
	LUT4 #(
		.INIT('haa3a)
	) name19277 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001 ,
		_w4155_,
		_w9925_,
		_w11602_,
		_w23325_
	);
	LUT4 #(
		.INIT('haaca)
	) name19278 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w9925_,
		_w11602_,
		_w23326_
	);
	LUT4 #(
		.INIT('haaca)
	) name19279 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w9925_,
		_w11602_,
		_w23327_
	);
	LUT4 #(
		.INIT('haaca)
	) name19280 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w9925_,
		_w11602_,
		_w23328_
	);
	LUT4 #(
		.INIT('haaca)
	) name19281 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w9925_,
		_w11602_,
		_w23329_
	);
	LUT4 #(
		.INIT('hccac)
	) name19282 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001 ,
		_w9925_,
		_w11602_,
		_w23330_
	);
	LUT4 #(
		.INIT('hccac)
	) name19283 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001 ,
		_w9925_,
		_w11602_,
		_w23331_
	);
	LUT4 #(
		.INIT('hccac)
	) name19284 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001 ,
		_w9925_,
		_w11602_,
		_w23332_
	);
	LUT4 #(
		.INIT('hccac)
	) name19285 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001 ,
		_w9925_,
		_w11602_,
		_w23333_
	);
	LUT4 #(
		.INIT('hccac)
	) name19286 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001 ,
		_w9925_,
		_w11602_,
		_w23334_
	);
	LUT4 #(
		.INIT('haaca)
	) name19287 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001 ,
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w9925_,
		_w11602_,
		_w23335_
	);
	LUT4 #(
		.INIT('hccac)
	) name19288 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001 ,
		_w9925_,
		_w11602_,
		_w23336_
	);
	LUT4 #(
		.INIT('hccac)
	) name19289 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001 ,
		_w9925_,
		_w11602_,
		_w23337_
	);
	LUT4 #(
		.INIT('hccac)
	) name19290 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001 ,
		_w9925_,
		_w11602_,
		_w23338_
	);
	LUT4 #(
		.INIT('hccac)
	) name19291 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001 ,
		_w9925_,
		_w11602_,
		_w23339_
	);
	LUT4 #(
		.INIT('hccac)
	) name19292 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001 ,
		_w9925_,
		_w11602_,
		_w23340_
	);
	LUT4 #(
		.INIT('hccac)
	) name19293 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001 ,
		_w9925_,
		_w11602_,
		_w23341_
	);
	LUT4 #(
		.INIT('hccac)
	) name19294 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001 ,
		_w9925_,
		_w11602_,
		_w23342_
	);
	LUT4 #(
		.INIT('hccac)
	) name19295 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001 ,
		_w9925_,
		_w11602_,
		_w23343_
	);
	LUT4 #(
		.INIT('hccac)
	) name19296 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001 ,
		_w9925_,
		_w11602_,
		_w23344_
	);
	LUT4 #(
		.INIT('hccac)
	) name19297 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001 ,
		_w9925_,
		_w11602_,
		_w23345_
	);
	LUT4 #(
		.INIT('haaca)
	) name19298 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w9925_,
		_w11602_,
		_w23346_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19299 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001 ,
		_w9908_,
		_w11602_,
		_w23347_
	);
	LUT4 #(
		.INIT('h0020)
	) name19300 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23348_
	);
	LUT2 #(
		.INIT('he)
	) name19301 (
		_w23347_,
		_w23348_,
		_w23349_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19302 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001 ,
		_w9908_,
		_w11602_,
		_w23350_
	);
	LUT4 #(
		.INIT('h0020)
	) name19303 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23351_
	);
	LUT2 #(
		.INIT('he)
	) name19304 (
		_w23350_,
		_w23351_,
		_w23352_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19305 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001 ,
		_w9908_,
		_w11602_,
		_w23353_
	);
	LUT4 #(
		.INIT('h0040)
	) name19306 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w9908_,
		_w11602_,
		_w23354_
	);
	LUT2 #(
		.INIT('he)
	) name19307 (
		_w23353_,
		_w23354_,
		_w23355_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19308 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001 ,
		_w9908_,
		_w11602_,
		_w23356_
	);
	LUT4 #(
		.INIT('h0010)
	) name19309 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w4155_,
		_w9908_,
		_w11602_,
		_w23357_
	);
	LUT2 #(
		.INIT('he)
	) name19310 (
		_w23356_,
		_w23357_,
		_w23358_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19311 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001 ,
		_w9908_,
		_w11602_,
		_w23359_
	);
	LUT4 #(
		.INIT('h0040)
	) name19312 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w9908_,
		_w11602_,
		_w23360_
	);
	LUT2 #(
		.INIT('he)
	) name19313 (
		_w23359_,
		_w23360_,
		_w23361_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19314 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001 ,
		_w9908_,
		_w11602_,
		_w23362_
	);
	LUT4 #(
		.INIT('h0040)
	) name19315 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w9908_,
		_w11602_,
		_w23363_
	);
	LUT2 #(
		.INIT('he)
	) name19316 (
		_w23362_,
		_w23363_,
		_w23364_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19317 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001 ,
		_w9908_,
		_w11602_,
		_w23365_
	);
	LUT4 #(
		.INIT('h0040)
	) name19318 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w9908_,
		_w11602_,
		_w23366_
	);
	LUT2 #(
		.INIT('he)
	) name19319 (
		_w23365_,
		_w23366_,
		_w23367_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19320 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001 ,
		_w9908_,
		_w11602_,
		_w23368_
	);
	LUT4 #(
		.INIT('h0040)
	) name19321 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w9908_,
		_w11602_,
		_w23369_
	);
	LUT2 #(
		.INIT('he)
	) name19322 (
		_w23368_,
		_w23369_,
		_w23370_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19323 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001 ,
		_w9908_,
		_w11602_,
		_w23371_
	);
	LUT4 #(
		.INIT('h0020)
	) name19324 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23372_
	);
	LUT2 #(
		.INIT('he)
	) name19325 (
		_w23371_,
		_w23372_,
		_w23373_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19326 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001 ,
		_w9908_,
		_w11602_,
		_w23374_
	);
	LUT4 #(
		.INIT('h0020)
	) name19327 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23375_
	);
	LUT2 #(
		.INIT('he)
	) name19328 (
		_w23374_,
		_w23375_,
		_w23376_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19329 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001 ,
		_w9908_,
		_w11602_,
		_w23377_
	);
	LUT4 #(
		.INIT('h0020)
	) name19330 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23378_
	);
	LUT2 #(
		.INIT('he)
	) name19331 (
		_w23377_,
		_w23378_,
		_w23379_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19332 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001 ,
		_w9908_,
		_w11602_,
		_w23380_
	);
	LUT4 #(
		.INIT('h0020)
	) name19333 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23381_
	);
	LUT2 #(
		.INIT('he)
	) name19334 (
		_w23380_,
		_w23381_,
		_w23382_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19335 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001 ,
		_w9908_,
		_w11602_,
		_w23383_
	);
	LUT4 #(
		.INIT('h0020)
	) name19336 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23384_
	);
	LUT2 #(
		.INIT('he)
	) name19337 (
		_w23383_,
		_w23384_,
		_w23385_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19338 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001 ,
		_w9908_,
		_w11602_,
		_w23386_
	);
	LUT4 #(
		.INIT('h0040)
	) name19339 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w9908_,
		_w11602_,
		_w23387_
	);
	LUT2 #(
		.INIT('he)
	) name19340 (
		_w23386_,
		_w23387_,
		_w23388_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19341 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001 ,
		_w9908_,
		_w11602_,
		_w23389_
	);
	LUT4 #(
		.INIT('h0020)
	) name19342 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23390_
	);
	LUT2 #(
		.INIT('he)
	) name19343 (
		_w23389_,
		_w23390_,
		_w23391_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19344 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001 ,
		_w9908_,
		_w11602_,
		_w23392_
	);
	LUT4 #(
		.INIT('h0020)
	) name19345 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23393_
	);
	LUT2 #(
		.INIT('he)
	) name19346 (
		_w23392_,
		_w23393_,
		_w23394_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19347 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001 ,
		_w9908_,
		_w11602_,
		_w23395_
	);
	LUT4 #(
		.INIT('h0020)
	) name19348 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23396_
	);
	LUT2 #(
		.INIT('he)
	) name19349 (
		_w23395_,
		_w23396_,
		_w23397_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19350 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001 ,
		_w9908_,
		_w11602_,
		_w23398_
	);
	LUT4 #(
		.INIT('h0020)
	) name19351 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23399_
	);
	LUT2 #(
		.INIT('he)
	) name19352 (
		_w23398_,
		_w23399_,
		_w23400_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19353 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001 ,
		_w9908_,
		_w11602_,
		_w23401_
	);
	LUT4 #(
		.INIT('h0020)
	) name19354 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23402_
	);
	LUT2 #(
		.INIT('he)
	) name19355 (
		_w23401_,
		_w23402_,
		_w23403_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19356 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001 ,
		_w9908_,
		_w11602_,
		_w23404_
	);
	LUT4 #(
		.INIT('h0020)
	) name19357 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23405_
	);
	LUT2 #(
		.INIT('he)
	) name19358 (
		_w23404_,
		_w23405_,
		_w23406_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19359 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001 ,
		_w9908_,
		_w11602_,
		_w23407_
	);
	LUT4 #(
		.INIT('h0020)
	) name19360 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23408_
	);
	LUT2 #(
		.INIT('he)
	) name19361 (
		_w23407_,
		_w23408_,
		_w23409_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19362 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001 ,
		_w9908_,
		_w11602_,
		_w23410_
	);
	LUT4 #(
		.INIT('h0020)
	) name19363 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23411_
	);
	LUT2 #(
		.INIT('he)
	) name19364 (
		_w23410_,
		_w23411_,
		_w23412_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19365 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001 ,
		_w9908_,
		_w11602_,
		_w23413_
	);
	LUT4 #(
		.INIT('h0020)
	) name19366 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23414_
	);
	LUT2 #(
		.INIT('he)
	) name19367 (
		_w23413_,
		_w23414_,
		_w23415_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19368 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001 ,
		_w9908_,
		_w11602_,
		_w23416_
	);
	LUT4 #(
		.INIT('h0020)
	) name19369 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w9908_,
		_w11602_,
		_w23417_
	);
	LUT2 #(
		.INIT('he)
	) name19370 (
		_w23416_,
		_w23417_,
		_w23418_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name19371 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001 ,
		_w9908_,
		_w11602_,
		_w23419_
	);
	LUT4 #(
		.INIT('h0040)
	) name19372 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w9908_,
		_w11602_,
		_w23420_
	);
	LUT2 #(
		.INIT('he)
	) name19373 (
		_w23419_,
		_w23420_,
		_w23421_
	);
	LUT4 #(
		.INIT('hccac)
	) name19374 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001 ,
		_w9912_,
		_w11602_,
		_w23422_
	);
	LUT4 #(
		.INIT('hccac)
	) name19375 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001 ,
		_w9912_,
		_w11602_,
		_w23423_
	);
	LUT4 #(
		.INIT('haaca)
	) name19376 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001 ,
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w9912_,
		_w11602_,
		_w23424_
	);
	LUT4 #(
		.INIT('haa3a)
	) name19377 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001 ,
		_w4155_,
		_w9912_,
		_w11602_,
		_w23425_
	);
	LUT4 #(
		.INIT('haaca)
	) name19378 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w9912_,
		_w11602_,
		_w23426_
	);
	LUT4 #(
		.INIT('haaca)
	) name19379 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w9912_,
		_w11602_,
		_w23427_
	);
	LUT4 #(
		.INIT('haaca)
	) name19380 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w9912_,
		_w11602_,
		_w23428_
	);
	LUT4 #(
		.INIT('haaca)
	) name19381 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w9912_,
		_w11602_,
		_w23429_
	);
	LUT4 #(
		.INIT('hccac)
	) name19382 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001 ,
		_w9912_,
		_w11602_,
		_w23430_
	);
	LUT4 #(
		.INIT('hccac)
	) name19383 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001 ,
		_w9912_,
		_w11602_,
		_w23431_
	);
	LUT4 #(
		.INIT('hccac)
	) name19384 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001 ,
		_w9912_,
		_w11602_,
		_w23432_
	);
	LUT4 #(
		.INIT('hccac)
	) name19385 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001 ,
		_w9912_,
		_w11602_,
		_w23433_
	);
	LUT4 #(
		.INIT('hccac)
	) name19386 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001 ,
		_w9912_,
		_w11602_,
		_w23434_
	);
	LUT4 #(
		.INIT('haaca)
	) name19387 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001 ,
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w9912_,
		_w11602_,
		_w23435_
	);
	LUT4 #(
		.INIT('hccac)
	) name19388 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001 ,
		_w9912_,
		_w11602_,
		_w23436_
	);
	LUT4 #(
		.INIT('h03aa)
	) name19389 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001 ,
		_w11332_,
		_w11598_,
		_w11830_,
		_w23437_
	);
	LUT4 #(
		.INIT('hccac)
	) name19390 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001 ,
		_w9912_,
		_w11602_,
		_w23438_
	);
	LUT4 #(
		.INIT('hccac)
	) name19391 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001 ,
		_w9912_,
		_w11602_,
		_w23439_
	);
	LUT2 #(
		.INIT('h8)
	) name19392 (
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w11610_,
		_w23440_
	);
	LUT3 #(
		.INIT('h08)
	) name19393 (
		_w5760_,
		_w11607_,
		_w11613_,
		_w23441_
	);
	LUT2 #(
		.INIT('he)
	) name19394 (
		_w23440_,
		_w23441_,
		_w23442_
	);
	LUT4 #(
		.INIT('hccac)
	) name19395 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001 ,
		_w9912_,
		_w11602_,
		_w23443_
	);
	LUT4 #(
		.INIT('hccac)
	) name19396 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001 ,
		_w9912_,
		_w11602_,
		_w23444_
	);
	LUT4 #(
		.INIT('hccac)
	) name19397 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001 ,
		_w9912_,
		_w11602_,
		_w23445_
	);
	LUT4 #(
		.INIT('hccac)
	) name19398 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001 ,
		_w9912_,
		_w11602_,
		_w23446_
	);
	LUT4 #(
		.INIT('hccac)
	) name19399 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001 ,
		_w9912_,
		_w11602_,
		_w23447_
	);
	LUT4 #(
		.INIT('hccac)
	) name19400 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001 ,
		_w9912_,
		_w11602_,
		_w23448_
	);
	LUT4 #(
		.INIT('hccac)
	) name19401 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001 ,
		_w9912_,
		_w11602_,
		_w23449_
	);
	LUT4 #(
		.INIT('hcddd)
	) name19402 (
		_w4065_,
		_w16153_,
		_w19997_,
		_w21216_,
		_w23450_
	);
	LUT2 #(
		.INIT('h8)
	) name19403 (
		\T_TMODE[1]_pad ,
		\core_c_dec_PPclr_reg/P0001 ,
		_w23451_
	);
	LUT3 #(
		.INIT('hf1)
	) name19404 (
		_w19773_,
		_w19774_,
		_w23451_,
		_w23452_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19405 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\T_PIOin[0]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23453_
	);
	LUT4 #(
		.INIT('h8000)
	) name19406 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[0]/P0001 ,
		_w23454_
	);
	LUT2 #(
		.INIT('he)
	) name19407 (
		_w23453_,
		_w23454_,
		_w23455_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19408 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\T_PIOin[10]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23456_
	);
	LUT4 #(
		.INIT('h8000)
	) name19409 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[10]/P0001 ,
		_w23457_
	);
	LUT2 #(
		.INIT('he)
	) name19410 (
		_w23456_,
		_w23457_,
		_w23458_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19411 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\T_PIOin[11]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23459_
	);
	LUT4 #(
		.INIT('h8000)
	) name19412 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[11]/P0001 ,
		_w23460_
	);
	LUT2 #(
		.INIT('he)
	) name19413 (
		_w23459_,
		_w23460_,
		_w23461_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19414 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\T_PIOin[1]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23462_
	);
	LUT4 #(
		.INIT('h8000)
	) name19415 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[1]/P0001 ,
		_w23463_
	);
	LUT2 #(
		.INIT('he)
	) name19416 (
		_w23462_,
		_w23463_,
		_w23464_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19417 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\T_PIOin[2]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23465_
	);
	LUT4 #(
		.INIT('h8000)
	) name19418 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[2]/P0001 ,
		_w23466_
	);
	LUT2 #(
		.INIT('he)
	) name19419 (
		_w23465_,
		_w23466_,
		_w23467_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19420 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\T_PIOin[3]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23468_
	);
	LUT4 #(
		.INIT('h8000)
	) name19421 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[3]/P0001 ,
		_w23469_
	);
	LUT2 #(
		.INIT('he)
	) name19422 (
		_w23468_,
		_w23469_,
		_w23470_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19423 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\T_PIOin[4]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23471_
	);
	LUT4 #(
		.INIT('h8000)
	) name19424 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[4]/P0001 ,
		_w23472_
	);
	LUT2 #(
		.INIT('he)
	) name19425 (
		_w23471_,
		_w23472_,
		_w23473_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19426 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\T_PIOin[5]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23474_
	);
	LUT4 #(
		.INIT('h8000)
	) name19427 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[5]/P0001 ,
		_w23475_
	);
	LUT2 #(
		.INIT('he)
	) name19428 (
		_w23474_,
		_w23475_,
		_w23476_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19429 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\T_PIOin[6]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23477_
	);
	LUT4 #(
		.INIT('h8000)
	) name19430 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[6]/P0001 ,
		_w23478_
	);
	LUT2 #(
		.INIT('he)
	) name19431 (
		_w23477_,
		_w23478_,
		_w23479_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19432 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\T_PIOin[7]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23480_
	);
	LUT4 #(
		.INIT('h8000)
	) name19433 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[7]/P0001 ,
		_w23481_
	);
	LUT2 #(
		.INIT('he)
	) name19434 (
		_w23480_,
		_w23481_,
		_w23482_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19435 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\T_PIOin[8]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23483_
	);
	LUT4 #(
		.INIT('h8000)
	) name19436 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[8]/P0001 ,
		_w23484_
	);
	LUT2 #(
		.INIT('he)
	) name19437 (
		_w23483_,
		_w23484_,
		_w23485_
	);
	LUT4 #(
		.INIT('h70f0)
	) name19438 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\T_PIOin[9]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		_w23486_
	);
	LUT4 #(
		.INIT('h8000)
	) name19439 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_IN_P_reg[9]/P0001 ,
		_w23487_
	);
	LUT2 #(
		.INIT('he)
	) name19440 (
		_w23486_,
		_w23487_,
		_w23488_
	);
	LUT4 #(
		.INIT('h7f00)
	) name19441 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[0]/NET0131 ,
		_w23489_
	);
	LUT4 #(
		.INIT('h8000)
	) name19442 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[0]/P0001 ,
		_w23490_
	);
	LUT2 #(
		.INIT('he)
	) name19443 (
		_w23489_,
		_w23490_,
		_w23491_
	);
	LUT4 #(
		.INIT('h7f00)
	) name19444 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[10]/NET0131 ,
		_w23492_
	);
	LUT4 #(
		.INIT('h8000)
	) name19445 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[10]/P0001 ,
		_w23493_
	);
	LUT2 #(
		.INIT('he)
	) name19446 (
		_w23492_,
		_w23493_,
		_w23494_
	);
	LUT4 #(
		.INIT('h7f00)
	) name19447 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[2]/NET0131 ,
		_w23495_
	);
	LUT4 #(
		.INIT('h8000)
	) name19448 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[2]/P0001 ,
		_w23496_
	);
	LUT2 #(
		.INIT('he)
	) name19449 (
		_w23495_,
		_w23496_,
		_w23497_
	);
	LUT4 #(
		.INIT('h7f00)
	) name19450 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[4]/NET0131 ,
		_w23498_
	);
	LUT4 #(
		.INIT('h8000)
	) name19451 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[4]/P0001 ,
		_w23499_
	);
	LUT2 #(
		.INIT('he)
	) name19452 (
		_w23498_,
		_w23499_,
		_w23500_
	);
	LUT4 #(
		.INIT('h7f00)
	) name19453 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_reg[6]/NET0131 ,
		_w23501_
	);
	LUT4 #(
		.INIT('h8000)
	) name19454 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		\memc_MMR_web_reg/NET0131 ,
		\pio_PIO_RES_OUT_reg[6]/P0001 ,
		_w23502_
	);
	LUT2 #(
		.INIT('he)
	) name19455 (
		_w23501_,
		_w23502_,
		_w23503_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name19456 (
		\sice_GO_NXi_reg/NET0131 ,
		\sice_SPC_reg[20]/P0001 ,
		_w14459_,
		_w14460_,
		_w23504_
	);
	LUT4 #(
		.INIT('h1d00)
	) name19457 (
		\T_RD0_pad ,
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w9377_,
		_w18895_,
		_w23505_
	);
	LUT4 #(
		.INIT('h3302)
	) name19458 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[0]/P0001 ,
		_w18892_,
		_w18894_,
		_w23506_
	);
	LUT2 #(
		.INIT('h1)
	) name19459 (
		_w23505_,
		_w23506_,
		_w23507_
	);
	LUT4 #(
		.INIT('hcc08)
	) name19460 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RXSHT_reg[1]/P0001 ,
		_w18892_,
		_w18894_,
		_w23508_
	);
	LUT2 #(
		.INIT('he)
	) name19461 (
		_w18896_,
		_w23508_,
		_w23509_
	);
	LUT4 #(
		.INIT('h1d00)
	) name19462 (
		\T_RD1_pad ,
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w9403_,
		_w18881_,
		_w23510_
	);
	LUT4 #(
		.INIT('h3302)
	) name19463 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[0]/P0001 ,
		_w18878_,
		_w18880_,
		_w23511_
	);
	LUT2 #(
		.INIT('h1)
	) name19464 (
		_w23510_,
		_w23511_,
		_w23512_
	);
	LUT4 #(
		.INIT('hcc08)
	) name19465 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RXSHT_reg[1]/P0001 ,
		_w18878_,
		_w18880_,
		_w23513_
	);
	LUT2 #(
		.INIT('he)
	) name19466 (
		_w18882_,
		_w23513_,
		_w23514_
	);
	assign CLKO_pad = _w4059_ ;
	assign \CMAinx[0]_pad  = _w4525_ ;
	assign \CMAinx[10]_pad  = _w4546_ ;
	assign \CMAinx[11]_pad  = _w4561_ ;
	assign \CMAinx[1]_pad  = _w4576_ ;
	assign \CMAinx[2]_pad  = _w4599_ ;
	assign \CMAinx[3]_pad  = _w4620_ ;
	assign \CMAinx[4]_pad  = _w4639_ ;
	assign \CMAinx[5]_pad  = _w4657_ ;
	assign \CMAinx[6]_pad  = _w4672_ ;
	assign \CMAinx[7]_pad  = _w4687_ ;
	assign \CMAinx[8]_pad  = _w4702_ ;
	assign \CMAinx[9]_pad  = _w4717_ ;
	assign CMSn_pad = _w4808_ ;
	assign CM_cs_pad = _w4883_ ;
	assign \CM_wd[0]_pad  = _w4889_ ;
	assign \CM_wd[10]_pad  = _w4891_ ;
	assign \CM_wd[11]_pad  = _w4893_ ;
	assign \CM_wd[12]_pad  = _w4895_ ;
	assign \CM_wd[13]_pad  = _w4897_ ;
	assign \CM_wd[14]_pad  = _w4899_ ;
	assign \CM_wd[15]_pad  = _w4901_ ;
	assign \CM_wd[16]_pad  = _w4903_ ;
	assign \CM_wd[17]_pad  = _w4905_ ;
	assign \CM_wd[18]_pad  = _w4907_ ;
	assign \CM_wd[19]_pad  = _w4909_ ;
	assign \CM_wd[1]_pad  = _w4911_ ;
	assign \CM_wd[20]_pad  = _w4913_ ;
	assign \CM_wd[21]_pad  = _w4915_ ;
	assign \CM_wd[22]_pad  = _w4917_ ;
	assign \CM_wd[23]_pad  = _w4919_ ;
	assign \CM_wd[2]_pad  = _w4921_ ;
	assign \CM_wd[3]_pad  = _w4923_ ;
	assign \CM_wd[4]_pad  = _w4925_ ;
	assign \CM_wd[5]_pad  = _w4927_ ;
	assign \CM_wd[6]_pad  = _w4929_ ;
	assign \CM_wd[7]_pad  = _w4931_ ;
	assign \CM_wd[8]_pad  = _w4933_ ;
	assign \CM_wd[9]_pad  = _w4935_ ;
	assign CM_web_pad = _w4945_ ;
	assign \CMo_cs0_pad  = _w4958_ ;
	assign \CMo_cs1_pad  = _w4959_ ;
	assign \CMo_cs2_pad  = _w4960_ ;
	assign \CMo_cs3_pad  = _w4961_ ;
	assign \CMo_cs4_pad  = _w4962_ ;
	assign \CMo_cs5_pad  = _w4963_ ;
	assign \CMo_cs6_pad  = _w4964_ ;
	assign \CMo_cs7_pad  = _w4965_ ;
	assign \DMAinx[0]_pad  = _w5917_ ;
	assign \DMAinx[10]_pad  = _w6242_ ;
	assign \DMAinx[11]_pad  = _w6571_ ;
	assign \DMAinx[12]_pad  = _w6902_ ;
	assign \DMAinx[13]_pad  = _w6945_ ;
	assign \DMAinx[1]_pad  = _w6986_ ;
	assign \DMAinx[2]_pad  = _w7024_ ;
	assign \DMAinx[3]_pad  = _w7061_ ;
	assign \DMAinx[4]_pad  = _w7382_ ;
	assign \DMAinx[5]_pad  = _w7714_ ;
	assign \DMAinx[6]_pad  = _w8048_ ;
	assign \DMAinx[7]_pad  = _w8087_ ;
	assign \DMAinx[8]_pad  = _w8125_ ;
	assign \DMAinx[9]_pad  = _w8166_ ;
	assign DMSn_pad = _w4802_ ;
	assign DM_cs_pad = _w8195_ ;
	assign \DM_wd[0]_pad  = _w8204_ ;
	assign \DM_wd[10]_pad  = _w8212_ ;
	assign \DM_wd[11]_pad  = _w8220_ ;
	assign \DM_wd[12]_pad  = _w8228_ ;
	assign \DM_wd[13]_pad  = _w8236_ ;
	assign \DM_wd[14]_pad  = _w8317_ ;
	assign \DM_wd[15]_pad  = _w8396_ ;
	assign \DM_wd[1]_pad  = _w8403_ ;
	assign \DM_wd[2]_pad  = _w8410_ ;
	assign \DM_wd[3]_pad  = _w8417_ ;
	assign \DM_wd[4]_pad  = _w8424_ ;
	assign \DM_wd[5]_pad  = _w8431_ ;
	assign \DM_wd[6]_pad  = _w8438_ ;
	assign \DM_wd[7]_pad  = _w8445_ ;
	assign \DM_wd[8]_pad  = _w8453_ ;
	assign \DM_wd[9]_pad  = _w8461_ ;
	assign \DMo_cs0_pad  = _w8471_ ;
	assign \DMo_cs1_pad  = _w8473_ ;
	assign \DMo_cs2_pad  = _w8474_ ;
	assign \DMo_cs3_pad  = _w8475_ ;
	assign \DMo_cs4_pad  = _w8477_ ;
	assign \DMo_cs5_pad  = _w8479_ ;
	assign \DMo_cs6_pad  = _w8480_ ;
	assign \DMo_cs7_pad  = _w8481_ ;
	assign \DSPCLK_cm1_pad  = _w8492_ ;
	assign \EA_do[0]_pad  = _w8499_ ;
	assign \EA_do[10]_pad  = _w8505_ ;
	assign \EA_do[12]_pad  = _w8518_ ;
	assign \EA_do[13]_pad  = _w8529_ ;
	assign \EA_do[14]_pad  = _w8539_ ;
	assign \EA_do[1]_pad  = _w8545_ ;
	assign \EA_do[2]_pad  = _w8551_ ;
	assign \EA_do[3]_pad  = _w8557_ ;
	assign \EA_do[4]_pad  = _w8563_ ;
	assign \EA_do[5]_pad  = _w8569_ ;
	assign \EA_do[6]_pad  = _w8575_ ;
	assign \EA_do[7]_pad  = _w8581_ ;
	assign \EA_do[8]_pad  = _w8587_ ;
	assign \EA_do[9]_pad  = _w8593_ ;
	assign EA_oe_pad = _w8600_ ;
	assign \ED_do[0]_pad  = _w8651_ ;
	assign \ED_do[10]_pad  = _w8674_ ;
	assign \ED_do[11]_pad  = _w8697_ ;
	assign \ED_do[12]_pad  = _w8720_ ;
	assign \ED_do[13]_pad  = _w8743_ ;
	assign \ED_do[14]_pad  = _w8784_ ;
	assign \ED_do[15]_pad  = _w8823_ ;
	assign \ED_do[1]_pad  = _w8845_ ;
	assign \ED_do[2]_pad  = _w8867_ ;
	assign \ED_do[3]_pad  = _w8889_ ;
	assign \ED_do[4]_pad  = _w8911_ ;
	assign \ED_do[5]_pad  = _w8933_ ;
	assign \ED_do[6]_pad  = _w8956_ ;
	assign \ED_do[7]_pad  = _w8978_ ;
	assign \ED_do[8]_pad  = _w9001_ ;
	assign \ED_do[9]_pad  = _w9024_ ;
	assign \ED_oe_14_8_pad  = _w9025_ ;
	assign \ED_oe_7_0_pad  = _w9026_ ;
	assign \IAD_do[0]_pad  = _w9029_ ;
	assign \IAD_do[10]_pad  = _w9030_ ;
	assign \IAD_do[11]_pad  = _w9031_ ;
	assign \IAD_do[12]_pad  = _w9032_ ;
	assign \IAD_do[13]_pad  = _w9033_ ;
	assign \IAD_do[14]_pad  = _w9034_ ;
	assign \IAD_do[15]_pad  = _w9035_ ;
	assign \IAD_do[1]_pad  = _w9038_ ;
	assign \IAD_do[2]_pad  = _w9041_ ;
	assign \IAD_do[3]_pad  = _w9044_ ;
	assign \IAD_do[4]_pad  = _w9047_ ;
	assign \IAD_do[5]_pad  = _w9050_ ;
	assign \IAD_do[6]_pad  = _w9053_ ;
	assign \IAD_do[7]_pad  = _w9056_ ;
	assign \IAD_do[8]_pad  = _w9057_ ;
	assign \IAD_do[9]_pad  = _w9058_ ;
	assign IAD_oe_pad = _w9059_ ;
	assign IDoe_pad = _w9060_ ;
	assign IOSn_pad = _w4800_ ;
	assign \PMAinx[0]_pad  = _w9095_ ;
	assign \PMAinx[10]_pad  = _w9108_ ;
	assign \PMAinx[11]_pad  = _w9121_ ;
	assign \PMAinx[1]_pad  = _w9134_ ;
	assign \PMAinx[2]_pad  = _w9147_ ;
	assign \PMAinx[3]_pad  = _w9159_ ;
	assign \PMAinx[4]_pad  = _w9171_ ;
	assign \PMAinx[5]_pad  = _w9183_ ;
	assign \PMAinx[6]_pad  = _w9195_ ;
	assign \PMAinx[7]_pad  = _w9207_ ;
	assign \PMAinx[8]_pad  = _w9220_ ;
	assign \PMAinx[9]_pad  = _w9233_ ;
	assign \PM_wd[0]_pad  = _w9238_ ;
	assign \PM_wd[10]_pad  = _w9241_ ;
	assign \PM_wd[11]_pad  = _w9244_ ;
	assign \PM_wd[12]_pad  = _w9247_ ;
	assign \PM_wd[13]_pad  = _w9250_ ;
	assign \PM_wd[14]_pad  = _w9253_ ;
	assign \PM_wd[15]_pad  = _w9256_ ;
	assign \PM_wd[1]_pad  = _w9259_ ;
	assign \PM_wd[2]_pad  = _w9262_ ;
	assign \PM_wd[3]_pad  = _w9265_ ;
	assign \PM_wd[4]_pad  = _w9268_ ;
	assign \PM_wd[5]_pad  = _w9271_ ;
	assign \PM_wd[6]_pad  = _w9274_ ;
	assign \PM_wd[7]_pad  = _w9277_ ;
	assign \PM_wd[8]_pad  = _w9280_ ;
	assign \PM_wd[9]_pad  = _w9283_ ;
	assign \PMo_cs0_pad  = _w9337_ ;
	assign \PMo_cs1_pad  = _w9340_ ;
	assign \PMo_cs2_pad  = _w9342_ ;
	assign \PMo_cs3_pad  = _w9344_ ;
	assign \PMo_cs4_pad  = _w9346_ ;
	assign \PMo_cs5_pad  = _w9347_ ;
	assign \PMo_cs6_pad  = _w9348_ ;
	assign \PMo_cs7_pad  = _w9349_ ;
	assign \PMo_oe0_pad  = 1'b1;
	assign \RFS0_pad  = _w9351_ ;
	assign \RFS1_pad  = _w9353_ ;
	assign \SCLK0_pad  = _w9354_ ;
	assign \SCLK1_pad  = _w9355_ ;
	assign \TD0_pad  = _w9378_ ;
	assign \TD1_pad  = _w9404_ ;
	assign \TFS0_pad  = _w9406_ ;
	assign \TFS1_pad  = _w9408_ ;
	assign \T_ISn_syn_2  = _w560_ ;
	assign WRn_pad = _w9409_ ;
	assign XTALoffn_pad = _w8487_ ;
	assign \_al_n0  = 1'b0;
	assign \bdma_BDMA_boot_reg/NET0131_reg_syn_3  = _w9425_ ;
	assign \bdma_BDMA_boot_reg/n0  = _w9410_ ;
	assign \bdma_BM_cyc_reg/P0000  = _w646_ ;
	assign \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_3  = _w9435_ ;
	assign \core_c_psq_MGNT_reg/P0001  = _w1137_ ;
	assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001_reg_syn_3  = _w9441_ ;
	assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001_reg_syn_3  = _w9444_ ;
	assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001_reg_syn_3  = _w9447_ ;
	assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001_reg_syn_3  = _w9450_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001_reg_syn_3  = _w9770_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001_reg_syn_3  = _w9837_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001_reg_syn_3  = _w9849_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001_reg_syn_3  = _w9856_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001_reg_syn_3  = _w9868_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001_reg_syn_3  = _w9880_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001_reg_syn_3  = _w9892_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001_reg_syn_3  = _w9896_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001_reg_syn_3  = _w9899_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001_reg_syn_3  = _w9900_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001_reg_syn_3  = _w9901_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001_reg_syn_3  = _w9902_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001_reg_syn_3  = _w9903_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001_reg_syn_3  = _w9904_ ;
	assign \core_eu_ec_cun_MVi_pre_C_reg/P0001_reg_syn_3  = _w9930_ ;
	assign \core_eu_em_mac_em_reg_Sq_E_reg/P0001_reg_syn_3  = _w9935_ ;
	assign \emc_DMDreg_reg[8]/P0001_reg_syn_3  = _w9941_ ;
	assign \emc_DMDreg_reg[9]/P0001_reg_syn_3  = _w9942_ ;
	assign \emc_ECMcs_reg/P0001  = _w2951_ ;
	assign \emc_PMDreg_reg[8]/P0001_reg_syn_3  = _w9944_ ;
	assign \emc_PMDreg_reg[9]/P0001_reg_syn_3  = _w9945_ ;
	assign \g10/_0_  = _w11327_ ;
	assign \g1000/_0_  = _w11599_ ;
	assign \g10000/_0_  = _w11603_ ;
	assign \g10001/_0_  = _w11616_ ;
	assign \g10002/_0_  = _w11617_ ;
	assign \g10003/_0_  = _w11618_ ;
	assign \g10004/_0_  = _w11619_ ;
	assign \g10005/_0_  = _w11620_ ;
	assign \g10007/_0_  = _w11621_ ;
	assign \g10008/_0_  = _w11622_ ;
	assign \g10009/_0_  = _w11623_ ;
	assign \g1001/_3_  = _w11642_ ;
	assign \g10010/_0_  = _w11643_ ;
	assign \g10011/_0_  = _w11644_ ;
	assign \g10012/_0_  = _w11645_ ;
	assign \g10013/_0_  = _w11646_ ;
	assign \g10014/_0_  = _w11647_ ;
	assign \g10015/_0_  = _w11648_ ;
	assign \g10016/_0_  = _w11649_ ;
	assign \g10017/_0_  = _w11650_ ;
	assign \g10018/_0_  = _w11651_ ;
	assign \g10019/_0_  = _w11652_ ;
	assign \g1002/_3_  = _w11662_ ;
	assign \g10020/_0_  = _w11663_ ;
	assign \g10021/_0_  = _w11664_ ;
	assign \g10022/_0_  = _w11665_ ;
	assign \g10023/_0_  = _w11666_ ;
	assign \g10024/_0_  = _w11667_ ;
	assign \g10025/_0_  = _w11668_ ;
	assign \g10026/_0_  = _w11669_ ;
	assign \g10027/_0_  = _w11670_ ;
	assign \g10028/_0_  = _w11671_ ;
	assign \g10029/_0_  = _w11672_ ;
	assign \g1003/_0_  = _w11744_ ;
	assign \g10030/_0_  = _w11745_ ;
	assign \g10031/_0_  = _w11746_ ;
	assign \g10032/_0_  = _w11747_ ;
	assign \g10033/_0_  = _w11748_ ;
	assign \g10034/_0_  = _w11749_ ;
	assign \g10035/_0_  = _w11750_ ;
	assign \g10036/_0_  = _w11751_ ;
	assign \g10037/_0_  = _w11752_ ;
	assign \g10038/_0_  = _w11753_ ;
	assign \g10039/_0_  = _w11754_ ;
	assign \g10040/_0_  = _w11755_ ;
	assign \g10041/_0_  = _w11756_ ;
	assign \g10042/_0_  = _w11757_ ;
	assign \g10043/_0_  = _w11758_ ;
	assign \g10044/_0_  = _w11759_ ;
	assign \g10045/_0_  = _w11760_ ;
	assign \g10046/_0_  = _w11761_ ;
	assign \g10047/_0_  = _w11762_ ;
	assign \g10048/_0_  = _w11763_ ;
	assign \g10049/_0_  = _w11764_ ;
	assign \g10050/_0_  = _w11765_ ;
	assign \g10051/_0_  = _w11766_ ;
	assign \g10052/_0_  = _w11767_ ;
	assign \g10053/_0_  = _w11768_ ;
	assign \g10054/_0_  = _w11769_ ;
	assign \g10055/_0_  = _w11770_ ;
	assign \g10056/_0_  = _w11771_ ;
	assign \g10057/_0_  = _w11772_ ;
	assign \g10058/_0_  = _w11773_ ;
	assign \g10059/_0_  = _w11774_ ;
	assign \g10060/_0_  = _w11775_ ;
	assign \g10061/_0_  = _w11776_ ;
	assign \g10062/_0_  = _w11777_ ;
	assign \g10063/_0_  = _w11778_ ;
	assign \g10064/_0_  = _w11779_ ;
	assign \g10065/_0_  = _w11780_ ;
	assign \g10066/_0_  = _w11781_ ;
	assign \g10067/_0_  = _w11782_ ;
	assign \g10068/_0_  = _w11783_ ;
	assign \g10069/_0_  = _w11784_ ;
	assign \g10070/_0_  = _w11785_ ;
	assign \g10071/_0_  = _w11786_ ;
	assign \g10072/_0_  = _w11791_ ;
	assign \g10073/_0_  = _w11792_ ;
	assign \g10074/_0_  = _w11793_ ;
	assign \g10075/_0_  = _w11794_ ;
	assign \g10076/_0_  = _w11795_ ;
	assign \g10077/_0_  = _w11798_ ;
	assign \g10078/_0_  = _w11799_ ;
	assign \g10080/_0_  = _w11800_ ;
	assign \g10081/_0_  = _w11805_ ;
	assign \g10083/_0_  = _w11808_ ;
	assign \g10089/_0_  = _w11811_ ;
	assign \g1009/_0_  = _w11814_ ;
	assign \g10090/_0_  = _w11817_ ;
	assign \g10091/_0_  = _w11820_ ;
	assign \g10092/_0_  = _w11823_ ;
	assign \g10093/_0_  = _w11826_ ;
	assign \g10094/_0_  = _w11829_ ;
	assign \g1010/_0_  = _w11916_ ;
	assign \g10108/_3_  = _w11929_ ;
	assign \g1011/_0_  = _w11930_ ;
	assign \g10110/_0_  = _w11933_ ;
	assign \g10111/_0_  = _w11937_ ;
	assign \g10113/_3_  = _w11939_ ;
	assign \g10115/_3_  = _w11941_ ;
	assign \g1013/_0_  = _w11944_ ;
	assign \g1014/_0_  = _w11983_ ;
	assign \g10152/_0_  = _w11988_ ;
	assign \g10153/_0_  = _w11991_ ;
	assign \g10154/_0_  = _w11994_ ;
	assign \g10155/_0_  = _w11995_ ;
	assign \g10156/_0_  = _w11998_ ;
	assign \g10157/_0_  = _w12001_ ;
	assign \g10158/_0_  = _w12004_ ;
	assign \g10159/_0_  = _w12005_ ;
	assign \g1016/_0_  = _w12029_ ;
	assign \g10160/_0_  = _w12033_ ;
	assign \g10161/_0_  = _w12036_ ;
	assign \g10162/_0_  = _w12039_ ;
	assign \g10163/_0_  = _w12041_ ;
	assign \g10164/_0_  = _w12044_ ;
	assign \g10165/_0_  = _w12047_ ;
	assign \g1017/_0_  = _w12049_ ;
	assign \g10170/_3_  = _w12063_ ;
	assign \g1018/_0_  = _w12064_ ;
	assign \g10190/_3_  = _w12065_ ;
	assign \g10194/_3_  = _w12066_ ;
	assign \g10198/_0_  = _w12088_ ;
	assign \g10199/_0_  = _w12110_ ;
	assign \g102/_0_  = _w12214_ ;
	assign \g103/_0_  = _w12229_ ;
	assign \g104/_0_  = _w12236_ ;
	assign \g105/_0_  = _w12240_ ;
	assign \g10598/_0_  = _w12242_ ;
	assign \g106/_0_  = _w12249_ ;
	assign \g10667/_0_  = _w12251_ ;
	assign \g10683/_0_  = _w12266_ ;
	assign \g10685/_0_  = _w12281_ ;
	assign \g107/_0_  = _w12295_ ;
	assign \g10721/_0_  = _w12300_ ;
	assign \g10758/_0_  = _w12303_ ;
	assign \g10765/_0_  = _w12305_ ;
	assign \g10778/_0_  = _w12313_ ;
	assign \g10791/_0_  = _w12314_ ;
	assign \g108/_0_  = _w12388_ ;
	assign \g10887/_0_  = _w12399_ ;
	assign \g1089/_0_  = _w12438_ ;
	assign \g109/_0_  = _w12445_ ;
	assign \g1090/_0_  = _w12484_ ;
	assign \g1091/_0_  = _w12521_ ;
	assign \g1092/_0_  = _w12524_ ;
	assign \g10923/_0_  = _w12526_ ;
	assign \g1093/_0_  = _w12527_ ;
	assign \g10930/_0_  = _w12531_ ;
	assign \g10931/_0_  = _w12532_ ;
	assign \g10936/_0_  = _w12536_ ;
	assign \g1097/_0_  = _w12539_ ;
	assign \g11/_0_  = _w12554_ ;
	assign \g110/_0_  = _w12559_ ;
	assign \g1101/_0_  = _w12603_ ;
	assign \g11013/_0_  = _w12607_ ;
	assign \g1102/_0_  = _w12614_ ;
	assign \g1103/_0_  = _w12617_ ;
	assign \g11032/_0_  = _w12625_ ;
	assign \g1104/_0_  = _w12671_ ;
	assign \g1105/_0_  = _w12699_ ;
	assign \g1107/_0_  = _w12702_ ;
	assign \g11074/_0_  = _w12712_ ;
	assign \g11077/_0_  = _w12714_ ;
	assign \g1108/_0_  = _w12717_ ;
	assign \g1109/_0_  = _w12720_ ;
	assign \g11112/_0_  = _w12726_ ;
	assign \g11115/_0_  = _w12728_ ;
	assign \g11116/_0_  = _w12730_ ;
	assign \g11119/_0_  = _w12734_ ;
	assign \g11120/_0_  = _w12735_ ;
	assign \g1113/_0_  = _w12759_ ;
	assign \g1115/_0_  = _w12782_ ;
	assign \g1116/_0_  = _w12783_ ;
	assign \g1117/_0_  = _w12786_ ;
	assign \g11267/_0_  = _w12787_ ;
	assign \g11281/_0_  = _w12795_ ;
	assign \g11287/_0_  = _w12806_ ;
	assign \g11300/_0_  = _w12810_ ;
	assign \g11323/_0_  = _w12815_ ;
	assign \g11325/_2__syn_2  = _w12822_ ;
	assign \g11345/_2_  = _w12823_ ;
	assign \g11470/_0_  = _w12827_ ;
	assign \g11471/_0_  = _w12835_ ;
	assign \g11472/_0_  = _w12839_ ;
	assign \g11473/_0_  = _w12847_ ;
	assign \g11474/_0_  = _w12851_ ;
	assign \g11476/_0_  = _w12852_ ;
	assign \g11477/_0_  = _w12859_ ;
	assign \g11496/_0_  = _w12864_ ;
	assign \g11497/_0_  = _w12866_ ;
	assign \g11498/_0_  = _w12869_ ;
	assign \g11499/_0_  = _w12871_ ;
	assign \g11500/_0_  = _w12874_ ;
	assign \g11501/_0_  = _w12876_ ;
	assign \g11502/_0_  = _w12879_ ;
	assign \g11503/_0_  = _w12881_ ;
	assign \g11504/_0_  = _w12884_ ;
	assign \g11505/_0_  = _w12887_ ;
	assign \g11506/_0_  = _w12889_ ;
	assign \g11507/_0_  = _w12891_ ;
	assign \g11509/_0_  = _w12892_ ;
	assign \g11510/_0_  = _w12893_ ;
	assign \g11515/_0_  = _w12904_ ;
	assign \g11516/_0_  = _w12905_ ;
	assign \g11520/_0_  = _w12907_ ;
	assign \g11521/_0_  = _w12911_ ;
	assign \g11576/_0_  = _w12921_ ;
	assign \g11577/_0_  = _w12929_ ;
	assign \g11578/_0_  = _w12937_ ;
	assign \g11579/_0_  = _w12945_ ;
	assign \g11580/_0_  = _w12953_ ;
	assign \g11581/_0_  = _w12959_ ;
	assign \g11582/_0_  = _w12967_ ;
	assign \g11583/_0_  = _w12975_ ;
	assign \g11584/_0_  = _w12982_ ;
	assign \g11585/_0_  = _w12989_ ;
	assign \g11586/_0_  = _w12998_ ;
	assign \g11587/_0_  = _w13006_ ;
	assign \g11588/_0_  = _w13014_ ;
	assign \g11589/_0_  = _w13020_ ;
	assign \g11591/_0_  = _w13028_ ;
	assign \g11593/_0_  = _w13035_ ;
	assign \g11595/_0_  = _w13039_ ;
	assign \g11596/_0_  = _w13040_ ;
	assign \g11597/_0_  = _w13041_ ;
	assign \g11605/_0_  = _w13046_ ;
	assign \g11606/_0_  = _w13049_ ;
	assign \g11607/_0_  = _w13052_ ;
	assign \g11608/_0_  = _w13055_ ;
	assign \g11609/_0_  = _w13058_ ;
	assign \g11610/_0_  = _w13061_ ;
	assign \g11611/_0_  = _w13064_ ;
	assign \g11612/_0_  = _w13067_ ;
	assign \g11613/_0_  = _w13068_ ;
	assign \g11615/_0_  = _w13071_ ;
	assign \g11616/_0_  = _w13079_ ;
	assign \g11617/_0_  = _w13080_ ;
	assign \g11651/_3_  = _w13083_ ;
	assign \g11704/_0_  = _w13084_ ;
	assign \g11705/_0_  = _w13085_ ;
	assign \g11709/_0_  = _w13086_ ;
	assign \g11722/_0_  = _w13089_ ;
	assign \g11723/_0_  = _w13090_ ;
	assign \g119/_0_  = _w13094_ ;
	assign \g1192/_0_  = _w13166_ ;
	assign \g11994/_0_  = _w13167_ ;
	assign \g120/_0_  = _w13171_ ;
	assign \g1200/_0_  = _w13203_ ;
	assign \g12003/_0_  = _w13205_ ;
	assign \g1201/_0_  = _w13208_ ;
	assign \g12019/_0_  = _w13210_ ;
	assign \g1203/_3_  = _w13216_ ;
	assign \g1204/_3_  = _w13221_ ;
	assign \g1207/_0_  = _w13252_ ;
	assign \g1208/_0_  = _w13255_ ;
	assign \g12092/_0_  = _w13260_ ;
	assign \g1210/_0_  = _w13284_ ;
	assign \g1211/_0_  = _w13317_ ;
	assign \g1212/_0_  = _w13318_ ;
	assign \g1213/_0_  = _w13321_ ;
	assign \g12145/_0_  = _w13331_ ;
	assign \g12155/_0_  = _w13336_ ;
	assign \g12186/_0_  = _w13341_ ;
	assign \g12187/_0_  = _w13343_ ;
	assign \g12192/_0_  = _w13345_ ;
	assign \g12201/_0_  = _w13352_ ;
	assign \g12202/_0_  = _w13356_ ;
	assign \g12203/_0_  = _w13360_ ;
	assign \g12204/_0_  = _w13363_ ;
	assign \g12207/_0_  = _w13365_ ;
	assign \g12229/_3_  = _w13370_ ;
	assign \g12267/_0_  = _w13371_ ;
	assign \g12276/_0_  = _w13373_ ;
	assign \g12278/_0_  = _w13375_ ;
	assign \g12279/_0_  = _w13377_ ;
	assign \g12280/_0_  = _w13379_ ;
	assign \g12302/_0_  = _w13381_ ;
	assign \g12316/_0_  = _w13387_ ;
	assign \g12317/_0_  = _w13390_ ;
	assign \g12319/_0_  = _w13394_ ;
	assign \g12328/_3_  = _w13398_ ;
	assign \g1233/_0_  = _w7378_ ;
	assign \g12348/_0_  = _w13400_ ;
	assign \g12351/_0_  = _w13403_ ;
	assign \g12352/_0_  = _w13406_ ;
	assign \g12353/_0_  = _w13409_ ;
	assign \g12354/_0_  = _w13412_ ;
	assign \g12355/_0_  = _w13415_ ;
	assign \g1237/_0_  = _w6176_ ;
	assign \g124/_0_  = _w13418_ ;
	assign \g12444/_0_  = _w13421_ ;
	assign \g125/_0_  = _w13424_ ;
	assign \g12637/_0_  = _w13427_ ;
	assign \g12639/_0_  = _w13430_ ;
	assign \g12658/_0_  = _w13435_ ;
	assign \g12659/_0_  = _w13440_ ;
	assign \g12660/_0_  = _w13445_ ;
	assign \g12663/_0_  = _w13449_ ;
	assign \g12664/_0_  = _w13453_ ;
	assign \g12665/_0_  = _w13457_ ;
	assign \g12672/_3_  = _w13462_ ;
	assign \g12673/_3_  = _w13467_ ;
	assign \g12674/_3_  = _w13471_ ;
	assign \g12675/_3_  = _w13476_ ;
	assign \g12676/_3_  = _w13480_ ;
	assign \g12677/_3_  = _w13485_ ;
	assign \g12678/_0_  = _w13488_ ;
	assign \g12679/_3_  = _w13493_ ;
	assign \g12697/_3_  = _w13498_ ;
	assign \g12701/_3_  = _w13503_ ;
	assign \g12711/_2_  = _w13509_ ;
	assign \g12713/_2_  = _w13513_ ;
	assign \g12715/_2_  = _w13518_ ;
	assign \g12717/_2_  = _w13522_ ;
	assign \g12718/_2__syn_2  = _w13527_ ;
	assign \g1272/_0_  = _w13535_ ;
	assign \g12728/_1__syn_2  = _w13537_ ;
	assign \g12730/_3_  = _w13542_ ;
	assign \g12741/_1__syn_2  = _w13547_ ;
	assign \g12746/_0__syn_2  = _w11807_ ;
	assign \g12748/_0_  = _w13552_ ;
	assign \g12749/_0_  = _w13553_ ;
	assign \g12759/_1__syn_2  = _w11611_ ;
	assign \g12760/_0_  = _w13555_ ;
	assign \g12762/_0_  = _w13558_ ;
	assign \g12763/_0_  = _w13561_ ;
	assign \g12764/_0_  = _w13564_ ;
	assign \g12765/_0_  = _w13567_ ;
	assign \g12766/_0_  = _w13570_ ;
	assign \g12767/_0_  = _w13573_ ;
	assign \g12768/_0_  = _w13576_ ;
	assign \g12769/_0_  = _w13579_ ;
	assign \g12770/_0_  = _w13582_ ;
	assign \g12771/_0_  = _w13585_ ;
	assign \g12772/_0_  = _w13588_ ;
	assign \g12773/_0_  = _w13591_ ;
	assign \g12774/_0_  = _w13594_ ;
	assign \g12775/_0_  = _w13597_ ;
	assign \g12776/_0_  = _w13600_ ;
	assign \g12777/_0_  = _w13603_ ;
	assign \g12778/_0_  = _w13606_ ;
	assign \g12779/_0_  = _w13609_ ;
	assign \g1278/_0_  = _w13633_ ;
	assign \g12780/_0_  = _w13636_ ;
	assign \g12781/_0_  = _w13639_ ;
	assign \g12782/_0_  = _w13642_ ;
	assign \g12783/_0_  = _w13645_ ;
	assign \g12784/_0_  = _w13648_ ;
	assign \g12785/_0_  = _w13651_ ;
	assign \g12786/_0_  = _w13654_ ;
	assign \g12787/_0_  = _w13657_ ;
	assign \g12788/_0_  = _w13660_ ;
	assign \g12789/_0_  = _w13663_ ;
	assign \g12790/_0_  = _w13666_ ;
	assign \g12791/_0_  = _w13669_ ;
	assign \g12792/_0_  = _w13672_ ;
	assign \g12793/_0_  = _w13675_ ;
	assign \g12794/_0_  = _w13678_ ;
	assign \g12795/_0_  = _w13681_ ;
	assign \g12796/_0_  = _w13684_ ;
	assign \g12797/_0_  = _w13687_ ;
	assign \g12798/_0_  = _w13688_ ;
	assign \g12799/_0_  = _w13689_ ;
	assign \g12800/_0_  = _w13690_ ;
	assign \g12801/_0_  = _w13691_ ;
	assign \g12802/_0_  = _w13692_ ;
	assign \g12803/_0_  = _w13693_ ;
	assign \g12804/_0_  = _w13694_ ;
	assign \g12805/_0_  = _w13695_ ;
	assign \g12806/_0_  = _w13696_ ;
	assign \g12807/_0_  = _w13697_ ;
	assign \g12808/_0_  = _w13698_ ;
	assign \g12809/_0_  = _w13699_ ;
	assign \g1281/_0_  = _w13702_ ;
	assign \g12810/_0_  = _w13703_ ;
	assign \g12811/_0_  = _w13704_ ;
	assign \g12812/_0_  = _w13705_ ;
	assign \g12813/_0_  = _w13706_ ;
	assign \g12814/_0_  = _w13707_ ;
	assign \g12815/_0_  = _w13710_ ;
	assign \g12816/_0_  = _w13713_ ;
	assign \g12817/_0_  = _w13716_ ;
	assign \g12818/_0_  = _w13719_ ;
	assign \g12819/_0_  = _w13722_ ;
	assign \g1282/_0_  = _w13723_ ;
	assign \g12820/_0_  = _w13726_ ;
	assign \g12821/_0_  = _w13729_ ;
	assign \g12822/_0_  = _w13732_ ;
	assign \g12823/_0_  = _w13735_ ;
	assign \g12824/_0_  = _w13738_ ;
	assign \g12825/_0_  = _w13741_ ;
	assign \g12826/_0_  = _w13744_ ;
	assign \g12827/_0_  = _w13747_ ;
	assign \g12828/_0_  = _w13750_ ;
	assign \g12829/_0_  = _w13753_ ;
	assign \g12830/_0_  = _w13756_ ;
	assign \g12831/_0_  = _w13758_ ;
	assign \g12832/_0_  = _w13762_ ;
	assign \g12833/_0_  = _w13763_ ;
	assign \g12835/_0_  = _w13766_ ;
	assign \g12836/_0_  = _w13767_ ;
	assign \g12838/_0_  = _w13770_ ;
	assign \g12848/_0_  = _w13772_ ;
	assign \g12849/_0_  = _w13774_ ;
	assign \g1285/_0_  = _w13775_ ;
	assign \g12850/_0_  = _w13776_ ;
	assign \g12857/_0_  = _w13778_ ;
	assign \g12858/_0_  = _w13779_ ;
	assign \g12859/_0_  = _w13780_ ;
	assign \g12861/_0_  = _w13781_ ;
	assign \g12862/_0_  = _w13782_ ;
	assign \g12868/_0_  = _w13785_ ;
	assign \g12869/_0_  = _w13786_ ;
	assign \g1287/_0_  = _w13807_ ;
	assign \g12870/_0_  = _w13808_ ;
	assign \g12871/_0_  = _w13809_ ;
	assign \g12872/_0_  = _w13810_ ;
	assign \g12873/_0_  = _w13811_ ;
	assign \g12874/_0_  = _w13813_ ;
	assign \g12875/_0_  = _w13814_ ;
	assign \g12876/_0_  = _w13815_ ;
	assign \g12877/_0_  = _w13816_ ;
	assign \g12878/_0_  = _w13824_ ;
	assign \g12879/_0_  = _w13829_ ;
	assign \g12880/_0_  = _w13834_ ;
	assign \g12881/_0_  = _w13839_ ;
	assign \g12882/_0_  = _w13844_ ;
	assign \g12883/_0_  = _w13849_ ;
	assign \g12884/_0_  = _w13854_ ;
	assign \g12885/_0_  = _w13859_ ;
	assign \g12886/_0_  = _w13864_ ;
	assign \g12887/_0_  = _w13869_ ;
	assign \g12888/_0_  = _w13872_ ;
	assign \g12889/_0_  = _w13875_ ;
	assign \g1289/_0_  = _w13876_ ;
	assign \g12890/_0_  = _w13881_ ;
	assign \g12891/_0_  = _w13886_ ;
	assign \g12894/_0_  = _w13887_ ;
	assign \g12898/_0_  = _w13889_ ;
	assign \g12899/_0_  = _w13890_ ;
	assign \g12900/_0_  = _w13891_ ;
	assign \g12901/_0_  = _w13892_ ;
	assign \g12902/_0_  = _w13893_ ;
	assign \g12903/_0_  = _w13894_ ;
	assign \g12906/_0_  = _w13895_ ;
	assign \g12907/_0_  = _w13896_ ;
	assign \g12908/_0_  = _w13901_ ;
	assign \g12912/_0_  = _w13905_ ;
	assign \g12913/_0_  = _w13908_ ;
	assign \g12914/_0_  = _w13909_ ;
	assign \g12915/_0_  = _w13910_ ;
	assign \g12916/_0_  = _w13911_ ;
	assign \g12917/_0_  = _w13912_ ;
	assign \g12918/_0_  = _w13913_ ;
	assign \g12919/_0_  = _w13914_ ;
	assign \g12920/_0_  = _w13915_ ;
	assign \g12921/_0_  = _w13918_ ;
	assign \g12922/_0_  = _w13921_ ;
	assign \g12923/_0_  = _w13922_ ;
	assign \g12924/_0_  = _w13923_ ;
	assign \g12925/_0_  = _w13926_ ;
	assign \g12926/_0_  = _w13929_ ;
	assign \g12932/_0_  = _w13930_ ;
	assign \g12933/_0_  = _w13933_ ;
	assign \g12936/_0_  = _w13936_ ;
	assign \g12955/_0_  = _w13937_ ;
	assign \g13015/_0_  = _w13940_ ;
	assign \g13016/_0_  = _w13943_ ;
	assign \g13017/_0_  = _w13946_ ;
	assign \g13018/_0_  = _w13947_ ;
	assign \g13019/_0_  = _w13948_ ;
	assign \g13020/_0_  = _w13951_ ;
	assign \g13021/_0_  = _w13954_ ;
	assign \g13024/_0_  = _w13957_ ;
	assign \g13025/_0_  = _w13960_ ;
	assign \g13027/_0_  = _w13963_ ;
	assign \g13028/_0_  = _w13966_ ;
	assign \g13030/_0_  = _w13969_ ;
	assign \g13031/_0_  = _w13970_ ;
	assign \g13033/_0_  = _w13973_ ;
	assign \g13047/_0_  = _w13974_ ;
	assign \g13060/_0_  = _w13977_ ;
	assign \g13062/_0_  = _w13980_ ;
	assign \g13063/_0_  = _w13983_ ;
	assign \g13064/_0_  = _w13986_ ;
	assign \g13067/_0_  = _w13989_ ;
	assign \g13068/_0_  = _w13992_ ;
	assign \g13069/_0_  = _w13993_ ;
	assign \g13070/_0_  = _w13994_ ;
	assign \g13072/_0_  = _w13997_ ;
	assign \g13094/_0_  = _w13999_ ;
	assign \g13104/_0_  = _w14003_ ;
	assign \g13110/_0_  = _w14006_ ;
	assign \g13114/_0_  = _w14010_ ;
	assign \g13115/_0_  = _w14013_ ;
	assign \g13116/_0_  = _w14016_ ;
	assign \g13117/_0_  = _w14019_ ;
	assign \g13118/_0_  = _w14022_ ;
	assign \g13119/_0_  = _w14025_ ;
	assign \g13120/_0_  = _w14028_ ;
	assign \g13121/_0_  = _w14031_ ;
	assign \g13124/_0_  = _w14034_ ;
	assign \g13125/_0_  = _w14037_ ;
	assign \g13127/_0_  = _w14040_ ;
	assign \g13128/_0_  = _w14043_ ;
	assign \g13129/_0_  = _w14046_ ;
	assign \g13130/_0_  = _w14049_ ;
	assign \g13131/_0_  = _w14052_ ;
	assign \g13132/_0_  = _w14053_ ;
	assign \g13133/_0_  = _w14054_ ;
	assign \g13134/_0_  = _w14057_ ;
	assign \g13138/_0_  = _w14060_ ;
	assign \g13139/_0_  = _w14063_ ;
	assign \g13140/_0_  = _w14066_ ;
	assign \g13141/_0_  = _w14069_ ;
	assign \g13142/_0_  = _w14072_ ;
	assign \g13143/_0_  = _w14075_ ;
	assign \g13144/_0_  = _w14078_ ;
	assign \g13146/_0_  = _w14081_ ;
	assign \g13150/_0_  = _w14084_ ;
	assign \g13152/_0_  = _w14087_ ;
	assign \g13154/_0_  = _w14090_ ;
	assign \g13155/_0_  = _w14093_ ;
	assign \g13156/_0_  = _w14096_ ;
	assign \g13157/_0_  = _w14099_ ;
	assign \g13158/_0_  = _w14100_ ;
	assign \g1320/_3_  = _w14118_ ;
	assign \g13266/_0_  = _w14121_ ;
	assign \g13269/_0_  = _w14124_ ;
	assign \g13274/_0_  = _w14127_ ;
	assign \g13277/_0_  = _w14130_ ;
	assign \g13280/_0_  = _w14133_ ;
	assign \g13283/_0_  = _w14134_ ;
	assign \g13294/_0_  = _w14137_ ;
	assign \g13330/_0_  = _w14139_ ;
	assign \g13333/_0_  = _w14142_ ;
	assign \g13334/_0_  = _w14143_ ;
	assign \g13335/_0_  = _w14144_ ;
	assign \g13336/_0_  = _w14145_ ;
	assign \g13337/_0_  = _w14146_ ;
	assign \g13338/_0_  = _w14147_ ;
	assign \g13345/_0_  = _w14149_ ;
	assign \g13346/_0_  = _w14150_ ;
	assign \g13347/_0_  = _w14152_ ;
	assign \g13348/_0_  = _w14153_ ;
	assign \g13349/_0_  = _w14154_ ;
	assign \g13350/_0_  = _w14155_ ;
	assign \g13351/_0_  = _w14156_ ;
	assign \g13352/_0_  = _w14157_ ;
	assign \g13486/_0_  = _w14158_ ;
	assign \g13488/_0_  = _w14159_ ;
	assign \g13508/_0_  = _w14160_ ;
	assign \g13509/_0_  = _w14161_ ;
	assign \g13510/_0_  = _w14162_ ;
	assign \g13511/_0_  = _w14163_ ;
	assign \g13512/_0_  = _w14164_ ;
	assign \g13513/_0_  = _w14165_ ;
	assign \g13514/_0_  = _w14166_ ;
	assign \g13515/_0_  = _w14167_ ;
	assign \g13516/_0_  = _w14168_ ;
	assign \g13517/_0_  = _w14169_ ;
	assign \g13518/_0_  = _w14170_ ;
	assign \g13519/_0_  = _w14171_ ;
	assign \g13520/_0_  = _w14172_ ;
	assign \g13521/_0_  = _w14173_ ;
	assign \g13540/_0_  = _w14176_ ;
	assign \g13541/_0_  = _w14179_ ;
	assign \g13542/_0_  = _w14182_ ;
	assign \g13543/_0_  = _w14185_ ;
	assign \g13544/_0_  = _w14188_ ;
	assign \g13545/_0_  = _w14191_ ;
	assign \g13546/_0_  = _w14194_ ;
	assign \g13547/_0_  = _w14195_ ;
	assign \g13548/_0_  = _w14196_ ;
	assign \g13549/_0_  = _w14199_ ;
	assign \g13550/_0_  = _w14200_ ;
	assign \g13551/_0_  = _w14203_ ;
	assign \g13552/_0_  = _w14204_ ;
	assign \g13553/_0_  = _w14205_ ;
	assign \g13554/_0_  = _w14208_ ;
	assign \g13555/_0_  = _w14211_ ;
	assign \g13556/_0_  = _w14214_ ;
	assign \g13557/_0_  = _w14217_ ;
	assign \g13558/_0_  = _w14220_ ;
	assign \g13559/_0_  = _w14223_ ;
	assign \g13560/_0_  = _w14226_ ;
	assign \g13561/_0_  = _w14227_ ;
	assign \g13562/_0_  = _w14228_ ;
	assign \g13563/_0_  = _w14231_ ;
	assign \g13564/_0_  = _w14234_ ;
	assign \g13565/_0_  = _w14237_ ;
	assign \g13566/_0_  = _w14240_ ;
	assign \g13567/_0_  = _w14243_ ;
	assign \g13568/_0_  = _w14246_ ;
	assign \g13569/_0_  = _w14249_ ;
	assign \g13570/_0_  = _w14252_ ;
	assign \g13571/_0_  = _w14253_ ;
	assign \g13572/_0_  = _w14256_ ;
	assign \g137/_3_  = _w14271_ ;
	assign \g1387/_3_  = _w14277_ ;
	assign \g1388/_3_  = _w14282_ ;
	assign \g1389/_0_  = _w14286_ ;
	assign \g139/_0_  = _w14368_ ;
	assign \g1390/_0_  = _w14388_ ;
	assign \g1393/_0_  = _w14389_ ;
	assign \g140/_0_  = _w14393_ ;
	assign \g141/_0_  = _w14394_ ;
	assign \g14173/_0_  = _w14396_ ;
	assign \g14176/_0_  = _w14398_ ;
	assign \g142/_3_  = _w14412_ ;
	assign \g14273/_1__syn_2  = _w12826_ ;
	assign \g14274/_0_  = _w14413_ ;
	assign \g14280/_0_  = _w14419_ ;
	assign \g14281/_0_  = _w14425_ ;
	assign \g143/_3_  = _w14436_ ;
	assign \g14354/_3__syn_2  = _w9440_ ;
	assign \g14370/_0_  = _w14438_ ;
	assign \g14385/_0_  = _w14441_ ;
	assign \g14386/_0_  = _w14443_ ;
	assign \g144/_3_  = _w14448_ ;
	assign \g14407/_0_  = _w14456_ ;
	assign \g14412/_0_  = _w14458_ ;
	assign \g14435/_0_  = _w14463_ ;
	assign \g14439/_0_  = _w14465_ ;
	assign \g145/_0_  = _w14495_ ;
	assign \g14522/_0_  = _w14497_ ;
	assign \g14528/_0_  = _w14498_ ;
	assign \g14533/_0_  = _w14507_ ;
	assign \g14581/_1_  = _w14508_ ;
	assign \g14582/_0_  = _w14509_ ;
	assign \g146/_3_  = _w14513_ ;
	assign \g14671/_0_  = _w14519_ ;
	assign \g14672/_0_  = _w14525_ ;
	assign \g147/_0_  = _w14545_ ;
	assign \g1473/_0_  = _w14554_ ;
	assign \g148/_0_  = _w14563_ ;
	assign \g14826/_0_  = _w12040_ ;
	assign \g149/_0_  = _w14568_ ;
	assign \g14908/_0_  = _w14572_ ;
	assign \g14911/_0_  = _w14575_ ;
	assign \g14936/_2_  = _w14577_ ;
	assign \g1494/_0_  = _w14586_ ;
	assign \g1495/_0_  = _w14589_ ;
	assign \g14950/_2_  = _w14595_ ;
	assign \g14953/_2_  = _w14601_ ;
	assign \g15003/_0_  = _w14605_ ;
	assign \g15004/_0_  = _w14608_ ;
	assign \g15006/_0_  = _w14611_ ;
	assign \g15007/_0_  = _w14614_ ;
	assign \g15008/_0_  = _w14617_ ;
	assign \g15009/_0_  = _w14620_ ;
	assign \g15010/_0_  = _w14623_ ;
	assign \g15011/_0_  = _w14626_ ;
	assign \g15012/_0_  = _w14629_ ;
	assign \g15013/_0_  = _w14632_ ;
	assign \g15014/_0_  = _w14635_ ;
	assign \g15015/_0_  = _w14638_ ;
	assign \g15016/_0_  = _w14641_ ;
	assign \g15017/_0_  = _w14644_ ;
	assign \g15018/_0_  = _w14647_ ;
	assign \g15019/_0_  = _w14648_ ;
	assign \g15035/_0_  = _w14650_ ;
	assign \g15036/_0_  = _w14653_ ;
	assign \g15038/_0_  = _w14658_ ;
	assign \g15039/_0_  = _w14662_ ;
	assign \g15040/_0_  = _w14666_ ;
	assign \g15041/_0_  = _w14670_ ;
	assign \g15042/_0_  = _w14674_ ;
	assign \g15043/_0_  = _w14678_ ;
	assign \g15044/_0_  = _w14682_ ;
	assign \g15045/_0_  = _w14686_ ;
	assign \g15046/_0_  = _w14690_ ;
	assign \g15056/_00_  = _w14693_ ;
	assign \g151/_0_  = _w14694_ ;
	assign \g15193/_0_  = _w14696_ ;
	assign \g152/_0_  = _w14697_ ;
	assign \g15256/_0_  = _w14701_ ;
	assign \g153/_0_  = _w14704_ ;
	assign \g15393/_0_  = _w14708_ ;
	assign \g15394/_0_  = _w14710_ ;
	assign \g15395/_0_  = _w14713_ ;
	assign \g15396/_0_  = _w14716_ ;
	assign \g15397/_0_  = _w14719_ ;
	assign \g15398/_0_  = _w14722_ ;
	assign \g15399/_0_  = _w14725_ ;
	assign \g154/_0_  = _w14728_ ;
	assign \g15400/_0_  = _w14731_ ;
	assign \g15401/_0_  = _w14734_ ;
	assign \g15402/_0_  = _w14736_ ;
	assign \g15403/_0_  = _w14738_ ;
	assign \g15404/_0_  = _w14741_ ;
	assign \g15405/_0_  = _w14744_ ;
	assign \g15406/_0_  = _w14746_ ;
	assign \g15407/_0_  = _w14748_ ;
	assign \g15408/_0_  = _w14751_ ;
	assign \g15473/_0_  = _w14754_ ;
	assign \g15650/_0_  = _w14755_ ;
	assign \g15651/_0_  = _w14756_ ;
	assign \g15652/_0_  = _w14757_ ;
	assign \g15653/_0_  = _w14758_ ;
	assign \g15662/_0_  = _w14759_ ;
	assign \g15663/_0_  = _w14760_ ;
	assign \g15664/_0_  = _w14761_ ;
	assign \g15665/_0_  = _w14762_ ;
	assign \g15666/_0_  = _w14763_ ;
	assign \g15667/_0_  = _w14764_ ;
	assign \g15668/_0_  = _w14765_ ;
	assign \g15669/_0_  = _w14766_ ;
	assign \g15670/_0_  = _w14767_ ;
	assign \g15671/_0_  = _w14768_ ;
	assign \g15672/_0_  = _w14769_ ;
	assign \g15673/_0_  = _w14770_ ;
	assign \g15674/_0_  = _w14771_ ;
	assign \g15675/_0_  = _w14772_ ;
	assign \g1569/_0_  = _w14808_ ;
	assign \g1570/_0_  = _w14812_ ;
	assign \g1575/_0_  = _w14815_ ;
	assign \g1576/_0_  = _w14816_ ;
	assign \g15922/_1_  = _w14817_ ;
	assign \g15970/_0_  = _w14818_ ;
	assign \g16059/_0_  = _w14820_ ;
	assign \g1606/_3_  = _w14826_ ;
	assign \g16124/_0_  = _w12898_ ;
	assign \g16144/_0_  = _w14828_ ;
	assign \g16202/_0_  = _w14831_ ;
	assign \g16214/_0_  = _w14833_ ;
	assign \g16247/_0_  = _w14837_ ;
	assign \g16257/_0_  = _w14841_ ;
	assign \g16274/_1_  = _w14842_ ;
	assign \g16324/_0_  = _w13042_ ;
	assign \g16343/_1__syn_2  = _w14002_ ;
	assign \g16381/_0_  = _w14844_ ;
	assign \g16383/_0_  = _w14851_ ;
	assign \g16386/_0_  = _w14853_ ;
	assign \g16414/_1__syn_2  = _w13777_ ;
	assign \g16416/_0__syn_2  = _w13091_ ;
	assign \g16448/_0_  = _w14854_ ;
	assign \g16460/_1_  = _w14855_ ;
	assign \g16625/_3_  = _w14461_ ;
	assign \g16662/_0_  = _w14862_ ;
	assign \g16668/_1__syn_2  = _w14148_ ;
	assign \g16692/_0_  = _w14863_ ;
	assign \g16721/_0_  = _w14867_ ;
	assign \g16723/_0_  = _w14870_ ;
	assign \g16725/_0_  = _w14872_ ;
	assign \g16726/_0_  = _w14873_ ;
	assign \g16727/_0_  = _w14876_ ;
	assign \g16728/_0_  = _w14879_ ;
	assign \g16729/_0_  = _w14880_ ;
	assign \g16730/_0_  = _w14882_ ;
	assign \g16731/_0_  = _w14885_ ;
	assign \g16732/_0_  = _w14888_ ;
	assign \g16733/_0_  = _w14889_ ;
	assign \g16734/_0_  = _w14890_ ;
	assign \g16735/_0_  = _w14892_ ;
	assign \g16736/_0_  = _w14893_ ;
	assign \g16737/_0_  = _w14896_ ;
	assign \g16738/_0_  = _w14897_ ;
	assign \g16739/_0_  = _w14898_ ;
	assign \g16740/_0_  = _w14900_ ;
	assign \g16741/_0_  = _w14901_ ;
	assign \g16742/_0_  = _w14904_ ;
	assign \g16743/_0_  = _w14905_ ;
	assign \g16747/_0_  = _w14907_ ;
	assign \g16748/_0_  = _w14908_ ;
	assign \g16749/_0_  = _w14909_ ;
	assign \g16750/_0_  = _w14910_ ;
	assign \g16753/_0_  = _w14911_ ;
	assign \g16754/_0_  = _w14912_ ;
	assign \g16755/_0_  = _w14913_ ;
	assign \g16756/_0_  = _w14914_ ;
	assign \g16757/_0_  = _w14915_ ;
	assign \g16758/_0_  = _w14916_ ;
	assign \g16761/_0_  = _w14919_ ;
	assign \g16765/_0_  = _w14922_ ;
	assign \g16766/_0_  = _w14923_ ;
	assign \g16767/_0_  = _w14924_ ;
	assign \g16768/_0_  = _w14925_ ;
	assign \g16769/_0_  = _w14926_ ;
	assign \g16772/_0_  = _w14927_ ;
	assign \g16785/_0_  = _w14930_ ;
	assign \g16786/_0_  = _w14932_ ;
	assign \g16787/_0_  = _w14933_ ;
	assign \g16788/_0_  = _w14936_ ;
	assign \g16789/_0_  = _w14939_ ;
	assign \g16790/_0_  = _w14940_ ;
	assign \g16791/_0_  = _w14941_ ;
	assign \g16804/_0_  = _w14943_ ;
	assign \g16805/_0_  = _w14944_ ;
	assign \g16806/_0_  = _w14947_ ;
	assign \g16807/_0_  = _w14952_ ;
	assign \g16808/_0_  = _w14953_ ;
	assign \g16809/_0_  = _w14954_ ;
	assign \g16810/_0_  = _w14956_ ;
	assign \g16811/_0_  = _w14957_ ;
	assign \g16812/_0_  = _w14960_ ;
	assign \g16813/_0_  = _w14963_ ;
	assign \g16814/_0_  = _w14964_ ;
	assign \g16815/_0_  = _w14965_ ;
	assign \g16816/_0_  = _w14966_ ;
	assign \g16817/_0_  = _w14969_ ;
	assign \g16819/_0_  = _w14975_ ;
	assign \g16822/_0_  = _w14977_ ;
	assign \g16823/_0_  = _w14979_ ;
	assign \g16824/_0_  = _w14981_ ;
	assign \g16825/_0_  = _w14983_ ;
	assign \g16828/_0_  = _w14984_ ;
	assign \g16829/_0_  = _w14985_ ;
	assign \g16830/_0_  = _w14986_ ;
	assign \g16831/_0_  = _w14987_ ;
	assign \g16832/_0_  = _w14988_ ;
	assign \g16833/_0_  = _w14989_ ;
	assign \g16834/_0_  = _w14990_ ;
	assign \g16835/_0_  = _w14991_ ;
	assign \g16836/_0_  = _w14992_ ;
	assign \g16837/_0_  = _w14998_ ;
	assign \g16840/_0_  = _w15000_ ;
	assign \g16841/_0_  = _w15002_ ;
	assign \g16842/_0_  = _w15004_ ;
	assign \g16843/_0_  = _w15006_ ;
	assign \g16846/_0_  = _w15012_ ;
	assign \g16847/_0_  = _w15013_ ;
	assign \g16848/_0_  = _w15014_ ;
	assign \g16849/_0_  = _w15016_ ;
	assign \g16850/_0_  = _w15018_ ;
	assign \g16851/_0_  = _w15020_ ;
	assign \g16852/_0_  = _w15022_ ;
	assign \g16853/_0_  = _w15023_ ;
	assign \g16854/_0_  = _w15024_ ;
	assign \g16855/_0_  = _w15025_ ;
	assign \g16856/_0_  = _w15028_ ;
	assign \g16857/_0_  = _w15031_ ;
	assign \g16859/_0_  = _w15034_ ;
	assign \g16862/_0_  = _w15037_ ;
	assign \g16865/_0_  = _w15040_ ;
	assign \g16866/_0_  = _w15043_ ;
	assign \g16867/_0_  = _w15046_ ;
	assign \g16868/_0_  = _w15049_ ;
	assign \g16869/_0_  = _w15050_ ;
	assign \g16870/_0_  = _w15054_ ;
	assign \g16871/_0_  = _w15056_ ;
	assign \g16872/_0_  = _w15060_ ;
	assign \g16873/_0_  = _w15064_ ;
	assign \g16874/_0_  = _w15066_ ;
	assign \g16875/_0_  = _w15070_ ;
	assign \g16876/_0_  = _w15074_ ;
	assign \g16877/_0_  = _w15077_ ;
	assign \g16878/_0_  = _w15078_ ;
	assign \g16879/_0_  = _w15079_ ;
	assign \g16880/_0_  = _w15080_ ;
	assign \g16881/_0_  = _w15081_ ;
	assign \g16882/_0_  = _w15086_ ;
	assign \g16884/_0_  = _w15088_ ;
	assign \g16887/_0_  = _w15091_ ;
	assign \g16891/_0_  = _w15093_ ;
	assign \g16892/_0_  = _w15094_ ;
	assign \g16893/_0_  = _w15095_ ;
	assign \g16894/_0_  = _w15096_ ;
	assign \g16895/_0_  = _w15097_ ;
	assign \g16897/_0_  = _w15098_ ;
	assign \g16898/_0_  = _w15101_ ;
	assign \g16899/_0_  = _w15104_ ;
	assign \g16900/_0_  = _w15105_ ;
	assign \g16901/_0_  = _w15107_ ;
	assign \g16902/_0_  = _w15108_ ;
	assign \g16903/_0_  = _w15109_ ;
	assign \g16904/_0_  = _w15112_ ;
	assign \g16905/_0_  = _w15114_ ;
	assign \g16906/_0_  = _w15115_ ;
	assign \g16907/_0_  = _w15116_ ;
	assign \g16908/_0_  = _w15117_ ;
	assign \g16909/_0_  = _w15118_ ;
	assign \g16910/_0_  = _w15120_ ;
	assign \g16912/_0_  = _w15121_ ;
	assign \g16914/_0_  = _w15124_ ;
	assign \g16915/_0_  = _w15125_ ;
	assign \g16950/_0_  = _w15127_ ;
	assign \g16951/_0_  = _w15129_ ;
	assign \g16952/_0_  = _w15131_ ;
	assign \g16953/_0_  = _w15133_ ;
	assign \g16954/_0_  = _w15135_ ;
	assign \g16955/_0_  = _w15136_ ;
	assign \g16956/_0_  = _w15137_ ;
	assign \g16957/_0_  = _w15138_ ;
	assign \g16958/_0_  = _w15139_ ;
	assign \g16959/_0_  = _w15140_ ;
	assign \g16960/_0_  = _w15142_ ;
	assign \g16961/_0_  = _w15144_ ;
	assign \g16962/_0_  = _w15146_ ;
	assign \g16963/_0_  = _w15148_ ;
	assign \g16964/_0_  = _w15150_ ;
	assign \g16965/_0_  = _w15152_ ;
	assign \g16966/_0_  = _w15154_ ;
	assign \g16967/_0_  = _w15156_ ;
	assign \g16968/_0_  = _w15158_ ;
	assign \g16970/_0_  = _w15160_ ;
	assign \g17102/_3_  = _w15163_ ;
	assign \g17106/_0_  = _w15167_ ;
	assign \g17107/_0_  = _w15168_ ;
	assign \g17109/_0_  = _w15169_ ;
	assign \g17110/_0_  = _w15170_ ;
	assign \g17111/_0_  = _w15171_ ;
	assign \g17112/_0_  = _w15172_ ;
	assign \g17115/_0_  = _w15173_ ;
	assign \g17116/_0_  = _w15174_ ;
	assign \g17119/_0_  = _w15175_ ;
	assign \g17120/_0_  = _w15176_ ;
	assign \g17122/_0_  = _w15177_ ;
	assign \g17123/_0_  = _w15178_ ;
	assign \g17124/_0_  = _w15179_ ;
	assign \g17125/_0_  = _w15180_ ;
	assign \g17126/_0_  = _w15181_ ;
	assign \g17127/_0_  = _w15182_ ;
	assign \g17128/_0_  = _w15183_ ;
	assign \g17130/_0_  = _w15184_ ;
	assign \g17131/_0_  = _w15185_ ;
	assign \g17132/_0_  = _w15186_ ;
	assign \g17133/_0_  = _w15187_ ;
	assign \g17134/_0_  = _w15188_ ;
	assign \g17135/_0_  = _w15189_ ;
	assign \g17136/_0_  = _w15190_ ;
	assign \g17137/_0_  = _w15191_ ;
	assign \g17138/_0_  = _w15192_ ;
	assign \g17140/_0_  = _w15193_ ;
	assign \g17141/_0_  = _w15194_ ;
	assign \g17142/_0_  = _w15195_ ;
	assign \g17143/_0_  = _w15196_ ;
	assign \g17144/_0_  = _w15197_ ;
	assign \g17145/_0_  = _w15198_ ;
	assign \g17146/_0_  = _w15199_ ;
	assign \g17147/_0_  = _w15200_ ;
	assign \g17148/_0_  = _w15201_ ;
	assign \g17149/_0_  = _w15202_ ;
	assign \g17150/_0_  = _w15203_ ;
	assign \g17151/_0_  = _w15204_ ;
	assign \g17152/_0_  = _w15205_ ;
	assign \g17153/_0_  = _w15206_ ;
	assign \g17154/_0_  = _w15207_ ;
	assign \g17155/_0_  = _w15208_ ;
	assign \g17157/_0_  = _w15209_ ;
	assign \g17159/_0_  = _w15213_ ;
	assign \g17160/_0_  = _w15215_ ;
	assign \g17161/_0_  = _w15216_ ;
	assign \g17162/_0_  = _w15217_ ;
	assign \g17163/_0_  = _w15220_ ;
	assign \g17164/_0_  = _w15221_ ;
	assign \g17165/_0_  = _w15223_ ;
	assign \g17166/_0_  = _w15224_ ;
	assign \g17168/_0_  = _w15225_ ;
	assign \g17171/_0_  = _w15226_ ;
	assign \g17173/_0_  = _w15230_ ;
	assign \g17177/_0_  = _w15231_ ;
	assign \g17178/_0_  = _w15232_ ;
	assign \g17179/_0_  = _w15233_ ;
	assign \g17180/_0_  = _w15234_ ;
	assign \g17182/_0_  = _w15235_ ;
	assign \g17183/_0_  = _w15236_ ;
	assign \g17184/_0_  = _w15237_ ;
	assign \g17185/_0_  = _w15238_ ;
	assign \g17186/_0_  = _w15239_ ;
	assign \g17188/_0_  = _w15240_ ;
	assign \g17189/_0_  = _w15241_ ;
	assign \g17190/_0_  = _w15242_ ;
	assign \g17191/_0_  = _w15243_ ;
	assign \g17193/_0_  = _w15244_ ;
	assign \g17194/_0_  = _w15245_ ;
	assign \g17195/_0_  = _w15246_ ;
	assign \g17196/_0_  = _w15247_ ;
	assign \g17197/_0_  = _w15248_ ;
	assign \g17198/_0_  = _w15249_ ;
	assign \g17199/_0_  = _w15250_ ;
	assign \g17200/_0_  = _w15251_ ;
	assign \g17201/_0_  = _w15252_ ;
	assign \g17202/_0_  = _w15253_ ;
	assign \g17203/_0_  = _w15256_ ;
	assign \g17204/_0_  = _w15257_ ;
	assign \g17205/_0_  = _w15258_ ;
	assign \g17206/_0_  = _w15259_ ;
	assign \g17207/_0_  = _w15260_ ;
	assign \g17208/_0_  = _w15261_ ;
	assign \g17209/_0_  = _w15262_ ;
	assign \g17210/_0_  = _w15263_ ;
	assign \g17211/_0_  = _w15264_ ;
	assign \g17212/_0_  = _w15267_ ;
	assign \g17213/_0_  = _w15270_ ;
	assign \g17214/_0_  = _w15273_ ;
	assign \g17215/_0_  = _w15276_ ;
	assign \g17216/_0_  = _w15279_ ;
	assign \g17217/_0_  = _w15282_ ;
	assign \g17218/_0_  = _w15285_ ;
	assign \g17219/_0_  = _w15288_ ;
	assign \g17223/_0_  = _w15291_ ;
	assign \g17224/_0_  = _w15294_ ;
	assign \g17225/_0_  = _w15297_ ;
	assign \g17226/_0_  = _w15298_ ;
	assign \g17227/_0_  = _w15299_ ;
	assign \g17228/_0_  = _w15302_ ;
	assign \g17229/_0_  = _w15303_ ;
	assign \g17231/_0_  = _w15304_ ;
	assign \g17232/_0_  = _w15305_ ;
	assign \g17233/_0_  = _w15306_ ;
	assign \g17234/_0_  = _w15307_ ;
	assign \g17237/_0_  = _w15308_ ;
	assign \g17239/_0_  = _w15309_ ;
	assign \g17240/_0_  = _w15310_ ;
	assign \g17243/_0_  = _w15311_ ;
	assign \g17246/_0_  = _w15312_ ;
	assign \g17247/_0_  = _w15313_ ;
	assign \g17248/_0_  = _w15314_ ;
	assign \g17249/_0_  = _w15315_ ;
	assign \g17250/_0_  = _w15316_ ;
	assign \g17251/_0_  = _w15317_ ;
	assign \g17252/_0_  = _w15318_ ;
	assign \g17253/_0_  = _w15319_ ;
	assign \g17254/_0_  = _w15320_ ;
	assign \g17258/_0_  = _w15321_ ;
	assign \g17261/_0_  = _w15329_ ;
	assign \g17262/_0_  = _w15330_ ;
	assign \g17269/_0_  = _w15331_ ;
	assign \g17271/_0_  = _w15332_ ;
	assign \g17274/_0_  = _w15335_ ;
	assign \g17275/_0_  = _w15336_ ;
	assign \g17276/_0_  = _w15339_ ;
	assign \g17277/_0_  = _w15342_ ;
	assign \g17278/_0_  = _w15345_ ;
	assign \g17279/_0_  = _w15348_ ;
	assign \g17280/_0_  = _w15351_ ;
	assign \g17281/_0_  = _w15354_ ;
	assign \g17282/_0_  = _w15355_ ;
	assign \g17283/_0_  = _w15356_ ;
	assign \g17285/_0_  = _w15359_ ;
	assign \g17290/_0_  = _w15360_ ;
	assign \g17292/_0_  = _w15361_ ;
	assign \g17293/_0_  = _w15362_ ;
	assign \g17296/_0_  = _w15363_ ;
	assign \g17297/_0_  = _w15364_ ;
	assign \g17298/_0_  = _w15366_ ;
	assign \g173/_0_  = _w15373_ ;
	assign \g17303/_0_  = _w15374_ ;
	assign \g17304/_0_  = _w15375_ ;
	assign \g17305/_0_  = _w15376_ ;
	assign \g17306/_0_  = _w15377_ ;
	assign \g17307/_0_  = _w15378_ ;
	assign \g17308/_0_  = _w15379_ ;
	assign \g17309/_0_  = _w15380_ ;
	assign \g17310/_0_  = _w15381_ ;
	assign \g17311/_0_  = _w15382_ ;
	assign \g17312/_0_  = _w15383_ ;
	assign \g17314/_0_  = _w15384_ ;
	assign \g17315/_0_  = _w15385_ ;
	assign \g17316/_0_  = _w15386_ ;
	assign \g17317/_0_  = _w15387_ ;
	assign \g17318/_0_  = _w15388_ ;
	assign \g17319/_0_  = _w15389_ ;
	assign \g17320/_0_  = _w15390_ ;
	assign \g17321/_0_  = _w15391_ ;
	assign \g17322/_0_  = _w15392_ ;
	assign \g17323/_0_  = _w15393_ ;
	assign \g17324/_0_  = _w15394_ ;
	assign \g17325/_0_  = _w15395_ ;
	assign \g17326/_0_  = _w15396_ ;
	assign \g17327/_0_  = _w15397_ ;
	assign \g17328/_0_  = _w15398_ ;
	assign \g17329/_0_  = _w15399_ ;
	assign \g17330/_0_  = _w15400_ ;
	assign \g17331/_0_  = _w15401_ ;
	assign \g17332/_0_  = _w15402_ ;
	assign \g17333/_0_  = _w15403_ ;
	assign \g17335/_0_  = _w15404_ ;
	assign \g17336/_0_  = _w15407_ ;
	assign \g17337/_0_  = _w15408_ ;
	assign \g17338/_0_  = _w15409_ ;
	assign \g17339/_0_  = _w15410_ ;
	assign \g17340/_0_  = _w15411_ ;
	assign \g17342/_0_  = _w15412_ ;
	assign \g17343/_0_  = _w15413_ ;
	assign \g17347/_0_  = _w15414_ ;
	assign \g17350/_0_  = _w15415_ ;
	assign \g17354/_0_  = _w15416_ ;
	assign \g17356/_0_  = _w15417_ ;
	assign \g17357/_0_  = _w15418_ ;
	assign \g17358/_0_  = _w15419_ ;
	assign \g17359/_0_  = _w15420_ ;
	assign \g17360/_0_  = _w15421_ ;
	assign \g17415/_0_  = _w15424_ ;
	assign \g17441/_0_  = _w15425_ ;
	assign \g17442/_0_  = _w15426_ ;
	assign \g17451/_0_  = _w15427_ ;
	assign \g17457/_0_  = _w15429_ ;
	assign \g17458/_0_  = _w15430_ ;
	assign \g17459/_0_  = _w15431_ ;
	assign \g17460/_0_  = _w15432_ ;
	assign \g17461/_0_  = _w15433_ ;
	assign \g17462/_0_  = _w15434_ ;
	assign \g17463/_0_  = _w15435_ ;
	assign \g17464/_0_  = _w15436_ ;
	assign \g17465/_0_  = _w15437_ ;
	assign \g17466/_0_  = _w15438_ ;
	assign \g17467/_0_  = _w15439_ ;
	assign \g17468/_0_  = _w15442_ ;
	assign \g17469/_0_  = _w15445_ ;
	assign \g17470/_0_  = _w15446_ ;
	assign \g17471/_0_  = _w15447_ ;
	assign \g17472/_0_  = _w15448_ ;
	assign \g175/_3_  = _w15457_ ;
	assign \g1750/_0_  = _w15465_ ;
	assign \g176/_3_  = _w15475_ ;
	assign \g17619/_0_  = _w15476_ ;
	assign \g17620/_0_  = _w15477_ ;
	assign \g1763/_3_  = _w15483_ ;
	assign \g1764/_3_  = _w15488_ ;
	assign \g1768/_0_  = _w15491_ ;
	assign \g1769/_0_  = _w15494_ ;
	assign \g177/_3_  = _w15503_ ;
	assign \g17737/_0_  = _w15507_ ;
	assign \g17747/_0_  = _w15509_ ;
	assign \g178/_3_  = _w15514_ ;
	assign \g17814/_1_  = _w13380_ ;
	assign \g17815/_0_  = _w15516_ ;
	assign \g17821/_1_  = _w15518_ ;
	assign \g17821/_1__syn_2  = _w15517_ ;
	assign \g17872/_0_  = _w15520_ ;
	assign \g179/_3_  = _w15526_ ;
	assign \g17902/_0_  = _w15528_ ;
	assign \g180/_3_  = _w15534_ ;
	assign \g18020/_1_  = _w15536_ ;
	assign \g18057/_0_  = _w15538_ ;
	assign \g18096/_0_  = _w15541_ ;
	assign \g18099/_0_  = _w15543_ ;
	assign \g18107/_0_  = _w15545_ ;
	assign \g18133/_0_  = _w15548_ ;
	assign \g18140/_1_  = _w14452_ ;
	assign \g18153/_0_  = _w15550_ ;
	assign \g182/_0_  = _w15555_ ;
	assign \g18218/_0_  = _w15558_ ;
	assign \g18244/_0_  = _w15560_ ;
	assign \g18262/_0_  = _w15563_ ;
	assign \g18267/_0_  = _w15566_ ;
	assign \g18387/_1__syn_2  = _w15569_ ;
	assign \g184/_0_  = _w15572_ ;
	assign \g18478/_1_  = _w14654_ ;
	assign \g18585/_3_  = _w14001_ ;
	assign \g18608/_0_  = _w15573_ ;
	assign \g18609/_0_  = _w15574_ ;
	assign \g18613/_0_  = _w15578_ ;
	assign \g18618/_0_  = _w15579_ ;
	assign \g18647/_0_  = _w15582_ ;
	assign \g18687/_2_  = _w13168_ ;
	assign \g18707/_0_  = _w15583_ ;
	assign \g18748/_0_  = _w15587_ ;
	assign \g18753/_0_  = _w15589_ ;
	assign \g18758/_0_  = _w15592_ ;
	assign \g18759/_0_  = _w15596_ ;
	assign \g18760/_0_  = _w15599_ ;
	assign \g18761/_0_  = _w15601_ ;
	assign \g18762/_0_  = _w15604_ ;
	assign \g18763/_0_  = _w15607_ ;
	assign \g18764/_0_  = _w15608_ ;
	assign \g18765/_0_  = _w15609_ ;
	assign \g18766/_0_  = _w15610_ ;
	assign \g18767/_0_  = _w15613_ ;
	assign \g18768/_0_  = _w15614_ ;
	assign \g18770/_0_  = _w15615_ ;
	assign \g18771/_0_  = _w15618_ ;
	assign \g18788/_0_  = _w15619_ ;
	assign \g18796/_0_  = _w15620_ ;
	assign \g18800/_0_  = _w15621_ ;
	assign \g18801/_0_  = _w15622_ ;
	assign \g18802/_0_  = _w15623_ ;
	assign \g18803/_0_  = _w15624_ ;
	assign \g18804/_0_  = _w15625_ ;
	assign \g18805/_0_  = _w15626_ ;
	assign \g18807/_0_  = _w15627_ ;
	assign \g18840/_0_  = _w15631_ ;
	assign \g18843/_0_  = _w15632_ ;
	assign \g18844/_0_  = _w15637_ ;
	assign \g18846/_0_  = _w15641_ ;
	assign \g18847/_0_  = _w15644_ ;
	assign \g18848/_0_  = _w15647_ ;
	assign \g18849/_0_  = _w15651_ ;
	assign \g18850/_0_  = _w15655_ ;
	assign \g18851/_0_  = _w15658_ ;
	assign \g18852/_0_  = _w15661_ ;
	assign \g18853/_0_  = _w15664_ ;
	assign \g18854/_0_  = _w15667_ ;
	assign \g18855/_0_  = _w15671_ ;
	assign \g18856/_0_  = _w13001_ ;
	assign \g18858/_0_  = _w12993_ ;
	assign \g18860/_0_  = _w15674_ ;
	assign \g18861/_0_  = _w15675_ ;
	assign \g18863/_0_  = _w15676_ ;
	assign \g18864/_0_  = _w15677_ ;
	assign \g18866/_0_  = _w15678_ ;
	assign \g18867/_0_  = _w15679_ ;
	assign \g18868/_0_  = _w15680_ ;
	assign \g18869/_0_  = _w15681_ ;
	assign \g18870/_0_  = _w15682_ ;
	assign \g18871/_0_  = _w15683_ ;
	assign \g18872/_0_  = _w15684_ ;
	assign \g18873/_0_  = _w15685_ ;
	assign \g18874/_0_  = _w15686_ ;
	assign \g18875/_0_  = _w15687_ ;
	assign \g18876/_0_  = _w15688_ ;
	assign \g18877/_0_  = _w15689_ ;
	assign \g18878/_0_  = _w15690_ ;
	assign \g18879/_0_  = _w15691_ ;
	assign \g18880/_0_  = _w15692_ ;
	assign \g18881/_0_  = _w15693_ ;
	assign \g18882/_0_  = _w15694_ ;
	assign \g18883/_0_  = _w15695_ ;
	assign \g18888/_0_  = _w15698_ ;
	assign \g18892/_0_  = _w15701_ ;
	assign \g18895/_0_  = _w15704_ ;
	assign \g18896/_0_  = _w15707_ ;
	assign \g18897/_0_  = _w15708_ ;
	assign \g18905/_0_  = _w15711_ ;
	assign \g18908/_0_  = _w15712_ ;
	assign \g18909/_0_  = _w15713_ ;
	assign \g18912/_0_  = _w15714_ ;
	assign \g18918/_0_  = _w15718_ ;
	assign \g18919/_0_  = _w15722_ ;
	assign \g18920/_0_  = _w15723_ ;
	assign \g18921/_0_  = _w15726_ ;
	assign \g18922/_0_  = _w15727_ ;
	assign \g18924/_0_  = _w15730_ ;
	assign \g18925/_0_  = _w15731_ ;
	assign \g18927/_0_  = _w15732_ ;
	assign \g18930/_0_  = _w15733_ ;
	assign \g18966/_0_  = _w15736_ ;
	assign \g18968/_0_  = _w15739_ ;
	assign \g18970/_0_  = _w15740_ ;
	assign \g18974/_0_  = _w15741_ ;
	assign \g18975/_0_  = _w15744_ ;
	assign \g18977/_0_  = _w15747_ ;
	assign \g18981/_0_  = _w13023_ ;
	assign \g18983/_0_  = _w12914_ ;
	assign \g18985/_0_  = _w12924_ ;
	assign \g18987/_0_  = _w12932_ ;
	assign \g18989/_0_  = _w12940_ ;
	assign \g18991/_0_  = _w15751_ ;
	assign \g18992/_0_  = _w15754_ ;
	assign \g18993/_0_  = _w15757_ ;
	assign \g18994/_0_  = _w15758_ ;
	assign \g18995/_0_  = _w15761_ ;
	assign \g18996/_0_  = _w15762_ ;
	assign \g18997/_0_  = _w15765_ ;
	assign \g18998/_0_  = _w15766_ ;
	assign \g18999/_0_  = _w15767_ ;
	assign \g19001/_0_  = _w15768_ ;
	assign \g19003/_0_  = _w15769_ ;
	assign \g19005/_0_  = _w15770_ ;
	assign \g19006/_0_  = _w15775_ ;
	assign \g19014/_0_  = _w12948_ ;
	assign \g19016/_0_  = _w12954_ ;
	assign \g19018/_0_  = _w12962_ ;
	assign \g19020/_0_  = _w12970_ ;
	assign \g19022/_0_  = _w13009_ ;
	assign \g19056/_3_  = _w15779_ ;
	assign \g19058/_3_  = _w15783_ ;
	assign \g19060/_3_  = _w15787_ ;
	assign \g19062/_3_  = _w15791_ ;
	assign \g1910/_0_  = _w15796_ ;
	assign \g19186/_0_  = _w13425_ ;
	assign \g19188/_0_  = _w13428_ ;
	assign \g19235/_0_  = _w15798_ ;
	assign \g19239/_0_  = _w15801_ ;
	assign \g19244/_0_  = _w15802_ ;
	assign \g19253/_0_  = _w15803_ ;
	assign \g19254/_0_  = _w15804_ ;
	assign \g19259/_0_  = _w15805_ ;
	assign \g19261/_0_  = _w15806_ ;
	assign \g19267/_0_  = _w15807_ ;
	assign \g19277/_0_  = _w15809_ ;
	assign \g19278/_0_  = _w15810_ ;
	assign \g19280/_0_  = _w15812_ ;
	assign \g19281/_0_  = _w15813_ ;
	assign \g19282/_0_  = _w15814_ ;
	assign \g19283/_0_  = _w15815_ ;
	assign \g19284/_0_  = _w15816_ ;
	assign \g19285/_0_  = _w15817_ ;
	assign \g19286/_0_  = _w15818_ ;
	assign \g19287/_0_  = _w15819_ ;
	assign \g19288/_0_  = _w15820_ ;
	assign \g19289/_0_  = _w15821_ ;
	assign \g19290/_0_  = _w15822_ ;
	assign \g19291/_0_  = _w15825_ ;
	assign \g19292/_0_  = _w15828_ ;
	assign \g19293/_0_  = _w15829_ ;
	assign \g19294/_0_  = _w15830_ ;
	assign \g19295/_0_  = _w15831_ ;
	assign \g19296/_0_  = _w15832_ ;
	assign \g19297/_0_  = _w15833_ ;
	assign \g19298/_0_  = _w15834_ ;
	assign \g19299/_0_  = _w15835_ ;
	assign \g19300/_0_  = _w15836_ ;
	assign \g19301/_0_  = _w15837_ ;
	assign \g19302/_0_  = _w15838_ ;
	assign \g19303/_0_  = _w15839_ ;
	assign \g19304/_0_  = _w15842_ ;
	assign \g19305/_0_  = _w15845_ ;
	assign \g19306/_0_  = _w15846_ ;
	assign \g19307/_0_  = _w15847_ ;
	assign \g19308/_0_  = _w15848_ ;
	assign \g19315/_0_  = _w15849_ ;
	assign \g19316/_0_  = _w15850_ ;
	assign \g19317/_0_  = _w15851_ ;
	assign \g19318/_0_  = _w15852_ ;
	assign \g19319/_0_  = _w15853_ ;
	assign \g19320/_0_  = _w15856_ ;
	assign \g19321/_0_  = _w15857_ ;
	assign \g19322/_0_  = _w15858_ ;
	assign \g19323/_0_  = _w15859_ ;
	assign \g19325/_3_  = _w15864_ ;
	assign \g19326/_3_  = _w15869_ ;
	assign \g19333/_3_  = _w15874_ ;
	assign \g19341/_3_  = _w15879_ ;
	assign \g19347/_3_  = _w15884_ ;
	assign \g19377/_3_  = _w15887_ ;
	assign \g19381/_3_  = _w15892_ ;
	assign \g19393/_0_  = _w15894_ ;
	assign \g19401/_0_  = _w15900_ ;
	assign \g19402/_0_  = _w15906_ ;
	assign \g195/_2_  = _w9296_ ;
	assign \g19513/_0_  = _w15907_ ;
	assign \g19514/_0_  = _w15908_ ;
	assign \g19515/_0_  = _w15909_ ;
	assign \g19516/_0_  = _w15910_ ;
	assign \g1952/_3_  = _w15915_ ;
	assign \g19529/_0_  = _w15916_ ;
	assign \g19530/_0_  = _w15917_ ;
	assign \g19531/_0_  = _w15918_ ;
	assign \g19532/_0_  = _w15919_ ;
	assign \g19533/_0_  = _w15920_ ;
	assign \g19534/_0_  = _w15921_ ;
	assign \g19535/_0_  = _w15922_ ;
	assign \g19536/_0_  = _w15923_ ;
	assign \g19537/_0_  = _w15924_ ;
	assign \g19539/_0_  = _w15925_ ;
	assign \g19546/_0_  = _w15926_ ;
	assign \g19552/_0_  = _w15927_ ;
	assign \g19553/_0_  = _w15928_ ;
	assign \g19562/_0_  = _w15931_ ;
	assign \g19563/_0_  = _w15934_ ;
	assign \g19564/_0_  = _w15937_ ;
	assign \g19572/_0_  = _w12391_ ;
	assign \g19575/_0_  = _w15938_ ;
	assign \g19615/_0_  = _w15939_ ;
	assign \g19686/_0_  = _w15940_ ;
	assign \g19688/_0_  = _w15941_ ;
	assign \g197/_0_  = _w15973_ ;
	assign \g19729/_0_  = _w15974_ ;
	assign \g19774/_0_  = _w15975_ ;
	assign \g19777/_0_  = _w15976_ ;
	assign \g19791/_0_  = _w15979_ ;
	assign \g19818/_0_  = _w15981_ ;
	assign \g19819/_0_  = _w15982_ ;
	assign \g19828/_0_  = _w15983_ ;
	assign \g19852/_1_  = _w5084_ ;
	assign \g19860/_0_  = _w15984_ ;
	assign \g19861/_0_  = _w15985_ ;
	assign \g19864/_0_  = _w15986_ ;
	assign \g19886/_0_  = _w15987_ ;
	assign \g19887/_0_  = _w15989_ ;
	assign \g199/_0_  = _w15999_ ;
	assign \g19908/_0_  = _w16000_ ;
	assign \g19918/_0_  = _w16003_ ;
	assign \g19927/_0_  = _w16004_ ;
	assign \g19933/_0_  = _w16005_ ;
	assign \g200/_0_  = _w14410_ ;
	assign \g20019/_0_  = _w16008_ ;
	assign \g20046/_0_  = _w16009_ ;
	assign \g20068/_1_  = _w14973_ ;
	assign \g20080/_1_  = _w14996_ ;
	assign \g201/_0_  = _w16027_ ;
	assign \g20137/_0_  = _w16028_ ;
	assign \g20139/_0_  = _w16033_ ;
	assign \g20141/_0_  = _w16034_ ;
	assign \g20152/_1_  = _w5092_ ;
	assign \g20154/_00_  = _w16038_ ;
	assign \g202/_0_  = _w16056_ ;
	assign \g20206/_0_  = _w16059_ ;
	assign \g20211/_2_  = _w16060_ ;
	assign \g20217/_2_  = _w16061_ ;
	assign \g20239/_0_  = _w16063_ ;
	assign \g20265/_2_  = _w16064_ ;
	assign \g20266/_0_  = _w16066_ ;
	assign \g20272/_2_  = _w16067_ ;
	assign \g20278/_2_  = _w16068_ ;
	assign \g20283/_0_  = _w11740_ ;
	assign \g20285/_2_  = _w16069_ ;
	assign \g20288/_2__syn_2  = _w14649_ ;
	assign \g20293/_0_  = _w16070_ ;
	assign \g20295/_2_  = _w13162_ ;
	assign \g203/_0_  = _w14435_ ;
	assign \g20302/_2_  = _w16071_ ;
	assign \g20303/_2_  = _w16072_ ;
	assign \g20304/_2_  = _w16073_ ;
	assign \g20311/_2_  = _w16074_ ;
	assign \g20326/_0_  = _w16078_ ;
	assign \g20330/_0_  = _w16080_ ;
	assign \g2034/_0_  = _w16083_ ;
	assign \g20345/_0_  = _w16087_ ;
	assign \g20346/_0_  = _w16090_ ;
	assign \g2035/_0_  = _w16091_ ;
	assign \g20363/_0_  = _w13326_ ;
	assign \g20364/_0_  = _w16095_ ;
	assign \g204/_0_  = _w16105_ ;
	assign \g2047/_0_  = _w16107_ ;
	assign \g20483/_0_  = _w16110_ ;
	assign \g20493/_00_  = _w16113_ ;
	assign \g205/_0_  = _w16117_ ;
	assign \g20569/_0_  = _w16118_ ;
	assign \g20570/_0_  = _w16119_ ;
	assign \g20571/_0_  = _w16120_ ;
	assign \g206/_0_  = _w16121_ ;
	assign \g20613/_0_  = _w16122_ ;
	assign \g20615/_0_  = _w16123_ ;
	assign \g20657/_1__syn_2  = _w16124_ ;
	assign \g20660/_0_  = _w16125_ ;
	assign \g20685/_0_  = _w16127_ ;
	assign \g207/_0_  = _w16128_ ;
	assign \g20713/_1_  = _w16129_ ;
	assign \g20747/_1_  = _w16130_ ;
	assign \g20784/_0_  = _w14454_ ;
	assign \g20820/_1_  = _w15535_ ;
	assign \g20859/_0_  = _w16132_ ;
	assign \g20873/_2_  = _w16133_ ;
	assign \g20886/_0_  = _w16134_ ;
	assign \g20887/_0_  = _w16135_ ;
	assign \g20891/_2__syn_2  = _w15876_ ;
	assign \g20907/_2_  = _w15557_ ;
	assign \g20936/_2__syn_2  = _w15871_ ;
	assign \g20937/_1_  = _w16136_ ;
	assign \g20955/_0_  = _w16137_ ;
	assign \g20959/_2__syn_2  = _w15866_ ;
	assign \g20967/_0_  = _w16138_ ;
	assign \g20971/_2__syn_2  = _w15889_ ;
	assign \g20974/_1__syn_2  = _w15893_ ;
	assign \g21015/_1_  = _w16139_ ;
	assign \g21051/_2_  = _w15547_ ;
	assign \g21079/_1_  = _w16140_ ;
	assign \g21081/_1_  = _w16141_ ;
	assign \g21087/_2__syn_2  = _w15881_ ;
	assign \g21114/_1_  = _w16142_ ;
	assign \g21116/_1_  = _w16143_ ;
	assign \g21120/_2__syn_2  = _w15861_ ;
	assign \g21147/_0_  = _w16144_ ;
	assign \g21179/_1_  = _w16145_ ;
	assign \g21185/_1_  = _w16146_ ;
	assign \g21223/_0_  = _w16147_ ;
	assign \g21242/_0_  = _w16148_ ;
	assign \g21253/_0_  = _w16149_ ;
	assign \g21257/_0_  = _w16151_ ;
	assign \g21323/_1_  = _w16152_ ;
	assign \g21324/_1_  = _w16153_ ;
	assign \g21366/_0_  = _w16155_ ;
	assign \g21385/_2_  = _w16157_ ;
	assign \g21464/_0_  = _w16159_ ;
	assign \g21475/_3_  = _w16160_ ;
	assign \g21481/_0_  = _w16163_ ;
	assign \g21482/_0_  = _w16165_ ;
	assign \g21494/_3_  = _w16166_ ;
	assign \g21500/_3_  = _w16167_ ;
	assign \g21507/_3_  = _w16168_ ;
	assign \g21511/_3_  = _w16169_ ;
	assign \g21537/_1_  = _w16171_ ;
	assign \g21568/_0_  = _w16172_ ;
	assign \g21591/_0_  = _w16173_ ;
	assign \g21604/_0_  = _w16175_ ;
	assign \g21605/_3_  = _w12913_ ;
	assign \g21606/_0_  = _w16176_ ;
	assign \g21607/_0_  = _w16177_ ;
	assign \g21608/_0_  = _w16178_ ;
	assign \g21609/_0_  = _w16179_ ;
	assign \g21610/_0_  = _w16180_ ;
	assign \g21611/_0_  = _w16181_ ;
	assign \g21612/_0_  = _w16182_ ;
	assign \g21613/_0_  = _w16183_ ;
	assign \g21614/_0_  = _w16184_ ;
	assign \g21615/_0_  = _w16185_ ;
	assign \g21616/_0_  = _w16186_ ;
	assign \g21617/_0_  = _w16187_ ;
	assign \g21618/_0_  = _w16188_ ;
	assign \g21621/_0_  = _w16190_ ;
	assign \g21640/_0_  = _w16191_ ;
	assign \g21678/_0_  = _w16192_ ;
	assign \g21679/_0_  = _w16193_ ;
	assign \g21686/_0_  = _w16194_ ;
	assign \g21692/_3_  = _w15053_ ;
	assign \g21696/_0_  = _w16197_ ;
	assign \g21698/_0_  = _w16200_ ;
	assign \g21702/_3_  = _w13000_ ;
	assign \g21707/_0_  = _w16201_ ;
	assign \g21709/_0_  = _w16202_ ;
	assign \g21728/_0_  = _w16205_ ;
	assign \g21729/_0_  = _w16208_ ;
	assign \g21731/_0_  = _w16211_ ;
	assign \g21732/_0_  = _w16214_ ;
	assign \g21733/_0_  = _w16217_ ;
	assign \g21736/_0_  = _w16218_ ;
	assign \g21744/_3_  = _w12992_ ;
	assign \g21753/_0_  = _w16219_ ;
	assign \g21754/_0_  = _w16220_ ;
	assign \g21755/_0_  = _w16221_ ;
	assign \g21756/_0_  = _w16222_ ;
	assign \g21757/_0_  = _w16223_ ;
	assign \g21759/_0_  = _w16224_ ;
	assign \g21761/_0_  = _w16225_ ;
	assign \g21763/_0_  = _w16226_ ;
	assign \g21764/_0_  = _w16227_ ;
	assign \g21766/_0_  = _w16228_ ;
	assign \g2180/_0_  = _w16237_ ;
	assign \g21853/_3_  = _w14929_ ;
	assign \g21861/_3_  = _w15063_ ;
	assign \g21863/_3_  = _w15069_ ;
	assign \g21869/_3_  = _w12923_ ;
	assign \g2187/_0_  = _w16250_ ;
	assign \g21875/_3_  = _w15072_ ;
	assign \g21877/_3_  = _w15083_ ;
	assign \g21879/_3_  = _w15058_ ;
	assign \g2188/_0_  = _w16251_ ;
	assign \g21900/_0_  = _w16252_ ;
	assign \g22080/_0_  = _w16253_ ;
	assign \g22082/_0_  = _w16254_ ;
	assign \g22135/_0_  = _w16255_ ;
	assign \g22145/_1_  = _w16256_ ;
	assign \g22225/_0_  = _w16257_ ;
	assign \g223/_0_  = _w15501_ ;
	assign \g22354/_0_  = _w16258_ ;
	assign \g224/_0_  = _w15455_ ;
	assign \g22412/_0_  = _w16261_ ;
	assign \g22415/_1__syn_2  = _w14450_ ;
	assign \g225/_0_  = _w15473_ ;
	assign \g2257/_0_  = _w4769_ ;
	assign \g226/_3_  = _w16271_ ;
	assign \g22624/_0_  = _w16272_ ;
	assign \g227/_3_  = _w16276_ ;
	assign \g22702/_0_  = _w16277_ ;
	assign \g22919/_1__syn_2  = _w16084_ ;
	assign \g22933/_0_  = _w16279_ ;
	assign \g22954/_0_  = _w16281_ ;
	assign \g22989/_1_  = _w16282_ ;
	assign \g23529/_0_  = _w556_ ;
	assign \g23539/_0_  = _w552_ ;
	assign \g2362/_2_  = _w16322_ ;
	assign \g23766/_0_  = _w576_ ;
	assign \g24/_3_  = _w16323_ ;
	assign \g24018/_0_  = _w548_ ;
	assign \g2416/_0_  = _w16502_ ;
	assign \g2420/_0_  = _w16505_ ;
	assign \g24213/_0_  = _w558_ ;
	assign \g24301/_0_  = _w550_ ;
	assign \g2479/_0_  = _w16552_ ;
	assign \g248/_3_  = _w16563_ ;
	assign \g2480/_0_  = _w16583_ ;
	assign \g2481/_0_  = _w16603_ ;
	assign \g2482/_0_  = _w16623_ ;
	assign \g2483/_0_  = _w16643_ ;
	assign \g2484/_0_  = _w16663_ ;
	assign \g2485/_0_  = _w16683_ ;
	assign \g2486/_0_  = _w16703_ ;
	assign \g2487/_0_  = _w16723_ ;
	assign \g2488/_0_  = _w16743_ ;
	assign \g249/_3_  = _w16747_ ;
	assign \g2490/_0_  = _w16767_ ;
	assign \g2491/_0_  = _w16787_ ;
	assign \g2492/_0_  = _w16807_ ;
	assign \g2493/_0_  = _w16827_ ;
	assign \g2494/_0_  = _w16847_ ;
	assign \g2495/_0_  = _w16867_ ;
	assign \g2496/_0_  = _w16872_ ;
	assign \g2497/_0_  = _w16873_ ;
	assign \g2507/_0_  = _w16882_ ;
	assign \g2508/_0_  = _w16889_ ;
	assign \g2509/_0_  = _w16897_ ;
	assign \g2510/_0_  = _w16905_ ;
	assign \g2511/_0_  = _w16913_ ;
	assign \g2512/_0_  = _w16921_ ;
	assign \g2513/_0_  = _w16929_ ;
	assign \g2514/_0_  = _w16946_ ;
	assign \g2515/_0_  = _w16963_ ;
	assign \g2516/_0_  = _w16971_ ;
	assign \g25237/_0_  = _w554_ ;
	assign \g2558/_0_  = _w16974_ ;
	assign \g2562/_0_  = _w16992_ ;
	assign \g2563/_0_  = _w17010_ ;
	assign \g2564/_0_  = _w17028_ ;
	assign \g2565/_0_  = _w17046_ ;
	assign \g2566/_0_  = _w17064_ ;
	assign \g2567/_0_  = _w17082_ ;
	assign \g2699/_0_  = _w16321_ ;
	assign \g27/_2_  = _w17086_ ;
	assign \g271/_0_  = _w16270_ ;
	assign \g272/_3_  = _w17096_ ;
	assign \g273/_3_  = _w17105_ ;
	assign \g274/_3_  = _w17109_ ;
	assign \g275/_3_  = _w17113_ ;
	assign \g276/_3_  = _w17119_ ;
	assign \g277/_3_  = _w17123_ ;
	assign \g2787/_3_  = _w17129_ ;
	assign \g2788/_3_  = _w17134_ ;
	assign \g279/_0_  = _w17140_ ;
	assign \g2795/_0_  = _w17143_ ;
	assign \g2796/_0_  = _w17144_ ;
	assign \g280/_0_  = _w17148_ ;
	assign \g2842/_3_  = _w17157_ ;
	assign \g29/_1_  = _w17159_ ;
	assign \g2927/_0_  = _w17295_ ;
	assign \g2978/_0_  = _w17301_ ;
	assign \g2979/_0_  = _w17304_ ;
	assign \g2980/_0_  = _w17307_ ;
	assign \g2981/_0_  = _w17310_ ;
	assign \g2982/_0_  = _w17313_ ;
	assign \g2983/_0_  = _w17316_ ;
	assign \g2984/_0_  = _w17319_ ;
	assign \g2985/_0_  = _w17322_ ;
	assign \g3021/_3_  = _w17326_ ;
	assign \g3022/_3_  = _w17329_ ;
	assign \g3023/_3_  = _w17332_ ;
	assign \g3024/_3_  = _w17335_ ;
	assign \g3025/_3_  = _w17338_ ;
	assign \g3026/_3_  = _w17341_ ;
	assign \g3027/_3_  = _w17344_ ;
	assign \g3028/_3_  = _w17347_ ;
	assign \g3029/_3_  = _w17352_ ;
	assign \g3030/_3_  = _w17357_ ;
	assign \g3031/_3_  = _w17362_ ;
	assign \g3032/_3_  = _w17367_ ;
	assign \g3033/_3_  = _w17372_ ;
	assign \g3034/_3_  = _w17377_ ;
	assign \g3035/_3_  = _w17382_ ;
	assign \g3036/_3_  = _w17387_ ;
	assign \g3037/_3_  = _w17390_ ;
	assign \g3038/_3_  = _w17393_ ;
	assign \g3039/_3_  = _w17396_ ;
	assign \g3040/_3_  = _w17399_ ;
	assign \g3041/_3_  = _w17402_ ;
	assign \g3042/_3_  = _w17405_ ;
	assign \g3049/_0_  = _w17407_ ;
	assign \g3050/_0_  = _w17409_ ;
	assign \g3051/_0_  = _w17411_ ;
	assign \g3052/_0_  = _w17413_ ;
	assign \g3053/_0_  = _w17415_ ;
	assign \g3054/_0_  = _w17417_ ;
	assign \g3058/_0_  = _w17419_ ;
	assign \g3059/_0_  = _w17421_ ;
	assign \g3088/_0_  = _w17426_ ;
	assign \g3089/_0_  = _w17430_ ;
	assign \g3090/_0_  = _w17434_ ;
	assign \g3091/_0_  = _w17438_ ;
	assign \g3092/_0_  = _w17443_ ;
	assign \g3093/_0_  = _w17448_ ;
	assign \g3094/_0_  = _w17452_ ;
	assign \g3095/_0_  = _w17456_ ;
	assign \g314/_0_  = _w16562_ ;
	assign \g3147/_3_  = _w17459_ ;
	assign \g3148/_3_  = _w17462_ ;
	assign \g3189/_0_  = _w17465_ ;
	assign \g3190/_0_  = _w17468_ ;
	assign \g3191/_0_  = _w17471_ ;
	assign \g3192/_0_  = _w17474_ ;
	assign \g3193/_0_  = _w17477_ ;
	assign \g3194/_0_  = _w17480_ ;
	assign \g3195/_0_  = _w17484_ ;
	assign \g3196/_0_  = _w17488_ ;
	assign \g3197/_0_  = _w17492_ ;
	assign \g3198/_0_  = _w17496_ ;
	assign \g3199/_0_  = _w17499_ ;
	assign \g32/_0_  = _w17510_ ;
	assign \g320/_3_  = _w17597_ ;
	assign \g3200/_0_  = _w17601_ ;
	assign \g3201/_0_  = _w17605_ ;
	assign \g3202/_0_  = _w17609_ ;
	assign \g3203/_0_  = _w17613_ ;
	assign \g3204/_0_  = _w17616_ ;
	assign \g321/_3_  = _w17646_ ;
	assign \g325/_3_  = _w17650_ ;
	assign \g3271/_2_  = _w16314_ ;
	assign \g33/_0_  = _w17656_ ;
	assign \g3363/_0_  = _w17663_ ;
	assign \g3413/_0_  = _w17699_ ;
	assign \g3414/_0_  = _w17735_ ;
	assign \g352/_0_  = _w17095_ ;
	assign \g355/_0_  = _w17104_ ;
	assign \g356/_3_  = _w17741_ ;
	assign \g357/_3_  = _w17746_ ;
	assign \g35_dup/_1_  = _w17747_ ;
	assign \g36/_3_  = _w17748_ ;
	assign \g365/_3_  = _w17786_ ;
	assign \g366/_3_  = _w17848_ ;
	assign \g367/_3_  = _w17886_ ;
	assign \g368/_3_  = _w17922_ ;
	assign \g3687/_0_  = _w17924_ ;
	assign \g369/_3_  = _w17990_ ;
	assign \g37/_3_  = _w17991_ ;
	assign \g370/_3_  = _w18004_ ;
	assign \g372/_3_  = _w18017_ ;
	assign \g374/_3_  = _w18030_ ;
	assign \g3740/_0_  = _w18032_ ;
	assign \g375/_3_  = _w18045_ ;
	assign \g376/_3_  = _w18057_ ;
	assign \g3878/_0_  = _w18061_ ;
	assign \g3879/_0_  = _w18063_ ;
	assign \g388/_3_  = _w18069_ ;
	assign \g3880/_0_  = _w18074_ ;
	assign \g3881/_0_  = _w18076_ ;
	assign \g3882/_0_  = _w18080_ ;
	assign \g389/_3_  = _w18085_ ;
	assign \g3894/_0_  = _w18086_ ;
	assign \g3895/_0_  = _w18087_ ;
	assign \g3896/_0_  = _w18088_ ;
	assign \g3897/_0_  = _w18089_ ;
	assign \g3898/_0_  = _w18090_ ;
	assign \g392/_3_  = _w18187_ ;
	assign \g393/_3_  = _w18228_ ;
	assign \g394/_3_  = _w18331_ ;
	assign \g395/_3_  = _w18397_ ;
	assign \g396/_3_  = _w18401_ ;
	assign \g397/_3_  = _w18405_ ;
	assign \g398/_3_  = _w18409_ ;
	assign \g399/_3_  = _w18413_ ;
	assign \g401/_3_  = _w18501_ ;
	assign \g402/_3_  = _w18505_ ;
	assign \g404/_3_  = _w18571_ ;
	assign \g4048/_0_  = _w18573_ ;
	assign \g405/_3_  = _w18614_ ;
	assign \g4050/_0_  = _w18616_ ;
	assign \g406/_3_  = _w18619_ ;
	assign \g407/_3_  = _w18623_ ;
	assign \g410/_3_  = _w18714_ ;
	assign \g411/_3_  = _w18718_ ;
	assign \g412/_3_  = _w18753_ ;
	assign \g413/_3_  = _w18821_ ;
	assign \g415/_3_  = _w18834_ ;
	assign \g416/_3_  = _w18847_ ;
	assign \g42/_0_  = _w18853_ ;
	assign \g4216/_3_  = _w18859_ ;
	assign \g4217/_3_  = _w18863_ ;
	assign \g4218/_3_  = _w18865_ ;
	assign \g4219/_3_  = _w18874_ ;
	assign \g4296/_0_  = _w18888_ ;
	assign \g4297/_0_  = _w18902_ ;
	assign \g4298/_0_  = _w18906_ ;
	assign \g4299/_0_  = _w18910_ ;
	assign \g43/_0_  = _w18915_ ;
	assign \g4300/_0_  = _w18919_ ;
	assign \g4301/_0_  = _w18923_ ;
	assign \g4302/_0_  = _w18927_ ;
	assign \g4303/_0_  = _w18931_ ;
	assign \g4304/_0_  = _w18935_ ;
	assign \g4305/_0_  = _w18939_ ;
	assign \g4306/_0_  = _w18943_ ;
	assign \g4307/_0_  = _w18947_ ;
	assign \g4308/_0_  = _w18951_ ;
	assign \g4309/_0_  = _w18955_ ;
	assign \g4310/_0_  = _w18959_ ;
	assign \g4311/_0_  = _w18963_ ;
	assign \g4312/_0_  = _w18967_ ;
	assign \g4313/_0_  = _w18971_ ;
	assign \g4314/_0_  = _w18975_ ;
	assign \g4315/_0_  = _w18979_ ;
	assign \g4316/_0_  = _w18983_ ;
	assign \g4317/_0_  = _w18987_ ;
	assign \g4318/_0_  = _w18991_ ;
	assign \g4319/_0_  = _w18995_ ;
	assign \g4320/_0_  = _w18999_ ;
	assign \g4321/_0_  = _w19003_ ;
	assign \g4322/_0_  = _w19007_ ;
	assign \g4323/_0_  = _w19011_ ;
	assign \g436/_0_  = _w19013_ ;
	assign \g44/_0_  = _w19019_ ;
	assign \g448/_3_  = _w19023_ ;
	assign \g45/_0_  = _w19030_ ;
	assign \g4587/_0_  = _w19069_ ;
	assign \g4588/_0_  = _w19071_ ;
	assign \g46/_0_  = _w11298_ ;
	assign \g4601/_0_  = _w19073_ ;
	assign \g4602/_0_  = _w19075_ ;
	assign \g4613/_3_  = _w19079_ ;
	assign \g4614/_3_  = _w19085_ ;
	assign \g4615/_3_  = _w19090_ ;
	assign \g463/_0_  = _w19110_ ;
	assign \g465/_0_  = _w19115_ ;
	assign \g4653/_0_  = _w19138_ ;
	assign \g4654/_0_  = _w19145_ ;
	assign \g4655/_0_  = _w19148_ ;
	assign \g4656/_0_  = _w19150_ ;
	assign \g4659/_0_  = _w19151_ ;
	assign \g466/_0_  = _w19155_ ;
	assign \g468/_3_  = _w19162_ ;
	assign \g469/_3_  = _w19167_ ;
	assign \g4697/_0_  = _w19168_ ;
	assign \g47/_3_  = _w19175_ ;
	assign \g470/_0_  = _w19181_ ;
	assign \g471/_0_  = _w19182_ ;
	assign \g4755/_0_  = _w19183_ ;
	assign \g476/_0_  = _w19204_ ;
	assign \g48/_3_  = _w19209_ ;
	assign \g480/_00_  = _w19227_ ;
	assign \g4839/_0_  = _w19243_ ;
	assign \g4840/_0_  = _w19245_ ;
	assign \g485/_3_  = _w19246_ ;
	assign \g4854/_0_  = _w19248_ ;
	assign \g4855/_0_  = _w19250_ ;
	assign \g4859/_0_  = _w19252_ ;
	assign \g486/_3_  = _w19253_ ;
	assign \g4860/_0_  = _w19255_ ;
	assign \g4880/_0_  = _w19286_ ;
	assign \g4881/_0_  = _w19295_ ;
	assign \g4882/_0_  = _w19305_ ;
	assign \g4883/_0_  = _w19315_ ;
	assign \g4884/_0_  = _w19338_ ;
	assign \g4885/_0_  = _w19348_ ;
	assign \g4886/_0_  = _w19357_ ;
	assign \g4887/_0_  = _w19367_ ;
	assign \g4888/_0_  = _w19377_ ;
	assign \g49/_0_  = _w19384_ ;
	assign \g494/_0_  = _w4844_ ;
	assign \g499/_1_  = _w4826_ ;
	assign \g50/_0_  = _w19389_ ;
	assign \g5002/_0_  = _w19407_ ;
	assign \g5003/_0_  = _w19412_ ;
	assign \g5009/_0_  = _w19419_ ;
	assign \g5010/_0_  = _w19425_ ;
	assign \g5011/_0_  = _w19433_ ;
	assign \g5014/_0_  = _w19434_ ;
	assign \g51/_0_  = _w19436_ ;
	assign \g5105/_0_  = _w19437_ ;
	assign \g5129/_2_  = _w19442_ ;
	assign \g5132/_0_  = _w19456_ ;
	assign \g5135/_0_  = _w19470_ ;
	assign \g5168/_0_  = _w19480_ ;
	assign \g5169/_0_  = _w19482_ ;
	assign \g5173/_0_  = _w19484_ ;
	assign \g5224/_0_  = _w19487_ ;
	assign \g5225/_0_  = _w19490_ ;
	assign \g5226/_0_  = _w19492_ ;
	assign \g5227/_0_  = _w19494_ ;
	assign \g5334/_0_  = _w19506_ ;
	assign \g5335/_0_  = _w19510_ ;
	assign \g5336/_0_  = _w19514_ ;
	assign \g5337/_0_  = _w19517_ ;
	assign \g5338/_0_  = _w19524_ ;
	assign \g5339/_0_  = _w19531_ ;
	assign \g5340/_0_  = _w19538_ ;
	assign \g5341/_0_  = _w19545_ ;
	assign \g5342/_0_  = _w19552_ ;
	assign \g5343/_0_  = _w19559_ ;
	assign \g5344/_0_  = _w19566_ ;
	assign \g5345/_0_  = _w19573_ ;
	assign \g5346/_0_  = _w19580_ ;
	assign \g5347/_0_  = _w19587_ ;
	assign \g5348/_0_  = _w19594_ ;
	assign \g5349/_0_  = _w19601_ ;
	assign \g5395/_0_  = _w19602_ ;
	assign \g54/_0_  = _w19605_ ;
	assign \g5434/_0_  = _w19612_ ;
	assign \g5447/_0_  = _w19616_ ;
	assign \g5450/_0_  = _w19628_ ;
	assign \g5451/_0_  = _w19632_ ;
	assign \g5452/_0_  = _w19636_ ;
	assign \g5453/_0_  = _w19640_ ;
	assign \g5454/_0_  = _w19643_ ;
	assign \g5461/_0_  = _w19644_ ;
	assign \g5483/_0_  = _w19649_ ;
	assign \g5484/_0_  = _w19659_ ;
	assign \g5492/_0_  = _w19660_ ;
	assign \g5493/_0_  = _w19662_ ;
	assign \g5496/_3_  = _w19668_ ;
	assign \g5497/_3_  = _w19673_ ;
	assign \g55/_0_  = _w19676_ ;
	assign \g5500/_0_  = _w19679_ ;
	assign \g5502/_0_  = _w19698_ ;
	assign \g5503/_0_  = _w19737_ ;
	assign \g5506/_0_  = _w19742_ ;
	assign \g5511/_0_  = _w19775_ ;
	assign \g5518/_0_  = _w19785_ ;
	assign \g5519/_0_  = _w19794_ ;
	assign \g5520/_0_  = _w19803_ ;
	assign \g5522/_0_  = _w19813_ ;
	assign \g5523/_0_  = _w19823_ ;
	assign \g5524/_0_  = _w19833_ ;
	assign \g5525/_0_  = _w19843_ ;
	assign \g5532/_0_  = _w19846_ ;
	assign \g5533/_0_  = _w19849_ ;
	assign \g5534/_0_  = _w19852_ ;
	assign \g5535/_0_  = _w19855_ ;
	assign \g5536/_0_  = _w19857_ ;
	assign \g5537/_0_  = _w19859_ ;
	assign \g5538/_0_  = _w19861_ ;
	assign \g5546/_0_  = _w19865_ ;
	assign \g5555/_00_  = _w19884_ ;
	assign \g5593/_0_  = _w4139_ ;
	assign \g5614/_2_  = _w5568_ ;
	assign \g567/_0_  = _w19886_ ;
	assign \g5677/_0_  = _w19887_ ;
	assign \g5678/_0_  = _w19888_ ;
	assign \g5682/_0_  = _w19890_ ;
	assign \g5683/_0_  = _w19893_ ;
	assign \g5684/_0_  = _w19895_ ;
	assign \g5686/_0_  = _w19898_ ;
	assign \g5687/_0_  = _w19900_ ;
	assign \g5689/_0_  = _w19903_ ;
	assign \g5690/_0_  = _w19905_ ;
	assign \g5691/_0_  = _w19908_ ;
	assign \g5692/_0_  = _w19910_ ;
	assign \g5698/_0_  = _w19912_ ;
	assign \g5699/_0_  = _w19914_ ;
	assign \g5700/_0_  = _w19916_ ;
	assign \g5701/_0_  = _w19918_ ;
	assign \g5702/_0_  = _w19920_ ;
	assign \g5703/_0_  = _w19921_ ;
	assign \g5704/_0_  = _w19928_ ;
	assign \g5709/_0_  = _w19929_ ;
	assign \g5711/_0_  = _w19930_ ;
	assign \g5714/_0_  = _w19931_ ;
	assign \g572/_0_  = _w19934_ ;
	assign \g5723/_0_  = _w19939_ ;
	assign \g5724/_0_  = _w19944_ ;
	assign \g5725/_0_  = _w19963_ ;
	assign \g573/_0_  = _w19964_ ;
	assign \g5739/_0_  = _w19974_ ;
	assign \g5740/_0_  = _w19981_ ;
	assign \g575/_0_  = _w19982_ ;
	assign \g5756/_0_  = _w19983_ ;
	assign \g5757/_0_  = _w19984_ ;
	assign \g5758/_0_  = _w19985_ ;
	assign \g5759/_0_  = _w19986_ ;
	assign \g576/_0_  = _w19987_ ;
	assign \g5760/_0_  = _w19988_ ;
	assign \g5761/_0_  = _w19989_ ;
	assign \g5762/_0_  = _w19990_ ;
	assign \g5763/_0_  = _w19991_ ;
	assign \g577/_0_  = _w19992_ ;
	assign \g5772/_0_  = _w20006_ ;
	assign \g5773/_0_  = _w20010_ ;
	assign \g5774/_0_  = _w20016_ ;
	assign \g5775/_0_  = _w20022_ ;
	assign \g5776/_0_  = _w20025_ ;
	assign \g5777/_0_  = _w20028_ ;
	assign \g578/_0_  = _w20029_ ;
	assign \g5781/_0_  = _w20036_ ;
	assign \g5783/_0_  = _w20040_ ;
	assign \g5784/_0_  = _w20045_ ;
	assign \g5785/_0_  = _w20049_ ;
	assign \g5786/_0_  = _w20054_ ;
	assign \g5787/_0_  = _w20059_ ;
	assign \g5788/_0_  = _w20064_ ;
	assign \g5789/_0_  = _w20069_ ;
	assign \g579/_0_  = _w20070_ ;
	assign \g5790/_0_  = _w20071_ ;
	assign \g5791/_0_  = _w20072_ ;
	assign \g5792/_0_  = _w20073_ ;
	assign \g5794/_0_  = _w20084_ ;
	assign \g5795/_0_  = _w20085_ ;
	assign \g5796/_0_  = _w20086_ ;
	assign \g580/_0_  = _w20087_ ;
	assign \g5801/_0_  = _w20090_ ;
	assign \g5802/_0_  = _w20093_ ;
	assign \g5803/_0_  = _w20096_ ;
	assign \g5804/_0_  = _w20099_ ;
	assign \g5805/_0_  = _w20102_ ;
	assign \g581/_0_  = _w20103_ ;
	assign \g5814/_0_  = _w20114_ ;
	assign \g582/_0_  = _w20115_ ;
	assign \g583/_0_  = _w20116_ ;
	assign \g5849/_3_  = _w20121_ ;
	assign \g585/_0_  = _w20122_ ;
	assign \g586/_0_  = _w20123_ ;
	assign \g587/_0_  = _w20124_ ;
	assign \g588/_0_  = _w20125_ ;
	assign \g589/_0_  = _w20126_ ;
	assign \g590/_0_  = _w20127_ ;
	assign \g591/_0_  = _w20128_ ;
	assign \g592/_0_  = _w20129_ ;
	assign \g593/_0_  = _w20130_ ;
	assign \g594/_0_  = _w20131_ ;
	assign \g595/_0_  = _w20132_ ;
	assign \g596/_0_  = _w20133_ ;
	assign \g597/_0_  = _w20134_ ;
	assign \g5971/_0_  = _w20135_ ;
	assign \g5972/_0_  = _w20136_ ;
	assign \g5976/_0_  = _w20137_ ;
	assign \g598/_0_  = _w20138_ ;
	assign \g5989/_0_  = _w20139_ ;
	assign \g599/_0_  = _w20140_ ;
	assign \g600/_0_  = _w20141_ ;
	assign \g601/_0_  = _w20142_ ;
	assign \g602/_0_  = _w20143_ ;
	assign \g603/_0_  = _w20144_ ;
	assign \g604/_0_  = _w20145_ ;
	assign \g605/_0_  = _w20146_ ;
	assign \g6092/_0_  = _w20149_ ;
	assign \g6093/_2_  = _w20259_ ;
	assign \g6094/_0_  = _w20261_ ;
	assign \g6114/_0_  = _w20262_ ;
	assign \g614/_3_  = _w20266_ ;
	assign \g6148/_0_  = _w20268_ ;
	assign \g6149/_0_  = _w20270_ ;
	assign \g6171/_0_  = _w20291_ ;
	assign \g6172/_0_  = _w20301_ ;
	assign \g6173/_0_  = _w20311_ ;
	assign \g6174/_0_  = _w20321_ ;
	assign \g6175/_0_  = _w20331_ ;
	assign \g6176/_0_  = _w20341_ ;
	assign \g6177/_0_  = _w20351_ ;
	assign \g6178/_0_  = _w20375_ ;
	assign \g6179/_0_  = _w20384_ ;
	assign \g6180/_0_  = _w20393_ ;
	assign \g6181/_0_  = _w20402_ ;
	assign \g6182/_0_  = _w20411_ ;
	assign \g6183/_0_  = _w20420_ ;
	assign \g6184/_0_  = _w20429_ ;
	assign \g6185/_0_  = _w20438_ ;
	assign \g6186/_0_  = _w20454_ ;
	assign \g6187/_0_  = _w20471_ ;
	assign \g6193/_0_  = _w20487_ ;
	assign \g6196/_0_  = _w20501_ ;
	assign \g6197/_0_  = _w20508_ ;
	assign \g6198/_3_  = _w20517_ ;
	assign \g6200/_2_  = _w19497_ ;
	assign \g6202/_2_  = _w19619_ ;
	assign \g6203/_3_  = _w20523_ ;
	assign \g6204/_3_  = _w20528_ ;
	assign \g6209/_0_  = _w20539_ ;
	assign \g6211/_0_  = _w20540_ ;
	assign \g6215/_0_  = _w20554_ ;
	assign \g6217/_0_  = _w20568_ ;
	assign \g6219/_0_  = _w20582_ ;
	assign \g6220/_0_  = _w20596_ ;
	assign \g6222/_0_  = _w20610_ ;
	assign \g6224/_0_  = _w20626_ ;
	assign \g6228/_0_  = _w20642_ ;
	assign \g6238/_0_  = _w20643_ ;
	assign \g6239/_0_  = _w20644_ ;
	assign \g6240/_0_  = _w20645_ ;
	assign \g6242/_0_  = _w20646_ ;
	assign \g6243/_0_  = _w20649_ ;
	assign \g6244/_0_  = _w20650_ ;
	assign \g6245/_0_  = _w20651_ ;
	assign \g6246/_0_  = _w20652_ ;
	assign \g6248/_0_  = _w20655_ ;
	assign \g6249/_0_  = _w20656_ ;
	assign \g6259/_0_  = _w20659_ ;
	assign \g6260/_0_  = _w20662_ ;
	assign \g6261/_0_  = _w20664_ ;
	assign \g6262/_0_  = _w20666_ ;
	assign \g6263/_0_  = _w20668_ ;
	assign \g6264/_0_  = _w20670_ ;
	assign \g6265/_0_  = _w20672_ ;
	assign \g6266/_0_  = _w20675_ ;
	assign \g6267/_0_  = _w20678_ ;
	assign \g6268/_0_  = _w20680_ ;
	assign \g6269/_0_  = _w20682_ ;
	assign \g6270/_0_  = _w20684_ ;
	assign \g6271/_0_  = _w20685_ ;
	assign \g6272/_0_  = _w20687_ ;
	assign \g6277/_0_  = _w20689_ ;
	assign \g6318/_0_  = _w20690_ ;
	assign \g6326/_0_  = _w20693_ ;
	assign \g6329/_0_  = _w20703_ ;
	assign \g6330/_0_  = _w20713_ ;
	assign \g6331/_0_  = _w20722_ ;
	assign \g6332/_0_  = _w20732_ ;
	assign \g6333/_0_  = _w20747_ ;
	assign \g6334/_0_  = _w20753_ ;
	assign \g6335/_0_  = _w20759_ ;
	assign \g6336/_0_  = _w20765_ ;
	assign \g6337/_0_  = _w20771_ ;
	assign \g6338/_0_  = _w20777_ ;
	assign \g6339/_0_  = _w20783_ ;
	assign \g6340/_0_  = _w20790_ ;
	assign \g6341/_0_  = _w20796_ ;
	assign \g6342/_0_  = _w20802_ ;
	assign \g6343/_0_  = _w20811_ ;
	assign \g6344/_0_  = _w20820_ ;
	assign \g6345/_0_  = _w20828_ ;
	assign \g6346/_0_  = _w20836_ ;
	assign \g6347/_0_  = _w20845_ ;
	assign \g6348/_0_  = _w20854_ ;
	assign \g6349/_0_  = _w20869_ ;
	assign \g6350/_0_  = _w20879_ ;
	assign \g6351/_0_  = _w20889_ ;
	assign \g6352/_0_  = _w20898_ ;
	assign \g6353/_0_  = _w20907_ ;
	assign \g6354/_0_  = _w20916_ ;
	assign \g6355/_0_  = _w20925_ ;
	assign \g6361/_0_  = _w20926_ ;
	assign \g637/_0_  = _w20929_ ;
	assign \g638/_0_  = _w20930_ ;
	assign \g639/_3_  = _w20937_ ;
	assign \g64/_3_  = _w20938_ ;
	assign \g640/_3_  = _w20943_ ;
	assign \g6419/_0_  = _w4877_ ;
	assign \g6442/_0_  = _w8483_ ;
	assign \g6442/_1_  = _w8482_ ;
	assign \g6489/_0_  = _w20944_ ;
	assign \g6490/_0_  = _w20945_ ;
	assign \g65/_3_  = _w20946_ ;
	assign \g6513/_0_  = _w20948_ ;
	assign \g6515/_0_  = _w20950_ ;
	assign \g6571/_0_  = _w20970_ ;
	assign \g6588/_0_  = _w20972_ ;
	assign \g6589/_0_  = _w20974_ ;
	assign \g6638/_0_  = _w20978_ ;
	assign \g6639/_0_  = _w20989_ ;
	assign \g6653/_0_  = _w20992_ ;
	assign \g6654/_3_  = _w21004_ ;
	assign \g6655/_0_  = _w21006_ ;
	assign \g6656/_0_  = _w21009_ ;
	assign \g6657/_0_  = _w21011_ ;
	assign \g6687/_0_  = _w21026_ ;
	assign \g6688/_0_  = _w21030_ ;
	assign \g6689/_0_  = _w21034_ ;
	assign \g6690/_0_  = _w21038_ ;
	assign \g6691/_0_  = _w21042_ ;
	assign \g6692/_0_  = _w21046_ ;
	assign \g6693/_0_  = _w21050_ ;
	assign \g6694/_0_  = _w21054_ ;
	assign \g6701/_0_  = _w21055_ ;
	assign \g6706/_0_  = _w21057_ ;
	assign \g6711/_0_  = _w21058_ ;
	assign \g6727/_0_  = _w21073_ ;
	assign \g6728/_0_  = _w21089_ ;
	assign \g6736/_0_  = _w21090_ ;
	assign \g6739/_0_  = _w21106_ ;
	assign \g6742/_0_  = _w21109_ ;
	assign \g6746/_0_  = _w21110_ ;
	assign \g6752/_0_  = _w21113_ ;
	assign \g6771/_0_  = _w21114_ ;
	assign \g684/_0_  = _w21137_ ;
	assign \g685/_0_  = _w21140_ ;
	assign \g686/_0_  = _w21144_ ;
	assign \g687/_0_  = _w21145_ ;
	assign \g688/_0_  = _w21149_ ;
	assign \g689/_0_  = _w21150_ ;
	assign \g690/_0_  = _w21154_ ;
	assign \g691/_0_  = _w21155_ ;
	assign \g692/_0_  = _w21156_ ;
	assign \g693/_0_  = _w21157_ ;
	assign \g696/_3_  = _w21163_ ;
	assign \g697/_3_  = _w21167_ ;
	assign \g699/_0_  = _w21188_ ;
	assign \g7/_0_  = _w21195_ ;
	assign \g700/_0_  = _w21211_ ;
	assign \g7005/_0_  = _w21217_ ;
	assign \g7056/_0_  = _w21219_ ;
	assign \g7057/_0_  = _w19502_ ;
	assign \g7058/_0_  = _w19624_ ;
	assign \g7060/_0_  = _w21221_ ;
	assign \g7075/_0_  = _w21235_ ;
	assign \g7086/_0_  = _w21240_ ;
	assign \g7087/_0_  = _w21243_ ;
	assign \g7089/_0_  = _w21251_ ;
	assign \g7108/_0_  = _w21255_ ;
	assign \g7109/_0_  = _w21259_ ;
	assign \g7112/_0_  = _w19771_ ;
	assign \g7172/_2_  = _w20534_ ;
	assign \g7210/_2_  = _w20110_ ;
	assign \g7211/_0_  = _w21261_ ;
	assign \g7212/_0_  = _w21264_ ;
	assign \g7213/_0_  = _w21266_ ;
	assign \g7214/_0_  = _w21268_ ;
	assign \g7215/_0_  = _w21271_ ;
	assign \g7216/_0_  = _w21273_ ;
	assign \g7217/_3_  = _w21276_ ;
	assign \g7218/_0_  = _w21278_ ;
	assign \g7219/_0_  = _w21281_ ;
	assign \g7220/_0_  = _w21283_ ;
	assign \g7222/_0_  = _w21285_ ;
	assign \g7227/_2_  = _w20080_ ;
	assign \g723/_3_  = _w21286_ ;
	assign \g7234/_0_  = _w21290_ ;
	assign \g7237/_3_  = _w21292_ ;
	assign \g7238/_3_  = _w21295_ ;
	assign \g7239/_3_  = _w9434_ ;
	assign \g724/_3_  = _w21296_ ;
	assign \g7240/_3_  = _w21300_ ;
	assign \g7241/_3_  = _w21303_ ;
	assign \g7242/_3_  = _w21305_ ;
	assign \g7243/_3_  = _w21308_ ;
	assign \g7244/_0_  = _w21311_ ;
	assign \g7245/_0_  = _w21313_ ;
	assign \g7246/_0_  = _w21315_ ;
	assign \g7247/_0_  = _w21317_ ;
	assign \g7248/_0_  = _w21320_ ;
	assign \g7249/_0_  = _w21322_ ;
	assign \g7250/_0_  = _w21324_ ;
	assign \g7251/_0_  = _w21327_ ;
	assign \g7253/_0_  = _w21328_ ;
	assign \g7254/_0_  = _w21329_ ;
	assign \g7255/_0_  = _w21330_ ;
	assign \g7256/_0_  = _w21331_ ;
	assign \g7257/_0_  = _w21332_ ;
	assign \g7258/_0_  = _w21333_ ;
	assign \g7261/_0_  = _w21334_ ;
	assign \g7264/_0_  = _w21343_ ;
	assign \g7265/_0_  = _w21353_ ;
	assign \g7266/_0_  = _w21359_ ;
	assign \g7267/_0_  = _w21365_ ;
	assign \g7268/_0_  = _w21371_ ;
	assign \g7269/_0_  = _w21380_ ;
	assign \g7278/_0_  = _w21390_ ;
	assign \g7279/_0_  = _w21396_ ;
	assign \g7280/_0_  = _w21406_ ;
	assign \g7281/_0_  = _w21415_ ;
	assign \g7282/_0_  = _w21424_ ;
	assign \g7283/_0_  = _w21433_ ;
	assign \g7284/_0_  = _w21443_ ;
	assign \g7285/_0_  = _w21453_ ;
	assign \g7286/_3_  = _w16512_ ;
	assign \g7288/_3_  = _w21456_ ;
	assign \g7291/_0_  = _w21457_ ;
	assign \g7296/_3_  = _w21475_ ;
	assign \g73/_0_  = _w21481_ ;
	assign \g7302/_3_  = _w21494_ ;
	assign \g7306/_3_  = _w21507_ ;
	assign \g7310/_3_  = _w21513_ ;
	assign \g7311/_3_  = _w21517_ ;
	assign \g7312/_3_  = _w21521_ ;
	assign \g7313/_3_  = _w21525_ ;
	assign \g7314/_3_  = _w21529_ ;
	assign \g7315/_3_  = _w21533_ ;
	assign \g7316/_3_  = _w21537_ ;
	assign \g7317/_3_  = _w21541_ ;
	assign \g7323/_3_  = _w21556_ ;
	assign \g7324/_3_  = _w21570_ ;
	assign \g7325/_3_  = _w21584_ ;
	assign \g7327/_0_  = _w21585_ ;
	assign \g7362/_0_  = _w21586_ ;
	assign \g74/_0_  = _w21592_ ;
	assign \g75/_0_  = _w21598_ ;
	assign \g7512/_0_  = _w9424_ ;
	assign \g7513/_0_  = _w21603_ ;
	assign \g7514/_0_  = _w21604_ ;
	assign \g7515/_0_  = _w21605_ ;
	assign \g7516/_0_  = _w21606_ ;
	assign \g7518/_0_  = _w21612_ ;
	assign \g7528/_0_  = _w21618_ ;
	assign \g7529/_0_  = _w21619_ ;
	assign \g7548/_0_  = _w21622_ ;
	assign \g7549/_0_  = _w21624_ ;
	assign \g7550/_0_  = _w21628_ ;
	assign \g7575/_0_  = _w21633_ ;
	assign \g7576/_0_  = _w21636_ ;
	assign \g7577/_0_  = _w21639_ ;
	assign \g7578/_0_  = _w21641_ ;
	assign \g7579/_0_  = _w21647_ ;
	assign \g7580/_0_  = _w21650_ ;
	assign \g7581/_0_  = _w21653_ ;
	assign \g7582/_0_  = _w21656_ ;
	assign \g7583/_0_  = _w21659_ ;
	assign \g7584/_0_  = _w21663_ ;
	assign \g7585/_0_  = _w21667_ ;
	assign \g7586/_0_  = _w21671_ ;
	assign \g7587/_0_  = _w21675_ ;
	assign \g7588/_0_  = _w21678_ ;
	assign \g7589/_0_  = _w21681_ ;
	assign \g7590/_0_  = _w21684_ ;
	assign \g7591/_0_  = _w21687_ ;
	assign \g7592/_0_  = _w21690_ ;
	assign \g7593/_0_  = _w21693_ ;
	assign \g7594/_0_  = _w21695_ ;
	assign \g7595/_0_  = _w21698_ ;
	assign \g7596/_0_  = _w21701_ ;
	assign \g7597/_0_  = _w21705_ ;
	assign \g7598/_0_  = _w21708_ ;
	assign \g7599/_0_  = _w21711_ ;
	assign \g76/_0_  = _w21717_ ;
	assign \g7600/_0_  = _w21720_ ;
	assign \g7601/_0_  = _w21723_ ;
	assign \g7602/_0_  = _w21725_ ;
	assign \g7603/_0_  = _w21728_ ;
	assign \g7604/_0_  = _w21731_ ;
	assign \g7614/_0_  = _w21733_ ;
	assign \g7618/_0_  = _w21734_ ;
	assign \g762/_0_  = _w21736_ ;
	assign \g7634/_0_  = _w20147_ ;
	assign \g766/_0_  = _w21739_ ;
	assign \g767/_0_  = _w21740_ ;
	assign \g768/_0_  = _w21743_ ;
	assign \g769/_0_  = _w21744_ ;
	assign \g77/_0_  = _w21750_ ;
	assign \g770/_3_  = _w21757_ ;
	assign \g771/_3_  = _w21762_ ;
	assign \g7715/_0_  = _w21773_ ;
	assign \g774/_0_  = _w21784_ ;
	assign \g7746/_0_  = _w21787_ ;
	assign \g7753/_0_  = _w21789_ ;
	assign \g7754/_0_  = _w21790_ ;
	assign \g7755/_0_  = _w21791_ ;
	assign \g7756/_0_  = _w21792_ ;
	assign \g7757/_0_  = _w21793_ ;
	assign \g7758/_0_  = _w21808_ ;
	assign \g7759/_0_  = _w21823_ ;
	assign \g7760/_0_  = _w21837_ ;
	assign \g7761/_0_  = _w21850_ ;
	assign \g7762/_0_  = _w21851_ ;
	assign \g7763/_0_  = _w21852_ ;
	assign \g7764/_0_  = _w21853_ ;
	assign \g7765/_0_  = _w21854_ ;
	assign \g7766/_0_  = _w21867_ ;
	assign \g7778/_0_  = _w21869_ ;
	assign \g7779/_0_  = _w21871_ ;
	assign \g7780/_0_  = _w21874_ ;
	assign \g7781/_0_  = _w21876_ ;
	assign \g7782/_0_  = _w21879_ ;
	assign \g7784/_0_  = _w21882_ ;
	assign \g78/_0_  = _w21888_ ;
	assign \g7800/_0_  = _w21889_ ;
	assign \g7823/_3_  = _w21891_ ;
	assign \g7837/_0_  = _w21894_ ;
	assign \g7841/_0_  = _w21897_ ;
	assign \g7842/_0_  = _w21900_ ;
	assign \g7843/_0_  = _w21903_ ;
	assign \g7844/_0_  = _w21905_ ;
	assign \g7845/_0_  = _w21908_ ;
	assign \g7846/_0_  = _w21911_ ;
	assign \g7847/_0_  = _w21914_ ;
	assign \g7849/_0_  = _w21915_ ;
	assign \g7850/_0_  = _w21917_ ;
	assign \g7852/_0_  = _w21918_ ;
	assign \g7854/_0_  = _w21919_ ;
	assign \g7855/_0_  = _w21922_ ;
	assign \g7857/_0_  = _w21924_ ;
	assign \g7858/_0_  = _w21926_ ;
	assign \g7859/_0_  = _w21928_ ;
	assign \g7860/_0_  = _w21930_ ;
	assign \g7861/_0_  = _w21932_ ;
	assign \g7862/_0_  = _w21934_ ;
	assign \g7863/_0_  = _w21936_ ;
	assign \g7864/_0_  = _w21938_ ;
	assign \g7865/_0_  = _w21940_ ;
	assign \g7866/_0_  = _w21942_ ;
	assign \g7867/_0_  = _w21944_ ;
	assign \g7868/_0_  = _w21946_ ;
	assign \g7869/_0_  = _w21948_ ;
	assign \g7870/_0_  = _w21950_ ;
	assign \g7871/_0_  = _w21954_ ;
	assign \g79211/_3_  = _w21955_ ;
	assign \g79258/_3_  = _w21956_ ;
	assign \g79299/_3_  = _w21957_ ;
	assign \g79316/_2_  = _w9311_ ;
	assign \g79342/_3_  = _w21958_ ;
	assign \g79401/_3_  = _w21959_ ;
	assign \g79452/_3_  = _w21960_ ;
	assign \g79457/_3_  = _w21961_ ;
	assign \g7951/_0_  = _w21962_ ;
	assign \g79541/_3_  = _w21963_ ;
	assign \g7958/_0_  = _w21964_ ;
	assign \g79598/_3_  = _w21965_ ;
	assign \g79654/_3_  = _w21966_ ;
	assign \g79675/_3_  = _w21967_ ;
	assign \g7971/_0_  = _w21968_ ;
	assign \g7972/_0_  = _w21977_ ;
	assign \g7973/_3_  = _w21989_ ;
	assign \g79753/_3_  = _w21990_ ;
	assign \g7976/_3_  = _w22002_ ;
	assign \g79855/_3_  = _w22003_ ;
	assign \g79858/_3_  = _w22004_ ;
	assign \g79997/_3_  = _w22005_ ;
	assign \g8/_0_  = _w22012_ ;
	assign \g80008/_3_  = _w8043_ ;
	assign \g80011/_0_  = _w22013_ ;
	assign \g80104/_0_  = _w12553_ ;
	assign \g80172/_1_  = _w8601_ ;
	assign \g80195/_3_  = _w6501_ ;
	assign \g80238/_3_  = _w22014_ ;
	assign \g80290/_2_  = _w5760_ ;
	assign \g80294/_0_  = _w7710_ ;
	assign \g80302/_0_  = _w7906_ ;
	assign \g80327/_0_  = _w22018_ ;
	assign \g80360/_3_  = _w7241_ ;
	assign \g80373/_0_  = _w22025_ ;
	assign \g80401/_0_  = _w5914_ ;
	assign \g80410/_0_  = _w6363_ ;
	assign \g80475/_0_  = _w6039_ ;
	assign \g80476/_0_  = _w7566_ ;
	assign \g80516/_3_  = _w22029_ ;
	assign \g80536/_0_  = _w22030_ ;
	assign \g80537/_0_  = _w6758_ ;
	assign \g80572/_0_  = _w22017_ ;
	assign \g80573/_0_  = _w22016_ ;
	assign \g80609/_2_  = _w8761_ ;
	assign \g80610/_2_  = _w8802_ ;
	assign \g80676/_0_  = _w14270_ ;
	assign \g80798/_0_  = _w22031_ ;
	assign \g80807/_0_  = _w16029_ ;
	assign \g80890/_2_  = _w4806_ ;
	assign \g80904/_0_  = _w16030_ ;
	assign \g81719/_2_  = _w12543_ ;
	assign \g81746/_0_  = _w4788_ ;
	assign \g81775/_0_  = _w4852_ ;
	assign \g81872/_0_  = _w22038_ ;
	assign \g81961/_0_  = _w4144_ ;
	assign \g81968/_0_  = _w4154_ ;
	assign \g82096/_0_  = _w4143_ ;
	assign \g82123/_0_  = _w4105_ ;
	assign \g82147/_0_  = _w4141_ ;
	assign \g82147/_1_  = _w4140_ ;
	assign \g82335/_0_  = _w4782_ ;
	assign \g82338/_2_  = _w4797_ ;
	assign \g82368/_0_  = _w4086_ ;
	assign \g82460/_2_  = _w14260_ ;
	assign \g82469/_0_  = _w12055_ ;
	assign \g82481/_0_  = _w4085_ ;
	assign \g82625/_1_  = _w8491_ ;
	assign \g82711/_0_  = _w4856_ ;
	assign \g82772/_0_  = _w4103_ ;
	assign \g82946/_0_  = _w14258_ ;
	assign \g82947/_0_  = _w12541_ ;
	assign \g82956/_0_  = _w4874_ ;
	assign \g83003/_0_  = _w4098_ ;
	assign \g83006/_1_  = _w8490_ ;
	assign \g83415/_0_  = _w4866_ ;
	assign \g83498/_0_  = _w4101_ ;
	assign \g837/_0_  = _w22041_ ;
	assign \g838/_0_  = _w22042_ ;
	assign \g83863/_0_  = _w8489_ ;
	assign \g839/_0_  = _w22048_ ;
	assign \g84049/_3_  = _w22049_ ;
	assign \g84050/_3_  = _w22050_ ;
	assign \g84077/_2_  = _w4858_ ;
	assign \g842/_0_  = _w22053_ ;
	assign \g84245/_0_  = _w4074_ ;
	assign \g843/_0_  = _w22056_ ;
	assign \g844/_0_  = _w22057_ ;
	assign \g84448/_0_  = _w5575_ ;
	assign \g84478/_3_  = _w22035_ ;
	assign \g845/_0_  = _w22060_ ;
	assign \g846/_0_  = _w22063_ ;
	assign \g847/_0_  = _w22066_ ;
	assign \g848/_0_  = _w22069_ ;
	assign \g8487/_0_  = _w22073_ ;
	assign \g8488/_0_  = _w22077_ ;
	assign \g8489/_0_  = _w22081_ ;
	assign \g849/_0_  = _w22082_ ;
	assign \g8490/_0_  = _w22086_ ;
	assign \g84904/_0_  = _w22087_ ;
	assign \g8491/_0_  = _w22090_ ;
	assign \g8492/_0_  = _w22094_ ;
	assign \g8493/_0_  = _w22097_ ;
	assign \g8494/_0_  = _w22101_ ;
	assign \g8496/_0_  = _w22102_ ;
	assign \g8517/_0_  = _w22104_ ;
	assign \g8534/_0_  = _w22106_ ;
	assign \g8538/_0_  = _w22113_ ;
	assign \g8540/_0_  = _w22115_ ;
	assign \g8576/_2_  = _w19740_ ;
	assign \g8597/_0_  = _w22118_ ;
	assign \g8598/_0_  = _w22123_ ;
	assign \g8599/_0_  = _w22126_ ;
	assign \g8600/_0_  = _w22130_ ;
	assign \g8601/_0_  = _w22133_ ;
	assign \g8602/_0_  = _w22136_ ;
	assign \g8603/_0_  = _w22140_ ;
	assign \g8605/_0_  = _w22143_ ;
	assign \g8606/_0_  = _w22146_ ;
	assign \g8607/_0_  = _w22148_ ;
	assign \g8608/_0_  = _w22153_ ;
	assign \g8609/_0_  = _w22157_ ;
	assign \g8610/_0_  = _w22161_ ;
	assign \g8611/_0_  = _w22165_ ;
	assign \g8612/_0_  = _w22169_ ;
	assign \g8613/_0_  = _w22173_ ;
	assign \g8614/_0_  = _w22177_ ;
	assign \g8615/_0_  = _w22181_ ;
	assign \g8617/_0_  = _w22183_ ;
	assign \g8643/_0_  = _w22186_ ;
	assign \g8644/_0_  = _w22189_ ;
	assign \g8645/_0_  = _w22193_ ;
	assign \g8646/_0_  = _w22196_ ;
	assign \g8647/_0_  = _w22199_ ;
	assign \g8648/_0_  = _w22203_ ;
	assign \g8650/_0_  = _w22206_ ;
	assign \g8651/_0_  = _w22209_ ;
	assign \g8652/_0_  = _w22211_ ;
	assign \g8653/_0_  = _w22215_ ;
	assign \g8654/_0_  = _w22219_ ;
	assign \g8655/_0_  = _w22223_ ;
	assign \g8656/_0_  = _w22227_ ;
	assign \g8657/_0_  = _w22231_ ;
	assign \g8658/_0_  = _w22235_ ;
	assign \g8659/_0_  = _w22239_ ;
	assign \g8660/_0_  = _w22243_ ;
	assign \g8665/_00_  = _w22248_ ;
	assign \g8666/_00_  = _w22252_ ;
	assign \g8667/_00_  = _w22256_ ;
	assign \g8668/_00_  = _w22259_ ;
	assign \g8669/_00_  = _w22263_ ;
	assign \g86715/_0_  = _w22264_ ;
	assign \g86745/_3_  = _w6897_ ;
	assign \g8691/_0_  = _w22265_ ;
	assign \g8700/_0_  = _w22269_ ;
	assign \g8701/_0_  = _w22272_ ;
	assign \g8702/_0_  = _w22275_ ;
	assign \g8703/_0_  = _w22278_ ;
	assign \g8704/_0_  = _w22281_ ;
	assign \g8705/_0_  = _w22284_ ;
	assign \g87063/_0_  = _w22298_ ;
	assign \g87114/_0_  = _w22312_ ;
	assign \g8712/_0_  = _w22314_ ;
	assign \g8713/_0_  = _w22316_ ;
	assign \g8714/_0_  = _w22320_ ;
	assign \g87171/_1_  = _w22324_ ;
	assign \g87252/_1_  = _w4089_ ;
	assign \g87298/_0_  = _w22325_ ;
	assign \g8730/_0_  = _w22327_ ;
	assign \g8741/_0_  = _w22331_ ;
	assign \g8747/_0_  = _w22332_ ;
	assign \g87480/_0_  = _w22333_ ;
	assign \g87484/_2_  = _w14460_ ;
	assign \g87488/_1__syn_2  = _w16259_ ;
	assign \g8761/_0_  = _w22338_ ;
	assign \g8762/_0_  = _w22340_ ;
	assign \g8763/_0_  = _w22345_ ;
	assign \g8764/_0_  = _w22347_ ;
	assign \g8765/_0_  = _w22349_ ;
	assign \g8775/_0_  = _w22360_ ;
	assign \g8776/_0_  = _w22364_ ;
	assign \g8777/_0_  = _w22366_ ;
	assign \g8778/_0_  = _w22367_ ;
	assign \g8784/_0_  = _w22371_ ;
	assign \g8804/_0_  = _w22376_ ;
	assign \g8807/_0_  = _w22378_ ;
	assign \g8808/_0_  = _w22380_ ;
	assign \g8809/_0_  = _w22383_ ;
	assign \g8810/_0_  = _w22385_ ;
	assign \g8811/_0_  = _w22388_ ;
	assign \g8812/_0_  = _w22390_ ;
	assign \g8813/_0_  = _w22391_ ;
	assign \g8814/_0_  = _w22393_ ;
	assign \g8815/_0_  = _w22395_ ;
	assign \g8816/_0_  = _w22397_ ;
	assign \g8817/_0_  = _w22399_ ;
	assign \g8818/_0_  = _w22404_ ;
	assign \g8819/_0_  = _w22408_ ;
	assign \g8820/_0_  = _w22412_ ;
	assign \g8821/_0_  = _w22415_ ;
	assign \g8822/_0_  = _w22417_ ;
	assign \g8823/_0_  = _w22418_ ;
	assign \g8824/_0_  = _w22420_ ;
	assign \g8825/_0_  = _w22421_ ;
	assign \g8826/_0_  = _w22423_ ;
	assign \g8827/_0_  = _w22424_ ;
	assign \g8828/_0_  = _w22425_ ;
	assign \g8829/_0_  = _w22426_ ;
	assign \g8830/_0_  = _w22428_ ;
	assign \g8831/_0_  = _w22430_ ;
	assign \g8832/_0_  = _w22432_ ;
	assign \g8833/_0_  = _w22434_ ;
	assign \g8834/_0_  = _w22437_ ;
	assign \g8835/_0_  = _w22439_ ;
	assign \g8836/_0_  = _w22442_ ;
	assign \g8837/_0_  = _w22444_ ;
	assign \g8838/_0_  = _w22445_ ;
	assign \g8839/_0_  = _w22446_ ;
	assign \g8840/_0_  = _w22448_ ;
	assign \g8842/_0_  = _w22450_ ;
	assign \g8843/_0_  = _w22453_ ;
	assign \g8846/_0_  = _w22455_ ;
	assign \g8848/_0_  = _w22459_ ;
	assign \g8857/_0_  = _w22460_ ;
	assign \g8895/_0_  = _w22462_ ;
	assign \g8902/_3_  = _w22479_ ;
	assign \g8903/_3_  = _w22496_ ;
	assign \g8904/_3_  = _w22513_ ;
	assign \g8905/_3_  = _w22530_ ;
	assign \g8906/_3_  = _w22547_ ;
	assign \g8909/_0_  = _w22549_ ;
	assign \g8910/_0_  = _w22550_ ;
	assign \g8911/_0_  = _w22552_ ;
	assign \g8924/_3_  = _w22565_ ;
	assign \g8926/_3_  = _w22578_ ;
	assign \g8927/_3_  = _w22591_ ;
	assign \g8943/_0_  = _w22592_ ;
	assign \g8944/_0_  = _w22593_ ;
	assign \g8958/_3_  = _w22606_ ;
	assign \g8960/_00_  = _w22610_ ;
	assign \g8961/_3_  = _w22623_ ;
	assign \g8965/_0_  = _w22631_ ;
	assign \g8966/_0_  = _w22639_ ;
	assign \g8967/_0_  = _w22647_ ;
	assign \g8968/_0_  = _w22655_ ;
	assign \g9/_0_  = _w22662_ ;
	assign \g9123/_0_  = _w19738_ ;
	assign \g9125/_0_  = _w22663_ ;
	assign \g9126/_0_  = _w22664_ ;
	assign \g913/_0_  = _w22675_ ;
	assign \g915/_0_  = _w22678_ ;
	assign \g916/_0_  = _w22681_ ;
	assign \g917/_0_  = _w22684_ ;
	assign \g918/_0_  = _w22687_ ;
	assign \g919/_0_  = _w22690_ ;
	assign \g920/_3_  = _w22695_ ;
	assign \g921/_3_  = _w22699_ ;
	assign \g925/_0_  = _w22707_ ;
	assign \g926/_0_  = _w22710_ ;
	assign \g927/_0_  = _w22713_ ;
	assign \g928/_0_  = _w22716_ ;
	assign \g929/_0_  = _w22717_ ;
	assign \g930/_0_  = _w22718_ ;
	assign \g9336/_0_  = _w22719_ ;
	assign \g9337/_0_  = _w22721_ ;
	assign \g939/_3_  = _w22725_ ;
	assign \g9396/_0_  = _w22728_ ;
	assign \g9397/_0_  = _w22729_ ;
	assign \g9399/_0_  = _w22730_ ;
	assign \g9400/_0_  = _w22731_ ;
	assign \g9401/_0_  = _w22732_ ;
	assign \g9402/_0_  = _w22733_ ;
	assign \g9403/_0_  = _w22734_ ;
	assign \g9404/_0_  = _w22735_ ;
	assign \g9415/_0_  = _w20081_ ;
	assign \g9418/_0_  = _w20111_ ;
	assign \g9419/_0_  = _w22740_ ;
	assign \g9420/_0_  = _w22742_ ;
	assign \g9446/_0_  = _w22743_ ;
	assign \g9465/_0_  = _w22744_ ;
	assign \g9493/_0_  = _w22745_ ;
	assign \g9536/_0_  = _w22747_ ;
	assign \g9537/_0_  = _w22752_ ;
	assign \g9538/_0_  = _w22754_ ;
	assign \g9539/_0_  = _w22756_ ;
	assign \g9540/_0_  = _w22758_ ;
	assign \g9541/_0_  = _w22760_ ;
	assign \g9542/_0_  = _w22763_ ;
	assign \g955/_2_  = _w22769_ ;
	assign \g9561/_0_  = _w22774_ ;
	assign \g9562/_0_  = _w22778_ ;
	assign \g9563/_0_  = _w22782_ ;
	assign \g9564/_0_  = _w22786_ ;
	assign \g9565/_0_  = _w22790_ ;
	assign \g9566/_0_  = _w22795_ ;
	assign \g9567/_0_  = _w22800_ ;
	assign \g9568/_0_  = _w22803_ ;
	assign \g9569/_0_  = _w22809_ ;
	assign \g9570/_0_  = _w22814_ ;
	assign \g9571/_0_  = _w22815_ ;
	assign \g9572/_0_  = _w22819_ ;
	assign \g9573/_0_  = _w22820_ ;
	assign \g9574/_0_  = _w22824_ ;
	assign \g9575/_0_  = _w22825_ ;
	assign \g9576/_0_  = _w22828_ ;
	assign \g9577/_0_  = _w22831_ ;
	assign \g9578/_0_  = _w22834_ ;
	assign \g9579/_0_  = _w22837_ ;
	assign \g9580/_0_  = _w22838_ ;
	assign \g9581/_0_  = _w22842_ ;
	assign \g9582/_0_  = _w22845_ ;
	assign \g9583/_0_  = _w22846_ ;
	assign \g9584/_0_  = _w22847_ ;
	assign \g9585/_0_  = _w22848_ ;
	assign \g9586/_0_  = _w22849_ ;
	assign \g9587/_0_  = _w22850_ ;
	assign \g9588/_0_  = _w22851_ ;
	assign \g9589/_0_  = _w22852_ ;
	assign \g9590/_0_  = _w22853_ ;
	assign \g9591/_0_  = _w22854_ ;
	assign \g9592/_0_  = _w22857_ ;
	assign \g9593/_0_  = _w22860_ ;
	assign \g9594/_0_  = _w22861_ ;
	assign \g9595/_0_  = _w22865_ ;
	assign \g9596/_0_  = _w22868_ ;
	assign \g9597/_0_  = _w22869_ ;
	assign \g9598/_0_  = _w22870_ ;
	assign \g9599/_0_  = _w22871_ ;
	assign \g9600/_0_  = _w22872_ ;
	assign \g9601/_0_  = _w22873_ ;
	assign \g9602/_0_  = _w22874_ ;
	assign \g9603/_0_  = _w22875_ ;
	assign \g9604/_0_  = _w22876_ ;
	assign \g9605/_0_  = _w22877_ ;
	assign \g9606/_0_  = _w22880_ ;
	assign \g9607/_0_  = _w22883_ ;
	assign \g9608/_0_  = _w22884_ ;
	assign \g9609/_0_  = _w22888_ ;
	assign \g9610/_0_  = _w22891_ ;
	assign \g9611/_0_  = _w22892_ ;
	assign \g9612/_0_  = _w22893_ ;
	assign \g9613/_0_  = _w22894_ ;
	assign \g9614/_0_  = _w22895_ ;
	assign \g9615/_0_  = _w22896_ ;
	assign \g9616/_0_  = _w22897_ ;
	assign \g9617/_0_  = _w22898_ ;
	assign \g9618/_0_  = _w22899_ ;
	assign \g9619/_0_  = _w22900_ ;
	assign \g9620/_0_  = _w22903_ ;
	assign \g9621/_0_  = _w22906_ ;
	assign \g9622/_0_  = _w22907_ ;
	assign \g9623/_0_  = _w22911_ ;
	assign \g9624/_0_  = _w22914_ ;
	assign \g9625/_0_  = _w22915_ ;
	assign \g9626/_0_  = _w22916_ ;
	assign \g9627/_0_  = _w22917_ ;
	assign \g9628/_0_  = _w22918_ ;
	assign \g9629/_0_  = _w22919_ ;
	assign \g9630/_0_  = _w22920_ ;
	assign \g9631/_0_  = _w22921_ ;
	assign \g9632/_0_  = _w22922_ ;
	assign \g9633/_0_  = _w22923_ ;
	assign \g9634/_0_  = _w22926_ ;
	assign \g9635/_0_  = _w22929_ ;
	assign \g9636/_0_  = _w22930_ ;
	assign \g9637/_0_  = _w22934_ ;
	assign \g9638/_0_  = _w22937_ ;
	assign \g9639/_0_  = _w22938_ ;
	assign \g9640/_0_  = _w22939_ ;
	assign \g9641/_0_  = _w22940_ ;
	assign \g9642/_0_  = _w22941_ ;
	assign \g9643/_0_  = _w22942_ ;
	assign \g9644/_0_  = _w22943_ ;
	assign \g9645/_0_  = _w22944_ ;
	assign \g9646/_0_  = _w22945_ ;
	assign \g9647/_0_  = _w22946_ ;
	assign \g9648/_0_  = _w22949_ ;
	assign \g9649/_0_  = _w22952_ ;
	assign \g9650/_0_  = _w22953_ ;
	assign \g9651/_0_  = _w22957_ ;
	assign \g9652/_0_  = _w22960_ ;
	assign \g9653/_0_  = _w22961_ ;
	assign \g9654/_0_  = _w22962_ ;
	assign \g9655/_0_  = _w22963_ ;
	assign \g9656/_0_  = _w22964_ ;
	assign \g9657/_0_  = _w22965_ ;
	assign \g9658/_0_  = _w22966_ ;
	assign \g9659/_0_  = _w22967_ ;
	assign \g9660/_0_  = _w22968_ ;
	assign \g9661/_0_  = _w22969_ ;
	assign \g9662/_0_  = _w22972_ ;
	assign \g9663/_0_  = _w22975_ ;
	assign \g9664/_0_  = _w22976_ ;
	assign \g9665/_0_  = _w22980_ ;
	assign \g9666/_0_  = _w22983_ ;
	assign \g9667/_0_  = _w22984_ ;
	assign \g9668/_0_  = _w22985_ ;
	assign \g9669/_0_  = _w22986_ ;
	assign \g9670/_0_  = _w22987_ ;
	assign \g9671/_0_  = _w22988_ ;
	assign \g9672/_0_  = _w22989_ ;
	assign \g9673/_0_  = _w22990_ ;
	assign \g9674/_0_  = _w22991_ ;
	assign \g9675/_0_  = _w22992_ ;
	assign \g9676/_0_  = _w22995_ ;
	assign \g9677/_0_  = _w22998_ ;
	assign \g9678/_0_  = _w22999_ ;
	assign \g9681/_0_  = _w23004_ ;
	assign \g9683/_0_  = _w23005_ ;
	assign \g9689/_0_  = _w23008_ ;
	assign \g9692/_0_  = _w23009_ ;
	assign \g9694/_0_  = _w23013_ ;
	assign \g9695/_0_  = _w23017_ ;
	assign \g9701/_0_  = _w23018_ ;
	assign \g9702/_0_  = _w23022_ ;
	assign \g9703/_0_  = _w23026_ ;
	assign \g9704/_0_  = _w23029_ ;
	assign \g9709/_0_  = _w23031_ ;
	assign \g9710/_0_  = _w23032_ ;
	assign \g9711/_0_  = _w23033_ ;
	assign \g9712/_0_  = _w23034_ ;
	assign \g9720/_0_  = _w23035_ ;
	assign \g9721/_0_  = _w23036_ ;
	assign \g9722/_0_  = _w23037_ ;
	assign \g9726/_0_  = _w23038_ ;
	assign \g9733/_0_  = _w23042_ ;
	assign \g9734/_0_  = _w23045_ ;
	assign \g9735/_0_  = _w23046_ ;
	assign \g9736/_0_  = _w23047_ ;
	assign \g9737/_0_  = _w23048_ ;
	assign \g9738/_0_  = _w23049_ ;
	assign \g9739/_0_  = _w23050_ ;
	assign \g9740/_0_  = _w23051_ ;
	assign \g9741/_0_  = _w23052_ ;
	assign \g9742/_0_  = _w23053_ ;
	assign \g9743/_0_  = _w23054_ ;
	assign \g9744/_0_  = _w23057_ ;
	assign \g9745/_0_  = _w23060_ ;
	assign \g9746/_0_  = _w23061_ ;
	assign \g9747/_0_  = _w23065_ ;
	assign \g9748/_0_  = _w23068_ ;
	assign \g9749/_0_  = _w23069_ ;
	assign \g9750/_0_  = _w23070_ ;
	assign \g9751/_0_  = _w23071_ ;
	assign \g9752/_0_  = _w23072_ ;
	assign \g9753/_0_  = _w23073_ ;
	assign \g9754/_0_  = _w23074_ ;
	assign \g9755/_0_  = _w23075_ ;
	assign \g9756/_0_  = _w23076_ ;
	assign \g9757/_0_  = _w23077_ ;
	assign \g9758/_0_  = _w23080_ ;
	assign \g9759/_0_  = _w23083_ ;
	assign \g9760/_0_  = _w23084_ ;
	assign \g9761/_0_  = _w23088_ ;
	assign \g9762/_0_  = _w23091_ ;
	assign \g9763/_0_  = _w23092_ ;
	assign \g9764/_0_  = _w23093_ ;
	assign \g9765/_0_  = _w23094_ ;
	assign \g9766/_0_  = _w23095_ ;
	assign \g9767/_0_  = _w23096_ ;
	assign \g9768/_0_  = _w23097_ ;
	assign \g9769/_0_  = _w23098_ ;
	assign \g9770/_0_  = _w23099_ ;
	assign \g9771/_0_  = _w23100_ ;
	assign \g9772/_0_  = _w23103_ ;
	assign \g9773/_0_  = _w23106_ ;
	assign \g9774/_0_  = _w23107_ ;
	assign \g9775/_0_  = _w23111_ ;
	assign \g9776/_0_  = _w23114_ ;
	assign \g9777/_0_  = _w23115_ ;
	assign \g9778/_0_  = _w23116_ ;
	assign \g9779/_0_  = _w23117_ ;
	assign \g9780/_0_  = _w23118_ ;
	assign \g9781/_0_  = _w23119_ ;
	assign \g9782/_0_  = _w23120_ ;
	assign \g9783/_0_  = _w23121_ ;
	assign \g9784/_0_  = _w23122_ ;
	assign \g9785/_0_  = _w23123_ ;
	assign \g9786/_0_  = _w23126_ ;
	assign \g9787/_0_  = _w23129_ ;
	assign \g9788/_0_  = _w23130_ ;
	assign \g9789/_0_  = _w23134_ ;
	assign \g9790/_0_  = _w23137_ ;
	assign \g9791/_0_  = _w23138_ ;
	assign \g9792/_0_  = _w23139_ ;
	assign \g9793/_0_  = _w23140_ ;
	assign \g9794/_0_  = _w23141_ ;
	assign \g9795/_0_  = _w23142_ ;
	assign \g9796/_0_  = _w23143_ ;
	assign \g9797/_0_  = _w23144_ ;
	assign \g9798/_0_  = _w23145_ ;
	assign \g9799/_0_  = _w23146_ ;
	assign \g9800/_0_  = _w23149_ ;
	assign \g9801/_0_  = _w23150_ ;
	assign \g9802/_0_  = _w23153_ ;
	assign \g9803/_0_  = _w23157_ ;
	assign \g9804/_0_  = _w23160_ ;
	assign \g9805/_0_  = _w23161_ ;
	assign \g9806/_0_  = _w23162_ ;
	assign \g9807/_0_  = _w23163_ ;
	assign \g9808/_0_  = _w23164_ ;
	assign \g9809/_0_  = _w23165_ ;
	assign \g9810/_0_  = _w23166_ ;
	assign \g9811/_0_  = _w23167_ ;
	assign \g9812/_0_  = _w23168_ ;
	assign \g9813/_0_  = _w23169_ ;
	assign \g9814/_0_  = _w23172_ ;
	assign \g9815/_0_  = _w23175_ ;
	assign \g9816/_0_  = _w23176_ ;
	assign \g9817/_0_  = _w23180_ ;
	assign \g9818/_0_  = _w23183_ ;
	assign \g9819/_0_  = _w23184_ ;
	assign \g9820/_0_  = _w23185_ ;
	assign \g9821/_0_  = _w23186_ ;
	assign \g9822/_0_  = _w23187_ ;
	assign \g9823/_0_  = _w23188_ ;
	assign \g9824/_0_  = _w23189_ ;
	assign \g9825/_0_  = _w23190_ ;
	assign \g9826/_0_  = _w23191_ ;
	assign \g9827/_0_  = _w23192_ ;
	assign \g9828/_0_  = _w23193_ ;
	assign \g9829/_0_  = _w23196_ ;
	assign \g9830/_0_  = _w23199_ ;
	assign \g9831/_0_  = _w23200_ ;
	assign \g9832/_0_  = _w23203_ ;
	assign \g9833/_0_  = _w23206_ ;
	assign \g9835/_0_  = _w23207_ ;
	assign \g9836/_0_  = _w23208_ ;
	assign \g9837/_0_  = _w23209_ ;
	assign \g9838/_0_  = _w23210_ ;
	assign \g9839/_0_  = _w23211_ ;
	assign \g9840/_0_  = _w23212_ ;
	assign \g9841/_0_  = _w23213_ ;
	assign \g9842/_0_  = _w23214_ ;
	assign \g9844/_0_  = _w23216_ ;
	assign \g9845/_0_  = _w23218_ ;
	assign \g9846/_0_  = _w23220_ ;
	assign \g9848/_0_  = _w23223_ ;
	assign \g9849/_0_  = _w23226_ ;
	assign \g9850/_0_  = _w23230_ ;
	assign \g9851/_0_  = _w23234_ ;
	assign \g9853/_0_  = _w23237_ ;
	assign \g9854/_0_  = _w23241_ ;
	assign \g9855/_0_  = _w23245_ ;
	assign \g9856/_0_  = _w23246_ ;
	assign \g9857/_0_  = _w23248_ ;
	assign \g9858/_0_  = _w23250_ ;
	assign \g9859/_0_  = _w23252_ ;
	assign \g9860/_0_  = _w23254_ ;
	assign \g9862/_0_  = _w23257_ ;
	assign \g9863/_0_  = _w23259_ ;
	assign \g9864/_0_  = _w23262_ ;
	assign \g9865/_0_  = _w23265_ ;
	assign \g9867/_0_  = _w23269_ ;
	assign \g9868/_0_  = _w23272_ ;
	assign \g9876/_0_  = _w23275_ ;
	assign \g9877/_0_  = _w23276_ ;
	assign \g9878/_0_  = _w23279_ ;
	assign \g9879/_0_  = _w23282_ ;
	assign \g9880/_0_  = _w23285_ ;
	assign \g9881/_0_  = _w23288_ ;
	assign \g9898/_0_  = _w23289_ ;
	assign \g9900/_0_  = _w23290_ ;
	assign \g9901/_0_  = _w23291_ ;
	assign \g9902/_0_  = _w23292_ ;
	assign \g9903/_0_  = _w23293_ ;
	assign \g9904/_0_  = _w23294_ ;
	assign \g9905/_0_  = _w23295_ ;
	assign \g9906/_0_  = _w23296_ ;
	assign \g9907/_0_  = _w23297_ ;
	assign \g9908/_0_  = _w23298_ ;
	assign \g9909/_0_  = _w23299_ ;
	assign \g9910/_0_  = _w23300_ ;
	assign \g9911/_0_  = _w23301_ ;
	assign \g9912/_0_  = _w23302_ ;
	assign \g9913/_0_  = _w23303_ ;
	assign \g9914/_0_  = _w23304_ ;
	assign \g9915/_0_  = _w23305_ ;
	assign \g9916/_0_  = _w23306_ ;
	assign \g9917/_0_  = _w23307_ ;
	assign \g9918/_0_  = _w23308_ ;
	assign \g9919/_0_  = _w23309_ ;
	assign \g992/_0_  = _w23317_ ;
	assign \g9920/_0_  = _w23318_ ;
	assign \g9921/_0_  = _w23319_ ;
	assign \g9922/_0_  = _w23320_ ;
	assign \g9923/_0_  = _w23321_ ;
	assign \g9924/_0_  = _w23322_ ;
	assign \g9925/_0_  = _w23323_ ;
	assign \g9926/_0_  = _w23324_ ;
	assign \g9927/_0_  = _w23325_ ;
	assign \g9928/_0_  = _w23326_ ;
	assign \g9929/_0_  = _w23327_ ;
	assign \g9930/_0_  = _w23328_ ;
	assign \g9931/_0_  = _w23329_ ;
	assign \g9932/_0_  = _w23330_ ;
	assign \g9933/_0_  = _w23331_ ;
	assign \g9934/_0_  = _w23332_ ;
	assign \g9935/_0_  = _w23333_ ;
	assign \g9936/_0_  = _w23334_ ;
	assign \g9937/_0_  = _w23335_ ;
	assign \g9938/_0_  = _w23336_ ;
	assign \g9939/_0_  = _w23337_ ;
	assign \g9940/_0_  = _w23338_ ;
	assign \g9941/_0_  = _w23339_ ;
	assign \g9942/_0_  = _w23340_ ;
	assign \g9943/_0_  = _w23341_ ;
	assign \g9944/_0_  = _w23342_ ;
	assign \g9945/_0_  = _w23343_ ;
	assign \g9946/_0_  = _w23344_ ;
	assign \g9947/_0_  = _w23345_ ;
	assign \g9948/_0_  = _w23346_ ;
	assign \g9949/_0_  = _w23349_ ;
	assign \g9950/_0_  = _w23352_ ;
	assign \g9951/_0_  = _w23355_ ;
	assign \g9952/_0_  = _w23358_ ;
	assign \g9953/_0_  = _w23361_ ;
	assign \g9954/_0_  = _w23364_ ;
	assign \g9955/_0_  = _w23367_ ;
	assign \g9956/_0_  = _w23370_ ;
	assign \g9957/_0_  = _w23373_ ;
	assign \g9958/_0_  = _w23376_ ;
	assign \g9959/_0_  = _w23379_ ;
	assign \g9960/_0_  = _w23382_ ;
	assign \g9961/_0_  = _w23385_ ;
	assign \g9962/_0_  = _w23388_ ;
	assign \g9963/_0_  = _w23391_ ;
	assign \g9964/_0_  = _w23394_ ;
	assign \g9965/_0_  = _w23397_ ;
	assign \g9966/_0_  = _w23400_ ;
	assign \g9967/_0_  = _w23403_ ;
	assign \g9968/_0_  = _w23406_ ;
	assign \g9969/_0_  = _w23409_ ;
	assign \g9970/_0_  = _w23412_ ;
	assign \g9971/_0_  = _w23415_ ;
	assign \g9972/_0_  = _w23418_ ;
	assign \g9973/_0_  = _w23421_ ;
	assign \g9974/_0_  = _w23422_ ;
	assign \g9975/_0_  = _w23423_ ;
	assign \g9976/_0_  = _w23424_ ;
	assign \g9977/_0_  = _w23425_ ;
	assign \g9978/_0_  = _w23426_ ;
	assign \g9979/_0_  = _w23427_ ;
	assign \g9980/_0_  = _w23428_ ;
	assign \g9981/_0_  = _w23429_ ;
	assign \g9982/_0_  = _w23430_ ;
	assign \g9983/_0_  = _w23431_ ;
	assign \g9984/_0_  = _w23432_ ;
	assign \g9985/_0_  = _w23433_ ;
	assign \g9987/_0_  = _w23434_ ;
	assign \g9988/_0_  = _w23435_ ;
	assign \g9989/_0_  = _w23436_ ;
	assign \g999/_0_  = _w23437_ ;
	assign \g9990/_0_  = _w23438_ ;
	assign \g9991/_0_  = _w23439_ ;
	assign \g9992/_0_  = _w23442_ ;
	assign \g9993/_0_  = _w23443_ ;
	assign \g9994/_0_  = _w23444_ ;
	assign \g9995/_0_  = _w23445_ ;
	assign \g9996/_0_  = _w23446_ ;
	assign \g9997/_0_  = _w23447_ ;
	assign \g9998/_0_  = _w23448_ ;
	assign \g9999/_0_  = _w23449_ ;
	assign \idma_IDMA_boot_reg/NET0131_reg_syn_3  = _w23450_ ;
	assign \memc_EXTC_Eg_reg/NET0131  = _w4070_ ;
	assign \memc_EXTC_Eg_reg/NET0131_reg_syn_3  = _w23452_ ;
	assign \memc_EXTC_Eg_reg/n0  = _w23451_ ;
	assign \pio_PIO_IN_P_reg[0]/P0001_reg_syn_3  = _w23455_ ;
	assign \pio_PIO_IN_P_reg[10]/P0001_reg_syn_3  = _w23458_ ;
	assign \pio_PIO_IN_P_reg[11]/P0001_reg_syn_3  = _w23461_ ;
	assign \pio_PIO_IN_P_reg[1]/P0001_reg_syn_3  = _w23464_ ;
	assign \pio_PIO_IN_P_reg[2]/P0001_reg_syn_3  = _w23467_ ;
	assign \pio_PIO_IN_P_reg[3]/P0001_reg_syn_3  = _w23470_ ;
	assign \pio_PIO_IN_P_reg[4]/P0001_reg_syn_3  = _w23473_ ;
	assign \pio_PIO_IN_P_reg[5]/P0001_reg_syn_3  = _w23476_ ;
	assign \pio_PIO_IN_P_reg[6]/P0001_reg_syn_3  = _w23479_ ;
	assign \pio_PIO_IN_P_reg[7]/P0001_reg_syn_3  = _w23482_ ;
	assign \pio_PIO_IN_P_reg[8]/P0001_reg_syn_3  = _w23485_ ;
	assign \pio_PIO_IN_P_reg[9]/P0001_reg_syn_3  = _w23488_ ;
	assign \pio_PIO_RES_OUT_reg[0]/P0001_reg_syn_3  = _w23491_ ;
	assign \pio_PIO_RES_OUT_reg[10]/P0001_reg_syn_3  = _w23494_ ;
	assign \pio_PIO_RES_OUT_reg[2]/P0001_reg_syn_3  = _w23497_ ;
	assign \pio_PIO_RES_OUT_reg[4]/P0001_reg_syn_3  = _w23500_ ;
	assign \pio_PIO_RES_OUT_reg[6]/P0001_reg_syn_3  = _w23503_ ;
	assign \sice_GO_NXi_reg/NET0131_reg_syn_3  = _w23504_ ;
	assign \sport0_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  = _w23507_ ;
	assign \sport0_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  = _w23509_ ;
	assign \sport1_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  = _w23512_ ;
	assign \sport1_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  = _w23514_ ;
endmodule;