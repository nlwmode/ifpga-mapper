module top (\data_i[0]_pad , \data_i[10]_pad , \data_i[11]_pad , \data_i[12]_pad , \data_i[13]_pad , \data_i[14]_pad , \data_i[15]_pad , \data_i[16]_pad , \data_i[17]_pad , \data_i[18]_pad , \data_i[19]_pad , \data_i[1]_pad , \data_i[20]_pad , \data_i[21]_pad , \data_i[22]_pad , \data_i[23]_pad , \data_i[24]_pad , \data_i[25]_pad , \data_i[26]_pad , \data_i[27]_pad , \data_i[28]_pad , \data_i[29]_pad , \data_i[2]_pad , \data_i[30]_pad , \data_i[31]_pad , \data_i[32]_pad , \data_i[33]_pad , \data_i[34]_pad , \data_i[35]_pad , \data_i[36]_pad , \data_i[37]_pad , \data_i[38]_pad , \data_i[39]_pad , \data_i[3]_pad , \data_i[40]_pad , \data_i[41]_pad , \data_i[42]_pad , \data_i[43]_pad , \data_i[44]_pad , \data_i[45]_pad , \data_i[46]_pad , \data_i[47]_pad , \data_i[48]_pad , \data_i[49]_pad , \data_i[4]_pad , \data_i[50]_pad , \data_i[51]_pad , \data_i[52]_pad , \data_i[53]_pad , \data_i[54]_pad , \data_i[55]_pad , \data_i[56]_pad , \data_i[57]_pad , \data_i[58]_pad , \data_i[59]_pad , \data_i[5]_pad , \data_i[60]_pad , \data_i[61]_pad , \data_i[62]_pad , \data_i[63]_pad , \data_i[6]_pad , \data_i[7]_pad , \data_i[8]_pad , \data_i[9]_pad , \data_ready_reg/NET0131 , decrypt_i_pad, \key_i[10]_pad , \key_i[11]_pad , \key_i[12]_pad , \key_i[13]_pad , \key_i[14]_pad , \key_i[15]_pad , \key_i[17]_pad , \key_i[18]_pad , \key_i[19]_pad , \key_i[1]_pad , \key_i[20]_pad , \key_i[21]_pad , \key_i[22]_pad , \key_i[23]_pad , \key_i[25]_pad , \key_i[26]_pad , \key_i[27]_pad , \key_i[28]_pad , \key_i[29]_pad , \key_i[2]_pad , \key_i[30]_pad , \key_i[31]_pad , \key_i[33]_pad , \key_i[34]_pad , \key_i[35]_pad , \key_i[36]_pad , \key_i[37]_pad , \key_i[38]_pad , \key_i[39]_pad , \key_i[3]_pad , \key_i[41]_pad , \key_i[42]_pad , \key_i[43]_pad , \key_i[44]_pad , \key_i[45]_pad , \key_i[46]_pad , \key_i[47]_pad , \key_i[49]_pad , \key_i[4]_pad , \key_i[50]_pad , \key_i[51]_pad , \key_i[52]_pad , \key_i[53]_pad , \key_i[54]_pad , \key_i[55]_pad , \key_i[57]_pad , \key_i[58]_pad , \key_i[59]_pad , \key_i[5]_pad , \key_i[60]_pad , \key_i[61]_pad , \key_i[62]_pad , \key_i[63]_pad , \key_i[6]_pad , \key_i[7]_pad , \key_i[9]_pad , load_i_pad, \rd1_Key_o_reg[0]/NET0131 , \rd1_Key_o_reg[10]/NET0131 , \rd1_Key_o_reg[11]/NET0131 , \rd1_Key_o_reg[12]/NET0131 , \rd1_Key_o_reg[13]/NET0131 , \rd1_Key_o_reg[14]/NET0131 , \rd1_Key_o_reg[15]/NET0131 , \rd1_Key_o_reg[16]/NET0131 , \rd1_Key_o_reg[17]/NET0131 , \rd1_Key_o_reg[18]/NET0131 , \rd1_Key_o_reg[19]/NET0131 , \rd1_Key_o_reg[1]/NET0131 , \rd1_Key_o_reg[20]/NET0131 , \rd1_Key_o_reg[21]/NET0131 , \rd1_Key_o_reg[22]/NET0131 , \rd1_Key_o_reg[23]/NET0131 , \rd1_Key_o_reg[24]/NET0131 , \rd1_Key_o_reg[25]/NET0131 , \rd1_Key_o_reg[26]/NET0131 , \rd1_Key_o_reg[27]/NET0131 , \rd1_Key_o_reg[28]/NET0131 , \rd1_Key_o_reg[29]/NET0131 , \rd1_Key_o_reg[2]/NET0131 , \rd1_Key_o_reg[30]/NET0131 , \rd1_Key_o_reg[31]/NET0131 , \rd1_Key_o_reg[32]/NET0131 , \rd1_Key_o_reg[33]/NET0131 , \rd1_Key_o_reg[34]/NET0131 , \rd1_Key_o_reg[35]/NET0131 , \rd1_Key_o_reg[36]/NET0131 , \rd1_Key_o_reg[37]/NET0131 , \rd1_Key_o_reg[38]/NET0131 , \rd1_Key_o_reg[39]/NET0131 , \rd1_Key_o_reg[3]/NET0131 , \rd1_Key_o_reg[40]/NET0131 , \rd1_Key_o_reg[41]/NET0131 , \rd1_Key_o_reg[42]/NET0131 , \rd1_Key_o_reg[43]/NET0131 , \rd1_Key_o_reg[44]/NET0131 , \rd1_Key_o_reg[45]/NET0131 , \rd1_Key_o_reg[46]/NET0131 , \rd1_Key_o_reg[47]/NET0131 , \rd1_Key_o_reg[48]/NET0131 , \rd1_Key_o_reg[49]/NET0131 , \rd1_Key_o_reg[4]/NET0131 , \rd1_Key_o_reg[50]/NET0131 , \rd1_Key_o_reg[51]/NET0131 , \rd1_Key_o_reg[52]/NET0131 , \rd1_Key_o_reg[53]/NET0131 , \rd1_Key_o_reg[54]/NET0131 , \rd1_Key_o_reg[55]/NET0131 , \rd1_Key_o_reg[5]/NET0131 , \rd1_Key_o_reg[6]/NET0131 , \rd1_Key_o_reg[7]/NET0131 , \rd1_Key_o_reg[8]/NET0131 , \rd1_Key_o_reg[9]/NET0131 , \rd1_L_o_reg[0]/NET0131 , \rd1_L_o_reg[10]/NET0131 , \rd1_L_o_reg[11]/NET0131 , \rd1_L_o_reg[12]/NET0131 , \rd1_L_o_reg[13]/NET0131 , \rd1_L_o_reg[14]/NET0131 , \rd1_L_o_reg[15]/NET0131 , \rd1_L_o_reg[16]/NET0131 , \rd1_L_o_reg[17]/NET0131 , \rd1_L_o_reg[18]/NET0131 , \rd1_L_o_reg[19]/NET0131 , \rd1_L_o_reg[1]/NET0131 , \rd1_L_o_reg[20]/NET0131 , \rd1_L_o_reg[21]/NET0131 , \rd1_L_o_reg[22]/NET0131 , \rd1_L_o_reg[23]/NET0131 , \rd1_L_o_reg[24]/NET0131 , \rd1_L_o_reg[25]/NET0131 , \rd1_L_o_reg[26]/NET0131 , \rd1_L_o_reg[27]/NET0131 , \rd1_L_o_reg[28]/NET0131 , \rd1_L_o_reg[29]/NET0131 , \rd1_L_o_reg[2]/NET0131 , \rd1_L_o_reg[30]/NET0131 , \rd1_L_o_reg[31]/NET0131 , \rd1_L_o_reg[3]/NET0131 , \rd1_L_o_reg[4]/NET0131 , \rd1_L_o_reg[5]/NET0131 , \rd1_L_o_reg[6]/NET0131 , \rd1_L_o_reg[7]/NET0131 , \rd1_L_o_reg[8]/NET0131 , \rd1_L_o_reg[9]/NET0131 , \rd1_R_o_reg[0]/NET0131 , \rd1_R_o_reg[10]/NET0131 , \rd1_R_o_reg[11]/NET0131 , \rd1_R_o_reg[12]/NET0131 , \rd1_R_o_reg[13]/NET0131 , \rd1_R_o_reg[14]/NET0131 , \rd1_R_o_reg[15]/NET0131 , \rd1_R_o_reg[16]/NET0131 , \rd1_R_o_reg[17]/NET0131 , \rd1_R_o_reg[18]/NET0131 , \rd1_R_o_reg[19]/NET0131 , \rd1_R_o_reg[1]/NET0131 , \rd1_R_o_reg[20]/NET0131 , \rd1_R_o_reg[21]/NET0131 , \rd1_R_o_reg[22]/NET0131 , \rd1_R_o_reg[23]/NET0131 , \rd1_R_o_reg[24]/NET0131 , \rd1_R_o_reg[25]/NET0131 , \rd1_R_o_reg[26]/NET0131 , \rd1_R_o_reg[27]/NET0131 , \rd1_R_o_reg[28]/NET0131 , \rd1_R_o_reg[29]/NET0131 , \rd1_R_o_reg[2]/NET0131 , \rd1_R_o_reg[30]/NET0131 , \rd1_R_o_reg[31]/NET0131 , \rd1_R_o_reg[3]/NET0131 , \rd1_R_o_reg[4]/NET0131 , \rd1_R_o_reg[5]/NET0131 , \rd1_R_o_reg[6]/NET0131 , \rd1_R_o_reg[7]/NET0131 , \rd1_R_o_reg[8]/NET0131 , \rd1_R_o_reg[9]/NET0131 , \stage1_iter_reg[0]/NET0131 , \stage1_iter_reg[1]/NET0131 , \stage1_iter_reg[2]/NET0131 , \stage1_iter_reg[3]/NET0131 , \_al_n0 , \_al_n1 , \g10087/_0_ , \g10220/_1_ , \g11117/_0_ , \g11124/_0_ , \g11125/_0_ , \g11170/_0_ , \g11182/_0_ , \g11184/_0_ , \g11378/_0_ , \g11393/_0_ , \g11415/_0_ , \g11432/_0_ , \g11433/_0_ , \g11453/_0_ , \g11500/_0_ , \g11588/_0_ , \g11607/_0_ , \g11616/_0_ , \g11625/_0_ , \g11641_dup/_0_ , \g11648/_0_ , \g11655/_0_ , \g11683/_0_ , \g11689/_2_ , \g11694/_0_ , \g11748/_0_ , \g11880/_0_ , \g11962/_1_ , \g12016/_0_ , \g12038/_0_ , \g12039/_0_ , \g12094/_0_ , \g12100/_0_ , \g12132/_0_ , \g12151/_0_ , \g12251/_0_ , \g12279/_0_ , \g12288/_0_ , \g12290/_0_ , \g12311/_0_ , \g12313/_0_ , \g12356/_0_ , \g12357/_0_ , \g12427/_0_ , \g12441/_0_ , \g12442/_0_ , \g12480/_0_ , \g12485/_0_ , \g12506/_0_ , \g12544/_0_ , \g12549/_2_ , \g12614/_0_ , \g12678/_0_ , \g12680/_0_ , \g12748/_0_ , \g15/_0_ , \g25/_0_ , \g31/_0_ , \g6843/_0_ , \g6861/_0_ , \g6863/_0_ , \g6865/_0_ , \g6887/_0_ , \g6888/_0_ , \g6889/_0_ , \g6890/_0_ , \g6891/_0_ , \g6892/_0_ , \g6893/_0_ , \g6894/_0_ , \g6922/_0_ , \g6923/_0_ , \g6924/_3_ , \g6926/_0_ , \g6927/_0_ , \g6928/_0_ , \g6931/_0_ , \g6933/_0_ , \g6967/_0_ , \g6968/_0_ , \g6969/_0_ , \g6974/_0_ , \g6975/_0_ , \g6976/_3_ , \g7006/_3_ , \g8882/_0_ , \g8883/_0_ , \g8884/_0_ , \g8895/_0_ , \g8896/_0_ , \g8898/_0_ , \g8900/_2_ , \g8902/_0_ , \g8907/_0_ , \g8911/_0_ , \g8924/_0_ , \g8927/_0_ , \g8929/_2_ , \g8967/_0_ , \g8969/_0_ , \g8973/_2_ , \g8987/_0_ , \g8989/_0_ , \g8991/_0_ , \g8996/_0_ , \g9099/_0_ , \g9543/_1_ , \g9751/_1_ , \g9755/_0_ , \g9786/_0_ , \g9794/_0_ , \g9817/_0_ , \g9836/_0_ , \g9859/_0_ , \g9862/_0_ , \g9867/_0_ , \g9869/_0_ , \g9876/_0_ , \g9887/_0_ , \g9895/_0_ , \g9897/_0_ , \g9908/_0_ , \g9910/_0_ , \g9915/_0_ , \g9938/_0_ , \g9970/_0_ );
	input \data_i[0]_pad  ;
	input \data_i[10]_pad  ;
	input \data_i[11]_pad  ;
	input \data_i[12]_pad  ;
	input \data_i[13]_pad  ;
	input \data_i[14]_pad  ;
	input \data_i[15]_pad  ;
	input \data_i[16]_pad  ;
	input \data_i[17]_pad  ;
	input \data_i[18]_pad  ;
	input \data_i[19]_pad  ;
	input \data_i[1]_pad  ;
	input \data_i[20]_pad  ;
	input \data_i[21]_pad  ;
	input \data_i[22]_pad  ;
	input \data_i[23]_pad  ;
	input \data_i[24]_pad  ;
	input \data_i[25]_pad  ;
	input \data_i[26]_pad  ;
	input \data_i[27]_pad  ;
	input \data_i[28]_pad  ;
	input \data_i[29]_pad  ;
	input \data_i[2]_pad  ;
	input \data_i[30]_pad  ;
	input \data_i[31]_pad  ;
	input \data_i[32]_pad  ;
	input \data_i[33]_pad  ;
	input \data_i[34]_pad  ;
	input \data_i[35]_pad  ;
	input \data_i[36]_pad  ;
	input \data_i[37]_pad  ;
	input \data_i[38]_pad  ;
	input \data_i[39]_pad  ;
	input \data_i[3]_pad  ;
	input \data_i[40]_pad  ;
	input \data_i[41]_pad  ;
	input \data_i[42]_pad  ;
	input \data_i[43]_pad  ;
	input \data_i[44]_pad  ;
	input \data_i[45]_pad  ;
	input \data_i[46]_pad  ;
	input \data_i[47]_pad  ;
	input \data_i[48]_pad  ;
	input \data_i[49]_pad  ;
	input \data_i[4]_pad  ;
	input \data_i[50]_pad  ;
	input \data_i[51]_pad  ;
	input \data_i[52]_pad  ;
	input \data_i[53]_pad  ;
	input \data_i[54]_pad  ;
	input \data_i[55]_pad  ;
	input \data_i[56]_pad  ;
	input \data_i[57]_pad  ;
	input \data_i[58]_pad  ;
	input \data_i[59]_pad  ;
	input \data_i[5]_pad  ;
	input \data_i[60]_pad  ;
	input \data_i[61]_pad  ;
	input \data_i[62]_pad  ;
	input \data_i[63]_pad  ;
	input \data_i[6]_pad  ;
	input \data_i[7]_pad  ;
	input \data_i[8]_pad  ;
	input \data_i[9]_pad  ;
	input \data_ready_reg/NET0131  ;
	input decrypt_i_pad ;
	input \key_i[10]_pad  ;
	input \key_i[11]_pad  ;
	input \key_i[12]_pad  ;
	input \key_i[13]_pad  ;
	input \key_i[14]_pad  ;
	input \key_i[15]_pad  ;
	input \key_i[17]_pad  ;
	input \key_i[18]_pad  ;
	input \key_i[19]_pad  ;
	input \key_i[1]_pad  ;
	input \key_i[20]_pad  ;
	input \key_i[21]_pad  ;
	input \key_i[22]_pad  ;
	input \key_i[23]_pad  ;
	input \key_i[25]_pad  ;
	input \key_i[26]_pad  ;
	input \key_i[27]_pad  ;
	input \key_i[28]_pad  ;
	input \key_i[29]_pad  ;
	input \key_i[2]_pad  ;
	input \key_i[30]_pad  ;
	input \key_i[31]_pad  ;
	input \key_i[33]_pad  ;
	input \key_i[34]_pad  ;
	input \key_i[35]_pad  ;
	input \key_i[36]_pad  ;
	input \key_i[37]_pad  ;
	input \key_i[38]_pad  ;
	input \key_i[39]_pad  ;
	input \key_i[3]_pad  ;
	input \key_i[41]_pad  ;
	input \key_i[42]_pad  ;
	input \key_i[43]_pad  ;
	input \key_i[44]_pad  ;
	input \key_i[45]_pad  ;
	input \key_i[46]_pad  ;
	input \key_i[47]_pad  ;
	input \key_i[49]_pad  ;
	input \key_i[4]_pad  ;
	input \key_i[50]_pad  ;
	input \key_i[51]_pad  ;
	input \key_i[52]_pad  ;
	input \key_i[53]_pad  ;
	input \key_i[54]_pad  ;
	input \key_i[55]_pad  ;
	input \key_i[57]_pad  ;
	input \key_i[58]_pad  ;
	input \key_i[59]_pad  ;
	input \key_i[5]_pad  ;
	input \key_i[60]_pad  ;
	input \key_i[61]_pad  ;
	input \key_i[62]_pad  ;
	input \key_i[63]_pad  ;
	input \key_i[6]_pad  ;
	input \key_i[7]_pad  ;
	input \key_i[9]_pad  ;
	input load_i_pad ;
	input \rd1_Key_o_reg[0]/NET0131  ;
	input \rd1_Key_o_reg[10]/NET0131  ;
	input \rd1_Key_o_reg[11]/NET0131  ;
	input \rd1_Key_o_reg[12]/NET0131  ;
	input \rd1_Key_o_reg[13]/NET0131  ;
	input \rd1_Key_o_reg[14]/NET0131  ;
	input \rd1_Key_o_reg[15]/NET0131  ;
	input \rd1_Key_o_reg[16]/NET0131  ;
	input \rd1_Key_o_reg[17]/NET0131  ;
	input \rd1_Key_o_reg[18]/NET0131  ;
	input \rd1_Key_o_reg[19]/NET0131  ;
	input \rd1_Key_o_reg[1]/NET0131  ;
	input \rd1_Key_o_reg[20]/NET0131  ;
	input \rd1_Key_o_reg[21]/NET0131  ;
	input \rd1_Key_o_reg[22]/NET0131  ;
	input \rd1_Key_o_reg[23]/NET0131  ;
	input \rd1_Key_o_reg[24]/NET0131  ;
	input \rd1_Key_o_reg[25]/NET0131  ;
	input \rd1_Key_o_reg[26]/NET0131  ;
	input \rd1_Key_o_reg[27]/NET0131  ;
	input \rd1_Key_o_reg[28]/NET0131  ;
	input \rd1_Key_o_reg[29]/NET0131  ;
	input \rd1_Key_o_reg[2]/NET0131  ;
	input \rd1_Key_o_reg[30]/NET0131  ;
	input \rd1_Key_o_reg[31]/NET0131  ;
	input \rd1_Key_o_reg[32]/NET0131  ;
	input \rd1_Key_o_reg[33]/NET0131  ;
	input \rd1_Key_o_reg[34]/NET0131  ;
	input \rd1_Key_o_reg[35]/NET0131  ;
	input \rd1_Key_o_reg[36]/NET0131  ;
	input \rd1_Key_o_reg[37]/NET0131  ;
	input \rd1_Key_o_reg[38]/NET0131  ;
	input \rd1_Key_o_reg[39]/NET0131  ;
	input \rd1_Key_o_reg[3]/NET0131  ;
	input \rd1_Key_o_reg[40]/NET0131  ;
	input \rd1_Key_o_reg[41]/NET0131  ;
	input \rd1_Key_o_reg[42]/NET0131  ;
	input \rd1_Key_o_reg[43]/NET0131  ;
	input \rd1_Key_o_reg[44]/NET0131  ;
	input \rd1_Key_o_reg[45]/NET0131  ;
	input \rd1_Key_o_reg[46]/NET0131  ;
	input \rd1_Key_o_reg[47]/NET0131  ;
	input \rd1_Key_o_reg[48]/NET0131  ;
	input \rd1_Key_o_reg[49]/NET0131  ;
	input \rd1_Key_o_reg[4]/NET0131  ;
	input \rd1_Key_o_reg[50]/NET0131  ;
	input \rd1_Key_o_reg[51]/NET0131  ;
	input \rd1_Key_o_reg[52]/NET0131  ;
	input \rd1_Key_o_reg[53]/NET0131  ;
	input \rd1_Key_o_reg[54]/NET0131  ;
	input \rd1_Key_o_reg[55]/NET0131  ;
	input \rd1_Key_o_reg[5]/NET0131  ;
	input \rd1_Key_o_reg[6]/NET0131  ;
	input \rd1_Key_o_reg[7]/NET0131  ;
	input \rd1_Key_o_reg[8]/NET0131  ;
	input \rd1_Key_o_reg[9]/NET0131  ;
	input \rd1_L_o_reg[0]/NET0131  ;
	input \rd1_L_o_reg[10]/NET0131  ;
	input \rd1_L_o_reg[11]/NET0131  ;
	input \rd1_L_o_reg[12]/NET0131  ;
	input \rd1_L_o_reg[13]/NET0131  ;
	input \rd1_L_o_reg[14]/NET0131  ;
	input \rd1_L_o_reg[15]/NET0131  ;
	input \rd1_L_o_reg[16]/NET0131  ;
	input \rd1_L_o_reg[17]/NET0131  ;
	input \rd1_L_o_reg[18]/NET0131  ;
	input \rd1_L_o_reg[19]/NET0131  ;
	input \rd1_L_o_reg[1]/NET0131  ;
	input \rd1_L_o_reg[20]/NET0131  ;
	input \rd1_L_o_reg[21]/NET0131  ;
	input \rd1_L_o_reg[22]/NET0131  ;
	input \rd1_L_o_reg[23]/NET0131  ;
	input \rd1_L_o_reg[24]/NET0131  ;
	input \rd1_L_o_reg[25]/NET0131  ;
	input \rd1_L_o_reg[26]/NET0131  ;
	input \rd1_L_o_reg[27]/NET0131  ;
	input \rd1_L_o_reg[28]/NET0131  ;
	input \rd1_L_o_reg[29]/NET0131  ;
	input \rd1_L_o_reg[2]/NET0131  ;
	input \rd1_L_o_reg[30]/NET0131  ;
	input \rd1_L_o_reg[31]/NET0131  ;
	input \rd1_L_o_reg[3]/NET0131  ;
	input \rd1_L_o_reg[4]/NET0131  ;
	input \rd1_L_o_reg[5]/NET0131  ;
	input \rd1_L_o_reg[6]/NET0131  ;
	input \rd1_L_o_reg[7]/NET0131  ;
	input \rd1_L_o_reg[8]/NET0131  ;
	input \rd1_L_o_reg[9]/NET0131  ;
	input \rd1_R_o_reg[0]/NET0131  ;
	input \rd1_R_o_reg[10]/NET0131  ;
	input \rd1_R_o_reg[11]/NET0131  ;
	input \rd1_R_o_reg[12]/NET0131  ;
	input \rd1_R_o_reg[13]/NET0131  ;
	input \rd1_R_o_reg[14]/NET0131  ;
	input \rd1_R_o_reg[15]/NET0131  ;
	input \rd1_R_o_reg[16]/NET0131  ;
	input \rd1_R_o_reg[17]/NET0131  ;
	input \rd1_R_o_reg[18]/NET0131  ;
	input \rd1_R_o_reg[19]/NET0131  ;
	input \rd1_R_o_reg[1]/NET0131  ;
	input \rd1_R_o_reg[20]/NET0131  ;
	input \rd1_R_o_reg[21]/NET0131  ;
	input \rd1_R_o_reg[22]/NET0131  ;
	input \rd1_R_o_reg[23]/NET0131  ;
	input \rd1_R_o_reg[24]/NET0131  ;
	input \rd1_R_o_reg[25]/NET0131  ;
	input \rd1_R_o_reg[26]/NET0131  ;
	input \rd1_R_o_reg[27]/NET0131  ;
	input \rd1_R_o_reg[28]/NET0131  ;
	input \rd1_R_o_reg[29]/NET0131  ;
	input \rd1_R_o_reg[2]/NET0131  ;
	input \rd1_R_o_reg[30]/NET0131  ;
	input \rd1_R_o_reg[31]/NET0131  ;
	input \rd1_R_o_reg[3]/NET0131  ;
	input \rd1_R_o_reg[4]/NET0131  ;
	input \rd1_R_o_reg[5]/NET0131  ;
	input \rd1_R_o_reg[6]/NET0131  ;
	input \rd1_R_o_reg[7]/NET0131  ;
	input \rd1_R_o_reg[8]/NET0131  ;
	input \rd1_R_o_reg[9]/NET0131  ;
	input \stage1_iter_reg[0]/NET0131  ;
	input \stage1_iter_reg[1]/NET0131  ;
	input \stage1_iter_reg[2]/NET0131  ;
	input \stage1_iter_reg[3]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g10087/_0_  ;
	output \g10220/_1_  ;
	output \g11117/_0_  ;
	output \g11124/_0_  ;
	output \g11125/_0_  ;
	output \g11170/_0_  ;
	output \g11182/_0_  ;
	output \g11184/_0_  ;
	output \g11378/_0_  ;
	output \g11393/_0_  ;
	output \g11415/_0_  ;
	output \g11432/_0_  ;
	output \g11433/_0_  ;
	output \g11453/_0_  ;
	output \g11500/_0_  ;
	output \g11588/_0_  ;
	output \g11607/_0_  ;
	output \g11616/_0_  ;
	output \g11625/_0_  ;
	output \g11641_dup/_0_  ;
	output \g11648/_0_  ;
	output \g11655/_0_  ;
	output \g11683/_0_  ;
	output \g11689/_2_  ;
	output \g11694/_0_  ;
	output \g11748/_0_  ;
	output \g11880/_0_  ;
	output \g11962/_1_  ;
	output \g12016/_0_  ;
	output \g12038/_0_  ;
	output \g12039/_0_  ;
	output \g12094/_0_  ;
	output \g12100/_0_  ;
	output \g12132/_0_  ;
	output \g12151/_0_  ;
	output \g12251/_0_  ;
	output \g12279/_0_  ;
	output \g12288/_0_  ;
	output \g12290/_0_  ;
	output \g12311/_0_  ;
	output \g12313/_0_  ;
	output \g12356/_0_  ;
	output \g12357/_0_  ;
	output \g12427/_0_  ;
	output \g12441/_0_  ;
	output \g12442/_0_  ;
	output \g12480/_0_  ;
	output \g12485/_0_  ;
	output \g12506/_0_  ;
	output \g12544/_0_  ;
	output \g12549/_2_  ;
	output \g12614/_0_  ;
	output \g12678/_0_  ;
	output \g12680/_0_  ;
	output \g12748/_0_  ;
	output \g15/_0_  ;
	output \g25/_0_  ;
	output \g31/_0_  ;
	output \g6843/_0_  ;
	output \g6861/_0_  ;
	output \g6863/_0_  ;
	output \g6865/_0_  ;
	output \g6887/_0_  ;
	output \g6888/_0_  ;
	output \g6889/_0_  ;
	output \g6890/_0_  ;
	output \g6891/_0_  ;
	output \g6892/_0_  ;
	output \g6893/_0_  ;
	output \g6894/_0_  ;
	output \g6922/_0_  ;
	output \g6923/_0_  ;
	output \g6924/_3_  ;
	output \g6926/_0_  ;
	output \g6927/_0_  ;
	output \g6928/_0_  ;
	output \g6931/_0_  ;
	output \g6933/_0_  ;
	output \g6967/_0_  ;
	output \g6968/_0_  ;
	output \g6969/_0_  ;
	output \g6974/_0_  ;
	output \g6975/_0_  ;
	output \g6976/_3_  ;
	output \g7006/_3_  ;
	output \g8882/_0_  ;
	output \g8883/_0_  ;
	output \g8884/_0_  ;
	output \g8895/_0_  ;
	output \g8896/_0_  ;
	output \g8898/_0_  ;
	output \g8900/_2_  ;
	output \g8902/_0_  ;
	output \g8907/_0_  ;
	output \g8911/_0_  ;
	output \g8924/_0_  ;
	output \g8927/_0_  ;
	output \g8929/_2_  ;
	output \g8967/_0_  ;
	output \g8969/_0_  ;
	output \g8973/_2_  ;
	output \g8987/_0_  ;
	output \g8989/_0_  ;
	output \g8991/_0_  ;
	output \g8996/_0_  ;
	output \g9099/_0_  ;
	output \g9543/_1_  ;
	output \g9751/_1_  ;
	output \g9755/_0_  ;
	output \g9786/_0_  ;
	output \g9794/_0_  ;
	output \g9817/_0_  ;
	output \g9836/_0_  ;
	output \g9859/_0_  ;
	output \g9862/_0_  ;
	output \g9867/_0_  ;
	output \g9869/_0_  ;
	output \g9876/_0_  ;
	output \g9887/_0_  ;
	output \g9895/_0_  ;
	output \g9897/_0_  ;
	output \g9908/_0_  ;
	output \g9910/_0_  ;
	output \g9915/_0_  ;
	output \g9938/_0_  ;
	output \g9970/_0_  ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\stage1_iter_reg[1]/NET0131 ,
		\stage1_iter_reg[2]/NET0131 ,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[3]/NET0131 ,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w248_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\data_ready_reg/NET0131 ,
		load_i_pad,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[1]/NET0131 ,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[1]/NET0131 ,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\rd1_Key_o_reg[26]/NET0131 ,
		_w250_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		load_i_pad,
		\rd1_Key_o_reg[26]/NET0131 ,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\key_i[9]_pad ,
		load_i_pad,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w257_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w250_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w256_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\stage1_iter_reg[2]/NET0131 ,
		_w254_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\stage1_iter_reg[3]/NET0131 ,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[3]/NET0131 ,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		_w248_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w263_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w261_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\rd1_Key_o_reg[25]/NET0131 ,
		_w250_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		load_i_pad,
		\rd1_Key_o_reg[25]/NET0131 ,
		_w269_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\key_i[17]_pad ,
		load_i_pad,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w269_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w250_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w268_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		_w266_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w267_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		decrypt_i_pad,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		load_i_pad,
		\rd1_Key_o_reg[27]/NET0131 ,
		_w277_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		\key_i[1]_pad ,
		load_i_pad,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w250_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		load_i_pad,
		_w250_,
		_w281_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\rd1_Key_o_reg[1]/NET0131 ,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\key_i[52]_pad ,
		_w281_,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w282_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		_w266_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		\rd1_Key_o_reg[0]/NET0131 ,
		_w250_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		load_i_pad,
		\rd1_Key_o_reg[0]/NET0131 ,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\key_i[60]_pad ,
		load_i_pad,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w287_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w250_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w286_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w249_,
		_w266_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		_w291_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w280_,
		_w285_,
		_w294_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w293_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		decrypt_i_pad,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w276_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		\rd1_R_o_reg[10]/NET0131 ,
		_w281_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\data_i[43]_pad ,
		_w281_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w298_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\rd1_Key_o_reg[3]/NET0131 ,
		_w281_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\key_i[36]_pad ,
		_w281_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w301_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		_w266_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\rd1_Key_o_reg[4]/NET0131 ,
		_w250_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		load_i_pad,
		\rd1_Key_o_reg[4]/NET0131 ,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		\key_i[59]_pad ,
		load_i_pad,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w250_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w305_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w266_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w304_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		decrypt_i_pad,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\rd1_Key_o_reg[5]/NET0131 ,
		_w281_,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\key_i[51]_pad ,
		_w281_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		_w250_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\rd1_Key_o_reg[7]/NET0131 ,
		_w250_,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		load_i_pad,
		\rd1_Key_o_reg[7]/NET0131 ,
		_w319_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		\key_i[35]_pad ,
		load_i_pad,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w319_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w250_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w318_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		_w266_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\rd1_Key_o_reg[6]/NET0131 ,
		_w250_,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		load_i_pad,
		\rd1_Key_o_reg[6]/NET0131 ,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\key_i[43]_pad ,
		load_i_pad,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w326_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w250_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w325_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		_w292_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w317_,
		_w324_,
		_w332_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w331_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		decrypt_i_pad,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w313_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		\rd1_Key_o_reg[28]/NET0131 ,
		_w250_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		load_i_pad,
		\rd1_Key_o_reg[28]/NET0131 ,
		_w337_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\key_i[28]_pad ,
		load_i_pad,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w337_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w250_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w336_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w266_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\rd1_Key_o_reg[55]/NET0131 ,
		_w250_,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		\key_i[7]_pad ,
		load_i_pad,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		load_i_pad,
		\rd1_Key_o_reg[55]/NET0131 ,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w344_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w250_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w343_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		_w266_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w342_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		decrypt_i_pad,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		load_i_pad,
		\rd1_Key_o_reg[29]/NET0131 ,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		\key_i[20]_pad ,
		load_i_pad,
		_w353_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w352_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w250_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		\rd1_Key_o_reg[31]/NET0131 ,
		_w250_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		load_i_pad,
		\rd1_Key_o_reg[31]/NET0131 ,
		_w357_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\key_i[4]_pad ,
		load_i_pad,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w357_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w250_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w356_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		_w266_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\rd1_Key_o_reg[30]/NET0131 ,
		_w250_,
		_w363_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		\key_i[12]_pad ,
		load_i_pad,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		load_i_pad,
		\rd1_Key_o_reg[30]/NET0131 ,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w364_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w250_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w363_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		_w292_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w355_,
		_w362_,
		_w370_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		_w369_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		decrypt_i_pad,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w351_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\rd1_R_o_reg[4]/NET0131 ,
		_w281_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\data_i[25]_pad ,
		_w281_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w374_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		\rd1_Key_o_reg[21]/NET0131 ,
		_w250_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		load_i_pad,
		\rd1_Key_o_reg[21]/NET0131 ,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		\key_i[49]_pad ,
		load_i_pad,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w250_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w377_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w266_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		\rd1_Key_o_reg[20]/NET0131 ,
		_w250_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		load_i_pad,
		\rd1_Key_o_reg[20]/NET0131 ,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		\key_i[57]_pad ,
		load_i_pad,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w385_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w250_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w384_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		_w266_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w383_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		decrypt_i_pad,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\rd1_Key_o_reg[24]/NET0131 ,
		_w250_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		load_i_pad,
		\rd1_Key_o_reg[24]/NET0131 ,
		_w394_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		\key_i[25]_pad ,
		load_i_pad,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w394_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w250_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w393_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		_w266_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		\rd1_Key_o_reg[23]/NET0131 ,
		_w281_,
		_w400_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		\key_i[33]_pad ,
		_w281_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w400_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		_w292_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		load_i_pad,
		\rd1_Key_o_reg[22]/NET0131 ,
		_w404_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		\key_i[41]_pad ,
		load_i_pad,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w404_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w250_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w399_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		_w403_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h2)
	) name162 (
		decrypt_i_pad,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w392_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w266_,
		_w330_,
		_w412_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		_w266_,
		_w316_,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w412_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		decrypt_i_pad,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		\rd1_Key_o_reg[9]/NET0131 ,
		_w281_,
		_w416_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\key_i[19]_pad ,
		_w281_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w416_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		_w266_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\rd1_Key_o_reg[8]/NET0131 ,
		_w281_,
		_w420_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		\key_i[27]_pad ,
		_w281_,
		_w421_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w420_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		_w292_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w322_,
		_w419_,
		_w424_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		_w423_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		decrypt_i_pad,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w415_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h2)
	) name180 (
		\rd1_Key_o_reg[10]/NET0131 ,
		_w250_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		load_i_pad,
		\rd1_Key_o_reg[10]/NET0131 ,
		_w429_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		\key_i[11]_pad ,
		load_i_pad,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w429_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w250_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w428_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w266_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w419_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		decrypt_i_pad,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		\rd1_Key_o_reg[12]/NET0131 ,
		_w281_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\key_i[58]_pad ,
		_w281_,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w437_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		_w292_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		\rd1_Key_o_reg[13]/NET0131 ,
		_w281_,
		_w441_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\key_i[50]_pad ,
		_w281_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w441_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h2)
	) name196 (
		_w266_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		load_i_pad,
		\rd1_Key_o_reg[11]/NET0131 ,
		_w445_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		\key_i[3]_pad ,
		load_i_pad,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		_w445_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w250_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w440_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h4)
	) name202 (
		_w444_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		decrypt_i_pad,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w436_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h2)
	) name205 (
		\rd1_Key_o_reg[29]/NET0131 ,
		_w250_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w355_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w266_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h2)
	) name208 (
		_w266_,
		_w341_,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		_w455_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		decrypt_i_pad,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\rd1_Key_o_reg[32]/NET0131 ,
		_w250_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		load_i_pad,
		\rd1_Key_o_reg[32]/NET0131 ,
		_w460_
	);
	LUT2 #(
		.INIT('h4)
	) name213 (
		\key_i[61]_pad ,
		load_i_pad,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w460_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		_w250_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w459_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h2)
	) name217 (
		_w266_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		_w292_,
		_w361_,
		_w466_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w367_,
		_w465_,
		_w467_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		_w466_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		decrypt_i_pad,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		_w458_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		_w266_,
		_w361_,
		_w471_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		_w266_,
		_w368_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w471_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		decrypt_i_pad,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h2)
	) name227 (
		\rd1_Key_o_reg[34]/NET0131 ,
		_w250_,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		load_i_pad,
		\rd1_Key_o_reg[34]/NET0131 ,
		_w476_
	);
	LUT2 #(
		.INIT('h4)
	) name229 (
		\key_i[45]_pad ,
		load_i_pad,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w476_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w250_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w475_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h2)
	) name233 (
		_w266_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		\rd1_Key_o_reg[33]/NET0131 ,
		_w281_,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\key_i[53]_pad ,
		_w281_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w482_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		_w292_,
		_w484_,
		_w485_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w463_,
		_w481_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w485_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		decrypt_i_pad,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		_w474_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h2)
	) name242 (
		\rd1_R_o_reg[29]/NET0131 ,
		_w281_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name243 (
		\data_i[23]_pad ,
		_w281_,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w490_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		_w292_,
		_w418_,
		_w493_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		_w266_,
		_w422_,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		_w250_,
		_w418_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		_w493_,
		_w494_,
		_w496_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		_w495_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		decrypt_i_pad,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		_w266_,
		_w439_,
		_w499_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		\rd1_Key_o_reg[11]/NET0131 ,
		_w250_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w448_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		_w292_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w432_,
		_w499_,
		_w503_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		_w502_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h2)
	) name257 (
		decrypt_i_pad,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w498_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w266_,
		_w464_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w362_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		decrypt_i_pad,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		_w250_,
		_w484_,
		_w510_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\rd1_Key_o_reg[35]/NET0131 ,
		_w250_,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		load_i_pad,
		\rd1_Key_o_reg[35]/NET0131 ,
		_w512_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		\key_i[37]_pad ,
		load_i_pad,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w512_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w250_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w511_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		_w266_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		_w292_,
		_w480_,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w510_,
		_w517_,
		_w519_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		_w518_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		decrypt_i_pad,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w509_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		\rd1_Key_o_reg[22]/NET0131 ,
		_w250_,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w407_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w266_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		_w266_,
		_w382_,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w525_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		decrypt_i_pad,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		_w250_,
		_w402_,
		_w529_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		_w292_,
		_w398_,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w274_,
		_w529_,
		_w531_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		_w530_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		decrypt_i_pad,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w528_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w266_,
		_w291_,
		_w535_
	);
	LUT2 #(
		.INIT('h2)
	) name288 (
		\rd1_Key_o_reg[27]/NET0131 ,
		_w250_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		_w266_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w535_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		decrypt_i_pad,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		_w250_,
		_w284_,
		_w540_
	);
	LUT2 #(
		.INIT('h2)
	) name293 (
		\rd1_Key_o_reg[2]/NET0131 ,
		_w250_,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		load_i_pad,
		\rd1_Key_o_reg[2]/NET0131 ,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		\key_i[44]_pad ,
		load_i_pad,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w542_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		_w250_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w541_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		_w292_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w304_,
		_w540_,
		_w548_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		_w547_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		decrypt_i_pad,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w539_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		load_i_pad,
		\rd1_Key_o_reg[48]/NET0131 ,
		_w552_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		\key_i[63]_pad ,
		load_i_pad,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w552_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w250_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h2)
	) name308 (
		\rd1_Key_o_reg[50]/NET0131 ,
		_w250_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		load_i_pad,
		\rd1_Key_o_reg[50]/NET0131 ,
		_w557_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		\key_i[47]_pad ,
		load_i_pad,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w557_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		_w250_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w556_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		_w266_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		\rd1_Key_o_reg[49]/NET0131 ,
		_w250_,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		load_i_pad,
		\rd1_Key_o_reg[49]/NET0131 ,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		\key_i[55]_pad ,
		load_i_pad,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w564_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w250_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w563_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		_w292_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w555_,
		_w562_,
		_w570_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		_w569_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h2)
	) name324 (
		decrypt_i_pad,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h2)
	) name325 (
		\rd1_Key_o_reg[47]/NET0131 ,
		_w281_,
		_w573_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		\key_i[6]_pad ,
		_w281_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w573_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h2)
	) name328 (
		_w250_,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		\rd1_Key_o_reg[46]/NET0131 ,
		_w281_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		\key_i[14]_pad ,
		_w281_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		_w577_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		_w266_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h2)
	) name333 (
		_w292_,
		_w575_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w576_,
		_w580_,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w581_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		decrypt_i_pad,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w572_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h2)
	) name338 (
		\rd1_R_o_reg[13]/NET0131 ,
		_w281_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\data_i[19]_pad ,
		_w281_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w266_,
		_w516_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w481_,
		_w589_,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		decrypt_i_pad,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		load_i_pad,
		\rd1_Key_o_reg[36]/NET0131 ,
		_w592_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		\key_i[29]_pad ,
		load_i_pad,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w592_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		_w250_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h2)
	) name348 (
		\rd1_Key_o_reg[38]/NET0131 ,
		_w281_,
		_w596_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		\key_i[13]_pad ,
		_w281_,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w596_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		_w266_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		\rd1_Key_o_reg[37]/NET0131 ,
		_w250_,
		_w600_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		load_i_pad,
		\rd1_Key_o_reg[37]/NET0131 ,
		_w601_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		\key_i[21]_pad ,
		load_i_pad,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		_w601_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w250_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w600_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		_w292_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w595_,
		_w599_,
		_w607_
	);
	LUT2 #(
		.INIT('h4)
	) name360 (
		_w606_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		decrypt_i_pad,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w591_,
		_w609_,
		_w610_
	);
	LUT2 #(
		.INIT('h2)
	) name363 (
		\rd1_Key_o_reg[48]/NET0131 ,
		_w250_,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w555_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w266_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		_w266_,
		_w575_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w613_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		decrypt_i_pad,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h2)
	) name369 (
		\rd1_Key_o_reg[51]/NET0131 ,
		_w250_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		load_i_pad,
		\rd1_Key_o_reg[51]/NET0131 ,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		\key_i[39]_pad ,
		load_i_pad,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w618_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		_w250_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w617_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		_w266_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		_w292_,
		_w561_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w567_,
		_w623_,
		_w625_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w624_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h2)
	) name379 (
		decrypt_i_pad,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w616_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h2)
	) name381 (
		\rd1_Key_o_reg[15]/NET0131 ,
		_w250_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		load_i_pad,
		\rd1_Key_o_reg[15]/NET0131 ,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		\key_i[34]_pad ,
		load_i_pad,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w630_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w250_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		_w629_,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		_w266_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h2)
	) name388 (
		\rd1_Key_o_reg[16]/NET0131 ,
		_w250_,
		_w636_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		load_i_pad,
		\rd1_Key_o_reg[16]/NET0131 ,
		_w637_
	);
	LUT2 #(
		.INIT('h4)
	) name390 (
		\key_i[26]_pad ,
		load_i_pad,
		_w638_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w637_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		_w250_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w636_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w266_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w635_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		decrypt_i_pad,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		load_i_pad,
		\rd1_Key_o_reg[17]/NET0131 ,
		_w645_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		\key_i[18]_pad ,
		load_i_pad,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		_w645_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		_w250_,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h2)
	) name401 (
		\rd1_Key_o_reg[19]/NET0131 ,
		_w281_,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name402 (
		\key_i[2]_pad ,
		_w281_,
		_w650_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w649_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h2)
	) name404 (
		_w266_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h2)
	) name405 (
		\rd1_Key_o_reg[18]/NET0131 ,
		_w250_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		load_i_pad,
		\rd1_Key_o_reg[18]/NET0131 ,
		_w654_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		\key_i[10]_pad ,
		load_i_pad,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w654_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w250_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w653_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		_w292_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		_w648_,
		_w652_,
		_w660_
	);
	LUT2 #(
		.INIT('h4)
	) name413 (
		_w659_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		decrypt_i_pad,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w644_,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h2)
	) name416 (
		\rd1_R_o_reg[0]/NET0131 ,
		_w281_,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		\data_i[57]_pad ,
		_w281_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		_w664_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		\rd1_R_o_reg[16]/NET0131 ,
		_w281_,
		_w667_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\data_i[61]_pad ,
		_w281_,
		_w668_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		_w667_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		\rd1_Key_o_reg[14]/NET0131 ,
		_w250_,
		_w670_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		load_i_pad,
		\rd1_Key_o_reg[14]/NET0131 ,
		_w671_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		\key_i[42]_pad ,
		load_i_pad,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w671_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		_w250_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		_w670_,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w266_,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w444_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		decrypt_i_pad,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h2)
	) name431 (
		\rd1_Key_o_reg[17]/NET0131 ,
		_w250_,
		_w679_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		_w266_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		_w292_,
		_w641_,
		_w681_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w633_,
		_w680_,
		_w682_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		_w681_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h2)
	) name436 (
		decrypt_i_pad,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w678_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		\rd1_R_o_reg[7]/NET0131 ,
		_w281_,
		_w686_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		\data_i[1]_pad ,
		_w281_,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		_w686_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h2)
	) name441 (
		_w266_,
		_w454_,
		_w689_
	);
	LUT2 #(
		.INIT('h2)
	) name442 (
		_w292_,
		_w341_,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		_w347_,
		_w689_,
		_w691_
	);
	LUT2 #(
		.INIT('h4)
	) name444 (
		_w690_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h2)
	) name445 (
		decrypt_i_pad,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		\rd1_Key_o_reg[54]/NET0131 ,
		_w281_,
		_w694_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		\key_i[15]_pad ,
		_w281_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		_w694_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h2)
	) name449 (
		_w250_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		_w292_,
		_w696_,
		_w698_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		\rd1_Key_o_reg[53]/NET0131 ,
		_w250_,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		load_i_pad,
		\rd1_Key_o_reg[53]/NET0131 ,
		_w700_
	);
	LUT2 #(
		.INIT('h4)
	) name453 (
		\key_i[23]_pad ,
		load_i_pad,
		_w701_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w700_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w250_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		_w699_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h2)
	) name457 (
		_w266_,
		_w704_,
		_w705_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w697_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h4)
	) name459 (
		_w698_,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		decrypt_i_pad,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w693_,
		_w708_,
		_w709_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		\rd1_Key_o_reg[44]/NET0131 ,
		_w250_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		load_i_pad,
		\rd1_Key_o_reg[44]/NET0131 ,
		_w711_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		\key_i[30]_pad ,
		load_i_pad,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w711_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h8)
	) name466 (
		_w250_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w710_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h2)
	) name468 (
		_w266_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h2)
	) name469 (
		\rd1_Key_o_reg[45]/NET0131 ,
		_w250_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		load_i_pad,
		\rd1_Key_o_reg[45]/NET0131 ,
		_w718_
	);
	LUT2 #(
		.INIT('h4)
	) name471 (
		\key_i[22]_pad ,
		load_i_pad,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w718_,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w250_,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w717_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w266_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		decrypt_i_pad,
		_w716_,
		_w724_
	);
	LUT2 #(
		.INIT('h4)
	) name477 (
		_w723_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		_w250_,
		_w579_,
		_w726_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		_w266_,
		_w612_,
		_w727_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		decrypt_i_pad,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		_w581_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		_w726_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		_w725_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		\rd1_Key_o_reg[36]/NET0131 ,
		_w250_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w595_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w266_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w517_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		decrypt_i_pad,
		_w735_,
		_w736_
	);
	LUT2 #(
		.INIT('h2)
	) name489 (
		\rd1_Key_o_reg[39]/NET0131 ,
		_w250_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		load_i_pad,
		\rd1_Key_o_reg[39]/NET0131 ,
		_w738_
	);
	LUT2 #(
		.INIT('h4)
	) name491 (
		\key_i[5]_pad ,
		load_i_pad,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w738_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h8)
	) name493 (
		_w250_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w737_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h2)
	) name495 (
		_w266_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h2)
	) name496 (
		_w292_,
		_w598_,
		_w744_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w604_,
		_w743_,
		_w745_
	);
	LUT2 #(
		.INIT('h4)
	) name498 (
		_w744_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h2)
	) name499 (
		decrypt_i_pad,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w736_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h2)
	) name501 (
		\rd1_R_o_reg[30]/NET0131 ,
		_w281_,
		_w749_
	);
	LUT2 #(
		.INIT('h8)
	) name502 (
		\data_i[15]_pad ,
		_w281_,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w749_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w266_,
		_w715_,
		_w752_
	);
	LUT2 #(
		.INIT('h2)
	) name505 (
		\rd1_Key_o_reg[43]/NET0131 ,
		_w250_,
		_w753_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		\key_i[38]_pad ,
		load_i_pad,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		load_i_pad,
		\rd1_Key_o_reg[43]/NET0131 ,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w754_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		_w250_,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h1)
	) name510 (
		_w753_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		_w266_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w752_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		decrypt_i_pad,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h2)
	) name514 (
		_w292_,
		_w579_,
		_w762_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w614_,
		_w721_,
		_w763_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w762_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		decrypt_i_pad,
		_w764_,
		_w765_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		_w761_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h2)
	) name519 (
		_w266_,
		_w641_,
		_w767_
	);
	LUT2 #(
		.INIT('h2)
	) name520 (
		_w292_,
		_w634_,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w674_,
		_w767_,
		_w769_
	);
	LUT2 #(
		.INIT('h4)
	) name522 (
		_w768_,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		decrypt_i_pad,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h2)
	) name524 (
		_w292_,
		_w443_,
		_w772_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		_w250_,
		_w443_,
		_w773_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		_w499_,
		_w772_,
		_w774_
	);
	LUT2 #(
		.INIT('h4)
	) name527 (
		_w773_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		decrypt_i_pad,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w771_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		\rd1_R_o_reg[3]/NET0131 ,
		_w281_,
		_w778_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		\data_i[33]_pad ,
		_w281_,
		_w779_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w778_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		_w777_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h2)
	) name534 (
		_w777_,
		_w780_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w781_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		_w292_,
		_w323_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		_w329_,
		_w494_,
		_w785_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		_w784_,
		_w785_,
		_w786_
	);
	LUT2 #(
		.INIT('h2)
	) name539 (
		decrypt_i_pad,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h2)
	) name540 (
		_w292_,
		_w316_,
		_w788_
	);
	LUT2 #(
		.INIT('h2)
	) name541 (
		_w266_,
		_w310_,
		_w789_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		_w317_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h4)
	) name543 (
		_w788_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		decrypt_i_pad,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		_w787_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h2)
	) name546 (
		\rd1_R_o_reg[2]/NET0131 ,
		_w281_,
		_w794_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		\data_i[41]_pad ,
		_w281_,
		_w795_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w794_,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h4)
	) name549 (
		_w793_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h2)
	) name550 (
		_w793_,
		_w796_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		_w797_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w783_,
		_w799_,
		_w800_
	);
	LUT2 #(
		.INIT('h2)
	) name553 (
		_w376_,
		_w506_,
		_w801_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w376_,
		_w506_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w801_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		_w800_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h2)
	) name557 (
		_w266_,
		_w524_,
		_w805_
	);
	LUT2 #(
		.INIT('h2)
	) name558 (
		_w292_,
		_w382_,
		_w806_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		_w388_,
		_w805_,
		_w807_
	);
	LUT2 #(
		.INIT('h4)
	) name560 (
		_w806_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		decrypt_i_pad,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		_w250_,
		_w651_,
		_w810_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		_w292_,
		_w651_,
		_w811_
	);
	LUT2 #(
		.INIT('h2)
	) name564 (
		_w266_,
		_w658_,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		_w810_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		_w811_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		decrypt_i_pad,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w809_,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h2)
	) name569 (
		\rd1_R_o_reg[1]/NET0131 ,
		_w281_,
		_w817_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		\data_i[49]_pad ,
		_w281_,
		_w818_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		_w817_,
		_w818_,
		_w819_
	);
	LUT2 #(
		.INIT('h4)
	) name572 (
		_w816_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h2)
	) name573 (
		_w816_,
		_w819_,
		_w821_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w820_,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		_w804_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h2)
	) name576 (
		_w783_,
		_w803_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name577 (
		_w799_,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h4)
	) name578 (
		_w822_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w823_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		_w799_,
		_w803_,
		_w828_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		_w783_,
		_w822_,
		_w829_
	);
	LUT2 #(
		.INIT('h4)
	) name582 (
		_w799_,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		_w783_,
		_w803_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w830_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		_w828_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		_w827_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h4)
	) name587 (
		_w297_,
		_w666_,
		_w835_
	);
	LUT2 #(
		.INIT('h2)
	) name588 (
		_w297_,
		_w666_,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		_w835_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		_w834_,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		_w799_,
		_w803_,
		_w839_
	);
	LUT2 #(
		.INIT('h4)
	) name592 (
		_w837_,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h2)
	) name593 (
		_w783_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h4)
	) name594 (
		_w803_,
		_w837_,
		_w842_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		_w822_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		_w841_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h4)
	) name597 (
		_w799_,
		_w837_,
		_w845_
	);
	LUT2 #(
		.INIT('h2)
	) name598 (
		_w822_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h4)
	) name599 (
		_w841_,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		_w403_,
		_w805_,
		_w848_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		_w529_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		decrypt_i_pad,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		_w261_,
		_w266_,
		_w851_
	);
	LUT2 #(
		.INIT('h4)
	) name604 (
		_w273_,
		_w292_,
		_w852_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		_w397_,
		_w851_,
		_w853_
	);
	LUT2 #(
		.INIT('h4)
	) name606 (
		_w852_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		decrypt_i_pad,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		_w850_,
		_w855_,
		_w856_
	);
	LUT2 #(
		.INIT('h2)
	) name609 (
		\rd1_R_o_reg[31]/NET0131 ,
		_w281_,
		_w857_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		\data_i[7]_pad ,
		_w281_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w857_,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('h4)
	) name612 (
		_w856_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h2)
	) name613 (
		_w856_,
		_w859_,
		_w861_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w860_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w844_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h4)
	) name616 (
		_w847_,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h4)
	) name617 (
		_w838_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h4)
	) name618 (
		_w822_,
		_w828_,
		_w866_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		_w783_,
		_w866_,
		_w867_
	);
	LUT2 #(
		.INIT('h4)
	) name620 (
		_w822_,
		_w824_,
		_w868_
	);
	LUT2 #(
		.INIT('h4)
	) name621 (
		_w825_,
		_w837_,
		_w869_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		_w803_,
		_w829_,
		_w870_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		_w800_,
		_w868_,
		_w871_
	);
	LUT2 #(
		.INIT('h4)
	) name624 (
		_w870_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h8)
	) name625 (
		_w869_,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		_w827_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h8)
	) name627 (
		_w803_,
		_w822_,
		_w875_
	);
	LUT2 #(
		.INIT('h2)
	) name628 (
		_w799_,
		_w824_,
		_w876_
	);
	LUT2 #(
		.INIT('h4)
	) name629 (
		_w875_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w830_,
		_w837_,
		_w878_
	);
	LUT2 #(
		.INIT('h4)
	) name631 (
		_w877_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		_w874_,
		_w879_,
		_w880_
	);
	LUT2 #(
		.INIT('h2)
	) name633 (
		_w862_,
		_w867_,
		_w881_
	);
	LUT2 #(
		.INIT('h4)
	) name634 (
		_w880_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w865_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h4)
	) name636 (
		\data_i[16]_pad ,
		_w281_,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		\rd1_L_o_reg[5]/NET0131 ,
		_w281_,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		_w884_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h2)
	) name639 (
		_w883_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h4)
	) name640 (
		_w883_,
		_w886_,
		_w888_
	);
	LUT2 #(
		.INIT('h1)
	) name641 (
		_w887_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h2)
	) name642 (
		\rd1_R_o_reg[18]/NET0131 ,
		_w281_,
		_w890_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		\data_i[45]_pad ,
		_w281_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w890_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h4)
	) name645 (
		_w373_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		_w373_,
		_w892_,
		_w894_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w893_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h2)
	) name648 (
		\rd1_R_o_reg[17]/NET0131 ,
		_w281_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		\data_i[53]_pad ,
		_w281_,
		_w897_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w896_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h4)
	) name651 (
		_w610_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		_w610_,
		_w898_,
		_w900_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w899_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		_w895_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		\rd1_R_o_reg[19]/NET0131 ,
		_w281_,
		_w903_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		\data_i[37]_pad ,
		_w281_,
		_w904_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w903_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w628_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		_w628_,
		_w905_,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		_w906_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w266_,
		_w742_,
		_w909_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w599_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		decrypt_i_pad,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		load_i_pad,
		\rd1_Key_o_reg[40]/NET0131 ,
		_w912_
	);
	LUT2 #(
		.INIT('h4)
	) name665 (
		\key_i[62]_pad ,
		load_i_pad,
		_w913_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w912_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h8)
	) name667 (
		_w250_,
		_w914_,
		_w915_
	);
	LUT2 #(
		.INIT('h2)
	) name668 (
		\rd1_Key_o_reg[42]/NET0131 ,
		_w281_,
		_w916_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		\key_i[46]_pad ,
		_w281_,
		_w917_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w916_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h2)
	) name671 (
		_w266_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h2)
	) name672 (
		\rd1_Key_o_reg[41]/NET0131 ,
		_w250_,
		_w920_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		load_i_pad,
		\rd1_Key_o_reg[41]/NET0131 ,
		_w921_
	);
	LUT2 #(
		.INIT('h4)
	) name674 (
		\key_i[54]_pad ,
		load_i_pad,
		_w922_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w921_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h8)
	) name676 (
		_w250_,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		_w920_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h2)
	) name678 (
		_w292_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w915_,
		_w919_,
		_w927_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		_w926_,
		_w927_,
		_w928_
	);
	LUT2 #(
		.INIT('h2)
	) name681 (
		decrypt_i_pad,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		_w911_,
		_w929_,
		_w930_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		\rd1_R_o_reg[20]/NET0131 ,
		_w281_,
		_w931_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		\data_i[29]_pad ,
		_w281_,
		_w932_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		_w931_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		_w930_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h2)
	) name687 (
		_w930_,
		_w933_,
		_w935_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		_w934_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w908_,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		_w908_,
		_w936_,
		_w938_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		_w937_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h2)
	) name692 (
		_w902_,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h8)
	) name693 (
		_w895_,
		_w939_,
		_w941_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		_w895_,
		_w937_,
		_w942_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w941_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		_w292_,
		_w918_,
		_w944_
	);
	LUT2 #(
		.INIT('h2)
	) name697 (
		_w250_,
		_w918_,
		_w945_
	);
	LUT2 #(
		.INIT('h2)
	) name698 (
		_w266_,
		_w925_,
		_w946_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w944_,
		_w946_,
		_w947_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w945_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		decrypt_i_pad,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h2)
	) name702 (
		_w266_,
		_w722_,
		_w950_
	);
	LUT2 #(
		.INIT('h2)
	) name703 (
		_w292_,
		_w715_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w757_,
		_w950_,
		_w952_
	);
	LUT2 #(
		.INIT('h4)
	) name705 (
		_w951_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h2)
	) name706 (
		decrypt_i_pad,
		_w953_,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w949_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h2)
	) name708 (
		_w669_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h4)
	) name709 (
		_w669_,
		_w955_,
		_w957_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w956_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w943_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		_w901_,
		_w938_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w895_,
		_w901_,
		_w961_
	);
	LUT2 #(
		.INIT('h8)
	) name714 (
		_w939_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w960_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h2)
	) name716 (
		_w958_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w940_,
		_w959_,
		_w965_
	);
	LUT2 #(
		.INIT('h4)
	) name718 (
		_w964_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		_w266_,
		_w704_,
		_w967_
	);
	LUT2 #(
		.INIT('h2)
	) name720 (
		\rd1_Key_o_reg[52]/NET0131 ,
		_w250_,
		_w968_
	);
	LUT2 #(
		.INIT('h4)
	) name721 (
		\key_i[31]_pad ,
		load_i_pad,
		_w969_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		load_i_pad,
		\rd1_Key_o_reg[52]/NET0131 ,
		_w970_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w969_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h8)
	) name724 (
		_w250_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name725 (
		_w968_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h2)
	) name726 (
		_w266_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		_w967_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		decrypt_i_pad,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h2)
	) name729 (
		_w292_,
		_w348_,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name730 (
		_w456_,
		_w697_,
		_w978_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		_w977_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h2)
	) name732 (
		decrypt_i_pad,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h1)
	) name733 (
		_w976_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h2)
	) name734 (
		\rd1_R_o_reg[15]/NET0131 ,
		_w281_,
		_w982_
	);
	LUT2 #(
		.INIT('h8)
	) name735 (
		\data_i[3]_pad ,
		_w281_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w982_,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h4)
	) name737 (
		_w981_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h2)
	) name738 (
		_w981_,
		_w984_,
		_w986_
	);
	LUT2 #(
		.INIT('h1)
	) name739 (
		_w985_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h4)
	) name740 (
		_w966_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h2)
	) name741 (
		_w902_,
		_w936_,
		_w989_
	);
	LUT2 #(
		.INIT('h4)
	) name742 (
		_w958_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		_w908_,
		_w936_,
		_w991_
	);
	LUT2 #(
		.INIT('h8)
	) name744 (
		_w901_,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		_w901_,
		_w936_,
		_w993_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		_w908_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w992_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h4)
	) name748 (
		_w941_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h2)
	) name749 (
		_w958_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name750 (
		_w938_,
		_w961_,
		_w998_
	);
	LUT2 #(
		.INIT('h1)
	) name751 (
		_w990_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		_w997_,
		_w999_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		_w987_,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h8)
	) name754 (
		_w895_,
		_w991_,
		_w1002_
	);
	LUT2 #(
		.INIT('h8)
	) name755 (
		_w901_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h4)
	) name756 (
		_w895_,
		_w938_,
		_w1004_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w994_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		_w958_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		_w961_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h2)
	) name760 (
		_w895_,
		_w901_,
		_w1008_
	);
	LUT2 #(
		.INIT('h8)
	) name761 (
		_w908_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h8)
	) name762 (
		_w901_,
		_w937_,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		_w1009_,
		_w1010_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w958_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w1003_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h4)
	) name766 (
		_w1007_,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h4)
	) name767 (
		_w1001_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h4)
	) name768 (
		_w988_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h4)
	) name769 (
		\data_i[8]_pad ,
		_w281_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		\rd1_L_o_reg[6]/NET0131 ,
		_w281_,
		_w1018_
	);
	LUT2 #(
		.INIT('h1)
	) name771 (
		_w1017_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h2)
	) name772 (
		_w1016_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h4)
	) name773 (
		_w1016_,
		_w1019_,
		_w1021_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		_w1020_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		_w266_,
		_w273_,
		_w1023_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		_w399_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		decrypt_i_pad,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h2)
	) name778 (
		_w266_,
		_w291_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		_w280_,
		_w536_,
		_w1027_
	);
	LUT2 #(
		.INIT('h2)
	) name780 (
		_w292_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h1)
	) name781 (
		_w260_,
		_w1026_,
		_w1029_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w1028_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h2)
	) name783 (
		decrypt_i_pad,
		_w1030_,
		_w1031_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w1025_,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w266_,
		_w561_,
		_w1033_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		_w266_,
		_w568_,
		_w1034_
	);
	LUT2 #(
		.INIT('h1)
	) name787 (
		_w1033_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		decrypt_i_pad,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h2)
	) name789 (
		_w292_,
		_w973_,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		_w621_,
		_w705_,
		_w1038_
	);
	LUT2 #(
		.INIT('h4)
	) name791 (
		_w1037_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h2)
	) name792 (
		decrypt_i_pad,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w1036_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		_w266_,
		_w658_,
		_w1042_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w680_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name796 (
		decrypt_i_pad,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h2)
	) name797 (
		_w292_,
		_w389_,
		_w1045_
	);
	LUT2 #(
		.INIT('h1)
	) name798 (
		_w526_,
		_w810_,
		_w1046_
	);
	LUT2 #(
		.INIT('h4)
	) name799 (
		_w1045_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h2)
	) name800 (
		decrypt_i_pad,
		_w1047_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		_w1044_,
		_w1048_,
		_w1049_
	);
	LUT2 #(
		.INIT('h2)
	) name802 (
		_w266_,
		_w330_,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		_w309_,
		_w1050_,
		_w1051_
	);
	LUT2 #(
		.INIT('h4)
	) name804 (
		_w788_,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h2)
	) name805 (
		decrypt_i_pad,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h2)
	) name806 (
		_w250_,
		_w303_,
		_w1054_
	);
	LUT2 #(
		.INIT('h2)
	) name807 (
		_w292_,
		_w303_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name808 (
		_w266_,
		_w546_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		_w1054_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h4)
	) name810 (
		_w1055_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		decrypt_i_pad,
		_w1058_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w1053_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h2)
	) name813 (
		\rd1_R_o_reg[28]/NET0131 ,
		_w281_,
		_w1061_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		\data_i[31]_pad ,
		_w281_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w1061_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w266_,
		_w973_,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w623_,
		_w1064_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		decrypt_i_pad,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		_w349_,
		_w703_,
		_w1067_
	);
	LUT2 #(
		.INIT('h4)
	) name820 (
		_w698_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h2)
	) name821 (
		decrypt_i_pad,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w1066_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h2)
	) name823 (
		\rd1_Key_o_reg[40]/NET0131 ,
		_w250_,
		_w1071_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w915_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h1)
	) name825 (
		_w266_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w743_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h1)
	) name827 (
		decrypt_i_pad,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w759_,
		_w924_,
		_w1076_
	);
	LUT2 #(
		.INIT('h4)
	) name829 (
		_w944_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h2)
	) name830 (
		decrypt_i_pad,
		_w1077_,
		_w1078_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		_w1075_,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		\rd1_R_o_reg[26]/NET0131 ,
		_w281_,
		_w1080_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		\data_i[47]_pad ,
		_w281_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name834 (
		_w1080_,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h2)
	) name835 (
		_w250_,
		_w422_,
		_w1083_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w324_,
		_w423_,
		_w1084_
	);
	LUT2 #(
		.INIT('h4)
	) name837 (
		_w1083_,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		decrypt_i_pad,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		_w266_,
		_w501_,
		_w1087_
	);
	LUT2 #(
		.INIT('h2)
	) name840 (
		_w292_,
		_w433_,
		_w1088_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		_w495_,
		_w1087_,
		_w1089_
	);
	LUT2 #(
		.INIT('h4)
	) name842 (
		_w1088_,
		_w1089_,
		_w1090_
	);
	LUT2 #(
		.INIT('h2)
	) name843 (
		decrypt_i_pad,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		_w1086_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h2)
	) name845 (
		\rd1_R_o_reg[12]/NET0131 ,
		_w281_,
		_w1093_
	);
	LUT2 #(
		.INIT('h8)
	) name846 (
		\data_i[27]_pad ,
		_w281_,
		_w1094_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		_w1093_,
		_w1094_,
		_w1095_
	);
	LUT2 #(
		.INIT('h4)
	) name848 (
		_w1092_,
		_w1095_,
		_w1096_
	);
	LUT2 #(
		.INIT('h2)
	) name849 (
		_w1092_,
		_w1095_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		_w1096_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h2)
	) name851 (
		_w669_,
		_w685_,
		_w1099_
	);
	LUT2 #(
		.INIT('h4)
	) name852 (
		_w669_,
		_w685_,
		_w1100_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w1099_,
		_w1100_,
		_w1101_
	);
	LUT2 #(
		.INIT('h2)
	) name854 (
		_w984_,
		_w1060_,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		_w984_,
		_w1060_,
		_w1103_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w1102_,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w1101_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		_w1101_,
		_w1104_,
		_w1106_
	);
	LUT2 #(
		.INIT('h2)
	) name859 (
		_w588_,
		_w1049_,
		_w1107_
	);
	LUT2 #(
		.INIT('h4)
	) name860 (
		_w588_,
		_w1049_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h2)
	) name862 (
		_w1106_,
		_w1109_,
		_w1110_
	);
	LUT2 #(
		.INIT('h1)
	) name863 (
		_w1105_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('h2)
	) name864 (
		_w266_,
		_w402_,
		_w1112_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		_w266_,
		_w398_,
		_w1113_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		_w1112_,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		decrypt_i_pad,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h4)
	) name868 (
		_w261_,
		_w292_,
		_w1116_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		_w272_,
		_w537_,
		_w1117_
	);
	LUT2 #(
		.INIT('h4)
	) name870 (
		_w1116_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h2)
	) name871 (
		decrypt_i_pad,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w1115_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h2)
	) name873 (
		\rd1_R_o_reg[14]/NET0131 ,
		_w281_,
		_w1121_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		\data_i[11]_pad ,
		_w281_,
		_w1122_
	);
	LUT2 #(
		.INIT('h1)
	) name875 (
		_w1121_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h4)
	) name876 (
		_w1120_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h2)
	) name877 (
		_w1120_,
		_w1123_,
		_w1125_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w1124_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h1)
	) name879 (
		_w1111_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h1)
	) name880 (
		_w1101_,
		_w1104_,
		_w1128_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		_w1109_,
		_w1128_,
		_w1129_
	);
	LUT2 #(
		.INIT('h2)
	) name882 (
		_w1104_,
		_w1109_,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		_w1126_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w1098_,
		_w1129_,
		_w1132_
	);
	LUT2 #(
		.INIT('h4)
	) name885 (
		_w1131_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w1127_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h2)
	) name887 (
		_w1104_,
		_w1126_,
		_w1135_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		_w1101_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h2)
	) name889 (
		_w1098_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h8)
	) name890 (
		_w1104_,
		_w1109_,
		_w1138_
	);
	LUT2 #(
		.INIT('h4)
	) name891 (
		_w1104_,
		_w1126_,
		_w1139_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w1138_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		_w1101_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h1)
	) name894 (
		_w1109_,
		_w1126_,
		_w1142_
	);
	LUT2 #(
		.INIT('h8)
	) name895 (
		_w1128_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		_w1137_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h4)
	) name897 (
		_w1141_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		_w1134_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name899 (
		_w1105_,
		_w1126_,
		_w1147_
	);
	LUT2 #(
		.INIT('h4)
	) name900 (
		_w1109_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h4)
	) name901 (
		_w1126_,
		_w1138_,
		_w1149_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		_w1101_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w1148_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h4)
	) name904 (
		_w1146_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		\rd1_R_o_reg[11]/NET0131 ,
		_w281_,
		_w1153_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		\data_i[35]_pad ,
		_w281_,
		_w1154_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w1153_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h4)
	) name908 (
		_w551_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h2)
	) name909 (
		_w551_,
		_w1155_,
		_w1157_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w1156_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w1152_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h8)
	) name912 (
		_w1101_,
		_w1126_,
		_w1160_
	);
	LUT2 #(
		.INIT('h1)
	) name913 (
		_w1101_,
		_w1109_,
		_w1161_
	);
	LUT2 #(
		.INIT('h1)
	) name914 (
		_w1160_,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w1130_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h8)
	) name916 (
		_w1101_,
		_w1142_,
		_w1164_
	);
	LUT2 #(
		.INIT('h8)
	) name917 (
		_w1104_,
		_w1164_,
		_w1165_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		_w1163_,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h2)
	) name919 (
		_w1158_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h4)
	) name920 (
		_w1101_,
		_w1138_,
		_w1168_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		_w1126_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w1167_,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h1)
	) name923 (
		_w1098_,
		_w1170_,
		_w1171_
	);
	LUT2 #(
		.INIT('h8)
	) name924 (
		_w1098_,
		_w1109_,
		_w1172_
	);
	LUT2 #(
		.INIT('h4)
	) name925 (
		_w1135_,
		_w1172_,
		_w1173_
	);
	LUT2 #(
		.INIT('h4)
	) name926 (
		_w1101_,
		_w1173_,
		_w1174_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w1101_,
		_w1135_,
		_w1175_
	);
	LUT2 #(
		.INIT('h2)
	) name928 (
		_w1140_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h8)
	) name929 (
		_w1137_,
		_w1176_,
		_w1177_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		_w1174_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h2)
	) name931 (
		_w1158_,
		_w1178_,
		_w1179_
	);
	LUT2 #(
		.INIT('h8)
	) name932 (
		_w1101_,
		_w1138_,
		_w1180_
	);
	LUT2 #(
		.INIT('h2)
	) name933 (
		_w1098_,
		_w1126_,
		_w1181_
	);
	LUT2 #(
		.INIT('h8)
	) name934 (
		_w1180_,
		_w1181_,
		_w1182_
	);
	LUT2 #(
		.INIT('h4)
	) name935 (
		_w1109_,
		_w1158_,
		_w1183_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w1172_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h8)
	) name937 (
		_w1126_,
		_w1128_,
		_w1185_
	);
	LUT2 #(
		.INIT('h4)
	) name938 (
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		_w1182_,
		_w1186_,
		_w1187_
	);
	LUT2 #(
		.INIT('h4)
	) name940 (
		_w1179_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w1171_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h4)
	) name942 (
		_w1159_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name943 (
		\data_i[44]_pad ,
		_w281_,
		_w1191_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		\rd1_L_o_reg[18]/NET0131 ,
		_w281_,
		_w1192_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		_w1191_,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h2)
	) name946 (
		_w1190_,
		_w1193_,
		_w1194_
	);
	LUT2 #(
		.INIT('h4)
	) name947 (
		_w1190_,
		_w1193_,
		_w1195_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		_w1194_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h2)
	) name949 (
		\rd1_R_o_reg[8]/NET0131 ,
		_w281_,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		\data_i[59]_pad ,
		_w281_,
		_w1198_
	);
	LUT2 #(
		.INIT('h1)
	) name951 (
		_w1197_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h1)
	) name952 (
		_w266_,
		_w501_,
		_w1200_
	);
	LUT2 #(
		.INIT('h2)
	) name953 (
		_w266_,
		_w433_,
		_w1201_
	);
	LUT2 #(
		.INIT('h1)
	) name954 (
		_w1200_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		decrypt_i_pad,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h2)
	) name956 (
		_w250_,
		_w439_,
		_w1204_
	);
	LUT2 #(
		.INIT('h2)
	) name957 (
		_w266_,
		_w675_,
		_w1205_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		_w772_,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name959 (
		_w1204_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name960 (
		decrypt_i_pad,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h1)
	) name961 (
		_w1203_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		_w266_,
		_w634_,
		_w1210_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w1205_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		decrypt_i_pad,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		_w648_,
		_w679_,
		_w1213_
	);
	LUT2 #(
		.INIT('h2)
	) name966 (
		_w292_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		_w640_,
		_w812_,
		_w1215_
	);
	LUT2 #(
		.INIT('h4)
	) name968 (
		_w1214_,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h2)
	) name969 (
		decrypt_i_pad,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		_w1212_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		_w266_,
		_w323_,
		_w1219_
	);
	LUT2 #(
		.INIT('h1)
	) name972 (
		_w1050_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		decrypt_i_pad,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		_w493_,
		_w1201_,
		_w1222_
	);
	LUT2 #(
		.INIT('h4)
	) name975 (
		_w1083_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h2)
	) name976 (
		decrypt_i_pad,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		_w1221_,
		_w1224_,
		_w1225_
	);
	LUT2 #(
		.INIT('h1)
	) name978 (
		_w266_,
		_w568_,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w727_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h1)
	) name980 (
		decrypt_i_pad,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h2)
	) name981 (
		_w292_,
		_w622_,
		_w1229_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		_w560_,
		_w974_,
		_w1230_
	);
	LUT2 #(
		.INIT('h4)
	) name983 (
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h2)
	) name984 (
		decrypt_i_pad,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w1228_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h2)
	) name986 (
		\rd1_R_o_reg[25]/NET0131 ,
		_w281_,
		_w1234_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		\data_i[55]_pad ,
		_w281_,
		_w1235_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		_w1234_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		_w1233_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h2)
	) name990 (
		_w1233_,
		_w1236_,
		_w1238_
	);
	LUT2 #(
		.INIT('h1)
	) name991 (
		_w1237_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h4)
	) name992 (
		_w1079_,
		_w1082_,
		_w1240_
	);
	LUT2 #(
		.INIT('h2)
	) name993 (
		_w1079_,
		_w1082_,
		_w1241_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w1240_,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w266_,
		_w348_,
		_w1243_
	);
	LUT2 #(
		.INIT('h2)
	) name996 (
		_w266_,
		_w696_,
		_w1244_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w1243_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		decrypt_i_pad,
		_w1245_,
		_w1246_
	);
	LUT2 #(
		.INIT('h2)
	) name999 (
		_w292_,
		_w454_,
		_w1247_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w340_,
		_w472_,
		_w1248_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		_w1247_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h2)
	) name1002 (
		decrypt_i_pad,
		_w1249_,
		_w1250_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w1246_,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h2)
	) name1004 (
		\rd1_R_o_reg[27]/NET0131 ,
		_w281_,
		_w1252_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		\data_i[39]_pad ,
		_w281_,
		_w1253_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		_w1252_,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h4)
	) name1007 (
		_w1251_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h2)
	) name1008 (
		_w1251_,
		_w1254_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w1255_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		_w1242_,
		_w1257_,
		_w1258_
	);
	LUT2 #(
		.INIT('h2)
	) name1011 (
		_w1063_,
		_w1070_,
		_w1259_
	);
	LUT2 #(
		.INIT('h4)
	) name1012 (
		_w1063_,
		_w1070_,
		_w1260_
	);
	LUT2 #(
		.INIT('h1)
	) name1013 (
		_w1259_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h8)
	) name1014 (
		_w1258_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h8)
	) name1015 (
		_w1239_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h2)
	) name1016 (
		\rd1_R_o_reg[23]/NET0131 ,
		_w281_,
		_w1264_
	);
	LUT2 #(
		.INIT('h8)
	) name1017 (
		\data_i[5]_pad ,
		_w281_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w1264_,
		_w1265_,
		_w1266_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		_w731_,
		_w1266_,
		_w1267_
	);
	LUT2 #(
		.INIT('h1)
	) name1020 (
		_w731_,
		_w1266_,
		_w1268_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		_w1267_,
		_w1268_,
		_w1269_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		_w1242_,
		_w1257_,
		_w1270_
	);
	LUT2 #(
		.INIT('h4)
	) name1023 (
		_w1261_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w1239_,
		_w1242_,
		_w1272_
	);
	LUT2 #(
		.INIT('h4)
	) name1025 (
		_w1257_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h1)
	) name1026 (
		_w1271_,
		_w1273_,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		_w1239_,
		_w1242_,
		_w1275_
	);
	LUT2 #(
		.INIT('h4)
	) name1028 (
		_w1261_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h2)
	) name1029 (
		_w1261_,
		_w1275_,
		_w1277_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		_w1257_,
		_w1276_,
		_w1278_
	);
	LUT2 #(
		.INIT('h4)
	) name1031 (
		_w1277_,
		_w1278_,
		_w1279_
	);
	LUT2 #(
		.INIT('h2)
	) name1032 (
		_w1274_,
		_w1279_,
		_w1280_
	);
	LUT2 #(
		.INIT('h2)
	) name1033 (
		_w1269_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h8)
	) name1034 (
		_w1261_,
		_w1270_,
		_w1282_
	);
	LUT2 #(
		.INIT('h4)
	) name1035 (
		_w1239_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h1)
	) name1036 (
		_w1281_,
		_w1283_,
		_w1284_
	);
	LUT2 #(
		.INIT('h2)
	) name1037 (
		_w266_,
		_w484_,
		_w1285_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		_w266_,
		_w480_,
		_w1286_
	);
	LUT2 #(
		.INIT('h1)
	) name1039 (
		_w1285_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		decrypt_i_pad,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h2)
	) name1041 (
		_w266_,
		_w605_,
		_w1289_
	);
	LUT2 #(
		.INIT('h2)
	) name1042 (
		_w292_,
		_w733_,
		_w1290_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		_w515_,
		_w1289_,
		_w1291_
	);
	LUT2 #(
		.INIT('h4)
	) name1044 (
		_w1290_,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h2)
	) name1045 (
		decrypt_i_pad,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h1)
	) name1046 (
		_w1288_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h2)
	) name1047 (
		\rd1_R_o_reg[24]/NET0131 ,
		_w281_,
		_w1295_
	);
	LUT2 #(
		.INIT('h8)
	) name1048 (
		\data_i[63]_pad ,
		_w281_,
		_w1296_
	);
	LUT2 #(
		.INIT('h1)
	) name1049 (
		_w1295_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h4)
	) name1050 (
		_w1294_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('h2)
	) name1051 (
		_w1294_,
		_w1297_,
		_w1299_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w1298_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h1)
	) name1053 (
		_w1284_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h2)
	) name1054 (
		_w1242_,
		_w1261_,
		_w1302_
	);
	LUT2 #(
		.INIT('h2)
	) name1055 (
		_w1239_,
		_w1257_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name1056 (
		_w1302_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h4)
	) name1057 (
		_w1257_,
		_w1300_,
		_w1305_
	);
	LUT2 #(
		.INIT('h4)
	) name1058 (
		_w1242_,
		_w1261_,
		_w1306_
	);
	LUT2 #(
		.INIT('h1)
	) name1059 (
		_w1302_,
		_w1306_,
		_w1307_
	);
	LUT2 #(
		.INIT('h2)
	) name1060 (
		_w1305_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		_w1242_,
		_w1257_,
		_w1309_
	);
	LUT2 #(
		.INIT('h1)
	) name1062 (
		_w1275_,
		_w1300_,
		_w1310_
	);
	LUT2 #(
		.INIT('h1)
	) name1063 (
		_w1302_,
		_w1309_,
		_w1311_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		_w1310_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('h1)
	) name1065 (
		_w1304_,
		_w1308_,
		_w1313_
	);
	LUT2 #(
		.INIT('h4)
	) name1066 (
		_w1312_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h1)
	) name1067 (
		_w1269_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h8)
	) name1068 (
		_w1262_,
		_w1300_,
		_w1316_
	);
	LUT2 #(
		.INIT('h4)
	) name1069 (
		_w1239_,
		_w1261_,
		_w1317_
	);
	LUT2 #(
		.INIT('h8)
	) name1070 (
		_w1305_,
		_w1317_,
		_w1318_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		_w1242_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w1316_,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h2)
	) name1073 (
		_w1269_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h4)
	) name1074 (
		_w1239_,
		_w1257_,
		_w1322_
	);
	LUT2 #(
		.INIT('h8)
	) name1075 (
		_w1302_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w1317_,
		_w1322_,
		_w1324_
	);
	LUT2 #(
		.INIT('h1)
	) name1077 (
		_w1302_,
		_w1303_,
		_w1325_
	);
	LUT2 #(
		.INIT('h8)
	) name1078 (
		_w1324_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w1323_,
		_w1326_,
		_w1327_
	);
	LUT2 #(
		.INIT('h2)
	) name1080 (
		_w1300_,
		_w1327_,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w1263_,
		_w1321_,
		_w1329_
	);
	LUT2 #(
		.INIT('h4)
	) name1082 (
		_w1328_,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h4)
	) name1083 (
		_w1315_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h4)
	) name1084 (
		_w1301_,
		_w1331_,
		_w1332_
	);
	LUT2 #(
		.INIT('h4)
	) name1085 (
		\data_i[14]_pad ,
		_w281_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name1086 (
		\rd1_L_o_reg[30]/NET0131 ,
		_w281_,
		_w1334_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		_w1333_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h2)
	) name1088 (
		_w1332_,
		_w1335_,
		_w1336_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w1332_,
		_w1335_,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name1090 (
		_w1336_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h2)
	) name1091 (
		_w266_,
		_w1072_,
		_w1339_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w266_,
		_w925_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name1093 (
		_w1339_,
		_w1340_,
		_w1341_
	);
	LUT2 #(
		.INIT('h1)
	) name1094 (
		decrypt_i_pad,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h2)
	) name1095 (
		_w292_,
		_w758_,
		_w1343_
	);
	LUT2 #(
		.INIT('h1)
	) name1096 (
		_w716_,
		_w945_,
		_w1344_
	);
	LUT2 #(
		.INIT('h4)
	) name1097 (
		_w1343_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h2)
	) name1098 (
		decrypt_i_pad,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h1)
	) name1099 (
		_w1342_,
		_w1346_,
		_w1347_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w266_,
		_w1027_,
		_w1348_
	);
	LUT2 #(
		.INIT('h1)
	) name1101 (
		_w851_,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h1)
	) name1102 (
		decrypt_i_pad,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h4)
	) name1103 (
		_w284_,
		_w292_,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name1104 (
		_w290_,
		_w1056_,
		_w1352_
	);
	LUT2 #(
		.INIT('h4)
	) name1105 (
		_w1351_,
		_w1352_,
		_w1353_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		decrypt_i_pad,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h1)
	) name1107 (
		_w1350_,
		_w1354_,
		_w1355_
	);
	LUT2 #(
		.INIT('h4)
	) name1108 (
		_w901_,
		_w938_,
		_w1356_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		_w895_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h8)
	) name1110 (
		_w908_,
		_w993_,
		_w1358_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w992_,
		_w1358_,
		_w1359_
	);
	LUT2 #(
		.INIT('h4)
	) name1112 (
		_w895_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w941_,
		_w958_,
		_w1361_
	);
	LUT2 #(
		.INIT('h4)
	) name1114 (
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h1)
	) name1115 (
		_w1357_,
		_w1362_,
		_w1363_
	);
	LUT2 #(
		.INIT('h2)
	) name1116 (
		_w987_,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('h4)
	) name1117 (
		_w901_,
		_w936_,
		_w1365_
	);
	LUT2 #(
		.INIT('h8)
	) name1118 (
		_w895_,
		_w958_,
		_w1366_
	);
	LUT2 #(
		.INIT('h8)
	) name1119 (
		_w1365_,
		_w1366_,
		_w1367_
	);
	LUT2 #(
		.INIT('h2)
	) name1120 (
		_w908_,
		_w936_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name1121 (
		_w895_,
		_w1368_,
		_w1369_
	);
	LUT2 #(
		.INIT('h8)
	) name1122 (
		_w901_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h1)
	) name1123 (
		_w1367_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h2)
	) name1124 (
		_w908_,
		_w1371_,
		_w1372_
	);
	LUT2 #(
		.INIT('h2)
	) name1125 (
		_w937_,
		_w958_,
		_w1373_
	);
	LUT2 #(
		.INIT('h8)
	) name1126 (
		_w1008_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h1)
	) name1127 (
		_w961_,
		_w1368_,
		_w1375_
	);
	LUT2 #(
		.INIT('h4)
	) name1128 (
		_w958_,
		_w987_,
		_w1376_
	);
	LUT2 #(
		.INIT('h4)
	) name1129 (
		_w993_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h4)
	) name1130 (
		_w1375_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h8)
	) name1131 (
		_w902_,
		_w937_,
		_w1379_
	);
	LUT2 #(
		.INIT('h1)
	) name1132 (
		_w1004_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h4)
	) name1133 (
		_w1003_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h1)
	) name1134 (
		_w958_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h1)
	) name1135 (
		_w992_,
		_w1369_,
		_w1383_
	);
	LUT2 #(
		.INIT('h1)
	) name1136 (
		_w958_,
		_w1383_,
		_w1384_
	);
	LUT2 #(
		.INIT('h8)
	) name1137 (
		_w937_,
		_w961_,
		_w1385_
	);
	LUT2 #(
		.INIT('h1)
	) name1138 (
		_w1384_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h2)
	) name1139 (
		_w901_,
		_w908_,
		_w1387_
	);
	LUT2 #(
		.INIT('h2)
	) name1140 (
		_w958_,
		_w1387_,
		_w1388_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w938_,
		_w993_,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		_w1388_,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h8)
	) name1143 (
		_w901_,
		_w1004_,
		_w1391_
	);
	LUT2 #(
		.INIT('h1)
	) name1144 (
		_w1390_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h8)
	) name1145 (
		_w1386_,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w987_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h1)
	) name1147 (
		_w1374_,
		_w1378_,
		_w1395_
	);
	LUT2 #(
		.INIT('h4)
	) name1148 (
		_w1372_,
		_w1395_,
		_w1396_
	);
	LUT2 #(
		.INIT('h4)
	) name1149 (
		_w1382_,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h4)
	) name1150 (
		_w1364_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h4)
	) name1151 (
		_w1394_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		\data_i[12]_pad ,
		_w281_,
		_w1400_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		\rd1_L_o_reg[22]/NET0131 ,
		_w281_,
		_w1401_
	);
	LUT2 #(
		.INIT('h1)
	) name1154 (
		_w1400_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h2)
	) name1155 (
		_w1399_,
		_w1402_,
		_w1403_
	);
	LUT2 #(
		.INIT('h4)
	) name1156 (
		_w1399_,
		_w1402_,
		_w1404_
	);
	LUT2 #(
		.INIT('h1)
	) name1157 (
		_w1403_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h1)
	) name1158 (
		_w266_,
		_w546_,
		_w1406_
	);
	LUT2 #(
		.INIT('h1)
	) name1159 (
		_w285_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h1)
	) name1160 (
		decrypt_i_pad,
		_w1407_,
		_w1408_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		_w292_,
		_w310_,
		_w1409_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		_w413_,
		_w1054_,
		_w1410_
	);
	LUT2 #(
		.INIT('h4)
	) name1163 (
		_w1409_,
		_w1410_,
		_w1411_
	);
	LUT2 #(
		.INIT('h2)
	) name1164 (
		decrypt_i_pad,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h1)
	) name1165 (
		_w1408_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h2)
	) name1166 (
		_w780_,
		_w1413_,
		_w1414_
	);
	LUT2 #(
		.INIT('h4)
	) name1167 (
		_w780_,
		_w1413_,
		_w1415_
	);
	LUT2 #(
		.INIT('h1)
	) name1168 (
		_w1414_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h2)
	) name1169 (
		_w376_,
		_w411_,
		_w1417_
	);
	LUT2 #(
		.INIT('h4)
	) name1170 (
		_w376_,
		_w411_,
		_w1418_
	);
	LUT2 #(
		.INIT('h1)
	) name1171 (
		_w1417_,
		_w1418_,
		_w1419_
	);
	LUT2 #(
		.INIT('h2)
	) name1172 (
		_w1199_,
		_w1209_,
		_w1420_
	);
	LUT2 #(
		.INIT('h4)
	) name1173 (
		_w1199_,
		_w1209_,
		_w1421_
	);
	LUT2 #(
		.INIT('h1)
	) name1174 (
		_w1420_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h4)
	) name1175 (
		_w427_,
		_w688_,
		_w1423_
	);
	LUT2 #(
		.INIT('h2)
	) name1176 (
		_w427_,
		_w688_,
		_w1424_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		_w1423_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		_w1422_,
		_w1425_,
		_w1426_
	);
	LUT2 #(
		.INIT('h2)
	) name1179 (
		\rd1_R_o_reg[6]/NET0131 ,
		_w281_,
		_w1427_
	);
	LUT2 #(
		.INIT('h8)
	) name1180 (
		\data_i[9]_pad ,
		_w281_,
		_w1428_
	);
	LUT2 #(
		.INIT('h1)
	) name1181 (
		_w1427_,
		_w1428_,
		_w1429_
	);
	LUT2 #(
		.INIT('h4)
	) name1182 (
		_w663_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h2)
	) name1183 (
		_w663_,
		_w1429_,
		_w1431_
	);
	LUT2 #(
		.INIT('h1)
	) name1184 (
		_w1430_,
		_w1431_,
		_w1432_
	);
	LUT2 #(
		.INIT('h2)
	) name1185 (
		_w1426_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h8)
	) name1186 (
		_w1419_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h2)
	) name1187 (
		\rd1_R_o_reg[5]/NET0131 ,
		_w281_,
		_w1435_
	);
	LUT2 #(
		.INIT('h8)
	) name1188 (
		\data_i[17]_pad ,
		_w281_,
		_w1436_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		_w1435_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h4)
	) name1190 (
		_w1355_,
		_w1437_,
		_w1438_
	);
	LUT2 #(
		.INIT('h2)
	) name1191 (
		_w1355_,
		_w1437_,
		_w1439_
	);
	LUT2 #(
		.INIT('h1)
	) name1192 (
		_w1438_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h4)
	) name1193 (
		_w1422_,
		_w1432_,
		_w1441_
	);
	LUT2 #(
		.INIT('h2)
	) name1194 (
		_w1425_,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h8)
	) name1195 (
		_w1426_,
		_w1432_,
		_w1443_
	);
	LUT2 #(
		.INIT('h2)
	) name1196 (
		_w1440_,
		_w1442_,
		_w1444_
	);
	LUT2 #(
		.INIT('h4)
	) name1197 (
		_w1443_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h1)
	) name1198 (
		_w1434_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h1)
	) name1199 (
		_w1416_,
		_w1446_,
		_w1447_
	);
	LUT2 #(
		.INIT('h2)
	) name1200 (
		_w1422_,
		_w1432_,
		_w1448_
	);
	LUT2 #(
		.INIT('h4)
	) name1201 (
		_w1425_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h4)
	) name1202 (
		_w1419_,
		_w1440_,
		_w1450_
	);
	LUT2 #(
		.INIT('h8)
	) name1203 (
		_w1449_,
		_w1450_,
		_w1451_
	);
	LUT2 #(
		.INIT('h8)
	) name1204 (
		_w1422_,
		_w1432_,
		_w1452_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		_w1425_,
		_w1440_,
		_w1453_
	);
	LUT2 #(
		.INIT('h2)
	) name1206 (
		_w1425_,
		_w1440_,
		_w1454_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		_w1453_,
		_w1454_,
		_w1455_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		_w1450_,
		_w1452_,
		_w1456_
	);
	LUT2 #(
		.INIT('h4)
	) name1209 (
		_w1455_,
		_w1456_,
		_w1457_
	);
	LUT2 #(
		.INIT('h1)
	) name1210 (
		_w1422_,
		_w1432_,
		_w1458_
	);
	LUT2 #(
		.INIT('h8)
	) name1211 (
		_w1454_,
		_w1458_,
		_w1459_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w1416_,
		_w1419_,
		_w1460_
	);
	LUT2 #(
		.INIT('h8)
	) name1213 (
		_w1422_,
		_w1454_,
		_w1461_
	);
	LUT2 #(
		.INIT('h4)
	) name1214 (
		_w1440_,
		_w1443_,
		_w1462_
	);
	LUT2 #(
		.INIT('h1)
	) name1215 (
		_w1449_,
		_w1461_,
		_w1463_
	);
	LUT2 #(
		.INIT('h4)
	) name1216 (
		_w1462_,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h2)
	) name1217 (
		_w1460_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h4)
	) name1218 (
		_w1422_,
		_w1453_,
		_w1466_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		_w1432_,
		_w1466_,
		_w1467_
	);
	LUT2 #(
		.INIT('h2)
	) name1220 (
		_w1425_,
		_w1432_,
		_w1468_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		_w1440_,
		_w1468_,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		_w1426_,
		_w1469_,
		_w1470_
	);
	LUT2 #(
		.INIT('h1)
	) name1223 (
		_w1458_,
		_w1470_,
		_w1471_
	);
	LUT2 #(
		.INIT('h8)
	) name1224 (
		_w1422_,
		_w1425_,
		_w1472_
	);
	LUT2 #(
		.INIT('h1)
	) name1225 (
		_w1426_,
		_w1472_,
		_w1473_
	);
	LUT2 #(
		.INIT('h1)
	) name1226 (
		_w1440_,
		_w1452_,
		_w1474_
	);
	LUT2 #(
		.INIT('h8)
	) name1227 (
		_w1473_,
		_w1474_,
		_w1475_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		_w1471_,
		_w1475_,
		_w1476_
	);
	LUT2 #(
		.INIT('h2)
	) name1229 (
		_w1419_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h1)
	) name1230 (
		_w1441_,
		_w1448_,
		_w1478_
	);
	LUT2 #(
		.INIT('h1)
	) name1231 (
		_w1419_,
		_w1453_,
		_w1479_
	);
	LUT2 #(
		.INIT('h8)
	) name1232 (
		_w1478_,
		_w1479_,
		_w1480_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		_w1467_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h4)
	) name1234 (
		_w1477_,
		_w1481_,
		_w1482_
	);
	LUT2 #(
		.INIT('h2)
	) name1235 (
		_w1416_,
		_w1482_,
		_w1483_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w1451_,
		_w1459_,
		_w1484_
	);
	LUT2 #(
		.INIT('h4)
	) name1237 (
		_w1457_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		_w1465_,
		_w1485_,
		_w1486_
	);
	LUT2 #(
		.INIT('h4)
	) name1239 (
		_w1447_,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h4)
	) name1240 (
		_w1483_,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		\data_i[42]_pad ,
		_w281_,
		_w1489_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		\rd1_L_o_reg[10]/NET0131 ,
		_w281_,
		_w1490_
	);
	LUT2 #(
		.INIT('h1)
	) name1243 (
		_w1489_,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h2)
	) name1244 (
		_w1488_,
		_w1491_,
		_w1492_
	);
	LUT2 #(
		.INIT('h4)
	) name1245 (
		_w1488_,
		_w1491_,
		_w1493_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		_w1492_,
		_w1493_,
		_w1494_
	);
	LUT2 #(
		.INIT('h4)
	) name1247 (
		_w1419_,
		_w1467_,
		_w1495_
	);
	LUT2 #(
		.INIT('h8)
	) name1248 (
		_w1425_,
		_w1452_,
		_w1496_
	);
	LUT2 #(
		.INIT('h4)
	) name1249 (
		_w1422_,
		_w1469_,
		_w1497_
	);
	LUT2 #(
		.INIT('h2)
	) name1250 (
		_w1419_,
		_w1496_,
		_w1498_
	);
	LUT2 #(
		.INIT('h4)
	) name1251 (
		_w1497_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		_w1419_,
		_w1443_,
		_w1500_
	);
	LUT2 #(
		.INIT('h4)
	) name1253 (
		_w1459_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h1)
	) name1254 (
		_w1499_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		_w1419_,
		_w1432_,
		_w1503_
	);
	LUT2 #(
		.INIT('h2)
	) name1256 (
		_w1461_,
		_w1503_,
		_w1504_
	);
	LUT2 #(
		.INIT('h2)
	) name1257 (
		_w1450_,
		_w1458_,
		_w1505_
	);
	LUT2 #(
		.INIT('h4)
	) name1258 (
		_w1496_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h1)
	) name1259 (
		_w1467_,
		_w1504_,
		_w1507_
	);
	LUT2 #(
		.INIT('h4)
	) name1260 (
		_w1506_,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h4)
	) name1261 (
		_w1502_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h1)
	) name1262 (
		_w1416_,
		_w1509_,
		_w1510_
	);
	LUT2 #(
		.INIT('h8)
	) name1263 (
		_w1432_,
		_w1473_,
		_w1511_
	);
	LUT2 #(
		.INIT('h4)
	) name1264 (
		_w1450_,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h2)
	) name1265 (
		_w1419_,
		_w1440_,
		_w1513_
	);
	LUT2 #(
		.INIT('h4)
	) name1266 (
		_w1422_,
		_w1425_,
		_w1514_
	);
	LUT2 #(
		.INIT('h8)
	) name1267 (
		_w1513_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h1)
	) name1268 (
		_w1448_,
		_w1450_,
		_w1516_
	);
	LUT2 #(
		.INIT('h1)
	) name1269 (
		_w1513_,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h4)
	) name1270 (
		_w1506_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h1)
	) name1271 (
		_w1512_,
		_w1515_,
		_w1519_
	);
	LUT2 #(
		.INIT('h4)
	) name1272 (
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h2)
	) name1273 (
		_w1416_,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h1)
	) name1274 (
		_w1433_,
		_w1511_,
		_w1522_
	);
	LUT2 #(
		.INIT('h2)
	) name1275 (
		_w1513_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('h1)
	) name1276 (
		_w1495_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h4)
	) name1277 (
		_w1510_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h4)
	) name1278 (
		_w1521_,
		_w1525_,
		_w1526_
	);
	LUT2 #(
		.INIT('h4)
	) name1279 (
		\data_i[54]_pad ,
		_w281_,
		_w1527_
	);
	LUT2 #(
		.INIT('h1)
	) name1280 (
		\rd1_L_o_reg[25]/NET0131 ,
		_w281_,
		_w1528_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w1527_,
		_w1528_,
		_w1529_
	);
	LUT2 #(
		.INIT('h2)
	) name1282 (
		_w1526_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		_w1526_,
		_w1529_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		_w1530_,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h4)
	) name1285 (
		_w489_,
		_w492_,
		_w1533_
	);
	LUT2 #(
		.INIT('h2)
	) name1286 (
		_w489_,
		_w492_,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name1287 (
		_w1533_,
		_w1534_,
		_w1535_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		_w751_,
		_w766_,
		_w1536_
	);
	LUT2 #(
		.INIT('h4)
	) name1289 (
		_w751_,
		_w766_,
		_w1537_
	);
	LUT2 #(
		.INIT('h1)
	) name1290 (
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h2)
	) name1291 (
		_w250_,
		_w598_,
		_w1539_
	);
	LUT2 #(
		.INIT('h1)
	) name1292 (
		_w744_,
		_w1289_,
		_w1540_
	);
	LUT2 #(
		.INIT('h4)
	) name1293 (
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		decrypt_i_pad,
		_w1541_,
		_w1542_
	);
	LUT2 #(
		.INIT('h2)
	) name1295 (
		_w292_,
		_w1072_,
		_w1543_
	);
	LUT2 #(
		.INIT('h1)
	) name1296 (
		_w741_,
		_w946_,
		_w1544_
	);
	LUT2 #(
		.INIT('h4)
	) name1297 (
		_w1543_,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h2)
	) name1298 (
		decrypt_i_pad,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name1299 (
		_w1542_,
		_w1546_,
		_w1547_
	);
	LUT2 #(
		.INIT('h2)
	) name1300 (
		_w859_,
		_w1547_,
		_w1548_
	);
	LUT2 #(
		.INIT('h4)
	) name1301 (
		_w859_,
		_w1547_,
		_w1549_
	);
	LUT2 #(
		.INIT('h1)
	) name1302 (
		_w1548_,
		_w1549_,
		_w1550_
	);
	LUT2 #(
		.INIT('h2)
	) name1303 (
		_w1538_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h2)
	) name1304 (
		_w666_,
		_w1347_,
		_w1552_
	);
	LUT2 #(
		.INIT('h4)
	) name1305 (
		_w666_,
		_w1347_,
		_w1553_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h2)
	) name1307 (
		_w1551_,
		_w1554_,
		_w1555_
	);
	LUT2 #(
		.INIT('h4)
	) name1308 (
		_w1535_,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('h1)
	) name1309 (
		_w1535_,
		_w1538_,
		_w1557_
	);
	LUT2 #(
		.INIT('h4)
	) name1310 (
		_w1550_,
		_w1557_,
		_w1558_
	);
	LUT2 #(
		.INIT('h2)
	) name1311 (
		_w1550_,
		_w1554_,
		_w1559_
	);
	LUT2 #(
		.INIT('h8)
	) name1312 (
		_w1535_,
		_w1559_,
		_w1560_
	);
	LUT2 #(
		.INIT('h8)
	) name1313 (
		_w1550_,
		_w1554_,
		_w1561_
	);
	LUT2 #(
		.INIT('h4)
	) name1314 (
		_w1535_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h1)
	) name1315 (
		_w1560_,
		_w1562_,
		_w1563_
	);
	LUT2 #(
		.INIT('h2)
	) name1316 (
		_w1538_,
		_w1563_,
		_w1564_
	);
	LUT2 #(
		.INIT('h1)
	) name1317 (
		_w1558_,
		_w1564_,
		_w1565_
	);
	LUT2 #(
		.INIT('h4)
	) name1318 (
		_w709_,
		_w1063_,
		_w1566_
	);
	LUT2 #(
		.INIT('h2)
	) name1319 (
		_w709_,
		_w1063_,
		_w1567_
	);
	LUT2 #(
		.INIT('h1)
	) name1320 (
		_w1566_,
		_w1567_,
		_w1568_
	);
	LUT2 #(
		.INIT('h4)
	) name1321 (
		_w1565_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h8)
	) name1322 (
		_w1535_,
		_w1561_,
		_w1570_
	);
	LUT2 #(
		.INIT('h4)
	) name1323 (
		_w1535_,
		_w1559_,
		_w1571_
	);
	LUT2 #(
		.INIT('h1)
	) name1324 (
		_w1551_,
		_w1570_,
		_w1572_
	);
	LUT2 #(
		.INIT('h4)
	) name1325 (
		_w1571_,
		_w1572_,
		_w1573_
	);
	LUT2 #(
		.INIT('h1)
	) name1326 (
		_w1568_,
		_w1573_,
		_w1574_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w1556_,
		_w1574_,
		_w1575_
	);
	LUT2 #(
		.INIT('h4)
	) name1328 (
		_w1569_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h4)
	) name1329 (
		_w1041_,
		_w1254_,
		_w1577_
	);
	LUT2 #(
		.INIT('h2)
	) name1330 (
		_w1041_,
		_w1254_,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name1331 (
		_w1577_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h1)
	) name1332 (
		_w1576_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h4)
	) name1333 (
		_w1538_,
		_w1561_,
		_w1581_
	);
	LUT2 #(
		.INIT('h4)
	) name1334 (
		_w1550_,
		_w1554_,
		_w1582_
	);
	LUT2 #(
		.INIT('h8)
	) name1335 (
		_w1538_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h1)
	) name1336 (
		_w1581_,
		_w1583_,
		_w1584_
	);
	LUT2 #(
		.INIT('h8)
	) name1337 (
		_w1535_,
		_w1582_,
		_w1585_
	);
	LUT2 #(
		.INIT('h1)
	) name1338 (
		_w1535_,
		_w1559_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name1339 (
		_w1560_,
		_w1585_,
		_w1587_
	);
	LUT2 #(
		.INIT('h4)
	) name1340 (
		_w1586_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h2)
	) name1341 (
		_w1584_,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h2)
	) name1342 (
		_w1568_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h1)
	) name1343 (
		_w1550_,
		_w1554_,
		_w1591_
	);
	LUT2 #(
		.INIT('h2)
	) name1344 (
		_w1535_,
		_w1538_,
		_w1592_
	);
	LUT2 #(
		.INIT('h8)
	) name1345 (
		_w1591_,
		_w1592_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name1346 (
		_w1590_,
		_w1593_,
		_w1594_
	);
	LUT2 #(
		.INIT('h2)
	) name1347 (
		_w1579_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h8)
	) name1348 (
		_w1568_,
		_w1593_,
		_w1596_
	);
	LUT2 #(
		.INIT('h2)
	) name1349 (
		_w1535_,
		_w1550_,
		_w1597_
	);
	LUT2 #(
		.INIT('h1)
	) name1350 (
		_w1568_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h1)
	) name1351 (
		_w1538_,
		_w1561_,
		_w1599_
	);
	LUT2 #(
		.INIT('h2)
	) name1352 (
		_w1579_,
		_w1591_,
		_w1600_
	);
	LUT2 #(
		.INIT('h8)
	) name1353 (
		_w1598_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h8)
	) name1354 (
		_w1599_,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h2)
	) name1355 (
		_w1535_,
		_w1584_,
		_w1603_
	);
	LUT2 #(
		.INIT('h2)
	) name1356 (
		_w1556_,
		_w1568_,
		_w1604_
	);
	LUT2 #(
		.INIT('h1)
	) name1357 (
		_w1596_,
		_w1602_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name1358 (
		_w1603_,
		_w1604_,
		_w1606_
	);
	LUT2 #(
		.INIT('h8)
	) name1359 (
		_w1605_,
		_w1606_,
		_w1607_
	);
	LUT2 #(
		.INIT('h4)
	) name1360 (
		_w1580_,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h4)
	) name1361 (
		_w1595_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h4)
	) name1362 (
		\data_i[50]_pad ,
		_w281_,
		_w1610_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		\rd1_L_o_reg[9]/NET0131 ,
		_w281_,
		_w1611_
	);
	LUT2 #(
		.INIT('h1)
	) name1364 (
		_w1610_,
		_w1611_,
		_w1612_
	);
	LUT2 #(
		.INIT('h2)
	) name1365 (
		_w1609_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h4)
	) name1366 (
		_w1609_,
		_w1612_,
		_w1614_
	);
	LUT2 #(
		.INIT('h1)
	) name1367 (
		_w1613_,
		_w1614_,
		_w1615_
	);
	LUT2 #(
		.INIT('h4)
	) name1368 (
		_w1032_,
		_w1095_,
		_w1616_
	);
	LUT2 #(
		.INIT('h2)
	) name1369 (
		_w1032_,
		_w1095_,
		_w1617_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		_w1616_,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('h2)
	) name1371 (
		_w1155_,
		_w1218_,
		_w1619_
	);
	LUT2 #(
		.INIT('h4)
	) name1372 (
		_w1155_,
		_w1218_,
		_w1620_
	);
	LUT2 #(
		.INIT('h1)
	) name1373 (
		_w1619_,
		_w1620_,
		_w1621_
	);
	LUT2 #(
		.INIT('h4)
	) name1374 (
		_w1618_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h2)
	) name1375 (
		_w1618_,
		_w1621_,
		_w1623_
	);
	LUT2 #(
		.INIT('h1)
	) name1376 (
		_w1622_,
		_w1623_,
		_w1624_
	);
	LUT2 #(
		.INIT('h2)
	) name1377 (
		_w300_,
		_w335_,
		_w1625_
	);
	LUT2 #(
		.INIT('h4)
	) name1378 (
		_w300_,
		_w335_,
		_w1626_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		_w1625_,
		_w1626_,
		_w1627_
	);
	LUT2 #(
		.INIT('h8)
	) name1380 (
		_w1624_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h2)
	) name1381 (
		_w1621_,
		_w1627_,
		_w1629_
	);
	LUT2 #(
		.INIT('h2)
	) name1382 (
		\rd1_R_o_reg[9]/NET0131 ,
		_w281_,
		_w1630_
	);
	LUT2 #(
		.INIT('h8)
	) name1383 (
		\data_i[51]_pad ,
		_w281_,
		_w1631_
	);
	LUT2 #(
		.INIT('h1)
	) name1384 (
		_w1630_,
		_w1631_,
		_w1632_
	);
	LUT2 #(
		.INIT('h4)
	) name1385 (
		_w452_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h2)
	) name1386 (
		_w452_,
		_w1632_,
		_w1634_
	);
	LUT2 #(
		.INIT('h1)
	) name1387 (
		_w1633_,
		_w1634_,
		_w1635_
	);
	LUT2 #(
		.INIT('h4)
	) name1388 (
		_w1629_,
		_w1635_,
		_w1636_
	);
	LUT2 #(
		.INIT('h4)
	) name1389 (
		_w1628_,
		_w1636_,
		_w1637_
	);
	LUT2 #(
		.INIT('h4)
	) name1390 (
		_w534_,
		_w1199_,
		_w1638_
	);
	LUT2 #(
		.INIT('h2)
	) name1391 (
		_w534_,
		_w1199_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name1392 (
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT2 #(
		.INIT('h8)
	) name1393 (
		_w1618_,
		_w1627_,
		_w1641_
	);
	LUT2 #(
		.INIT('h4)
	) name1394 (
		_w1635_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h8)
	) name1395 (
		_w1621_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h1)
	) name1396 (
		_w1637_,
		_w1640_,
		_w1644_
	);
	LUT2 #(
		.INIT('h4)
	) name1397 (
		_w1643_,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h2)
	) name1398 (
		_w1621_,
		_w1635_,
		_w1646_
	);
	LUT2 #(
		.INIT('h2)
	) name1399 (
		_w1628_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h1)
	) name1400 (
		_w1618_,
		_w1627_,
		_w1648_
	);
	LUT2 #(
		.INIT('h1)
	) name1401 (
		_w1635_,
		_w1648_,
		_w1649_
	);
	LUT2 #(
		.INIT('h4)
	) name1402 (
		_w1641_,
		_w1649_,
		_w1650_
	);
	LUT2 #(
		.INIT('h2)
	) name1403 (
		_w1640_,
		_w1647_,
		_w1651_
	);
	LUT2 #(
		.INIT('h4)
	) name1404 (
		_w1650_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h1)
	) name1405 (
		_w1645_,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h2)
	) name1406 (
		_w1623_,
		_w1627_,
		_w1654_
	);
	LUT2 #(
		.INIT('h1)
	) name1407 (
		_w1653_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h2)
	) name1408 (
		_w688_,
		_w1225_,
		_w1656_
	);
	LUT2 #(
		.INIT('h4)
	) name1409 (
		_w688_,
		_w1225_,
		_w1657_
	);
	LUT2 #(
		.INIT('h1)
	) name1410 (
		_w1656_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h1)
	) name1411 (
		_w1655_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h8)
	) name1412 (
		_w1622_,
		_w1635_,
		_w1660_
	);
	LUT2 #(
		.INIT('h8)
	) name1413 (
		_w1623_,
		_w1627_,
		_w1661_
	);
	LUT2 #(
		.INIT('h1)
	) name1414 (
		_w1618_,
		_w1621_,
		_w1662_
	);
	LUT2 #(
		.INIT('h4)
	) name1415 (
		_w1627_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h1)
	) name1416 (
		_w1660_,
		_w1661_,
		_w1664_
	);
	LUT2 #(
		.INIT('h4)
	) name1417 (
		_w1663_,
		_w1664_,
		_w1665_
	);
	LUT2 #(
		.INIT('h4)
	) name1418 (
		_w1642_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h2)
	) name1419 (
		_w1640_,
		_w1666_,
		_w1667_
	);
	LUT2 #(
		.INIT('h8)
	) name1420 (
		_w1629_,
		_w1635_,
		_w1668_
	);
	LUT2 #(
		.INIT('h2)
	) name1421 (
		_w1640_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h8)
	) name1422 (
		_w1618_,
		_w1635_,
		_w1670_
	);
	LUT2 #(
		.INIT('h8)
	) name1423 (
		_w1621_,
		_w1670_,
		_w1671_
	);
	LUT2 #(
		.INIT('h8)
	) name1424 (
		_w1627_,
		_w1662_,
		_w1672_
	);
	LUT2 #(
		.INIT('h1)
	) name1425 (
		_w1629_,
		_w1672_,
		_w1673_
	);
	LUT2 #(
		.INIT('h4)
	) name1426 (
		_w1671_,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w1669_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name1428 (
		_w1667_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h2)
	) name1429 (
		_w1658_,
		_w1676_,
		_w1677_
	);
	LUT2 #(
		.INIT('h1)
	) name1430 (
		_w1627_,
		_w1635_,
		_w1678_
	);
	LUT2 #(
		.INIT('h4)
	) name1431 (
		_w1624_,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h4)
	) name1432 (
		_w1640_,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h4)
	) name1433 (
		_w1635_,
		_w1662_,
		_w1681_
	);
	LUT2 #(
		.INIT('h1)
	) name1434 (
		_w1660_,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w1627_,
		_w1682_,
		_w1683_
	);
	LUT2 #(
		.INIT('h8)
	) name1436 (
		_w1640_,
		_w1683_,
		_w1684_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		_w1680_,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h4)
	) name1438 (
		_w1677_,
		_w1685_,
		_w1686_
	);
	LUT2 #(
		.INIT('h4)
	) name1439 (
		_w1659_,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name1440 (
		\data_i[32]_pad ,
		_w281_,
		_w1688_
	);
	LUT2 #(
		.INIT('h1)
	) name1441 (
		\rd1_L_o_reg[3]/NET0131 ,
		_w281_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		_w1688_,
		_w1689_,
		_w1690_
	);
	LUT2 #(
		.INIT('h2)
	) name1443 (
		_w1687_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h4)
	) name1444 (
		_w1687_,
		_w1690_,
		_w1692_
	);
	LUT2 #(
		.INIT('h1)
	) name1445 (
		_w1691_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h4)
	) name1446 (
		_w1535_,
		_w1582_,
		_w1694_
	);
	LUT2 #(
		.INIT('h8)
	) name1447 (
		_w1538_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h4)
	) name1448 (
		_w1538_,
		_w1559_,
		_w1696_
	);
	LUT2 #(
		.INIT('h4)
	) name1449 (
		_w1554_,
		_w1557_,
		_w1697_
	);
	LUT2 #(
		.INIT('h8)
	) name1450 (
		_w1538_,
		_w1570_,
		_w1698_
	);
	LUT2 #(
		.INIT('h1)
	) name1451 (
		_w1696_,
		_w1697_,
		_w1699_
	);
	LUT2 #(
		.INIT('h4)
	) name1452 (
		_w1695_,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		_w1698_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		_w1568_,
		_w1701_,
		_w1702_
	);
	LUT2 #(
		.INIT('h2)
	) name1455 (
		_w1538_,
		_w1554_,
		_w1703_
	);
	LUT2 #(
		.INIT('h8)
	) name1456 (
		_w1597_,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h4)
	) name1457 (
		_w1538_,
		_w1582_,
		_w1705_
	);
	LUT2 #(
		.INIT('h8)
	) name1458 (
		_w1535_,
		_w1538_,
		_w1706_
	);
	LUT2 #(
		.INIT('h4)
	) name1459 (
		_w1554_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w1705_,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h2)
	) name1461 (
		_w1568_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h8)
	) name1462 (
		_w1550_,
		_w1557_,
		_w1710_
	);
	LUT2 #(
		.INIT('h1)
	) name1463 (
		_w1704_,
		_w1710_,
		_w1711_
	);
	LUT2 #(
		.INIT('h4)
	) name1464 (
		_w1709_,
		_w1711_,
		_w1712_
	);
	LUT2 #(
		.INIT('h4)
	) name1465 (
		_w1702_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('h1)
	) name1466 (
		_w1579_,
		_w1713_,
		_w1714_
	);
	LUT2 #(
		.INIT('h2)
	) name1467 (
		_w1538_,
		_w1559_,
		_w1715_
	);
	LUT2 #(
		.INIT('h4)
	) name1468 (
		_w1582_,
		_w1715_,
		_w1716_
	);
	LUT2 #(
		.INIT('h4)
	) name1469 (
		_w1535_,
		_w1716_,
		_w1717_
	);
	LUT2 #(
		.INIT('h8)
	) name1470 (
		_w1538_,
		_w1560_,
		_w1718_
	);
	LUT2 #(
		.INIT('h8)
	) name1471 (
		_w1554_,
		_w1592_,
		_w1719_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		_w1568_,
		_w1705_,
		_w1720_
	);
	LUT2 #(
		.INIT('h4)
	) name1473 (
		_w1719_,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('h4)
	) name1474 (
		_w1718_,
		_w1721_,
		_w1722_
	);
	LUT2 #(
		.INIT('h4)
	) name1475 (
		_w1554_,
		_w1592_,
		_w1723_
	);
	LUT2 #(
		.INIT('h2)
	) name1476 (
		_w1568_,
		_w1591_,
		_w1724_
	);
	LUT2 #(
		.INIT('h4)
	) name1477 (
		_w1597_,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h4)
	) name1478 (
		_w1723_,
		_w1725_,
		_w1726_
	);
	LUT2 #(
		.INIT('h1)
	) name1479 (
		_w1722_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h1)
	) name1480 (
		_w1717_,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h2)
	) name1481 (
		_w1579_,
		_w1728_,
		_w1729_
	);
	LUT2 #(
		.INIT('h8)
	) name1482 (
		_w1535_,
		_w1705_,
		_w1730_
	);
	LUT2 #(
		.INIT('h1)
	) name1483 (
		_w1555_,
		_w1562_,
		_w1731_
	);
	LUT2 #(
		.INIT('h2)
	) name1484 (
		_w1568_,
		_w1731_,
		_w1732_
	);
	LUT2 #(
		.INIT('h1)
	) name1485 (
		_w1535_,
		_w1568_,
		_w1733_
	);
	LUT2 #(
		.INIT('h8)
	) name1486 (
		_w1696_,
		_w1733_,
		_w1734_
	);
	LUT2 #(
		.INIT('h1)
	) name1487 (
		_w1730_,
		_w1734_,
		_w1735_
	);
	LUT2 #(
		.INIT('h4)
	) name1488 (
		_w1732_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h4)
	) name1489 (
		_w1714_,
		_w1736_,
		_w1737_
	);
	LUT2 #(
		.INIT('h4)
	) name1490 (
		_w1729_,
		_w1737_,
		_w1738_
	);
	LUT2 #(
		.INIT('h4)
	) name1491 (
		\data_i[48]_pad ,
		_w281_,
		_w1739_
	);
	LUT2 #(
		.INIT('h1)
	) name1492 (
		\rd1_L_o_reg[1]/NET0131 ,
		_w281_,
		_w1740_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		_w1739_,
		_w1740_,
		_w1741_
	);
	LUT2 #(
		.INIT('h2)
	) name1494 (
		_w1738_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h4)
	) name1495 (
		_w1738_,
		_w1741_,
		_w1743_
	);
	LUT2 #(
		.INIT('h1)
	) name1496 (
		_w1742_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h2)
	) name1497 (
		_w1105_,
		_w1109_,
		_w1745_
	);
	LUT2 #(
		.INIT('h2)
	) name1498 (
		_w1137_,
		_w1745_,
		_w1746_
	);
	LUT2 #(
		.INIT('h2)
	) name1499 (
		_w1109_,
		_w1126_,
		_w1747_
	);
	LUT2 #(
		.INIT('h4)
	) name1500 (
		_w1101_,
		_w1747_,
		_w1748_
	);
	LUT2 #(
		.INIT('h2)
	) name1501 (
		_w1126_,
		_w1138_,
		_w1749_
	);
	LUT2 #(
		.INIT('h1)
	) name1502 (
		_w1098_,
		_w1110_,
		_w1750_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		_w1748_,
		_w1749_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name1504 (
		_w1750_,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		_w1746_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		_w1126_,
		_w1129_,
		_w1754_
	);
	LUT2 #(
		.INIT('h1)
	) name1507 (
		_w1753_,
		_w1754_,
		_w1755_
	);
	LUT2 #(
		.INIT('h2)
	) name1508 (
		_w1158_,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h4)
	) name1509 (
		_w1098_,
		_w1180_,
		_w1757_
	);
	LUT2 #(
		.INIT('h4)
	) name1510 (
		_w1098_,
		_w1161_,
		_w1758_
	);
	LUT2 #(
		.INIT('h8)
	) name1511 (
		_w1106_,
		_w1747_,
		_w1759_
	);
	LUT2 #(
		.INIT('h1)
	) name1512 (
		_w1143_,
		_w1758_,
		_w1760_
	);
	LUT2 #(
		.INIT('h4)
	) name1513 (
		_w1759_,
		_w1760_,
		_w1761_
	);
	LUT2 #(
		.INIT('h1)
	) name1514 (
		_w1165_,
		_w1757_,
		_w1762_
	);
	LUT2 #(
		.INIT('h8)
	) name1515 (
		_w1761_,
		_w1762_,
		_w1763_
	);
	LUT2 #(
		.INIT('h1)
	) name1516 (
		_w1158_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h4)
	) name1517 (
		_w1098_,
		_w1185_,
		_w1765_
	);
	LUT2 #(
		.INIT('h8)
	) name1518 (
		_w1101_,
		_w1139_,
		_w1766_
	);
	LUT2 #(
		.INIT('h1)
	) name1519 (
		_w1168_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h1)
	) name1520 (
		_w1158_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h4)
	) name1521 (
		_w1109_,
		_w1766_,
		_w1769_
	);
	LUT2 #(
		.INIT('h1)
	) name1522 (
		_w1759_,
		_w1769_,
		_w1770_
	);
	LUT2 #(
		.INIT('h4)
	) name1523 (
		_w1768_,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h2)
	) name1524 (
		_w1098_,
		_w1771_,
		_w1772_
	);
	LUT2 #(
		.INIT('h1)
	) name1525 (
		_w1764_,
		_w1765_,
		_w1773_
	);
	LUT2 #(
		.INIT('h4)
	) name1526 (
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h4)
	) name1527 (
		_w1756_,
		_w1774_,
		_w1775_
	);
	LUT2 #(
		.INIT('h4)
	) name1528 (
		\data_i[22]_pad ,
		_w281_,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name1529 (
		\rd1_L_o_reg[29]/NET0131 ,
		_w281_,
		_w1777_
	);
	LUT2 #(
		.INIT('h1)
	) name1530 (
		_w1776_,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h2)
	) name1531 (
		_w1775_,
		_w1778_,
		_w1779_
	);
	LUT2 #(
		.INIT('h4)
	) name1532 (
		_w1775_,
		_w1778_,
		_w1780_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		_w1779_,
		_w1780_,
		_w1781_
	);
	LUT2 #(
		.INIT('h1)
	) name1534 (
		_w1419_,
		_w1440_,
		_w1782_
	);
	LUT2 #(
		.INIT('h1)
	) name1535 (
		_w1454_,
		_w1782_,
		_w1783_
	);
	LUT2 #(
		.INIT('h2)
	) name1536 (
		_w1441_,
		_w1783_,
		_w1784_
	);
	LUT2 #(
		.INIT('h2)
	) name1537 (
		_w1419_,
		_w1448_,
		_w1785_
	);
	LUT2 #(
		.INIT('h1)
	) name1538 (
		_w1425_,
		_w1440_,
		_w1786_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		_w1514_,
		_w1786_,
		_w1787_
	);
	LUT2 #(
		.INIT('h8)
	) name1540 (
		_w1785_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h1)
	) name1541 (
		_w1416_,
		_w1788_,
		_w1789_
	);
	LUT2 #(
		.INIT('h8)
	) name1542 (
		_w1425_,
		_w1478_,
		_w1790_
	);
	LUT2 #(
		.INIT('h1)
	) name1543 (
		_w1449_,
		_w1453_,
		_w1791_
	);
	LUT2 #(
		.INIT('h4)
	) name1544 (
		_w1790_,
		_w1791_,
		_w1792_
	);
	LUT2 #(
		.INIT('h2)
	) name1545 (
		_w1789_,
		_w1792_,
		_w1793_
	);
	LUT2 #(
		.INIT('h2)
	) name1546 (
		_w1454_,
		_w1785_,
		_w1794_
	);
	LUT2 #(
		.INIT('h2)
	) name1547 (
		_w1416_,
		_w1467_,
		_w1795_
	);
	LUT2 #(
		.INIT('h4)
	) name1548 (
		_w1794_,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('h2)
	) name1549 (
		_w1422_,
		_w1468_,
		_w1797_
	);
	LUT2 #(
		.INIT('h4)
	) name1550 (
		_w1786_,
		_w1797_,
		_w1798_
	);
	LUT2 #(
		.INIT('h2)
	) name1551 (
		_w1796_,
		_w1798_,
		_w1799_
	);
	LUT2 #(
		.INIT('h1)
	) name1552 (
		_w1419_,
		_w1793_,
		_w1800_
	);
	LUT2 #(
		.INIT('h4)
	) name1553 (
		_w1799_,
		_w1800_,
		_w1801_
	);
	LUT2 #(
		.INIT('h4)
	) name1554 (
		_w1475_,
		_w1789_,
		_w1802_
	);
	LUT2 #(
		.INIT('h8)
	) name1555 (
		_w1478_,
		_w1786_,
		_w1803_
	);
	LUT2 #(
		.INIT('h1)
	) name1556 (
		_w1469_,
		_w1803_,
		_w1804_
	);
	LUT2 #(
		.INIT('h8)
	) name1557 (
		_w1796_,
		_w1804_,
		_w1805_
	);
	LUT2 #(
		.INIT('h2)
	) name1558 (
		_w1419_,
		_w1802_,
		_w1806_
	);
	LUT2 #(
		.INIT('h4)
	) name1559 (
		_w1805_,
		_w1806_,
		_w1807_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w1451_,
		_w1784_,
		_w1808_
	);
	LUT2 #(
		.INIT('h4)
	) name1561 (
		_w1801_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h4)
	) name1562 (
		_w1807_,
		_w1809_,
		_w1810_
	);
	LUT2 #(
		.INIT('h4)
	) name1563 (
		\data_i[56]_pad ,
		_w281_,
		_w1811_
	);
	LUT2 #(
		.INIT('h1)
	) name1564 (
		\rd1_L_o_reg[0]/NET0131 ,
		_w281_,
		_w1812_
	);
	LUT2 #(
		.INIT('h1)
	) name1565 (
		_w1811_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h2)
	) name1566 (
		_w1810_,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h4)
	) name1567 (
		_w1810_,
		_w1813_,
		_w1815_
	);
	LUT2 #(
		.INIT('h1)
	) name1568 (
		_w1814_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h4)
	) name1569 (
		_w1126_,
		_w1129_,
		_w1817_
	);
	LUT2 #(
		.INIT('h2)
	) name1570 (
		_w1098_,
		_w1147_,
		_w1818_
	);
	LUT2 #(
		.INIT('h4)
	) name1571 (
		_w1817_,
		_w1818_,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1572 (
		_w1104_,
		_w1160_,
		_w1820_
	);
	LUT2 #(
		.INIT('h1)
	) name1573 (
		_w1098_,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('h4)
	) name1574 (
		_w1759_,
		_w1821_,
		_w1822_
	);
	LUT2 #(
		.INIT('h1)
	) name1575 (
		_w1819_,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h1)
	) name1576 (
		_w1110_,
		_w1138_,
		_w1824_
	);
	LUT2 #(
		.INIT('h2)
	) name1577 (
		_w1126_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h1)
	) name1578 (
		_w1158_,
		_w1765_,
		_w1826_
	);
	LUT2 #(
		.INIT('h4)
	) name1579 (
		_w1825_,
		_w1826_,
		_w1827_
	);
	LUT2 #(
		.INIT('h4)
	) name1580 (
		_w1823_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h8)
	) name1581 (
		_w1098_,
		_w1185_,
		_w1829_
	);
	LUT2 #(
		.INIT('h1)
	) name1582 (
		_w1142_,
		_w1172_,
		_w1830_
	);
	LUT2 #(
		.INIT('h2)
	) name1583 (
		_w1106_,
		_w1830_,
		_w1831_
	);
	LUT2 #(
		.INIT('h4)
	) name1584 (
		_w1139_,
		_w1758_,
		_w1832_
	);
	LUT2 #(
		.INIT('h2)
	) name1585 (
		_w1158_,
		_w1169_,
		_w1833_
	);
	LUT2 #(
		.INIT('h1)
	) name1586 (
		_w1757_,
		_w1829_,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name1587 (
		_w1831_,
		_w1832_,
		_w1835_
	);
	LUT2 #(
		.INIT('h8)
	) name1588 (
		_w1834_,
		_w1835_,
		_w1836_
	);
	LUT2 #(
		.INIT('h8)
	) name1589 (
		_w1833_,
		_w1836_,
		_w1837_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w1828_,
		_w1837_,
		_w1838_
	);
	LUT2 #(
		.INIT('h2)
	) name1591 (
		_w1098_,
		_w1164_,
		_w1839_
	);
	LUT2 #(
		.INIT('h4)
	) name1592 (
		_w1101_,
		_w1135_,
		_w1840_
	);
	LUT2 #(
		.INIT('h1)
	) name1593 (
		_w1098_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h4)
	) name1594 (
		_w1754_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h4)
	) name1595 (
		_w1769_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h1)
	) name1596 (
		_w1839_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('h1)
	) name1597 (
		_w1838_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h4)
	) name1598 (
		\data_i[62]_pad ,
		_w281_,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name1599 (
		\rd1_L_o_reg[24]/NET0131 ,
		_w281_,
		_w1847_
	);
	LUT2 #(
		.INIT('h1)
	) name1600 (
		_w1846_,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h2)
	) name1601 (
		_w1845_,
		_w1848_,
		_w1849_
	);
	LUT2 #(
		.INIT('h4)
	) name1602 (
		_w1845_,
		_w1848_,
		_w1850_
	);
	LUT2 #(
		.INIT('h1)
	) name1603 (
		_w1849_,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h1)
	) name1604 (
		_w266_,
		_w622_,
		_w1852_
	);
	LUT2 #(
		.INIT('h1)
	) name1605 (
		_w562_,
		_w1852_,
		_w1853_
	);
	LUT2 #(
		.INIT('h1)
	) name1606 (
		decrypt_i_pad,
		_w1853_,
		_w1854_
	);
	LUT2 #(
		.INIT('h2)
	) name1607 (
		_w292_,
		_w704_,
		_w1855_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w972_,
		_w1244_,
		_w1856_
	);
	LUT2 #(
		.INIT('h4)
	) name1609 (
		_w1855_,
		_w1856_,
		_w1857_
	);
	LUT2 #(
		.INIT('h2)
	) name1610 (
		decrypt_i_pad,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h1)
	) name1611 (
		_w1854_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h2)
	) name1612 (
		\rd1_R_o_reg[21]/NET0131 ,
		_w281_,
		_w1860_
	);
	LUT2 #(
		.INIT('h8)
	) name1613 (
		\data_i[21]_pad ,
		_w281_,
		_w1861_
	);
	LUT2 #(
		.INIT('h1)
	) name1614 (
		_w1860_,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h4)
	) name1615 (
		_w1859_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('h2)
	) name1616 (
		_w1859_,
		_w1862_,
		_w1864_
	);
	LUT2 #(
		.INIT('h1)
	) name1617 (
		_w1863_,
		_w1864_,
		_w1865_
	);
	LUT2 #(
		.INIT('h4)
	) name1618 (
		_w470_,
		_w933_,
		_w1866_
	);
	LUT2 #(
		.INIT('h2)
	) name1619 (
		_w470_,
		_w933_,
		_w1867_
	);
	LUT2 #(
		.INIT('h1)
	) name1620 (
		_w1866_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h4)
	) name1621 (
		_w1865_,
		_w1868_,
		_w1869_
	);
	LUT2 #(
		.INIT('h4)
	) name1622 (
		_w522_,
		_w1297_,
		_w1870_
	);
	LUT2 #(
		.INIT('h2)
	) name1623 (
		_w522_,
		_w1297_,
		_w1871_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		_w1870_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h1)
	) name1625 (
		_w266_,
		_w758_,
		_w1873_
	);
	LUT2 #(
		.INIT('h1)
	) name1626 (
		_w919_,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h1)
	) name1627 (
		decrypt_i_pad,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h2)
	) name1628 (
		_w292_,
		_w722_,
		_w1876_
	);
	LUT2 #(
		.INIT('h1)
	) name1629 (
		_w580_,
		_w714_,
		_w1877_
	);
	LUT2 #(
		.INIT('h4)
	) name1630 (
		_w1876_,
		_w1877_,
		_w1878_
	);
	LUT2 #(
		.INIT('h2)
	) name1631 (
		decrypt_i_pad,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('h1)
	) name1632 (
		_w1875_,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		\rd1_R_o_reg[22]/NET0131 ,
		_w281_,
		_w1881_
	);
	LUT2 #(
		.INIT('h8)
	) name1634 (
		\data_i[13]_pad ,
		_w281_,
		_w1882_
	);
	LUT2 #(
		.INIT('h1)
	) name1635 (
		_w1881_,
		_w1882_,
		_w1883_
	);
	LUT2 #(
		.INIT('h4)
	) name1636 (
		_w1880_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h2)
	) name1637 (
		_w1880_,
		_w1883_,
		_w1885_
	);
	LUT2 #(
		.INIT('h1)
	) name1638 (
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h8)
	) name1639 (
		_w1872_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h4)
	) name1640 (
		_w748_,
		_w1266_,
		_w1888_
	);
	LUT2 #(
		.INIT('h2)
	) name1641 (
		_w748_,
		_w1266_,
		_w1889_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		_w1888_,
		_w1889_,
		_w1890_
	);
	LUT2 #(
		.INIT('h2)
	) name1643 (
		_w1872_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('h4)
	) name1644 (
		_w1872_,
		_w1890_,
		_w1892_
	);
	LUT2 #(
		.INIT('h1)
	) name1645 (
		_w1891_,
		_w1892_,
		_w1893_
	);
	LUT2 #(
		.INIT('h4)
	) name1646 (
		_w1886_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('h1)
	) name1647 (
		_w1887_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h2)
	) name1648 (
		_w1869_,
		_w1895_,
		_w1896_
	);
	LUT2 #(
		.INIT('h1)
	) name1649 (
		_w1865_,
		_w1886_,
		_w1897_
	);
	LUT2 #(
		.INIT('h8)
	) name1650 (
		_w1865_,
		_w1886_,
		_w1898_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		_w1897_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h1)
	) name1652 (
		_w1891_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h2)
	) name1653 (
		_w1872_,
		_w1897_,
		_w1901_
	);
	LUT2 #(
		.INIT('h1)
	) name1654 (
		_w1868_,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h4)
	) name1655 (
		_w1900_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h4)
	) name1656 (
		_w585_,
		_w905_,
		_w1904_
	);
	LUT2 #(
		.INIT('h2)
	) name1657 (
		_w585_,
		_w905_,
		_w1905_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		_w1904_,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		_w1865_,
		_w1872_,
		_w1907_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		_w1890_,
		_w1907_,
		_w1908_
	);
	LUT2 #(
		.INIT('h4)
	) name1661 (
		_w1886_,
		_w1908_,
		_w1909_
	);
	LUT2 #(
		.INIT('h8)
	) name1662 (
		_w1886_,
		_w1907_,
		_w1910_
	);
	LUT2 #(
		.INIT('h8)
	) name1663 (
		_w1868_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h2)
	) name1664 (
		_w1906_,
		_w1909_,
		_w1912_
	);
	LUT2 #(
		.INIT('h4)
	) name1665 (
		_w1911_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h4)
	) name1666 (
		_w1903_,
		_w1913_,
		_w1914_
	);
	LUT2 #(
		.INIT('h4)
	) name1667 (
		_w1896_,
		_w1914_,
		_w1915_
	);
	LUT2 #(
		.INIT('h2)
	) name1668 (
		_w1865_,
		_w1890_,
		_w1916_
	);
	LUT2 #(
		.INIT('h4)
	) name1669 (
		_w1886_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h8)
	) name1670 (
		_w1872_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name1671 (
		_w1872_,
		_w1886_,
		_w1919_
	);
	LUT2 #(
		.INIT('h1)
	) name1672 (
		_w1887_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h1)
	) name1673 (
		_w1890_,
		_w1907_,
		_w1921_
	);
	LUT2 #(
		.INIT('h4)
	) name1674 (
		_w1920_,
		_w1921_,
		_w1922_
	);
	LUT2 #(
		.INIT('h8)
	) name1675 (
		_w1872_,
		_w1890_,
		_w1923_
	);
	LUT2 #(
		.INIT('h4)
	) name1676 (
		_w1865_,
		_w1923_,
		_w1924_
	);
	LUT2 #(
		.INIT('h1)
	) name1677 (
		_w1910_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h4)
	) name1678 (
		_w1922_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h1)
	) name1679 (
		_w1868_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h1)
	) name1680 (
		_w1906_,
		_w1918_,
		_w1928_
	);
	LUT2 #(
		.INIT('h4)
	) name1681 (
		_w1927_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		_w1915_,
		_w1929_,
		_w1930_
	);
	LUT2 #(
		.INIT('h2)
	) name1683 (
		_w1906_,
		_w1918_,
		_w1931_
	);
	LUT2 #(
		.INIT('h4)
	) name1684 (
		_w1865_,
		_w1892_,
		_w1932_
	);
	LUT2 #(
		.INIT('h1)
	) name1685 (
		_w1907_,
		_w1923_,
		_w1933_
	);
	LUT2 #(
		.INIT('h8)
	) name1686 (
		_w1920_,
		_w1933_,
		_w1934_
	);
	LUT2 #(
		.INIT('h1)
	) name1687 (
		_w1917_,
		_w1932_,
		_w1935_
	);
	LUT2 #(
		.INIT('h4)
	) name1688 (
		_w1934_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		_w1931_,
		_w1936_,
		_w1937_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		_w1898_,
		_w1923_,
		_w1938_
	);
	LUT2 #(
		.INIT('h2)
	) name1691 (
		_w1868_,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h4)
	) name1692 (
		_w1937_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h4)
	) name1693 (
		_w1865_,
		_w1890_,
		_w1941_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w1916_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h2)
	) name1695 (
		_w1887_,
		_w1942_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w1868_,
		_w1909_,
		_w1944_
	);
	LUT2 #(
		.INIT('h4)
	) name1697 (
		_w1943_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h1)
	) name1698 (
		_w1940_,
		_w1945_,
		_w1946_
	);
	LUT2 #(
		.INIT('h1)
	) name1699 (
		_w1930_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h4)
	) name1700 (
		\data_i[58]_pad ,
		_w281_,
		_w1948_
	);
	LUT2 #(
		.INIT('h1)
	) name1701 (
		\rd1_L_o_reg[8]/NET0131 ,
		_w281_,
		_w1949_
	);
	LUT2 #(
		.INIT('h1)
	) name1702 (
		_w1948_,
		_w1949_,
		_w1950_
	);
	LUT2 #(
		.INIT('h2)
	) name1703 (
		_w1947_,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('h4)
	) name1704 (
		_w1947_,
		_w1950_,
		_w1952_
	);
	LUT2 #(
		.INIT('h1)
	) name1705 (
		_w1951_,
		_w1952_,
		_w1953_
	);
	LUT2 #(
		.INIT('h2)
	) name1706 (
		_w1239_,
		_w1300_,
		_w1954_
	);
	LUT2 #(
		.INIT('h4)
	) name1707 (
		_w1257_,
		_w1307_,
		_w1955_
	);
	LUT2 #(
		.INIT('h8)
	) name1708 (
		_w1954_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w1239_,
		_w1257_,
		_w1957_
	);
	LUT2 #(
		.INIT('h8)
	) name1710 (
		_w1302_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h8)
	) name1711 (
		_w1239_,
		_w1261_,
		_w1959_
	);
	LUT2 #(
		.INIT('h1)
	) name1712 (
		_w1258_,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		_w1263_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('h1)
	) name1714 (
		_w1300_,
		_w1958_,
		_w1962_
	);
	LUT2 #(
		.INIT('h4)
	) name1715 (
		_w1961_,
		_w1962_,
		_w1963_
	);
	LUT2 #(
		.INIT('h4)
	) name1716 (
		_w1262_,
		_w1300_,
		_w1964_
	);
	LUT2 #(
		.INIT('h4)
	) name1717 (
		_w1276_,
		_w1964_,
		_w1965_
	);
	LUT2 #(
		.INIT('h8)
	) name1718 (
		_w1274_,
		_w1965_,
		_w1966_
	);
	LUT2 #(
		.INIT('h1)
	) name1719 (
		_w1963_,
		_w1966_,
		_w1967_
	);
	LUT2 #(
		.INIT('h2)
	) name1720 (
		_w1269_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h2)
	) name1721 (
		_w1282_,
		_w1954_,
		_w1969_
	);
	LUT2 #(
		.INIT('h4)
	) name1722 (
		_w1261_,
		_w1303_,
		_w1970_
	);
	LUT2 #(
		.INIT('h1)
	) name1723 (
		_w1300_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h2)
	) name1724 (
		_w1261_,
		_w1309_,
		_w1972_
	);
	LUT2 #(
		.INIT('h1)
	) name1725 (
		_w1324_,
		_w1972_,
		_w1973_
	);
	LUT2 #(
		.INIT('h4)
	) name1726 (
		_w1263_,
		_w1971_,
		_w1974_
	);
	LUT2 #(
		.INIT('h4)
	) name1727 (
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h2)
	) name1728 (
		_w1258_,
		_w1261_,
		_w1976_
	);
	LUT2 #(
		.INIT('h1)
	) name1729 (
		_w1257_,
		_w1272_,
		_w1977_
	);
	LUT2 #(
		.INIT('h4)
	) name1730 (
		_w1275_,
		_w1977_,
		_w1978_
	);
	LUT2 #(
		.INIT('h2)
	) name1731 (
		_w1300_,
		_w1976_,
		_w1979_
	);
	LUT2 #(
		.INIT('h4)
	) name1732 (
		_w1978_,
		_w1979_,
		_w1980_
	);
	LUT2 #(
		.INIT('h1)
	) name1733 (
		_w1975_,
		_w1980_,
		_w1981_
	);
	LUT2 #(
		.INIT('h1)
	) name1734 (
		_w1269_,
		_w1969_,
		_w1982_
	);
	LUT2 #(
		.INIT('h4)
	) name1735 (
		_w1981_,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('h1)
	) name1736 (
		_w1968_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h1)
	) name1737 (
		_w1319_,
		_w1956_,
		_w1985_
	);
	LUT2 #(
		.INIT('h4)
	) name1738 (
		_w1984_,
		_w1985_,
		_w1986_
	);
	LUT2 #(
		.INIT('h4)
	) name1739 (
		\data_i[36]_pad ,
		_w281_,
		_w1987_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		\rd1_L_o_reg[19]/NET0131 ,
		_w281_,
		_w1988_
	);
	LUT2 #(
		.INIT('h1)
	) name1741 (
		_w1987_,
		_w1988_,
		_w1989_
	);
	LUT2 #(
		.INIT('h2)
	) name1742 (
		_w1986_,
		_w1989_,
		_w1990_
	);
	LUT2 #(
		.INIT('h4)
	) name1743 (
		_w1986_,
		_w1989_,
		_w1991_
	);
	LUT2 #(
		.INIT('h1)
	) name1744 (
		_w1990_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h8)
	) name1745 (
		_w1635_,
		_w1641_,
		_w1993_
	);
	LUT2 #(
		.INIT('h1)
	) name1746 (
		_w1671_,
		_w1679_,
		_w1994_
	);
	LUT2 #(
		.INIT('h2)
	) name1747 (
		_w1640_,
		_w1994_,
		_w1995_
	);
	LUT2 #(
		.INIT('h8)
	) name1748 (
		_w1635_,
		_w1662_,
		_w1996_
	);
	LUT2 #(
		.INIT('h1)
	) name1749 (
		_w1661_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h1)
	) name1750 (
		_w1640_,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h8)
	) name1751 (
		_w1635_,
		_w1663_,
		_w1999_
	);
	LUT2 #(
		.INIT('h1)
	) name1752 (
		_w1993_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h4)
	) name1753 (
		_w1998_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h4)
	) name1754 (
		_w1995_,
		_w2001_,
		_w2002_
	);
	LUT2 #(
		.INIT('h2)
	) name1755 (
		_w1658_,
		_w2002_,
		_w2003_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		_w1618_,
		_w1629_,
		_w2004_
	);
	LUT2 #(
		.INIT('h4)
	) name1757 (
		_w1635_,
		_w2004_,
		_w2005_
	);
	LUT2 #(
		.INIT('h1)
	) name1758 (
		_w1648_,
		_w1661_,
		_w2006_
	);
	LUT2 #(
		.INIT('h2)
	) name1759 (
		_w1635_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h8)
	) name1760 (
		_w1622_,
		_w1627_,
		_w2008_
	);
	LUT2 #(
		.INIT('h4)
	) name1761 (
		_w1635_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h1)
	) name1762 (
		_w2005_,
		_w2009_,
		_w2010_
	);
	LUT2 #(
		.INIT('h4)
	) name1763 (
		_w2007_,
		_w2010_,
		_w2011_
	);
	LUT2 #(
		.INIT('h1)
	) name1764 (
		_w1640_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		_w1627_,
		_w1640_,
		_w2013_
	);
	LUT2 #(
		.INIT('h4)
	) name1766 (
		_w1682_,
		_w2013_,
		_w2014_
	);
	LUT2 #(
		.INIT('h4)
	) name1767 (
		_w1627_,
		_w1670_,
		_w2015_
	);
	LUT2 #(
		.INIT('h4)
	) name1768 (
		_w1621_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h2)
	) name1769 (
		_w1640_,
		_w1642_,
		_w2017_
	);
	LUT2 #(
		.INIT('h4)
	) name1770 (
		_w2016_,
		_w2017_,
		_w2018_
	);
	LUT2 #(
		.INIT('h8)
	) name1771 (
		_w1618_,
		_w1678_,
		_w2019_
	);
	LUT2 #(
		.INIT('h1)
	) name1772 (
		_w1640_,
		_w2004_,
		_w2020_
	);
	LUT2 #(
		.INIT('h4)
	) name1773 (
		_w2019_,
		_w2020_,
		_w2021_
	);
	LUT2 #(
		.INIT('h1)
	) name1774 (
		_w2018_,
		_w2021_,
		_w2022_
	);
	LUT2 #(
		.INIT('h1)
	) name1775 (
		_w1683_,
		_w2005_,
		_w2023_
	);
	LUT2 #(
		.INIT('h4)
	) name1776 (
		_w2022_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h1)
	) name1777 (
		_w1658_,
		_w2024_,
		_w2025_
	);
	LUT2 #(
		.INIT('h1)
	) name1778 (
		_w2003_,
		_w2014_,
		_w2026_
	);
	LUT2 #(
		.INIT('h4)
	) name1779 (
		_w2012_,
		_w2026_,
		_w2027_
	);
	LUT2 #(
		.INIT('h4)
	) name1780 (
		_w2025_,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h4)
	) name1781 (
		\data_i[20]_pad ,
		_w281_,
		_w2029_
	);
	LUT2 #(
		.INIT('h1)
	) name1782 (
		\rd1_L_o_reg[21]/NET0131 ,
		_w281_,
		_w2030_
	);
	LUT2 #(
		.INIT('h1)
	) name1783 (
		_w2029_,
		_w2030_,
		_w2031_
	);
	LUT2 #(
		.INIT('h2)
	) name1784 (
		_w2028_,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h4)
	) name1785 (
		_w2028_,
		_w2031_,
		_w2033_
	);
	LUT2 #(
		.INIT('h1)
	) name1786 (
		_w2032_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h1)
	) name1787 (
		_w895_,
		_w995_,
		_w2035_
	);
	LUT2 #(
		.INIT('h8)
	) name1788 (
		_w895_,
		_w901_,
		_w2036_
	);
	LUT2 #(
		.INIT('h4)
	) name1789 (
		_w936_,
		_w2036_,
		_w2037_
	);
	LUT2 #(
		.INIT('h1)
	) name1790 (
		_w1356_,
		_w2037_,
		_w2038_
	);
	LUT2 #(
		.INIT('h1)
	) name1791 (
		_w987_,
		_w2038_,
		_w2039_
	);
	LUT2 #(
		.INIT('h2)
	) name1792 (
		_w941_,
		_w1387_,
		_w2040_
	);
	LUT2 #(
		.INIT('h1)
	) name1793 (
		_w2035_,
		_w2039_,
		_w2041_
	);
	LUT2 #(
		.INIT('h4)
	) name1794 (
		_w2040_,
		_w2041_,
		_w2042_
	);
	LUT2 #(
		.INIT('h2)
	) name1795 (
		_w958_,
		_w2042_,
		_w2043_
	);
	LUT2 #(
		.INIT('h8)
	) name1796 (
		_w908_,
		_w989_,
		_w2044_
	);
	LUT2 #(
		.INIT('h2)
	) name1797 (
		_w895_,
		_w960_,
		_w2045_
	);
	LUT2 #(
		.INIT('h1)
	) name1798 (
		_w942_,
		_w1004_,
		_w2046_
	);
	LUT2 #(
		.INIT('h1)
	) name1799 (
		_w958_,
		_w2045_,
		_w2047_
	);
	LUT2 #(
		.INIT('h8)
	) name1800 (
		_w2046_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h1)
	) name1801 (
		_w987_,
		_w1374_,
		_w2049_
	);
	LUT2 #(
		.INIT('h4)
	) name1802 (
		_w2044_,
		_w2049_,
		_w2050_
	);
	LUT2 #(
		.INIT('h4)
	) name1803 (
		_w2048_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h2)
	) name1804 (
		_w895_,
		_w1359_,
		_w2052_
	);
	LUT2 #(
		.INIT('h1)
	) name1805 (
		_w1010_,
		_w1356_,
		_w2053_
	);
	LUT2 #(
		.INIT('h1)
	) name1806 (
		_w958_,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('h2)
	) name1807 (
		_w987_,
		_w1006_,
		_w2055_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w2052_,
		_w2054_,
		_w2056_
	);
	LUT2 #(
		.INIT('h8)
	) name1809 (
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT2 #(
		.INIT('h1)
	) name1810 (
		_w2051_,
		_w2057_,
		_w2058_
	);
	LUT2 #(
		.INIT('h4)
	) name1811 (
		_w895_,
		_w1365_,
		_w2059_
	);
	LUT2 #(
		.INIT('h1)
	) name1812 (
		_w990_,
		_w2059_,
		_w2060_
	);
	LUT2 #(
		.INIT('h2)
	) name1813 (
		_w908_,
		_w2060_,
		_w2061_
	);
	LUT2 #(
		.INIT('h1)
	) name1814 (
		_w2043_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h4)
	) name1815 (
		_w2058_,
		_w2062_,
		_w2063_
	);
	LUT2 #(
		.INIT('h4)
	) name1816 (
		\data_i[26]_pad ,
		_w281_,
		_w2064_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		\rd1_L_o_reg[12]/NET0131 ,
		_w281_,
		_w2065_
	);
	LUT2 #(
		.INIT('h1)
	) name1818 (
		_w2064_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h2)
	) name1819 (
		_w2063_,
		_w2066_,
		_w2067_
	);
	LUT2 #(
		.INIT('h4)
	) name1820 (
		_w2063_,
		_w2066_,
		_w2068_
	);
	LUT2 #(
		.INIT('h1)
	) name1821 (
		_w2067_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h8)
	) name1822 (
		_w1893_,
		_w1898_,
		_w2070_
	);
	LUT2 #(
		.INIT('h4)
	) name1823 (
		_w1890_,
		_w1920_,
		_w2071_
	);
	LUT2 #(
		.INIT('h1)
	) name1824 (
		_w1909_,
		_w2071_,
		_w2072_
	);
	LUT2 #(
		.INIT('h2)
	) name1825 (
		_w1868_,
		_w2072_,
		_w2073_
	);
	LUT2 #(
		.INIT('h8)
	) name1826 (
		_w1865_,
		_w1923_,
		_w2074_
	);
	LUT2 #(
		.INIT('h4)
	) name1827 (
		_w1890_,
		_w1919_,
		_w2075_
	);
	LUT2 #(
		.INIT('h4)
	) name1828 (
		_w1872_,
		_w1897_,
		_w2076_
	);
	LUT2 #(
		.INIT('h1)
	) name1829 (
		_w2074_,
		_w2075_,
		_w2077_
	);
	LUT2 #(
		.INIT('h4)
	) name1830 (
		_w2076_,
		_w2077_,
		_w2078_
	);
	LUT2 #(
		.INIT('h1)
	) name1831 (
		_w1868_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h1)
	) name1832 (
		_w2070_,
		_w2073_,
		_w2080_
	);
	LUT2 #(
		.INIT('h4)
	) name1833 (
		_w2079_,
		_w2080_,
		_w2081_
	);
	LUT2 #(
		.INIT('h1)
	) name1834 (
		_w1906_,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h8)
	) name1835 (
		_w1886_,
		_w1892_,
		_w2083_
	);
	LUT2 #(
		.INIT('h8)
	) name1836 (
		_w1865_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h8)
	) name1837 (
		_w1868_,
		_w1894_,
		_w2085_
	);
	LUT2 #(
		.INIT('h8)
	) name1838 (
		_w1872_,
		_w1942_,
		_w2086_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w1872_,
		_w1942_,
		_w2087_
	);
	LUT2 #(
		.INIT('h1)
	) name1840 (
		_w1868_,
		_w2086_,
		_w2088_
	);
	LUT2 #(
		.INIT('h4)
	) name1841 (
		_w2087_,
		_w2088_,
		_w2089_
	);
	LUT2 #(
		.INIT('h1)
	) name1842 (
		_w2084_,
		_w2085_,
		_w2090_
	);
	LUT2 #(
		.INIT('h4)
	) name1843 (
		_w2089_,
		_w2090_,
		_w2091_
	);
	LUT2 #(
		.INIT('h2)
	) name1844 (
		_w1906_,
		_w2091_,
		_w2092_
	);
	LUT2 #(
		.INIT('h4)
	) name1845 (
		_w1865_,
		_w1887_,
		_w2093_
	);
	LUT2 #(
		.INIT('h4)
	) name1846 (
		_w1890_,
		_w2093_,
		_w2094_
	);
	LUT2 #(
		.INIT('h8)
	) name1847 (
		_w1869_,
		_w1890_,
		_w2095_
	);
	LUT2 #(
		.INIT('h8)
	) name1848 (
		_w1920_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('h1)
	) name1849 (
		_w2094_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h4)
	) name1850 (
		_w2092_,
		_w2097_,
		_w2098_
	);
	LUT2 #(
		.INIT('h4)
	) name1851 (
		_w2082_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h4)
	) name1852 (
		\data_i[60]_pad ,
		_w281_,
		_w2100_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		\rd1_L_o_reg[16]/NET0131 ,
		_w281_,
		_w2101_
	);
	LUT2 #(
		.INIT('h1)
	) name1854 (
		_w2100_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('h2)
	) name1855 (
		_w2099_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h4)
	) name1856 (
		_w2099_,
		_w2102_,
		_w2104_
	);
	LUT2 #(
		.INIT('h1)
	) name1857 (
		_w2103_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h8)
	) name1858 (
		_w804_,
		_w822_,
		_w2106_
	);
	LUT2 #(
		.INIT('h8)
	) name1859 (
		_w822_,
		_w825_,
		_w2107_
	);
	LUT2 #(
		.INIT('h1)
	) name1860 (
		_w2106_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h8)
	) name1861 (
		_w783_,
		_w828_,
		_w2109_
	);
	LUT2 #(
		.INIT('h2)
	) name1862 (
		_w837_,
		_w2109_,
		_w2110_
	);
	LUT2 #(
		.INIT('h8)
	) name1863 (
		_w2108_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('h4)
	) name1864 (
		_w822_,
		_w831_,
		_w2112_
	);
	LUT2 #(
		.INIT('h1)
	) name1865 (
		_w837_,
		_w870_,
		_w2113_
	);
	LUT2 #(
		.INIT('h4)
	) name1866 (
		_w2112_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h1)
	) name1867 (
		_w2111_,
		_w2114_,
		_w2115_
	);
	LUT2 #(
		.INIT('h2)
	) name1868 (
		_w799_,
		_w822_,
		_w2116_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w839_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h4)
	) name1870 (
		_w783_,
		_w837_,
		_w2118_
	);
	LUT2 #(
		.INIT('h4)
	) name1871 (
		_w2117_,
		_w2118_,
		_w2119_
	);
	LUT2 #(
		.INIT('h4)
	) name1872 (
		_w799_,
		_w868_,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name1873 (
		_w783_,
		_w803_,
		_w2121_
	);
	LUT2 #(
		.INIT('h1)
	) name1874 (
		_w825_,
		_w2121_,
		_w2122_
	);
	LUT2 #(
		.INIT('h2)
	) name1875 (
		_w822_,
		_w869_,
		_w2123_
	);
	LUT2 #(
		.INIT('h4)
	) name1876 (
		_w2122_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h2)
	) name1877 (
		_w862_,
		_w2119_,
		_w2125_
	);
	LUT2 #(
		.INIT('h4)
	) name1878 (
		_w2120_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h4)
	) name1879 (
		_w2124_,
		_w2126_,
		_w2127_
	);
	LUT2 #(
		.INIT('h1)
	) name1880 (
		_w829_,
		_w831_,
		_w2128_
	);
	LUT2 #(
		.INIT('h1)
	) name1881 (
		_w799_,
		_w837_,
		_w2129_
	);
	LUT2 #(
		.INIT('h4)
	) name1882 (
		_w2128_,
		_w2129_,
		_w2130_
	);
	LUT2 #(
		.INIT('h8)
	) name1883 (
		_w822_,
		_w837_,
		_w2131_
	);
	LUT2 #(
		.INIT('h8)
	) name1884 (
		_w2121_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h1)
	) name1885 (
		_w862_,
		_w2132_,
		_w2133_
	);
	LUT2 #(
		.INIT('h4)
	) name1886 (
		_w2130_,
		_w2133_,
		_w2134_
	);
	LUT2 #(
		.INIT('h8)
	) name1887 (
		_w827_,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h1)
	) name1888 (
		_w2127_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h4)
	) name1889 (
		_w783_,
		_w839_,
		_w2137_
	);
	LUT2 #(
		.INIT('h4)
	) name1890 (
		_w822_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h1)
	) name1891 (
		_w2115_,
		_w2138_,
		_w2139_
	);
	LUT2 #(
		.INIT('h4)
	) name1892 (
		_w2136_,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h4)
	) name1893 (
		\data_i[52]_pad ,
		_w281_,
		_w2141_
	);
	LUT2 #(
		.INIT('h1)
	) name1894 (
		\rd1_L_o_reg[17]/NET0131 ,
		_w281_,
		_w2142_
	);
	LUT2 #(
		.INIT('h1)
	) name1895 (
		_w2141_,
		_w2142_,
		_w2143_
	);
	LUT2 #(
		.INIT('h2)
	) name1896 (
		_w2140_,
		_w2143_,
		_w2144_
	);
	LUT2 #(
		.INIT('h4)
	) name1897 (
		_w2140_,
		_w2143_,
		_w2145_
	);
	LUT2 #(
		.INIT('h1)
	) name1898 (
		_w2144_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h4)
	) name1899 (
		_w1432_,
		_w1466_,
		_w2147_
	);
	LUT2 #(
		.INIT('h1)
	) name1900 (
		_w1419_,
		_w1454_,
		_w2148_
	);
	LUT2 #(
		.INIT('h4)
	) name1901 (
		_w1466_,
		_w2148_,
		_w2149_
	);
	LUT2 #(
		.INIT('h2)
	) name1902 (
		_w1416_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		_w1460_,
		_w1511_,
		_w2151_
	);
	LUT2 #(
		.INIT('h4)
	) name1904 (
		_w2147_,
		_w2151_,
		_w2152_
	);
	LUT2 #(
		.INIT('h4)
	) name1905 (
		_w2150_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h1)
	) name1906 (
		_w1416_,
		_w1786_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name1907 (
		_w1419_,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h4)
	) name1908 (
		_w1432_,
		_w1473_,
		_w2156_
	);
	LUT2 #(
		.INIT('h4)
	) name1909 (
		_w1416_,
		_w1419_,
		_w2157_
	);
	LUT2 #(
		.INIT('h1)
	) name1910 (
		_w1462_,
		_w2157_,
		_w2158_
	);
	LUT2 #(
		.INIT('h1)
	) name1911 (
		_w2155_,
		_w2156_,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1912 (
		_w2158_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h1)
	) name1913 (
		_w2153_,
		_w2160_,
		_w2161_
	);
	LUT2 #(
		.INIT('h8)
	) name1914 (
		_w1419_,
		_w1440_,
		_w2162_
	);
	LUT2 #(
		.INIT('h8)
	) name1915 (
		_w1472_,
		_w2162_,
		_w2163_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		_w1452_,
		_w1782_,
		_w2164_
	);
	LUT2 #(
		.INIT('h1)
	) name1917 (
		_w2163_,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('h4)
	) name1918 (
		_w1495_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h4)
	) name1919 (
		_w2161_,
		_w2166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h4)
	) name1920 (
		\data_i[28]_pad ,
		_w281_,
		_w2168_
	);
	LUT2 #(
		.INIT('h1)
	) name1921 (
		\rd1_L_o_reg[20]/NET0131 ,
		_w281_,
		_w2169_
	);
	LUT2 #(
		.INIT('h1)
	) name1922 (
		_w2168_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h2)
	) name1923 (
		_w2167_,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h4)
	) name1924 (
		_w2167_,
		_w2170_,
		_w2172_
	);
	LUT2 #(
		.INIT('h1)
	) name1925 (
		_w2171_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h1)
	) name1926 (
		_w1571_,
		_w1581_,
		_w2174_
	);
	LUT2 #(
		.INIT('h8)
	) name1927 (
		_w1598_,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h8)
	) name1928 (
		_w1535_,
		_w1696_,
		_w2176_
	);
	LUT2 #(
		.INIT('h2)
	) name1929 (
		_w1568_,
		_w1716_,
		_w2177_
	);
	LUT2 #(
		.INIT('h4)
	) name1930 (
		_w2176_,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h1)
	) name1931 (
		_w2175_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h2)
	) name1932 (
		_w1579_,
		_w2179_,
		_w2180_
	);
	LUT2 #(
		.INIT('h8)
	) name1933 (
		_w1550_,
		_w1706_,
		_w2181_
	);
	LUT2 #(
		.INIT('h1)
	) name1934 (
		_w1560_,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w1568_,
		_w2182_,
		_w2183_
	);
	LUT2 #(
		.INIT('h8)
	) name1936 (
		_w1568_,
		_w1592_,
		_w2184_
	);
	LUT2 #(
		.INIT('h1)
	) name1937 (
		_w1733_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h1)
	) name1938 (
		_w1550_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h2)
	) name1939 (
		_w1568_,
		_w1584_,
		_w2187_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w1579_,
		_w1718_,
		_w2188_
	);
	LUT2 #(
		.INIT('h4)
	) name1941 (
		_w2183_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h1)
	) name1942 (
		_w2186_,
		_w2187_,
		_w2190_
	);
	LUT2 #(
		.INIT('h8)
	) name1943 (
		_w2189_,
		_w2190_,
		_w2191_
	);
	LUT2 #(
		.INIT('h1)
	) name1944 (
		_w2180_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h1)
	) name1945 (
		_w1695_,
		_w1704_,
		_w2193_
	);
	LUT2 #(
		.INIT('h1)
	) name1946 (
		_w1568_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h4)
	) name1947 (
		_w1535_,
		_w1568_,
		_w2195_
	);
	LUT2 #(
		.INIT('h4)
	) name1948 (
		_w1599_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h4)
	) name1949 (
		_w1715_,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h1)
	) name1950 (
		_w2194_,
		_w2197_,
		_w2198_
	);
	LUT2 #(
		.INIT('h4)
	) name1951 (
		_w2192_,
		_w2198_,
		_w2199_
	);
	LUT2 #(
		.INIT('h4)
	) name1952 (
		\data_i[4]_pad ,
		_w281_,
		_w2200_
	);
	LUT2 #(
		.INIT('h1)
	) name1953 (
		\rd1_L_o_reg[23]/NET0131 ,
		_w281_,
		_w2201_
	);
	LUT2 #(
		.INIT('h1)
	) name1954 (
		_w2200_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h2)
	) name1955 (
		_w2199_,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h4)
	) name1956 (
		_w2199_,
		_w2202_,
		_w2204_
	);
	LUT2 #(
		.INIT('h1)
	) name1957 (
		_w2203_,
		_w2204_,
		_w2205_
	);
	LUT2 #(
		.INIT('h8)
	) name1958 (
		_w1624_,
		_w1649_,
		_w2206_
	);
	LUT2 #(
		.INIT('h1)
	) name1959 (
		_w2007_,
		_w2206_,
		_w2207_
	);
	LUT2 #(
		.INIT('h2)
	) name1960 (
		_w1658_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h4)
	) name1961 (
		_w1635_,
		_w1654_,
		_w2209_
	);
	LUT2 #(
		.INIT('h1)
	) name1962 (
		_w2208_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h1)
	) name1963 (
		_w1640_,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h2)
	) name1964 (
		_w1622_,
		_w1635_,
		_w2212_
	);
	LUT2 #(
		.INIT('h1)
	) name1965 (
		_w1654_,
		_w2212_,
		_w2213_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		_w1671_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h1)
	) name1967 (
		_w1640_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h8)
	) name1968 (
		_w1629_,
		_w1640_,
		_w2216_
	);
	LUT2 #(
		.INIT('h4)
	) name1969 (
		_w1670_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h8)
	) name1970 (
		_w1635_,
		_w1672_,
		_w2218_
	);
	LUT2 #(
		.INIT('h1)
	) name1971 (
		_w1635_,
		_w2006_,
		_w2219_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		_w2217_,
		_w2218_,
		_w2220_
	);
	LUT2 #(
		.INIT('h4)
	) name1973 (
		_w2219_,
		_w2220_,
		_w2221_
	);
	LUT2 #(
		.INIT('h4)
	) name1974 (
		_w2215_,
		_w2221_,
		_w2222_
	);
	LUT2 #(
		.INIT('h1)
	) name1975 (
		_w1658_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h8)
	) name1976 (
		_w1621_,
		_w1627_,
		_w2224_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		_w2015_,
		_w2224_,
		_w2225_
	);
	LUT2 #(
		.INIT('h2)
	) name1978 (
		_w1640_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		_w1635_,
		_w2008_,
		_w2227_
	);
	LUT2 #(
		.INIT('h1)
	) name1980 (
		_w2226_,
		_w2227_,
		_w2228_
	);
	LUT2 #(
		.INIT('h2)
	) name1981 (
		_w1658_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h8)
	) name1982 (
		_w1618_,
		_w2224_,
		_w2230_
	);
	LUT2 #(
		.INIT('h2)
	) name1983 (
		_w1635_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h2)
	) name1984 (
		_w1640_,
		_w1649_,
		_w2232_
	);
	LUT2 #(
		.INIT('h4)
	) name1985 (
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('h1)
	) name1986 (
		_w2229_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h4)
	) name1987 (
		_w2211_,
		_w2234_,
		_w2235_
	);
	LUT2 #(
		.INIT('h4)
	) name1988 (
		_w2223_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h4)
	) name1989 (
		\data_i[30]_pad ,
		_w281_,
		_w2237_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		\rd1_L_o_reg[28]/NET0131 ,
		_w281_,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		_w2237_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h2)
	) name1992 (
		_w2236_,
		_w2239_,
		_w2240_
	);
	LUT2 #(
		.INIT('h4)
	) name1993 (
		_w2236_,
		_w2239_,
		_w2241_
	);
	LUT2 #(
		.INIT('h1)
	) name1994 (
		_w2240_,
		_w2241_,
		_w2242_
	);
	LUT2 #(
		.INIT('h1)
	) name1995 (
		_w1570_,
		_w1694_,
		_w2243_
	);
	LUT2 #(
		.INIT('h2)
	) name1996 (
		_w1579_,
		_w2243_,
		_w2244_
	);
	LUT2 #(
		.INIT('h1)
	) name1997 (
		_w1698_,
		_w2244_,
		_w2245_
	);
	LUT2 #(
		.INIT('h1)
	) name1998 (
		_w1568_,
		_w2245_,
		_w2246_
	);
	LUT2 #(
		.INIT('h1)
	) name1999 (
		_w1538_,
		_w1585_,
		_w2247_
	);
	LUT2 #(
		.INIT('h4)
	) name2000 (
		_w1551_,
		_w1568_,
		_w2248_
	);
	LUT2 #(
		.INIT('h4)
	) name2001 (
		_w2247_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h1)
	) name2002 (
		_w1704_,
		_w2176_,
		_w2250_
	);
	LUT2 #(
		.INIT('h4)
	) name2003 (
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h2)
	) name2004 (
		_w1579_,
		_w2251_,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name2005 (
		_w1560_,
		_w1707_,
		_w2253_
	);
	LUT2 #(
		.INIT('h2)
	) name2006 (
		_w1568_,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h1)
	) name2007 (
		_w1538_,
		_w1591_,
		_w2255_
	);
	LUT2 #(
		.INIT('h4)
	) name2008 (
		_w1703_,
		_w2195_,
		_w2256_
	);
	LUT2 #(
		.INIT('h4)
	) name2009 (
		_w2255_,
		_w2256_,
		_w2257_
	);
	LUT2 #(
		.INIT('h1)
	) name2010 (
		_w1585_,
		_w1697_,
		_w2258_
	);
	LUT2 #(
		.INIT('h1)
	) name2011 (
		_w1568_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		_w1568_,
		_w1581_,
		_w2260_
	);
	LUT2 #(
		.INIT('h1)
	) name2013 (
		_w1564_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h4)
	) name2014 (
		_w2259_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h1)
	) name2015 (
		_w1579_,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		_w1604_,
		_w2257_,
		_w2264_
	);
	LUT2 #(
		.INIT('h4)
	) name2017 (
		_w2254_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h4)
	) name2018 (
		_w2246_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h4)
	) name2019 (
		_w2252_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h4)
	) name2020 (
		_w2263_,
		_w2267_,
		_w2268_
	);
	LUT2 #(
		.INIT('h4)
	) name2021 (
		\data_i[2]_pad ,
		_w281_,
		_w2269_
	);
	LUT2 #(
		.INIT('h1)
	) name2022 (
		\rd1_L_o_reg[15]/NET0131 ,
		_w281_,
		_w2270_
	);
	LUT2 #(
		.INIT('h1)
	) name2023 (
		_w2269_,
		_w2270_,
		_w2271_
	);
	LUT2 #(
		.INIT('h2)
	) name2024 (
		_w2268_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h4)
	) name2025 (
		_w2268_,
		_w2271_,
		_w2273_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		_w2272_,
		_w2273_,
		_w2274_
	);
	LUT2 #(
		.INIT('h1)
	) name2027 (
		_w1261_,
		_w1322_,
		_w2275_
	);
	LUT2 #(
		.INIT('h2)
	) name2028 (
		_w1300_,
		_w1317_,
		_w2276_
	);
	LUT2 #(
		.INIT('h4)
	) name2029 (
		_w2275_,
		_w2276_,
		_w2277_
	);
	LUT2 #(
		.INIT('h4)
	) name2030 (
		_w1242_,
		_w2277_,
		_w2278_
	);
	LUT2 #(
		.INIT('h4)
	) name2031 (
		_w1303_,
		_w2275_,
		_w2279_
	);
	LUT2 #(
		.INIT('h4)
	) name2032 (
		_w1257_,
		_w1261_,
		_w2280_
	);
	LUT2 #(
		.INIT('h8)
	) name2033 (
		_w1242_,
		_w2280_,
		_w2281_
	);
	LUT2 #(
		.INIT('h1)
	) name2034 (
		_w2279_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w1300_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h8)
	) name2036 (
		_w1257_,
		_w2277_,
		_w2284_
	);
	LUT2 #(
		.INIT('h1)
	) name2037 (
		_w1308_,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('h4)
	) name2038 (
		_w2283_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h2)
	) name2039 (
		_w1269_,
		_w2286_,
		_w2287_
	);
	LUT2 #(
		.INIT('h4)
	) name2040 (
		_w1242_,
		_w1317_,
		_w2288_
	);
	LUT2 #(
		.INIT('h1)
	) name2041 (
		_w1282_,
		_w2288_,
		_w2289_
	);
	LUT2 #(
		.INIT('h8)
	) name2042 (
		_w1971_,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h1)
	) name2043 (
		_w1282_,
		_w1324_,
		_w2291_
	);
	LUT2 #(
		.INIT('h2)
	) name2044 (
		_w1239_,
		_w2280_,
		_w2292_
	);
	LUT2 #(
		.INIT('h4)
	) name2045 (
		_w1271_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h1)
	) name2046 (
		_w2291_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name2047 (
		_w1300_,
		_w2294_,
		_w2295_
	);
	LUT2 #(
		.INIT('h1)
	) name2048 (
		_w1269_,
		_w2290_,
		_w2296_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		_w2295_,
		_w2296_,
		_w2297_
	);
	LUT2 #(
		.INIT('h8)
	) name2050 (
		_w1239_,
		_w1976_,
		_w2298_
	);
	LUT2 #(
		.INIT('h8)
	) name2051 (
		_w1261_,
		_w1322_,
		_w2299_
	);
	LUT2 #(
		.INIT('h1)
	) name2052 (
		_w2298_,
		_w2299_,
		_w2300_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		_w1300_,
		_w2300_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name2054 (
		_w1958_,
		_w2278_,
		_w2302_
	);
	LUT2 #(
		.INIT('h4)
	) name2055 (
		_w2301_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h4)
	) name2056 (
		_w2297_,
		_w2303_,
		_w2304_
	);
	LUT2 #(
		.INIT('h4)
	) name2057 (
		_w2287_,
		_w2304_,
		_w2305_
	);
	LUT2 #(
		.INIT('h4)
	) name2058 (
		\data_i[24]_pad ,
		_w281_,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name2059 (
		\rd1_L_o_reg[4]/NET0131 ,
		_w281_,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name2060 (
		_w2306_,
		_w2307_,
		_w2308_
	);
	LUT2 #(
		.INIT('h2)
	) name2061 (
		_w2305_,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('h4)
	) name2062 (
		_w2305_,
		_w2308_,
		_w2310_
	);
	LUT2 #(
		.INIT('h1)
	) name2063 (
		_w2309_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h4)
	) name2064 (
		_w1160_,
		_w1173_,
		_w2312_
	);
	LUT2 #(
		.INIT('h1)
	) name2065 (
		_w1098_,
		_w1109_,
		_w2313_
	);
	LUT2 #(
		.INIT('h2)
	) name2066 (
		_w1820_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h1)
	) name2067 (
		_w1158_,
		_w2314_,
		_w2315_
	);
	LUT2 #(
		.INIT('h4)
	) name2068 (
		_w1754_,
		_w2315_,
		_w2316_
	);
	LUT2 #(
		.INIT('h4)
	) name2069 (
		_w2312_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('h4)
	) name2070 (
		_w1098_,
		_w1147_,
		_w2318_
	);
	LUT2 #(
		.INIT('h1)
	) name2071 (
		_w1110_,
		_w1135_,
		_w2319_
	);
	LUT2 #(
		.INIT('h2)
	) name2072 (
		_w1098_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h4)
	) name2073 (
		_w1136_,
		_w1158_,
		_w2321_
	);
	LUT2 #(
		.INIT('h4)
	) name2074 (
		_w1817_,
		_w2321_,
		_w2322_
	);
	LUT2 #(
		.INIT('h4)
	) name2075 (
		_w2318_,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h4)
	) name2076 (
		_w2320_,
		_w2323_,
		_w2324_
	);
	LUT2 #(
		.INIT('h1)
	) name2077 (
		_w2317_,
		_w2324_,
		_w2325_
	);
	LUT2 #(
		.INIT('h1)
	) name2078 (
		_w1143_,
		_w1148_,
		_w2326_
	);
	LUT2 #(
		.INIT('h1)
	) name2079 (
		_w1098_,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h8)
	) name2080 (
		_w1181_,
		_w1745_,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w1105_,
		_w1106_,
		_w2329_
	);
	LUT2 #(
		.INIT('h8)
	) name2082 (
		_w1173_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h1)
	) name2083 (
		_w1110_,
		_w1149_,
		_w2331_
	);
	LUT2 #(
		.INIT('h1)
	) name2084 (
		_w1098_,
		_w1158_,
		_w2332_
	);
	LUT2 #(
		.INIT('h4)
	) name2085 (
		_w2331_,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h1)
	) name2086 (
		_w1769_,
		_w2328_,
		_w2334_
	);
	LUT2 #(
		.INIT('h4)
	) name2087 (
		_w2330_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h4)
	) name2088 (
		_w2333_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h4)
	) name2089 (
		_w2327_,
		_w2336_,
		_w2337_
	);
	LUT2 #(
		.INIT('h4)
	) name2090 (
		_w2325_,
		_w2337_,
		_w2338_
	);
	LUT2 #(
		.INIT('h4)
	) name2091 (
		\data_i[0]_pad ,
		_w281_,
		_w2339_
	);
	LUT2 #(
		.INIT('h1)
	) name2092 (
		\rd1_L_o_reg[7]/NET0131 ,
		_w281_,
		_w2340_
	);
	LUT2 #(
		.INIT('h1)
	) name2093 (
		_w2339_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('h2)
	) name2094 (
		_w2338_,
		_w2341_,
		_w2342_
	);
	LUT2 #(
		.INIT('h4)
	) name2095 (
		_w2338_,
		_w2341_,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name2096 (
		_w2342_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h2)
	) name2097 (
		_w1886_,
		_w1893_,
		_w2345_
	);
	LUT2 #(
		.INIT('h1)
	) name2098 (
		_w1894_,
		_w2345_,
		_w2346_
	);
	LUT2 #(
		.INIT('h2)
	) name2099 (
		_w1906_,
		_w1907_,
		_w2347_
	);
	LUT2 #(
		.INIT('h4)
	) name2100 (
		_w2346_,
		_w2347_,
		_w2348_
	);
	LUT2 #(
		.INIT('h4)
	) name2101 (
		_w1906_,
		_w2346_,
		_w2349_
	);
	LUT2 #(
		.INIT('h4)
	) name2102 (
		_w1890_,
		_w1910_,
		_w2350_
	);
	LUT2 #(
		.INIT('h1)
	) name2103 (
		_w1909_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h4)
	) name2104 (
		_w2348_,
		_w2351_,
		_w2352_
	);
	LUT2 #(
		.INIT('h4)
	) name2105 (
		_w2349_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('h1)
	) name2106 (
		_w1868_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		_w2083_,
		_w2086_,
		_w2355_
	);
	LUT2 #(
		.INIT('h2)
	) name2108 (
		_w1868_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h8)
	) name2109 (
		_w1865_,
		_w2075_,
		_w2357_
	);
	LUT2 #(
		.INIT('h1)
	) name2110 (
		_w2356_,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('h1)
	) name2111 (
		_w1906_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h2)
	) name2112 (
		_w1906_,
		_w1942_,
		_w2360_
	);
	LUT2 #(
		.INIT('h4)
	) name2113 (
		_w2083_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w2084_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h2)
	) name2115 (
		_w1868_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h1)
	) name2116 (
		_w2359_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('h4)
	) name2117 (
		_w2354_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h4)
	) name2118 (
		\data_i[46]_pad ,
		_w281_,
		_w2366_
	);
	LUT2 #(
		.INIT('h1)
	) name2119 (
		\rd1_L_o_reg[26]/NET0131 ,
		_w281_,
		_w2367_
	);
	LUT2 #(
		.INIT('h1)
	) name2120 (
		_w2366_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h2)
	) name2121 (
		_w2365_,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h4)
	) name2122 (
		_w2365_,
		_w2368_,
		_w2370_
	);
	LUT2 #(
		.INIT('h1)
	) name2123 (
		_w2369_,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('h4)
	) name2124 (
		_w1886_,
		_w2074_,
		_w2372_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w1897_,
		_w2074_,
		_w2373_
	);
	LUT2 #(
		.INIT('h4)
	) name2126 (
		_w2071_,
		_w2373_,
		_w2374_
	);
	LUT2 #(
		.INIT('h2)
	) name2127 (
		_w1868_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h1)
	) name2128 (
		_w1908_,
		_w2075_,
		_w2376_
	);
	LUT2 #(
		.INIT('h4)
	) name2129 (
		_w2093_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h1)
	) name2130 (
		_w1868_,
		_w2377_,
		_w2378_
	);
	LUT2 #(
		.INIT('h1)
	) name2131 (
		_w2372_,
		_w2375_,
		_w2379_
	);
	LUT2 #(
		.INIT('h4)
	) name2132 (
		_w2378_,
		_w2379_,
		_w2380_
	);
	LUT2 #(
		.INIT('h2)
	) name2133 (
		_w1906_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		_w1887_,
		_w1892_,
		_w2382_
	);
	LUT2 #(
		.INIT('h4)
	) name2135 (
		_w1916_,
		_w2382_,
		_w2383_
	);
	LUT2 #(
		.INIT('h2)
	) name2136 (
		_w1865_,
		_w1906_,
		_w2384_
	);
	LUT2 #(
		.INIT('h4)
	) name2137 (
		_w1923_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h4)
	) name2138 (
		_w1920_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h2)
	) name2139 (
		_w1868_,
		_w2383_,
		_w2387_
	);
	LUT2 #(
		.INIT('h4)
	) name2140 (
		_w2386_,
		_w2387_,
		_w2388_
	);
	LUT2 #(
		.INIT('h2)
	) name2141 (
		_w1890_,
		_w1899_,
		_w2389_
	);
	LUT2 #(
		.INIT('h4)
	) name2142 (
		_w1897_,
		_w2071_,
		_w2390_
	);
	LUT2 #(
		.INIT('h1)
	) name2143 (
		_w2389_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name2144 (
		_w1906_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h1)
	) name2145 (
		_w1868_,
		_w2094_,
		_w2393_
	);
	LUT2 #(
		.INIT('h4)
	) name2146 (
		_w2392_,
		_w2393_,
		_w2394_
	);
	LUT2 #(
		.INIT('h1)
	) name2147 (
		_w2388_,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h1)
	) name2148 (
		_w2381_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h4)
	) name2149 (
		\data_i[40]_pad ,
		_w281_,
		_w2397_
	);
	LUT2 #(
		.INIT('h1)
	) name2150 (
		\rd1_L_o_reg[2]/NET0131 ,
		_w281_,
		_w2398_
	);
	LUT2 #(
		.INIT('h1)
	) name2151 (
		_w2397_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		_w2396_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h4)
	) name2153 (
		_w2396_,
		_w2399_,
		_w2401_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		_w2400_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h1)
	) name2155 (
		_w1277_,
		_w2275_,
		_w2403_
	);
	LUT2 #(
		.INIT('h4)
	) name2156 (
		_w1242_,
		_w1970_,
		_w2404_
	);
	LUT2 #(
		.INIT('h8)
	) name2157 (
		_w1257_,
		_w1959_,
		_w2405_
	);
	LUT2 #(
		.INIT('h1)
	) name2158 (
		_w1300_,
		_w1323_,
		_w2406_
	);
	LUT2 #(
		.INIT('h1)
	) name2159 (
		_w1955_,
		_w2405_,
		_w2407_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		_w2406_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h2)
	) name2161 (
		_w1300_,
		_w1304_,
		_w2409_
	);
	LUT2 #(
		.INIT('h4)
	) name2162 (
		_w2288_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h1)
	) name2163 (
		_w2408_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h2)
	) name2164 (
		_w1269_,
		_w2403_,
		_w2412_
	);
	LUT2 #(
		.INIT('h4)
	) name2165 (
		_w2404_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h4)
	) name2166 (
		_w2411_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h1)
	) name2167 (
		_w1309_,
		_w1322_,
		_w2415_
	);
	LUT2 #(
		.INIT('h4)
	) name2168 (
		_w2280_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h2)
	) name2169 (
		_w1300_,
		_w2416_,
		_w2417_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w1282_,
		_w1309_,
		_w2418_
	);
	LUT2 #(
		.INIT('h8)
	) name2171 (
		_w2406_,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		_w2417_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h1)
	) name2173 (
		_w1269_,
		_w1318_,
		_w2421_
	);
	LUT2 #(
		.INIT('h4)
	) name2174 (
		_w2298_,
		_w2421_,
		_w2422_
	);
	LUT2 #(
		.INIT('h4)
	) name2175 (
		_w2420_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h1)
	) name2176 (
		_w2414_,
		_w2423_,
		_w2424_
	);
	LUT2 #(
		.INIT('h4)
	) name2177 (
		\data_i[10]_pad ,
		_w281_,
		_w2425_
	);
	LUT2 #(
		.INIT('h1)
	) name2178 (
		\rd1_L_o_reg[14]/NET0131 ,
		_w281_,
		_w2426_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w2425_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h2)
	) name2180 (
		_w2424_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h4)
	) name2181 (
		_w2424_,
		_w2427_,
		_w2429_
	);
	LUT2 #(
		.INIT('h1)
	) name2182 (
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h8)
	) name2183 (
		_w995_,
		_w2046_,
		_w2431_
	);
	LUT2 #(
		.INIT('h1)
	) name2184 (
		_w958_,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h2)
	) name2185 (
		_w1371_,
		_w2432_,
		_w2433_
	);
	LUT2 #(
		.INIT('h2)
	) name2186 (
		_w987_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h4)
	) name2187 (
		_w901_,
		_w941_,
		_w2435_
	);
	LUT2 #(
		.INIT('h4)
	) name2188 (
		_w939_,
		_w2036_,
		_w2436_
	);
	LUT2 #(
		.INIT('h1)
	) name2189 (
		_w1358_,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h1)
	) name2190 (
		_w958_,
		_w2437_,
		_w2438_
	);
	LUT2 #(
		.INIT('h4)
	) name2191 (
		_w1002_,
		_w2046_,
		_w2439_
	);
	LUT2 #(
		.INIT('h2)
	) name2192 (
		_w958_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h1)
	) name2193 (
		_w2435_,
		_w2438_,
		_w2441_
	);
	LUT2 #(
		.INIT('h4)
	) name2194 (
		_w2440_,
		_w2441_,
		_w2442_
	);
	LUT2 #(
		.INIT('h1)
	) name2195 (
		_w987_,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('h1)
	) name2196 (
		_w1386_,
		_w2036_,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name2197 (
		_w902_,
		_w991_,
		_w2445_
	);
	LUT2 #(
		.INIT('h2)
	) name2198 (
		_w1388_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h1)
	) name2199 (
		_w2444_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('h4)
	) name2200 (
		_w2434_,
		_w2447_,
		_w2448_
	);
	LUT2 #(
		.INIT('h4)
	) name2201 (
		_w2443_,
		_w2448_,
		_w2449_
	);
	LUT2 #(
		.INIT('h4)
	) name2202 (
		\data_i[6]_pad ,
		_w281_,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		\rd1_L_o_reg[31]/NET0131 ,
		_w281_,
		_w2451_
	);
	LUT2 #(
		.INIT('h1)
	) name2204 (
		_w2450_,
		_w2451_,
		_w2452_
	);
	LUT2 #(
		.INIT('h2)
	) name2205 (
		_w2449_,
		_w2452_,
		_w2453_
	);
	LUT2 #(
		.INIT('h4)
	) name2206 (
		_w2449_,
		_w2452_,
		_w2454_
	);
	LUT2 #(
		.INIT('h1)
	) name2207 (
		_w2453_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h8)
	) name2208 (
		_w799_,
		_w870_,
		_w2456_
	);
	LUT2 #(
		.INIT('h4)
	) name2209 (
		_w862_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h1)
	) name2210 (
		_w800_,
		_w824_,
		_w2458_
	);
	LUT2 #(
		.INIT('h1)
	) name2211 (
		_w804_,
		_w822_,
		_w2459_
	);
	LUT2 #(
		.INIT('h1)
	) name2212 (
		_w2458_,
		_w2459_,
		_w2460_
	);
	LUT2 #(
		.INIT('h1)
	) name2213 (
		_w2138_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('h8)
	) name2214 (
		_w837_,
		_w862_,
		_w2462_
	);
	LUT2 #(
		.INIT('h4)
	) name2215 (
		_w2461_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h1)
	) name2216 (
		_w804_,
		_w868_,
		_w2464_
	);
	LUT2 #(
		.INIT('h4)
	) name2217 (
		_w2137_,
		_w2464_,
		_w2465_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		_w837_,
		_w862_,
		_w2466_
	);
	LUT2 #(
		.INIT('h4)
	) name2219 (
		_w2465_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		_w783_,
		_w866_,
		_w2468_
	);
	LUT2 #(
		.INIT('h2)
	) name2221 (
		_w837_,
		_w2456_,
		_w2469_
	);
	LUT2 #(
		.INIT('h4)
	) name2222 (
		_w2468_,
		_w2469_,
		_w2470_
	);
	LUT2 #(
		.INIT('h1)
	) name2223 (
		_w2109_,
		_w2137_,
		_w2471_
	);
	LUT2 #(
		.INIT('h2)
	) name2224 (
		_w822_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h1)
	) name2225 (
		_w825_,
		_w837_,
		_w2473_
	);
	LUT2 #(
		.INIT('h4)
	) name2226 (
		_w2472_,
		_w2473_,
		_w2474_
	);
	LUT2 #(
		.INIT('h1)
	) name2227 (
		_w2470_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h4)
	) name2228 (
		_w803_,
		_w2116_,
		_w2476_
	);
	LUT2 #(
		.INIT('h1)
	) name2229 (
		_w866_,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h2)
	) name2230 (
		_w862_,
		_w2477_,
		_w2478_
	);
	LUT2 #(
		.INIT('h4)
	) name2231 (
		_w831_,
		_w876_,
		_w2479_
	);
	LUT2 #(
		.INIT('h1)
	) name2232 (
		_w866_,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name2233 (
		_w837_,
		_w2480_,
		_w2481_
	);
	LUT2 #(
		.INIT('h1)
	) name2234 (
		_w2478_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('h1)
	) name2235 (
		_w2462_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h1)
	) name2236 (
		_w2106_,
		_w2457_,
		_w2484_
	);
	LUT2 #(
		.INIT('h4)
	) name2237 (
		_w2467_,
		_w2484_,
		_w2485_
	);
	LUT2 #(
		.INIT('h4)
	) name2238 (
		_w2463_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('h4)
	) name2239 (
		_w2475_,
		_w2486_,
		_w2487_
	);
	LUT2 #(
		.INIT('h4)
	) name2240 (
		_w2483_,
		_w2487_,
		_w2488_
	);
	LUT2 #(
		.INIT('h4)
	) name2241 (
		\data_i[34]_pad ,
		_w281_,
		_w2489_
	);
	LUT2 #(
		.INIT('h1)
	) name2242 (
		\rd1_L_o_reg[11]/NET0131 ,
		_w281_,
		_w2490_
	);
	LUT2 #(
		.INIT('h1)
	) name2243 (
		_w2489_,
		_w2490_,
		_w2491_
	);
	LUT2 #(
		.INIT('h2)
	) name2244 (
		_w2488_,
		_w2491_,
		_w2492_
	);
	LUT2 #(
		.INIT('h4)
	) name2245 (
		_w2488_,
		_w2491_,
		_w2493_
	);
	LUT2 #(
		.INIT('h1)
	) name2246 (
		_w2492_,
		_w2493_,
		_w2494_
	);
	LUT2 #(
		.INIT('h8)
	) name2247 (
		_w800_,
		_w875_,
		_w2495_
	);
	LUT2 #(
		.INIT('h2)
	) name2248 (
		_w837_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h4)
	) name2249 (
		_w823_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name2250 (
		_w2107_,
		_w2138_,
		_w2498_
	);
	LUT2 #(
		.INIT('h8)
	) name2251 (
		_w2497_,
		_w2498_,
		_w2499_
	);
	LUT2 #(
		.INIT('h1)
	) name2252 (
		_w837_,
		_w866_,
		_w2500_
	);
	LUT2 #(
		.INIT('h4)
	) name2253 (
		_w2106_,
		_w2500_,
		_w2501_
	);
	LUT2 #(
		.INIT('h1)
	) name2254 (
		_w2499_,
		_w2501_,
		_w2502_
	);
	LUT2 #(
		.INIT('h2)
	) name2255 (
		_w783_,
		_w828_,
		_w2503_
	);
	LUT2 #(
		.INIT('h8)
	) name2256 (
		_w2131_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('h8)
	) name2257 (
		_w822_,
		_w2137_,
		_w2505_
	);
	LUT2 #(
		.INIT('h1)
	) name2258 (
		_w2109_,
		_w2476_,
		_w2506_
	);
	LUT2 #(
		.INIT('h4)
	) name2259 (
		_w2505_,
		_w2506_,
		_w2507_
	);
	LUT2 #(
		.INIT('h1)
	) name2260 (
		_w837_,
		_w2507_,
		_w2508_
	);
	LUT2 #(
		.INIT('h1)
	) name2261 (
		_w862_,
		_w2468_,
		_w2509_
	);
	LUT2 #(
		.INIT('h4)
	) name2262 (
		_w2504_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h8)
	) name2263 (
		_w2108_,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h4)
	) name2264 (
		_w2508_,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h8)
	) name2265 (
		_w799_,
		_w822_,
		_w2513_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		_w2121_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h2)
	) name2267 (
		_w783_,
		_w837_,
		_w2515_
	);
	LUT2 #(
		.INIT('h2)
	) name2268 (
		_w822_,
		_w839_,
		_w2516_
	);
	LUT2 #(
		.INIT('h2)
	) name2269 (
		_w2515_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h8)
	) name2270 (
		_w822_,
		_w828_,
		_w2518_
	);
	LUT2 #(
		.INIT('h4)
	) name2271 (
		_w2515_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h2)
	) name2272 (
		_w862_,
		_w2514_,
		_w2520_
	);
	LUT2 #(
		.INIT('h4)
	) name2273 (
		_w826_,
		_w2520_,
		_w2521_
	);
	LUT2 #(
		.INIT('h1)
	) name2274 (
		_w2517_,
		_w2519_,
		_w2522_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		_w2521_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h1)
	) name2276 (
		_w2512_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h1)
	) name2277 (
		_w2502_,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h4)
	) name2278 (
		\data_i[38]_pad ,
		_w281_,
		_w2526_
	);
	LUT2 #(
		.INIT('h1)
	) name2279 (
		\rd1_L_o_reg[27]/NET0131 ,
		_w281_,
		_w2527_
	);
	LUT2 #(
		.INIT('h1)
	) name2280 (
		_w2526_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h2)
	) name2281 (
		_w2525_,
		_w2528_,
		_w2529_
	);
	LUT2 #(
		.INIT('h4)
	) name2282 (
		_w2525_,
		_w2528_,
		_w2530_
	);
	LUT2 #(
		.INIT('h1)
	) name2283 (
		_w2529_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h1)
	) name2284 (
		_w1672_,
		_w2004_,
		_w2532_
	);
	LUT2 #(
		.INIT('h8)
	) name2285 (
		_w1635_,
		_w1640_,
		_w2533_
	);
	LUT2 #(
		.INIT('h4)
	) name2286 (
		_w2532_,
		_w2533_,
		_w2534_
	);
	LUT2 #(
		.INIT('h1)
	) name2287 (
		_w1663_,
		_w2008_,
		_w2535_
	);
	LUT2 #(
		.INIT('h2)
	) name2288 (
		_w1640_,
		_w2535_,
		_w2536_
	);
	LUT2 #(
		.INIT('h1)
	) name2289 (
		_w2212_,
		_w2230_,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name2290 (
		_w1640_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w1999_,
		_w2209_,
		_w2539_
	);
	LUT2 #(
		.INIT('h4)
	) name2292 (
		_w2536_,
		_w2539_,
		_w2540_
	);
	LUT2 #(
		.INIT('h4)
	) name2293 (
		_w2538_,
		_w2540_,
		_w2541_
	);
	LUT2 #(
		.INIT('h2)
	) name2294 (
		_w1658_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w1635_,
		_w2532_,
		_w2543_
	);
	LUT2 #(
		.INIT('h1)
	) name2296 (
		_w1640_,
		_w1682_,
		_w2544_
	);
	LUT2 #(
		.INIT('h1)
	) name2297 (
		_w2216_,
		_w2544_,
		_w2545_
	);
	LUT2 #(
		.INIT('h4)
	) name2298 (
		_w2543_,
		_w2545_,
		_w2546_
	);
	LUT2 #(
		.INIT('h1)
	) name2299 (
		_w1658_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h1)
	) name2300 (
		_w1623_,
		_w1993_,
		_w2548_
	);
	LUT2 #(
		.INIT('h1)
	) name2301 (
		_w1635_,
		_w1640_,
		_w2549_
	);
	LUT2 #(
		.INIT('h1)
	) name2302 (
		_w2533_,
		_w2549_,
		_w2550_
	);
	LUT2 #(
		.INIT('h4)
	) name2303 (
		_w2548_,
		_w2550_,
		_w2551_
	);
	LUT2 #(
		.INIT('h1)
	) name2304 (
		_w2534_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('h4)
	) name2305 (
		_w2542_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h4)
	) name2306 (
		_w2547_,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h4)
	) name2307 (
		\data_i[18]_pad ,
		_w281_,
		_w2555_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		\rd1_L_o_reg[13]/NET0131 ,
		_w281_,
		_w2556_
	);
	LUT2 #(
		.INIT('h1)
	) name2309 (
		_w2555_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name2310 (
		_w2554_,
		_w2557_,
		_w2558_
	);
	LUT2 #(
		.INIT('h4)
	) name2311 (
		_w2554_,
		_w2557_,
		_w2559_
	);
	LUT2 #(
		.INIT('h1)
	) name2312 (
		_w2558_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h1)
	) name2313 (
		_w440_,
		_w1087_,
		_w2561_
	);
	LUT2 #(
		.INIT('h4)
	) name2314 (
		_w1204_,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		decrypt_i_pad,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h2)
	) name2316 (
		_w292_,
		_w675_,
		_w2564_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		_w635_,
		_w773_,
		_w2565_
	);
	LUT2 #(
		.INIT('h4)
	) name2318 (
		_w2564_,
		_w2565_,
		_w2566_
	);
	LUT2 #(
		.INIT('h2)
	) name2319 (
		decrypt_i_pad,
		_w2566_,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name2320 (
		_w2563_,
		_w2567_,
		_w2568_
	);
	LUT2 #(
		.INIT('h1)
	) name2321 (
		_w266_,
		_w389_,
		_w2569_
	);
	LUT2 #(
		.INIT('h1)
	) name2322 (
		_w652_,
		_w2569_,
		_w2570_
	);
	LUT2 #(
		.INIT('h1)
	) name2323 (
		decrypt_i_pad,
		_w2570_,
		_w2571_
	);
	LUT2 #(
		.INIT('h2)
	) name2324 (
		_w292_,
		_w524_,
		_w2572_
	);
	LUT2 #(
		.INIT('h1)
	) name2325 (
		_w381_,
		_w1112_,
		_w2573_
	);
	LUT2 #(
		.INIT('h4)
	) name2326 (
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h2)
	) name2327 (
		decrypt_i_pad,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h1)
	) name2328 (
		_w2571_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		_w266_,
		_w368_,
		_w2577_
	);
	LUT2 #(
		.INIT('h1)
	) name2330 (
		_w689_,
		_w2577_,
		_w2578_
	);
	LUT2 #(
		.INIT('h1)
	) name2331 (
		decrypt_i_pad,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h2)
	) name2332 (
		_w292_,
		_w464_,
		_w2580_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		_w360_,
		_w1285_,
		_w2581_
	);
	LUT2 #(
		.INIT('h4)
	) name2334 (
		_w2580_,
		_w2581_,
		_w2582_
	);
	LUT2 #(
		.INIT('h2)
	) name2335 (
		decrypt_i_pad,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h1)
	) name2336 (
		_w2579_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h1)
	) name2337 (
		_w726_,
		_w950_,
		_w2585_
	);
	LUT2 #(
		.INIT('h4)
	) name2338 (
		_w762_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h1)
	) name2339 (
		decrypt_i_pad,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('h2)
	) name2340 (
		_w292_,
		_w612_,
		_w2588_
	);
	LUT2 #(
		.INIT('h1)
	) name2341 (
		_w576_,
		_w1034_,
		_w2589_
	);
	LUT2 #(
		.INIT('h4)
	) name2342 (
		_w2588_,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h2)
	) name2343 (
		decrypt_i_pad,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('h1)
	) name2344 (
		_w2587_,
		_w2591_,
		_w2592_
	);
	LUT2 #(
		.INIT('h1)
	) name2345 (
		_w540_,
		_w1026_,
		_w2593_
	);
	LUT2 #(
		.INIT('h4)
	) name2346 (
		_w1351_,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h1)
	) name2347 (
		decrypt_i_pad,
		_w2594_,
		_w2595_
	);
	LUT2 #(
		.INIT('h1)
	) name2348 (
		_w545_,
		_w789_,
		_w2596_
	);
	LUT2 #(
		.INIT('h4)
	) name2349 (
		_w1055_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h2)
	) name2350 (
		decrypt_i_pad,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name2351 (
		_w2595_,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h1)
	) name2352 (
		_w266_,
		_w605_,
		_w2600_
	);
	LUT2 #(
		.INIT('h2)
	) name2353 (
		_w266_,
		_w733_,
		_w2601_
	);
	LUT2 #(
		.INIT('h1)
	) name2354 (
		_w2600_,
		_w2601_,
		_w2602_
	);
	LUT2 #(
		.INIT('h1)
	) name2355 (
		decrypt_i_pad,
		_w2602_,
		_w2603_
	);
	LUT2 #(
		.INIT('h2)
	) name2356 (
		_w292_,
		_w742_,
		_w2604_
	);
	LUT2 #(
		.INIT('h1)
	) name2357 (
		_w1339_,
		_w1539_,
		_w2605_
	);
	LUT2 #(
		.INIT('h4)
	) name2358 (
		_w2604_,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('h2)
	) name2359 (
		decrypt_i_pad,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h1)
	) name2360 (
		_w2603_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h1)
	) name2361 (
		_w465_,
		_w485_,
		_w2609_
	);
	LUT2 #(
		.INIT('h4)
	) name2362 (
		_w510_,
		_w2609_,
		_w2610_
	);
	LUT2 #(
		.INIT('h1)
	) name2363 (
		decrypt_i_pad,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h2)
	) name2364 (
		_w292_,
		_w516_,
		_w2612_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		_w479_,
		_w2601_,
		_w2613_
	);
	LUT2 #(
		.INIT('h4)
	) name2366 (
		_w2612_,
		_w2613_,
		_w2614_
	);
	LUT2 #(
		.INIT('h2)
	) name2367 (
		decrypt_i_pad,
		_w2614_,
		_w2615_
	);
	LUT2 #(
		.INIT('h1)
	) name2368 (
		_w2611_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h1)
	) name2369 (
		_w266_,
		_w1213_,
		_w2617_
	);
	LUT2 #(
		.INIT('h1)
	) name2370 (
		_w767_,
		_w2617_,
		_w2618_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		decrypt_i_pad,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h1)
	) name2372 (
		_w390_,
		_w657_,
		_w2620_
	);
	LUT2 #(
		.INIT('h4)
	) name2373 (
		_w811_,
		_w2620_,
		_w2621_
	);
	LUT2 #(
		.INIT('h2)
	) name2374 (
		decrypt_i_pad,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h1)
	) name2375 (
		_w2619_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h8)
	) name2376 (
		\data_ready_reg/NET0131 ,
		\stage1_iter_reg[0]/NET0131 ,
		_w2624_
	);
	LUT2 #(
		.INIT('h1)
	) name2377 (
		load_i_pad,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h2)
	) name2378 (
		_w250_,
		_w2625_,
		_w2626_
	);
	LUT2 #(
		.INIT('h1)
	) name2379 (
		\stage1_iter_reg[0]/NET0131 ,
		_w250_,
		_w2627_
	);
	LUT2 #(
		.INIT('h4)
	) name2380 (
		_w263_,
		_w2627_,
		_w2628_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		_w2626_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h1)
	) name2382 (
		\stage1_iter_reg[3]/NET0131 ,
		_w262_,
		_w2630_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w263_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h1)
	) name2384 (
		\stage1_iter_reg[2]/NET0131 ,
		_w254_,
		_w2632_
	);
	LUT2 #(
		.INIT('h1)
	) name2385 (
		_w262_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		\data_ready_reg/NET0131 ,
		_w250_,
		_w2634_
	);
	LUT2 #(
		.INIT('h1)
	) name2387 (
		_w281_,
		_w2634_,
		_w2635_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g10087/_0_  = _w252_ ;
	assign \g10220/_1_  = _w255_ ;
	assign \g11117/_0_  = _w297_ ;
	assign \g11124/_0_  = _w300_ ;
	assign \g11125/_0_  = _w335_ ;
	assign \g11170/_0_  = _w373_ ;
	assign \g11182/_0_  = _w376_ ;
	assign \g11184/_0_  = _w411_ ;
	assign \g11378/_0_  = _w427_ ;
	assign \g11393/_0_  = _w452_ ;
	assign \g11415/_0_  = _w470_ ;
	assign \g11432/_0_  = _w489_ ;
	assign \g11433/_0_  = _w492_ ;
	assign \g11453/_0_  = _w506_ ;
	assign \g11500/_0_  = _w522_ ;
	assign \g11588/_0_  = _w534_ ;
	assign \g11607/_0_  = _w551_ ;
	assign \g11616/_0_  = _w585_ ;
	assign \g11625/_0_  = _w588_ ;
	assign \g11641_dup/_0_  = _w610_ ;
	assign \g11648/_0_  = _w628_ ;
	assign \g11655/_0_  = _w663_ ;
	assign \g11683/_0_  = _w666_ ;
	assign \g11689/_2_  = _w669_ ;
	assign \g11694/_0_  = _w685_ ;
	assign \g11748/_0_  = _w688_ ;
	assign \g11880/_0_  = _w709_ ;
	assign \g11962/_1_  = _w731_ ;
	assign \g12016/_0_  = _w748_ ;
	assign \g12038/_0_  = _w751_ ;
	assign \g12039/_0_  = _w766_ ;
	assign \g12094/_0_  = _w889_ ;
	assign \g12100/_0_  = _w777_ ;
	assign \g12132/_0_  = _w1022_ ;
	assign \g12151/_0_  = _w1032_ ;
	assign \g12251/_0_  = _w1041_ ;
	assign \g12279/_0_  = _w1049_ ;
	assign \g12288/_0_  = _w984_ ;
	assign \g12290/_0_  = _w1060_ ;
	assign \g12311/_0_  = _w1063_ ;
	assign \g12313/_0_  = _w1070_ ;
	assign \g12356/_0_  = _w1079_ ;
	assign \g12357/_0_  = _w1082_ ;
	assign \g12427/_0_  = _w1196_ ;
	assign \g12441/_0_  = _w1199_ ;
	assign \g12442/_0_  = _w1209_ ;
	assign \g12480/_0_  = _w1092_ ;
	assign \g12485/_0_  = _w1095_ ;
	assign \g12506/_0_  = _w892_ ;
	assign \g12544/_0_  = _w1218_ ;
	assign \g12549/_2_  = _w1225_ ;
	assign \g12614/_0_  = _w1338_ ;
	assign \g12678/_0_  = _w1123_ ;
	assign \g12680/_0_  = _w1120_ ;
	assign \g12748/_0_  = _w1347_ ;
	assign \g15/_0_  = _w1355_ ;
	assign \g25/_0_  = _w1294_ ;
	assign \g31/_0_  = _w1405_ ;
	assign \g6843/_0_  = _w1494_ ;
	assign \g6861/_0_  = _w1532_ ;
	assign \g6863/_0_  = _w1615_ ;
	assign \g6865/_0_  = _w1693_ ;
	assign \g6887/_0_  = _w1744_ ;
	assign \g6888/_0_  = _w1781_ ;
	assign \g6889/_0_  = _w1816_ ;
	assign \g6890/_0_  = _w1851_ ;
	assign \g6891/_0_  = _w1953_ ;
	assign \g6892/_0_  = _w1992_ ;
	assign \g6893/_0_  = _w2034_ ;
	assign \g6894/_0_  = _w2069_ ;
	assign \g6922/_0_  = _w2105_ ;
	assign \g6923/_0_  = _w2146_ ;
	assign \g6924/_3_  = _w2173_ ;
	assign \g6926/_0_  = _w2205_ ;
	assign \g6927/_0_  = _w2242_ ;
	assign \g6928/_0_  = _w2274_ ;
	assign \g6931/_0_  = _w2311_ ;
	assign \g6933/_0_  = _w2344_ ;
	assign \g6967/_0_  = _w2371_ ;
	assign \g6968/_0_  = _w2402_ ;
	assign \g6969/_0_  = _w2430_ ;
	assign \g6974/_0_  = _w2455_ ;
	assign \g6975/_0_  = _w2494_ ;
	assign \g6976/_3_  = _w2531_ ;
	assign \g7006/_3_  = _w2560_ ;
	assign \g8882/_0_  = _w1859_ ;
	assign \g8883/_0_  = _w2568_ ;
	assign \g8884/_0_  = _w2576_ ;
	assign \g8895/_0_  = _w856_ ;
	assign \g8896/_0_  = _w2584_ ;
	assign \g8898/_0_  = _w793_ ;
	assign \g8900/_2_  = _w981_ ;
	assign \g8902/_0_  = _w2592_ ;
	assign \g8907/_0_  = _w1251_ ;
	assign \g8911/_0_  = _w2599_ ;
	assign \g8924/_0_  = _w2608_ ;
	assign \g8927/_0_  = _w1547_ ;
	assign \g8929/_2_  = _w1413_ ;
	assign \g8967/_0_  = _w955_ ;
	assign \g8969/_0_  = _w1880_ ;
	assign \g8973/_2_  = _w816_ ;
	assign \g8987/_0_  = _w1233_ ;
	assign \g8989/_0_  = _w2616_ ;
	assign \g8991/_0_  = _w930_ ;
	assign \g8996/_0_  = _w2623_ ;
	assign \g9099/_0_  = _w2629_ ;
	assign \g9543/_1_  = _w2631_ ;
	assign \g9751/_1_  = _w2633_ ;
	assign \g9755/_0_  = _w2635_ ;
	assign \g9786/_0_  = _w1437_ ;
	assign \g9794/_0_  = _w933_ ;
	assign \g9817/_0_  = _w1266_ ;
	assign \g9836/_0_  = _w1155_ ;
	assign \g9859/_0_  = _w905_ ;
	assign \g9862/_0_  = _w819_ ;
	assign \g9867/_0_  = _w1429_ ;
	assign \g9869/_0_  = _w1883_ ;
	assign \g9876/_0_  = _w1297_ ;
	assign \g9887/_0_  = _w796_ ;
	assign \g9895/_0_  = _w859_ ;
	assign \g9897/_0_  = _w780_ ;
	assign \g9908/_0_  = _w1236_ ;
	assign \g9910/_0_  = _w1632_ ;
	assign \g9915/_0_  = _w1254_ ;
	assign \g9938/_0_  = _w898_ ;
	assign \g9970/_0_  = _w1862_ ;
endmodule;