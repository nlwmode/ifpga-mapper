module top (\G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G18_pad , \G19_pad , \G20_pad , \G22_pad , \G23_pad , \G24_pad , \G25_pad , \G26_pad , \G28_pad , \G2_pad , \G30_pad , \G31_pad , \G32_pad , \G33_pad , \G34_pad , \G35_pad , \G3_pad , \G4_pad , \G5_pad , \G64_reg/NET0131 , \G65_reg/NET0131 , \G66_reg/NET0131 , \G69_reg/NET0131 , \G6_pad , \G70_reg/NET0131 , \G71_reg/NET0131 , \G72_reg/NET0131 , \G73_reg/NET0131 , \G74_reg/NET0131 , \G75_reg/NET0131 , \G76_reg/NET0131 , \G77_reg/NET0131 , \G79_reg/NET0131 , \G81_reg/NET0131 , \G8_pad , \G9_pad , \G100BF_pad , \G103BF_pad , \G104BF_pad , \G105BF_pad , \G107_pad , \G83_pad , \G84_pad , \G86BF_pad , \G87BF_pad , \G88BF_pad , \G89BF_pad , \G90_pad , \G95BF_pad , \G96BF_pad , \G97BF_pad , \G98BF_pad , \G99BF_pad , \_al_n0 , \_al_n1 , \g1049/_0_ , \g1081/_0_ , \g1115/_0_ , \g13/_1_ , \g809/_0_ , \g810/_0_ , \g814/_0_ , \g825/_2_ , \g834/_0_ , \g863/_0_ , \g870/_0_ , \g871/_0_ , \g916/_0_ , \g917/_0_ , \g940/_3_ );
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G18_pad  ;
	input \G19_pad  ;
	input \G20_pad  ;
	input \G22_pad  ;
	input \G23_pad  ;
	input \G24_pad  ;
	input \G25_pad  ;
	input \G26_pad  ;
	input \G28_pad  ;
	input \G2_pad  ;
	input \G30_pad  ;
	input \G31_pad  ;
	input \G32_pad  ;
	input \G33_pad  ;
	input \G34_pad  ;
	input \G35_pad  ;
	input \G3_pad  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G64_reg/NET0131  ;
	input \G65_reg/NET0131  ;
	input \G66_reg/NET0131  ;
	input \G69_reg/NET0131  ;
	input \G6_pad  ;
	input \G70_reg/NET0131  ;
	input \G71_reg/NET0131  ;
	input \G72_reg/NET0131  ;
	input \G73_reg/NET0131  ;
	input \G74_reg/NET0131  ;
	input \G75_reg/NET0131  ;
	input \G76_reg/NET0131  ;
	input \G77_reg/NET0131  ;
	input \G79_reg/NET0131  ;
	input \G81_reg/NET0131  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G100BF_pad  ;
	output \G103BF_pad  ;
	output \G104BF_pad  ;
	output \G105BF_pad  ;
	output \G107_pad  ;
	output \G83_pad  ;
	output \G84_pad  ;
	output \G86BF_pad  ;
	output \G87BF_pad  ;
	output \G88BF_pad  ;
	output \G89BF_pad  ;
	output \G90_pad  ;
	output \G95BF_pad  ;
	output \G96BF_pad  ;
	output \G97BF_pad  ;
	output \G98BF_pad  ;
	output \G99BF_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1049/_0_  ;
	output \g1081/_0_  ;
	output \g1115/_0_  ;
	output \g13/_1_  ;
	output \g809/_0_  ;
	output \g810/_0_  ;
	output \g814/_0_  ;
	output \g825/_2_  ;
	output \g834/_0_  ;
	output \g863/_0_  ;
	output \g870/_0_  ;
	output \g871/_0_  ;
	output \g916/_0_  ;
	output \g917/_0_  ;
	output \g940/_3_  ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\G4_pad ,
		\G69_reg/NET0131 ,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\G35_pad ,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\G2_pad ,
		\G66_reg/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\G10_pad ,
		\G13_pad ,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\G3_pad ,
		\G9_pad ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\G11_pad ,
		\G3_pad ,
		_w50_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\G24_pad ,
		_w46_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w49_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\G3_pad ,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\G77_reg/NET0131 ,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\G10_pad ,
		\G13_pad ,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\G3_pad ,
		\G9_pad ,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w56_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\G23_pad ,
		\G65_reg/NET0131 ,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w50_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w58_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\G3_pad ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\G76_reg/NET0131 ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\G2_pad ,
		\G64_reg/NET0131 ,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w63_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w55_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		\G9_pad ,
		_w47_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\G11_pad ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\G3_pad ,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\G22_pad ,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w66_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\G3_pad ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\G75_reg/NET0131 ,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\G14_pad ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\G15_pad ,
		_w63_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\G16_pad ,
		_w55_,
		_w76_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\G18_pad ,
		\G4_pad ,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\G79_reg/NET0131 ,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		\G19_pad ,
		\G4_pad ,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		\G65_reg/NET0131 ,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		\G20_pad ,
		\G4_pad ,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\G81_reg/NET0131 ,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w48_,
		_w56_,
		_w83_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\G25_pad ,
		_w50_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		\G4_pad ,
		\G71_reg/NET0131 ,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\G72_reg/NET0131 ,
		_w61_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		\G9_pad ,
		_w56_,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w86_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w87_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\G70_reg/NET0131 ,
		_w53_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\G9_pad ,
		_w44_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w47_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w91_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\G74_reg/NET0131 ,
		_w71_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		\G4_pad ,
		\G73_reg/NET0131 ,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w67_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w95_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\G12_pad ,
		\G26_pad ,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w90_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		_w94_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w98_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\G30_pad ,
		_w95_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\G31_pad ,
		_w96_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\G32_pad ,
		_w87_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\G33_pad ,
		_w86_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\G34_pad ,
		_w91_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\G2_pad ,
		_w55_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w63_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w71_,
		_w96_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w95_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\G2_pad ,
		\G5_pad ,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		_w63_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\G5_pad ,
		_w86_,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w87_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w55_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w73_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w113_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		\G2_pad ,
		\G6_pad ,
		_w119_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		_w55_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\G6_pad ,
		_w44_,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		_w63_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w91_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w73_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w120_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\G2_pad ,
		\G8_pad ,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		_w73_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\G8_pad ,
		_w96_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w63_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w55_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w95_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w127_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w63_,
		_w108_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w73_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w95_,
		_w96_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\G2_pad ,
		_w55_,
		_w136_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		_w44_,
		_w53_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w91_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w44_,
		_w91_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		_w86_,
		_w87_,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w61_,
		_w86_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w87_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\G11_pad ,
		\G12_pad ,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\G13_pad ,
		\G28_pad ,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w143_,
		_w144_,
		_w145_
	);
	assign \G100BF_pad  = _w45_ ;
	assign \G103BF_pad  = _w74_ ;
	assign \G104BF_pad  = _w75_ ;
	assign \G105BF_pad  = _w76_ ;
	assign \G107_pad  = _w78_ ;
	assign \G83_pad  = _w80_ ;
	assign \G84_pad  = _w82_ ;
	assign \G86BF_pad  = _w71_ ;
	assign \G87BF_pad  = _w61_ ;
	assign \G88BF_pad  = _w53_ ;
	assign \G89BF_pad  = _w85_ ;
	assign \G90_pad  = _w102_ ;
	assign \G95BF_pad  = _w103_ ;
	assign \G96BF_pad  = _w104_ ;
	assign \G97BF_pad  = _w105_ ;
	assign \G98BF_pad  = _w106_ ;
	assign \G99BF_pad  = _w107_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1049/_0_  = _w109_ ;
	assign \g1081/_0_  = _w73_ ;
	assign \g1115/_0_  = _w111_ ;
	assign \g13/_1_  = _w55_ ;
	assign \g809/_0_  = _w118_ ;
	assign \g810/_0_  = _w125_ ;
	assign \g814/_0_  = _w132_ ;
	assign \g825/_2_  = _w134_ ;
	assign \g834/_0_  = _w135_ ;
	assign \g863/_0_  = _w136_ ;
	assign \g870/_0_  = _w138_ ;
	assign \g871/_0_  = _w139_ ;
	assign \g916/_0_  = _w140_ ;
	assign \g917/_0_  = _w142_ ;
	assign \g940/_3_  = _w145_ ;
endmodule;