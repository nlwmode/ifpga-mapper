module top (\a0_pad , a_pad, \b0_pad , b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, \l0_pad , l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \d0_pad , \e0_pad , \f0_pad , \g0_pad , \h0_pad , \i0_pad , \j0_pad , \k0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , \u0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input \l0_pad  ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \d0_pad  ;
	output \e0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \h0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output \u0_pad  ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\l0_pad ,
		u_pad,
		_w29_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		i_pad,
		\l0_pad ,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w29_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\l0_pad ,
		v_pad,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		j_pad,
		\l0_pad ,
		_w33_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w32_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\l0_pad ,
		w_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		k_pad,
		\l0_pad ,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\l0_pad ,
		x_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		\l0_pad ,
		l_pad,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w38_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\l0_pad ,
		y_pad,
		_w41_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\l0_pad ,
		m_pad,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w41_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\l0_pad ,
		z_pad,
		_w44_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\l0_pad ,
		n_pad,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\a0_pad ,
		\l0_pad ,
		_w47_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\l0_pad ,
		o_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\b0_pad ,
		\l0_pad ,
		_w50_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\l0_pad ,
		p_pad,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		q_pad,
		s_pad,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		i_pad,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		r_pad,
		u_pad,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		q_pad,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		q_pad,
		s_pad,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		a_pad,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		q_pad,
		r_pad,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		u_pad,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w54_,
		_w56_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w58_,
		_w60_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w61_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		j_pad,
		_w53_,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		b_pad,
		_w57_,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		v_pad,
		_w55_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		v_pad,
		_w55_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		q_pad,
		_w66_,
		_w68_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w64_,
		_w65_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w69_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		k_pad,
		s_pad,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		c_pad,
		s_pad,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		q_pad,
		_w72_,
		_w74_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		w_pad,
		_w66_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		v_pad,
		w_pad,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w55_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		q_pad,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w76_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w75_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		x_pad,
		_w78_,
		_w82_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		x_pad,
		_w78_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		q_pad,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		l_pad,
		s_pad,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		d_pad,
		s_pad,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		q_pad,
		_w86_,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w87_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w85_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		m_pad,
		s_pad,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		e_pad,
		s_pad,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		q_pad,
		_w91_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w92_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		y_pad,
		_w82_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		y_pad,
		_w82_,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		q_pad,
		_w95_,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w94_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		n_pad,
		s_pad,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		f_pad,
		s_pad,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		q_pad,
		_w100_,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		_w101_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		z_pad,
		_w96_,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		x_pad,
		y_pad,
		_w105_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		z_pad,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w78_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		q_pad,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w104_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w103_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\a0_pad ,
		_w107_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		\a0_pad ,
		_w107_,
		_w112_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w111_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		q_pad,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		o_pad,
		s_pad,
		_w115_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		g_pad,
		s_pad,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		q_pad,
		_w115_,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w116_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w114_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		\a0_pad ,
		\b0_pad ,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		y_pad,
		z_pad,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w82_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		\b0_pad ,
		_w112_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		q_pad,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		p_pad,
		s_pad,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		h_pad,
		s_pad,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		q_pad,
		_w127_,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w128_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w126_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		\l0_pad ,
		r_pad,
		_w132_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\a0_pad ,
		u_pad,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w77_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w106_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		_w122_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		r_pad,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		q_pad,
		_w132_,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w137_,
		_w138_,
		_w139_
	);
	assign \d0_pad  = _w31_ ;
	assign \e0_pad  = _w34_ ;
	assign \f0_pad  = _w37_ ;
	assign \g0_pad  = _w40_ ;
	assign \h0_pad  = _w43_ ;
	assign \i0_pad  = _w46_ ;
	assign \j0_pad  = _w49_ ;
	assign \k0_pad  = _w52_ ;
	assign \m0_pad  = _w63_ ;
	assign \n0_pad  = _w71_ ;
	assign \o0_pad  = _w81_ ;
	assign \p0_pad  = _w90_ ;
	assign \q0_pad  = _w99_ ;
	assign \r0_pad  = _w110_ ;
	assign \s0_pad  = _w119_ ;
	assign \t0_pad  = _w131_ ;
	assign \u0_pad  = _w139_ ;
endmodule;