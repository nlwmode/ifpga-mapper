module top( decrypt_pad , \key1[0]_pad  , \key1[10]_pad  , \key1[11]_pad  , \key1[12]_pad  , \key1[13]_pad  , \key1[14]_pad  , \key1[15]_pad  , \key1[16]_pad  , \key1[17]_pad  , \key1[18]_pad  , \key1[19]_pad  , \key1[1]_pad  , \key1[20]_pad  , \key1[21]_pad  , \key1[22]_pad  , \key1[23]_pad  , \key1[24]_pad  , \key1[25]_pad  , \key1[26]_pad  , \key1[27]_pad  , \key1[28]_pad  , \key1[29]_pad  , \key1[2]_pad  , \key1[30]_pad  , \key1[31]_pad  , \key1[32]_pad  , \key1[33]_pad  , \key1[34]_pad  , \key1[35]_pad  , \key1[36]_pad  , \key1[37]_pad  , \key1[38]_pad  , \key1[39]_pad  , \key1[3]_pad  , \key1[40]_pad  , \key1[41]_pad  , \key1[42]_pad  , \key1[43]_pad  , \key1[44]_pad  , \key1[45]_pad  , \key1[46]_pad  , \key1[47]_pad  , \key1[48]_pad  , \key1[49]_pad  , \key1[4]_pad  , \key1[50]_pad  , \key1[51]_pad  , \key1[52]_pad  , \key1[53]_pad  , \key1[54]_pad  , \key1[55]_pad  , \key1[5]_pad  , \key1[6]_pad  , \key1[7]_pad  , \key1[8]_pad  , \key1[9]_pad  , \key3[0]_pad  , \key3[10]_pad  , \key3[11]_pad  , \key3[12]_pad  , \key3[13]_pad  , \key3[14]_pad  , \key3[15]_pad  , \key3[16]_pad  , \key3[17]_pad  , \key3[18]_pad  , \key3[19]_pad  , \key3[1]_pad  , \key3[20]_pad  , \key3[21]_pad  , \key3[22]_pad  , \key3[23]_pad  , \key3[24]_pad  , \key3[25]_pad  , \key3[26]_pad  , \key3[27]_pad  , \key3[28]_pad  , \key3[29]_pad  , \key3[2]_pad  , \key3[30]_pad  , \key3[31]_pad  , \key3[32]_pad  , \key3[33]_pad  , \key3[34]_pad  , \key3[35]_pad  , \key3[36]_pad  , \key3[37]_pad  , \key3[38]_pad  , \key3[39]_pad  , \key3[3]_pad  , \key3[40]_pad  , \key3[41]_pad  , \key3[42]_pad  , \key3[43]_pad  , \key3[44]_pad  , \key3[45]_pad  , \key3[46]_pad  , \key3[47]_pad  , \key3[48]_pad  , \key3[49]_pad  , \key3[4]_pad  , \key3[50]_pad  , \key3[51]_pad  , \key3[52]_pad  , \key3[53]_pad  , \key3[54]_pad  , \key3[55]_pad  , \key3[5]_pad  , \key3[6]_pad  , \key3[7]_pad  , \key3[8]_pad  , \key3[9]_pad  , \u0_L0_reg[10]/NET0131  , \u0_L0_reg[11]/NET0131  , \u0_L0_reg[12]/NET0131  , \u0_L0_reg[13]/NET0131  , \u0_L0_reg[14]/NET0131  , \u0_L0_reg[15]/P0001  , \u0_L0_reg[16]/NET0131  , \u0_L0_reg[17]/NET0131  , \u0_L0_reg[18]/NET0131  , \u0_L0_reg[19]/P0001  , \u0_L0_reg[1]/NET0131  , \u0_L0_reg[20]/NET0131  , \u0_L0_reg[21]/NET0131  , \u0_L0_reg[22]/NET0131  , \u0_L0_reg[23]/NET0131  , \u0_L0_reg[24]/NET0131  , \u0_L0_reg[25]/NET0131  , \u0_L0_reg[26]/NET0131  , \u0_L0_reg[27]/NET0131  , \u0_L0_reg[28]/NET0131  , \u0_L0_reg[29]/NET0131  , \u0_L0_reg[2]/NET0131  , \u0_L0_reg[30]/P0001  , \u0_L0_reg[31]/NET0131  , \u0_L0_reg[32]/NET0131  , \u0_L0_reg[3]/NET0131  , \u0_L0_reg[4]/NET0131  , \u0_L0_reg[5]/NET0131  , \u0_L0_reg[6]/NET0131  , \u0_L0_reg[7]/NET0131  , \u0_L0_reg[8]/NET0131  , \u0_L0_reg[9]/NET0131  , \u0_L10_reg[10]/NET0131  , \u0_L10_reg[11]/NET0131  , \u0_L10_reg[12]/NET0131  , \u0_L10_reg[13]/NET0131  , \u0_L10_reg[14]/NET0131  , \u0_L10_reg[15]/P0001  , \u0_L10_reg[16]/NET0131  , \u0_L10_reg[17]/NET0131  , \u0_L10_reg[18]/NET0131  , \u0_L10_reg[19]/NET0131  , \u0_L10_reg[1]/NET0131  , \u0_L10_reg[20]/NET0131  , \u0_L10_reg[21]/NET0131  , \u0_L10_reg[22]/NET0131  , \u0_L10_reg[23]/NET0131  , \u0_L10_reg[24]/NET0131  , \u0_L10_reg[25]/NET0131  , \u0_L10_reg[26]/NET0131  , \u0_L10_reg[27]/NET0131  , \u0_L10_reg[28]/NET0131  , \u0_L10_reg[29]/NET0131  , \u0_L10_reg[2]/NET0131  , \u0_L10_reg[30]/NET0131  , \u0_L10_reg[31]/NET0131  , \u0_L10_reg[32]/NET0131  , \u0_L10_reg[3]/NET0131  , \u0_L10_reg[4]/NET0131  , \u0_L10_reg[5]/NET0131  , \u0_L10_reg[6]/NET0131  , \u0_L10_reg[7]/NET0131  , \u0_L10_reg[8]/NET0131  , \u0_L10_reg[9]/NET0131  , \u0_L11_reg[10]/NET0131  , \u0_L11_reg[11]/P0001  , \u0_L11_reg[12]/NET0131  , \u0_L11_reg[13]/NET0131  , \u0_L11_reg[14]/NET0131  , \u0_L11_reg[15]/P0001  , \u0_L11_reg[16]/NET0131  , \u0_L11_reg[17]/NET0131  , \u0_L11_reg[18]/NET0131  , \u0_L11_reg[19]/NET0131  , \u0_L11_reg[1]/NET0131  , \u0_L11_reg[20]/NET0131  , \u0_L11_reg[21]/NET0131  , \u0_L11_reg[22]/NET0131  , \u0_L11_reg[23]/NET0131  , \u0_L11_reg[24]/NET0131  , \u0_L11_reg[25]/NET0131  , \u0_L11_reg[26]/NET0131  , \u0_L11_reg[27]/NET0131  , \u0_L11_reg[28]/NET0131  , \u0_L11_reg[29]/NET0131  , \u0_L11_reg[2]/NET0131  , \u0_L11_reg[30]/NET0131  , \u0_L11_reg[31]/NET0131  , \u0_L11_reg[32]/NET0131  , \u0_L11_reg[3]/NET0131  , \u0_L11_reg[4]/NET0131  , \u0_L11_reg[5]/NET0131  , \u0_L11_reg[6]/NET0131  , \u0_L11_reg[7]/NET0131  , \u0_L11_reg[8]/NET0131  , \u0_L11_reg[9]/NET0131  , \u0_L12_reg[10]/NET0131  , \u0_L12_reg[11]/NET0131  , \u0_L12_reg[12]/NET0131  , \u0_L12_reg[13]/NET0131  , \u0_L12_reg[14]/NET0131  , \u0_L12_reg[15]/P0001  , \u0_L12_reg[16]/NET0131  , \u0_L12_reg[17]/NET0131  , \u0_L12_reg[18]/NET0131  , \u0_L12_reg[19]/P0001  , \u0_L12_reg[1]/NET0131  , \u0_L12_reg[20]/NET0131  , \u0_L12_reg[21]/NET0131  , \u0_L12_reg[22]/NET0131  , \u0_L12_reg[23]/NET0131  , \u0_L12_reg[24]/NET0131  , \u0_L12_reg[25]/NET0131  , \u0_L12_reg[26]/NET0131  , \u0_L12_reg[27]/NET0131  , \u0_L12_reg[28]/NET0131  , \u0_L12_reg[29]/NET0131  , \u0_L12_reg[2]/NET0131  , \u0_L12_reg[30]/NET0131  , \u0_L12_reg[31]/NET0131  , \u0_L12_reg[32]/NET0131  , \u0_L12_reg[3]/NET0131  , \u0_L12_reg[4]/NET0131  , \u0_L12_reg[5]/NET0131  , \u0_L12_reg[6]/NET0131  , \u0_L12_reg[7]/NET0131  , \u0_L12_reg[8]/NET0131  , \u0_L12_reg[9]/NET0131  , \u0_L13_reg[10]/NET0131  , \u0_L13_reg[11]/NET0131  , \u0_L13_reg[12]/NET0131  , \u0_L13_reg[13]/NET0131  , \u0_L13_reg[14]/NET0131  , \u0_L13_reg[15]/P0001  , \u0_L13_reg[16]/NET0131  , \u0_L13_reg[17]/NET0131  , \u0_L13_reg[18]/NET0131  , \u0_L13_reg[19]/NET0131  , \u0_L13_reg[1]/NET0131  , \u0_L13_reg[20]/NET0131  , \u0_L13_reg[21]/NET0131  , \u0_L13_reg[22]/NET0131  , \u0_L13_reg[23]/NET0131  , \u0_L13_reg[24]/NET0131  , \u0_L13_reg[25]/NET0131  , \u0_L13_reg[26]/NET0131  , \u0_L13_reg[27]/NET0131  , \u0_L13_reg[28]/NET0131  , \u0_L13_reg[29]/NET0131  , \u0_L13_reg[2]/NET0131  , \u0_L13_reg[30]/NET0131  , \u0_L13_reg[31]/NET0131  , \u0_L13_reg[32]/NET0131  , \u0_L13_reg[3]/NET0131  , \u0_L13_reg[4]/NET0131  , \u0_L13_reg[5]/NET0131  , \u0_L13_reg[6]/NET0131  , \u0_L13_reg[7]/NET0131  , \u0_L13_reg[8]/NET0131  , \u0_L13_reg[9]/NET0131  , \u0_L14_reg[10]/P0001  , \u0_L14_reg[11]/P0001  , \u0_L14_reg[12]/P0001  , \u0_L14_reg[13]/P0001  , \u0_L14_reg[14]/P0001  , \u0_L14_reg[15]/P0001  , \u0_L14_reg[16]/P0001  , \u0_L14_reg[17]/P0001  , \u0_L14_reg[18]/P0001  , \u0_L14_reg[19]/P0001  , \u0_L14_reg[1]/P0001  , \u0_L14_reg[20]/P0001  , \u0_L14_reg[21]/P0001  , \u0_L14_reg[22]/P0001  , \u0_L14_reg[23]/P0001  , \u0_L14_reg[24]/P0001  , \u0_L14_reg[25]/P0001  , \u0_L14_reg[26]/P0001  , \u0_L14_reg[27]/P0001  , \u0_L14_reg[28]/P0001  , \u0_L14_reg[29]/P0001  , \u0_L14_reg[2]/P0001  , \u0_L14_reg[30]/P0001  , \u0_L14_reg[31]/P0001  , \u0_L14_reg[32]/P0001  , \u0_L14_reg[3]/P0001  , \u0_L14_reg[4]/P0001  , \u0_L14_reg[5]/P0001  , \u0_L14_reg[6]/P0001  , \u0_L14_reg[7]/P0001  , \u0_L14_reg[8]/P0001  , \u0_L14_reg[9]/P0001  , \u0_L1_reg[10]/NET0131  , \u0_L1_reg[11]/NET0131  , \u0_L1_reg[12]/NET0131  , \u0_L1_reg[13]/NET0131  , \u0_L1_reg[14]/NET0131  , \u0_L1_reg[15]/P0001  , \u0_L1_reg[16]/NET0131  , \u0_L1_reg[17]/NET0131  , \u0_L1_reg[18]/NET0131  , \u0_L1_reg[19]/NET0131  , \u0_L1_reg[1]/NET0131  , \u0_L1_reg[20]/NET0131  , \u0_L1_reg[21]/NET0131  , \u0_L1_reg[22]/NET0131  , \u0_L1_reg[23]/NET0131  , \u0_L1_reg[24]/NET0131  , \u0_L1_reg[25]/NET0131  , \u0_L1_reg[26]/NET0131  , \u0_L1_reg[27]/NET0131  , \u0_L1_reg[28]/NET0131  , \u0_L1_reg[29]/NET0131  , \u0_L1_reg[2]/NET0131  , \u0_L1_reg[30]/NET0131  , \u0_L1_reg[31]/NET0131  , \u0_L1_reg[32]/NET0131  , \u0_L1_reg[3]/NET0131  , \u0_L1_reg[4]/NET0131  , \u0_L1_reg[5]/NET0131  , \u0_L1_reg[6]/NET0131  , \u0_L1_reg[7]/NET0131  , \u0_L1_reg[8]/NET0131  , \u0_L1_reg[9]/NET0131  , \u0_L2_reg[10]/NET0131  , \u0_L2_reg[11]/NET0131  , \u0_L2_reg[12]/NET0131  , \u0_L2_reg[13]/NET0131  , \u0_L2_reg[14]/NET0131  , \u0_L2_reg[15]/P0001  , \u0_L2_reg[16]/NET0131  , \u0_L2_reg[17]/NET0131  , \u0_L2_reg[18]/NET0131  , \u0_L2_reg[19]/P0001  , \u0_L2_reg[1]/NET0131  , \u0_L2_reg[20]/NET0131  , \u0_L2_reg[21]/NET0131  , \u0_L2_reg[22]/NET0131  , \u0_L2_reg[23]/NET0131  , \u0_L2_reg[24]/NET0131  , \u0_L2_reg[25]/NET0131  , \u0_L2_reg[26]/NET0131  , \u0_L2_reg[27]/NET0131  , \u0_L2_reg[28]/NET0131  , \u0_L2_reg[29]/NET0131  , \u0_L2_reg[2]/NET0131  , \u0_L2_reg[30]/NET0131  , \u0_L2_reg[31]/NET0131  , \u0_L2_reg[32]/NET0131  , \u0_L2_reg[3]/NET0131  , \u0_L2_reg[4]/NET0131  , \u0_L2_reg[5]/NET0131  , \u0_L2_reg[6]/NET0131  , \u0_L2_reg[7]/NET0131  , \u0_L2_reg[8]/NET0131  , \u0_L2_reg[9]/NET0131  , \u0_L3_reg[10]/NET0131  , \u0_L3_reg[11]/NET0131  , \u0_L3_reg[12]/NET0131  , \u0_L3_reg[13]/NET0131  , \u0_L3_reg[14]/NET0131  , \u0_L3_reg[15]/P0001  , \u0_L3_reg[16]/NET0131  , \u0_L3_reg[17]/NET0131  , \u0_L3_reg[18]/NET0131  , \u0_L3_reg[19]/P0001  , \u0_L3_reg[1]/NET0131  , \u0_L3_reg[20]/NET0131  , \u0_L3_reg[21]/NET0131  , \u0_L3_reg[22]/NET0131  , \u0_L3_reg[23]/NET0131  , \u0_L3_reg[24]/NET0131  , \u0_L3_reg[25]/NET0131  , \u0_L3_reg[26]/NET0131  , \u0_L3_reg[27]/NET0131  , \u0_L3_reg[28]/NET0131  , \u0_L3_reg[29]/NET0131  , \u0_L3_reg[2]/NET0131  , \u0_L3_reg[30]/NET0131  , \u0_L3_reg[31]/NET0131  , \u0_L3_reg[32]/NET0131  , \u0_L3_reg[3]/NET0131  , \u0_L3_reg[4]/NET0131  , \u0_L3_reg[5]/NET0131  , \u0_L3_reg[6]/NET0131  , \u0_L3_reg[7]/NET0131  , \u0_L3_reg[8]/NET0131  , \u0_L3_reg[9]/NET0131  , \u0_L4_reg[10]/NET0131  , \u0_L4_reg[11]/NET0131  , \u0_L4_reg[12]/NET0131  , \u0_L4_reg[13]/NET0131  , \u0_L4_reg[14]/NET0131  , \u0_L4_reg[15]/P0001  , \u0_L4_reg[16]/NET0131  , \u0_L4_reg[17]/NET0131  , \u0_L4_reg[18]/NET0131  , \u0_L4_reg[19]/NET0131  , \u0_L4_reg[1]/NET0131  , \u0_L4_reg[20]/NET0131  , \u0_L4_reg[21]/NET0131  , \u0_L4_reg[22]/NET0131  , \u0_L4_reg[23]/NET0131  , \u0_L4_reg[24]/NET0131  , \u0_L4_reg[25]/NET0131  , \u0_L4_reg[26]/NET0131  , \u0_L4_reg[27]/NET0131  , \u0_L4_reg[28]/NET0131  , \u0_L4_reg[29]/NET0131  , \u0_L4_reg[2]/NET0131  , \u0_L4_reg[30]/NET0131  , \u0_L4_reg[31]/NET0131  , \u0_L4_reg[32]/NET0131  , \u0_L4_reg[3]/NET0131  , \u0_L4_reg[4]/NET0131  , \u0_L4_reg[5]/NET0131  , \u0_L4_reg[6]/NET0131  , \u0_L4_reg[7]/NET0131  , \u0_L4_reg[8]/NET0131  , \u0_L4_reg[9]/NET0131  , \u0_L5_reg[10]/NET0131  , \u0_L5_reg[11]/NET0131  , \u0_L5_reg[12]/NET0131  , \u0_L5_reg[13]/NET0131  , \u0_L5_reg[14]/NET0131  , \u0_L5_reg[15]/P0001  , \u0_L5_reg[16]/NET0131  , \u0_L5_reg[17]/NET0131  , \u0_L5_reg[18]/NET0131  , \u0_L5_reg[19]/P0001  , \u0_L5_reg[1]/NET0131  , \u0_L5_reg[20]/NET0131  , \u0_L5_reg[21]/NET0131  , \u0_L5_reg[22]/NET0131  , \u0_L5_reg[23]/NET0131  , \u0_L5_reg[24]/NET0131  , \u0_L5_reg[25]/NET0131  , \u0_L5_reg[26]/NET0131  , \u0_L5_reg[27]/NET0131  , \u0_L5_reg[28]/NET0131  , \u0_L5_reg[29]/NET0131  , \u0_L5_reg[2]/NET0131  , \u0_L5_reg[30]/NET0131  , \u0_L5_reg[31]/NET0131  , \u0_L5_reg[32]/NET0131  , \u0_L5_reg[3]/NET0131  , \u0_L5_reg[4]/NET0131  , \u0_L5_reg[5]/NET0131  , \u0_L5_reg[6]/NET0131  , \u0_L5_reg[7]/NET0131  , \u0_L5_reg[8]/NET0131  , \u0_L5_reg[9]/NET0131  , \u0_L6_reg[10]/NET0131  , \u0_L6_reg[11]/NET0131  , \u0_L6_reg[12]/NET0131  , \u0_L6_reg[13]/NET0131  , \u0_L6_reg[14]/NET0131  , \u0_L6_reg[15]/P0001  , \u0_L6_reg[16]/NET0131  , \u0_L6_reg[17]/NET0131  , \u0_L6_reg[18]/NET0131  , \u0_L6_reg[19]/P0001  , \u0_L6_reg[1]/NET0131  , \u0_L6_reg[20]/NET0131  , \u0_L6_reg[21]/NET0131  , \u0_L6_reg[22]/NET0131  , \u0_L6_reg[23]/NET0131  , \u0_L6_reg[24]/NET0131  , \u0_L6_reg[25]/NET0131  , \u0_L6_reg[26]/NET0131  , \u0_L6_reg[27]/NET0131  , \u0_L6_reg[28]/NET0131  , \u0_L6_reg[29]/NET0131  , \u0_L6_reg[2]/NET0131  , \u0_L6_reg[30]/NET0131  , \u0_L6_reg[31]/NET0131  , \u0_L6_reg[32]/NET0131  , \u0_L6_reg[3]/NET0131  , \u0_L6_reg[4]/NET0131  , \u0_L6_reg[5]/NET0131  , \u0_L6_reg[6]/NET0131  , \u0_L6_reg[7]/NET0131  , \u0_L6_reg[8]/NET0131  , \u0_L6_reg[9]/NET0131  , \u0_L7_reg[10]/NET0131  , \u0_L7_reg[11]/NET0131  , \u0_L7_reg[12]/NET0131  , \u0_L7_reg[13]/NET0131  , \u0_L7_reg[14]/NET0131  , \u0_L7_reg[15]/P0001  , \u0_L7_reg[16]/NET0131  , \u0_L7_reg[17]/NET0131  , \u0_L7_reg[18]/NET0131  , \u0_L7_reg[19]/NET0131  , \u0_L7_reg[1]/NET0131  , \u0_L7_reg[20]/NET0131  , \u0_L7_reg[21]/NET0131  , \u0_L7_reg[22]/NET0131  , \u0_L7_reg[23]/NET0131  , \u0_L7_reg[24]/NET0131  , \u0_L7_reg[25]/NET0131  , \u0_L7_reg[26]/NET0131  , \u0_L7_reg[27]/NET0131  , \u0_L7_reg[28]/NET0131  , \u0_L7_reg[29]/NET0131  , \u0_L7_reg[2]/NET0131  , \u0_L7_reg[30]/NET0131  , \u0_L7_reg[31]/NET0131  , \u0_L7_reg[32]/NET0131  , \u0_L7_reg[3]/NET0131  , \u0_L7_reg[4]/NET0131  , \u0_L7_reg[5]/NET0131  , \u0_L7_reg[6]/NET0131  , \u0_L7_reg[7]/NET0131  , \u0_L7_reg[8]/NET0131  , \u0_L7_reg[9]/NET0131  , \u0_L8_reg[10]/NET0131  , \u0_L8_reg[11]/NET0131  , \u0_L8_reg[12]/NET0131  , \u0_L8_reg[13]/NET0131  , \u0_L8_reg[14]/NET0131  , \u0_L8_reg[15]/P0001  , \u0_L8_reg[16]/NET0131  , \u0_L8_reg[17]/NET0131  , \u0_L8_reg[18]/NET0131  , \u0_L8_reg[19]/NET0131  , \u0_L8_reg[1]/NET0131  , \u0_L8_reg[20]/NET0131  , \u0_L8_reg[21]/NET0131  , \u0_L8_reg[22]/NET0131  , \u0_L8_reg[23]/NET0131  , \u0_L8_reg[24]/NET0131  , \u0_L8_reg[25]/NET0131  , \u0_L8_reg[26]/NET0131  , \u0_L8_reg[27]/NET0131  , \u0_L8_reg[28]/NET0131  , \u0_L8_reg[29]/NET0131  , \u0_L8_reg[2]/NET0131  , \u0_L8_reg[30]/NET0131  , \u0_L8_reg[31]/NET0131  , \u0_L8_reg[32]/NET0131  , \u0_L8_reg[3]/NET0131  , \u0_L8_reg[4]/NET0131  , \u0_L8_reg[5]/NET0131  , \u0_L8_reg[6]/NET0131  , \u0_L8_reg[7]/NET0131  , \u0_L8_reg[8]/NET0131  , \u0_L8_reg[9]/NET0131  , \u0_L9_reg[10]/NET0131  , \u0_L9_reg[11]/NET0131  , \u0_L9_reg[12]/NET0131  , \u0_L9_reg[13]/NET0131  , \u0_L9_reg[14]/NET0131  , \u0_L9_reg[15]/P0001  , \u0_L9_reg[16]/NET0131  , \u0_L9_reg[17]/NET0131  , \u0_L9_reg[18]/NET0131  , \u0_L9_reg[19]/P0001  , \u0_L9_reg[1]/NET0131  , \u0_L9_reg[20]/NET0131  , \u0_L9_reg[21]/NET0131  , \u0_L9_reg[22]/NET0131  , \u0_L9_reg[23]/NET0131  , \u0_L9_reg[24]/NET0131  , \u0_L9_reg[25]/NET0131  , \u0_L9_reg[26]/NET0131  , \u0_L9_reg[27]/NET0131  , \u0_L9_reg[28]/NET0131  , \u0_L9_reg[29]/NET0131  , \u0_L9_reg[2]/NET0131  , \u0_L9_reg[30]/NET0131  , \u0_L9_reg[31]/NET0131  , \u0_L9_reg[32]/NET0131  , \u0_L9_reg[3]/NET0131  , \u0_L9_reg[4]/NET0131  , \u0_L9_reg[5]/NET0131  , \u0_L9_reg[6]/NET0131  , \u0_L9_reg[7]/NET0131  , \u0_L9_reg[8]/NET0131  , \u0_L9_reg[9]/NET0131  , \u0_R0_reg[10]/NET0131  , \u0_R0_reg[11]/NET0131  , \u0_R0_reg[12]/NET0131  , \u0_R0_reg[13]/NET0131  , \u0_R0_reg[14]/NET0131  , \u0_R0_reg[15]/NET0131  , \u0_R0_reg[16]/NET0131  , \u0_R0_reg[17]/NET0131  , \u0_R0_reg[18]/NET0131  , \u0_R0_reg[19]/NET0131  , \u0_R0_reg[1]/NET0131  , \u0_R0_reg[20]/NET0131  , \u0_R0_reg[21]/NET0131  , \u0_R0_reg[22]/NET0131  , \u0_R0_reg[23]/NET0131  , \u0_R0_reg[24]/NET0131  , \u0_R0_reg[25]/NET0131  , \u0_R0_reg[26]/NET0131  , \u0_R0_reg[27]/NET0131  , \u0_R0_reg[28]/NET0131  , \u0_R0_reg[29]/NET0131  , \u0_R0_reg[2]/NET0131  , \u0_R0_reg[30]/NET0131  , \u0_R0_reg[31]/NET0131  , \u0_R0_reg[32]/NET0131  , \u0_R0_reg[3]/NET0131  , \u0_R0_reg[4]/NET0131  , \u0_R0_reg[5]/NET0131  , \u0_R0_reg[6]/NET0131  , \u0_R0_reg[7]/NET0131  , \u0_R0_reg[8]/NET0131  , \u0_R0_reg[9]/NET0131  , \u0_R10_reg[10]/NET0131  , \u0_R10_reg[11]/NET0131  , \u0_R10_reg[12]/NET0131  , \u0_R10_reg[13]/NET0131  , \u0_R10_reg[14]/NET0131  , \u0_R10_reg[15]/NET0131  , \u0_R10_reg[16]/NET0131  , \u0_R10_reg[17]/NET0131  , \u0_R10_reg[18]/NET0131  , \u0_R10_reg[19]/NET0131  , \u0_R10_reg[1]/NET0131  , \u0_R10_reg[20]/NET0131  , \u0_R10_reg[21]/NET0131  , \u0_R10_reg[22]/NET0131  , \u0_R10_reg[23]/NET0131  , \u0_R10_reg[24]/NET0131  , \u0_R10_reg[25]/NET0131  , \u0_R10_reg[26]/NET0131  , \u0_R10_reg[27]/NET0131  , \u0_R10_reg[28]/NET0131  , \u0_R10_reg[29]/NET0131  , \u0_R10_reg[2]/NET0131  , \u0_R10_reg[30]/NET0131  , \u0_R10_reg[31]/P0001  , \u0_R10_reg[32]/NET0131  , \u0_R10_reg[3]/NET0131  , \u0_R10_reg[4]/NET0131  , \u0_R10_reg[5]/NET0131  , \u0_R10_reg[6]/NET0131  , \u0_R10_reg[7]/NET0131  , \u0_R10_reg[8]/NET0131  , \u0_R10_reg[9]/NET0131  , \u0_R11_reg[10]/NET0131  , \u0_R11_reg[11]/P0001  , \u0_R11_reg[12]/NET0131  , \u0_R11_reg[13]/NET0131  , \u0_R11_reg[14]/NET0131  , \u0_R11_reg[15]/NET0131  , \u0_R11_reg[16]/NET0131  , \u0_R11_reg[17]/NET0131  , \u0_R11_reg[18]/NET0131  , \u0_R11_reg[19]/NET0131  , \u0_R11_reg[1]/NET0131  , \u0_R11_reg[20]/NET0131  , \u0_R11_reg[21]/NET0131  , \u0_R11_reg[22]/NET0131  , \u0_R11_reg[23]/NET0131  , \u0_R11_reg[24]/NET0131  , \u0_R11_reg[25]/NET0131  , \u0_R11_reg[26]/NET0131  , \u0_R11_reg[27]/NET0131  , \u0_R11_reg[28]/NET0131  , \u0_R11_reg[29]/NET0131  , \u0_R11_reg[2]/NET0131  , \u0_R11_reg[30]/NET0131  , \u0_R11_reg[31]/P0001  , \u0_R11_reg[32]/NET0131  , \u0_R11_reg[3]/NET0131  , \u0_R11_reg[4]/NET0131  , \u0_R11_reg[5]/NET0131  , \u0_R11_reg[6]/NET0131  , \u0_R11_reg[7]/NET0131  , \u0_R11_reg[8]/NET0131  , \u0_R11_reg[9]/NET0131  , \u0_R12_reg[10]/NET0131  , \u0_R12_reg[11]/NET0131  , \u0_R12_reg[12]/NET0131  , \u0_R12_reg[13]/NET0131  , \u0_R12_reg[14]/NET0131  , \u0_R12_reg[15]/NET0131  , \u0_R12_reg[16]/NET0131  , \u0_R12_reg[17]/NET0131  , \u0_R12_reg[18]/NET0131  , \u0_R12_reg[19]/NET0131  , \u0_R12_reg[1]/NET0131  , \u0_R12_reg[20]/NET0131  , \u0_R12_reg[21]/NET0131  , \u0_R12_reg[22]/NET0131  , \u0_R12_reg[23]/NET0131  , \u0_R12_reg[24]/NET0131  , \u0_R12_reg[25]/NET0131  , \u0_R12_reg[26]/NET0131  , \u0_R12_reg[27]/NET0131  , \u0_R12_reg[28]/NET0131  , \u0_R12_reg[29]/NET0131  , \u0_R12_reg[2]/NET0131  , \u0_R12_reg[30]/NET0131  , \u0_R12_reg[31]/P0001  , \u0_R12_reg[32]/NET0131  , \u0_R12_reg[3]/NET0131  , \u0_R12_reg[4]/NET0131  , \u0_R12_reg[5]/NET0131  , \u0_R12_reg[6]/NET0131  , \u0_R12_reg[7]/NET0131  , \u0_R12_reg[8]/NET0131  , \u0_R12_reg[9]/NET0131  , \u0_R13_reg[10]/NET0131  , \u0_R13_reg[11]/NET0131  , \u0_R13_reg[12]/NET0131  , \u0_R13_reg[13]/NET0131  , \u0_R13_reg[14]/NET0131  , \u0_R13_reg[15]/NET0131  , \u0_R13_reg[16]/NET0131  , \u0_R13_reg[17]/NET0131  , \u0_R13_reg[18]/NET0131  , \u0_R13_reg[19]/NET0131  , \u0_R13_reg[1]/NET0131  , \u0_R13_reg[20]/NET0131  , \u0_R13_reg[21]/NET0131  , \u0_R13_reg[22]/P0001  , \u0_R13_reg[23]/NET0131  , \u0_R13_reg[24]/NET0131  , \u0_R13_reg[25]/NET0131  , \u0_R13_reg[26]/NET0131  , \u0_R13_reg[27]/P0001  , \u0_R13_reg[28]/NET0131  , \u0_R13_reg[29]/NET0131  , \u0_R13_reg[2]/NET0131  , \u0_R13_reg[30]/NET0131  , \u0_R13_reg[31]/NET0131  , \u0_R13_reg[32]/NET0131  , \u0_R13_reg[3]/NET0131  , \u0_R13_reg[4]/NET0131  , \u0_R13_reg[5]/NET0131  , \u0_R13_reg[6]/NET0131  , \u0_R13_reg[7]/NET0131  , \u0_R13_reg[8]/NET0131  , \u0_R13_reg[9]/NET0131  , \u0_R14_reg[10]/NET0131  , \u0_R14_reg[11]/P0001  , \u0_R14_reg[12]/NET0131  , \u0_R14_reg[13]/NET0131  , \u0_R14_reg[14]/NET0131  , \u0_R14_reg[15]/NET0131  , \u0_R14_reg[16]/NET0131  , \u0_R14_reg[17]/NET0131  , \u0_R14_reg[18]/NET0131  , \u0_R14_reg[19]/NET0131  , \u0_R14_reg[1]/NET0131  , \u0_R14_reg[20]/NET0131  , \u0_R14_reg[21]/NET0131  , \u0_R14_reg[22]/P0001  , \u0_R14_reg[23]/NET0131  , \u0_R14_reg[24]/NET0131  , \u0_R14_reg[25]/NET0131  , \u0_R14_reg[26]/P0001  , \u0_R14_reg[27]/P0001  , \u0_R14_reg[28]/NET0131  , \u0_R14_reg[29]/NET0131  , \u0_R14_reg[2]/NET0131  , \u0_R14_reg[30]/NET0131  , \u0_R14_reg[31]/P0001  , \u0_R14_reg[32]/NET0131  , \u0_R14_reg[3]/NET0131  , \u0_R14_reg[4]/NET0131  , \u0_R14_reg[5]/NET0131  , \u0_R14_reg[6]/NET0131  , \u0_R14_reg[7]/NET0131  , \u0_R14_reg[8]/NET0131  , \u0_R14_reg[9]/NET0131  , \u0_R1_reg[10]/NET0131  , \u0_R1_reg[11]/NET0131  , \u0_R1_reg[12]/NET0131  , \u0_R1_reg[13]/NET0131  , \u0_R1_reg[14]/NET0131  , \u0_R1_reg[15]/NET0131  , \u0_R1_reg[16]/NET0131  , \u0_R1_reg[17]/NET0131  , \u0_R1_reg[18]/NET0131  , \u0_R1_reg[19]/NET0131  , \u0_R1_reg[1]/NET0131  , \u0_R1_reg[20]/NET0131  , \u0_R1_reg[21]/NET0131  , \u0_R1_reg[22]/NET0131  , \u0_R1_reg[23]/NET0131  , \u0_R1_reg[24]/NET0131  , \u0_R1_reg[25]/NET0131  , \u0_R1_reg[26]/NET0131  , \u0_R1_reg[27]/NET0131  , \u0_R1_reg[28]/NET0131  , \u0_R1_reg[29]/NET0131  , \u0_R1_reg[2]/NET0131  , \u0_R1_reg[30]/NET0131  , \u0_R1_reg[31]/NET0131  , \u0_R1_reg[32]/NET0131  , \u0_R1_reg[3]/NET0131  , \u0_R1_reg[4]/NET0131  , \u0_R1_reg[5]/NET0131  , \u0_R1_reg[6]/NET0131  , \u0_R1_reg[7]/NET0131  , \u0_R1_reg[8]/NET0131  , \u0_R1_reg[9]/NET0131  , \u0_R2_reg[10]/NET0131  , \u0_R2_reg[11]/NET0131  , \u0_R2_reg[12]/NET0131  , \u0_R2_reg[13]/NET0131  , \u0_R2_reg[14]/NET0131  , \u0_R2_reg[15]/NET0131  , \u0_R2_reg[16]/NET0131  , \u0_R2_reg[17]/NET0131  , \u0_R2_reg[18]/NET0131  , \u0_R2_reg[19]/NET0131  , \u0_R2_reg[1]/NET0131  , \u0_R2_reg[20]/NET0131  , \u0_R2_reg[21]/NET0131  , \u0_R2_reg[22]/NET0131  , \u0_R2_reg[23]/NET0131  , \u0_R2_reg[24]/NET0131  , \u0_R2_reg[25]/NET0131  , \u0_R2_reg[26]/NET0131  , \u0_R2_reg[27]/NET0131  , \u0_R2_reg[28]/NET0131  , \u0_R2_reg[29]/NET0131  , \u0_R2_reg[2]/NET0131  , \u0_R2_reg[30]/NET0131  , \u0_R2_reg[31]/NET0131  , \u0_R2_reg[32]/NET0131  , \u0_R2_reg[3]/NET0131  , \u0_R2_reg[4]/NET0131  , \u0_R2_reg[5]/NET0131  , \u0_R2_reg[6]/NET0131  , \u0_R2_reg[7]/NET0131  , \u0_R2_reg[8]/NET0131  , \u0_R2_reg[9]/NET0131  , \u0_R3_reg[10]/NET0131  , \u0_R3_reg[11]/NET0131  , \u0_R3_reg[12]/NET0131  , \u0_R3_reg[13]/NET0131  , \u0_R3_reg[14]/NET0131  , \u0_R3_reg[15]/NET0131  , \u0_R3_reg[16]/NET0131  , \u0_R3_reg[17]/NET0131  , \u0_R3_reg[18]/NET0131  , \u0_R3_reg[19]/NET0131  , \u0_R3_reg[1]/NET0131  , \u0_R3_reg[20]/NET0131  , \u0_R3_reg[21]/NET0131  , \u0_R3_reg[22]/NET0131  , \u0_R3_reg[23]/NET0131  , \u0_R3_reg[24]/NET0131  , \u0_R3_reg[25]/NET0131  , \u0_R3_reg[26]/NET0131  , \u0_R3_reg[27]/NET0131  , \u0_R3_reg[28]/NET0131  , \u0_R3_reg[29]/NET0131  , \u0_R3_reg[2]/NET0131  , \u0_R3_reg[30]/NET0131  , \u0_R3_reg[31]/P0001  , \u0_R3_reg[32]/NET0131  , \u0_R3_reg[3]/NET0131  , \u0_R3_reg[4]/NET0131  , \u0_R3_reg[5]/NET0131  , \u0_R3_reg[6]/NET0131  , \u0_R3_reg[7]/NET0131  , \u0_R3_reg[8]/NET0131  , \u0_R3_reg[9]/NET0131  , \u0_R4_reg[10]/NET0131  , \u0_R4_reg[11]/NET0131  , \u0_R4_reg[12]/NET0131  , \u0_R4_reg[13]/NET0131  , \u0_R4_reg[14]/NET0131  , \u0_R4_reg[15]/NET0131  , \u0_R4_reg[16]/NET0131  , \u0_R4_reg[17]/NET0131  , \u0_R4_reg[18]/NET0131  , \u0_R4_reg[19]/NET0131  , \u0_R4_reg[1]/NET0131  , \u0_R4_reg[20]/NET0131  , \u0_R4_reg[21]/NET0131  , \u0_R4_reg[22]/NET0131  , \u0_R4_reg[23]/NET0131  , \u0_R4_reg[24]/NET0131  , \u0_R4_reg[25]/NET0131  , \u0_R4_reg[26]/NET0131  , \u0_R4_reg[27]/NET0131  , \u0_R4_reg[28]/NET0131  , \u0_R4_reg[29]/NET0131  , \u0_R4_reg[2]/NET0131  , \u0_R4_reg[30]/NET0131  , \u0_R4_reg[31]/P0001  , \u0_R4_reg[32]/NET0131  , \u0_R4_reg[3]/NET0131  , \u0_R4_reg[4]/NET0131  , \u0_R4_reg[5]/NET0131  , \u0_R4_reg[6]/NET0131  , \u0_R4_reg[7]/NET0131  , \u0_R4_reg[8]/NET0131  , \u0_R4_reg[9]/NET0131  , \u0_R5_reg[10]/NET0131  , \u0_R5_reg[11]/P0001  , \u0_R5_reg[12]/NET0131  , \u0_R5_reg[13]/NET0131  , \u0_R5_reg[14]/NET0131  , \u0_R5_reg[15]/NET0131  , \u0_R5_reg[16]/NET0131  , \u0_R5_reg[17]/NET0131  , \u0_R5_reg[18]/NET0131  , \u0_R5_reg[19]/NET0131  , \u0_R5_reg[1]/NET0131  , \u0_R5_reg[20]/NET0131  , \u0_R5_reg[21]/NET0131  , \u0_R5_reg[22]/NET0131  , \u0_R5_reg[23]/NET0131  , \u0_R5_reg[24]/NET0131  , \u0_R5_reg[25]/NET0131  , \u0_R5_reg[26]/NET0131  , \u0_R5_reg[27]/NET0131  , \u0_R5_reg[28]/NET0131  , \u0_R5_reg[29]/NET0131  , \u0_R5_reg[2]/NET0131  , \u0_R5_reg[30]/NET0131  , \u0_R5_reg[31]/P0001  , \u0_R5_reg[32]/NET0131  , \u0_R5_reg[3]/NET0131  , \u0_R5_reg[4]/NET0131  , \u0_R5_reg[5]/NET0131  , \u0_R5_reg[6]/NET0131  , \u0_R5_reg[7]/NET0131  , \u0_R5_reg[8]/NET0131  , \u0_R5_reg[9]/NET0131  , \u0_R6_reg[10]/NET0131  , \u0_R6_reg[11]/NET0131  , \u0_R6_reg[12]/NET0131  , \u0_R6_reg[13]/NET0131  , \u0_R6_reg[14]/NET0131  , \u0_R6_reg[15]/NET0131  , \u0_R6_reg[16]/NET0131  , \u0_R6_reg[17]/NET0131  , \u0_R6_reg[18]/NET0131  , \u0_R6_reg[19]/NET0131  , \u0_R6_reg[1]/NET0131  , \u0_R6_reg[20]/NET0131  , \u0_R6_reg[21]/NET0131  , \u0_R6_reg[22]/NET0131  , \u0_R6_reg[23]/NET0131  , \u0_R6_reg[24]/NET0131  , \u0_R6_reg[25]/NET0131  , \u0_R6_reg[26]/NET0131  , \u0_R6_reg[27]/NET0131  , \u0_R6_reg[28]/NET0131  , \u0_R6_reg[29]/NET0131  , \u0_R6_reg[2]/NET0131  , \u0_R6_reg[30]/NET0131  , \u0_R6_reg[31]/P0001  , \u0_R6_reg[32]/NET0131  , \u0_R6_reg[3]/NET0131  , \u0_R6_reg[4]/NET0131  , \u0_R6_reg[5]/NET0131  , \u0_R6_reg[6]/NET0131  , \u0_R6_reg[7]/NET0131  , \u0_R6_reg[8]/NET0131  , \u0_R6_reg[9]/NET0131  , \u0_R7_reg[10]/NET0131  , \u0_R7_reg[11]/P0001  , \u0_R7_reg[12]/NET0131  , \u0_R7_reg[13]/NET0131  , \u0_R7_reg[14]/NET0131  , \u0_R7_reg[15]/NET0131  , \u0_R7_reg[16]/NET0131  , \u0_R7_reg[17]/NET0131  , \u0_R7_reg[18]/NET0131  , \u0_R7_reg[19]/NET0131  , \u0_R7_reg[1]/NET0131  , \u0_R7_reg[20]/NET0131  , \u0_R7_reg[21]/NET0131  , \u0_R7_reg[22]/NET0131  , \u0_R7_reg[23]/NET0131  , \u0_R7_reg[24]/NET0131  , \u0_R7_reg[25]/NET0131  , \u0_R7_reg[26]/NET0131  , \u0_R7_reg[27]/NET0131  , \u0_R7_reg[28]/NET0131  , \u0_R7_reg[29]/NET0131  , \u0_R7_reg[2]/NET0131  , \u0_R7_reg[30]/NET0131  , \u0_R7_reg[31]/P0001  , \u0_R7_reg[32]/NET0131  , \u0_R7_reg[3]/NET0131  , \u0_R7_reg[4]/NET0131  , \u0_R7_reg[5]/NET0131  , \u0_R7_reg[6]/NET0131  , \u0_R7_reg[7]/NET0131  , \u0_R7_reg[8]/NET0131  , \u0_R7_reg[9]/NET0131  , \u0_R8_reg[10]/NET0131  , \u0_R8_reg[11]/NET0131  , \u0_R8_reg[12]/NET0131  , \u0_R8_reg[13]/NET0131  , \u0_R8_reg[14]/NET0131  , \u0_R8_reg[15]/NET0131  , \u0_R8_reg[16]/NET0131  , \u0_R8_reg[17]/NET0131  , \u0_R8_reg[18]/NET0131  , \u0_R8_reg[19]/NET0131  , \u0_R8_reg[1]/NET0131  , \u0_R8_reg[20]/NET0131  , \u0_R8_reg[21]/NET0131  , \u0_R8_reg[22]/NET0131  , \u0_R8_reg[23]/NET0131  , \u0_R8_reg[24]/NET0131  , \u0_R8_reg[25]/NET0131  , \u0_R8_reg[26]/NET0131  , \u0_R8_reg[27]/NET0131  , \u0_R8_reg[28]/NET0131  , \u0_R8_reg[29]/NET0131  , \u0_R8_reg[2]/NET0131  , \u0_R8_reg[30]/NET0131  , \u0_R8_reg[31]/P0001  , \u0_R8_reg[32]/NET0131  , \u0_R8_reg[3]/NET0131  , \u0_R8_reg[4]/NET0131  , \u0_R8_reg[5]/NET0131  , \u0_R8_reg[6]/NET0131  , \u0_R8_reg[7]/NET0131  , \u0_R8_reg[8]/NET0131  , \u0_R8_reg[9]/NET0131  , \u0_R9_reg[10]/NET0131  , \u0_R9_reg[11]/P0001  , \u0_R9_reg[12]/NET0131  , \u0_R9_reg[13]/NET0131  , \u0_R9_reg[14]/NET0131  , \u0_R9_reg[15]/NET0131  , \u0_R9_reg[16]/NET0131  , \u0_R9_reg[17]/NET0131  , \u0_R9_reg[18]/NET0131  , \u0_R9_reg[19]/NET0131  , \u0_R9_reg[1]/NET0131  , \u0_R9_reg[20]/NET0131  , \u0_R9_reg[21]/NET0131  , \u0_R9_reg[22]/NET0131  , \u0_R9_reg[23]/NET0131  , \u0_R9_reg[24]/NET0131  , \u0_R9_reg[25]/NET0131  , \u0_R9_reg[26]/NET0131  , \u0_R9_reg[27]/NET0131  , \u0_R9_reg[28]/NET0131  , \u0_R9_reg[29]/NET0131  , \u0_R9_reg[2]/NET0131  , \u0_R9_reg[30]/NET0131  , \u0_R9_reg[31]/P0001  , \u0_R9_reg[32]/NET0131  , \u0_R9_reg[3]/NET0131  , \u0_R9_reg[4]/NET0131  , \u0_R9_reg[5]/NET0131  , \u0_R9_reg[6]/NET0131  , \u0_R9_reg[7]/NET0131  , \u0_R9_reg[8]/NET0131  , \u0_R9_reg[9]/NET0131  , \u0_desIn_r_reg[0]/NET0131  , \u0_desIn_r_reg[10]/NET0131  , \u0_desIn_r_reg[11]/NET0131  , \u0_desIn_r_reg[12]/NET0131  , \u0_desIn_r_reg[13]/NET0131  , \u0_desIn_r_reg[14]/NET0131  , \u0_desIn_r_reg[15]/NET0131  , \u0_desIn_r_reg[16]/NET0131  , \u0_desIn_r_reg[17]/NET0131  , \u0_desIn_r_reg[18]/NET0131  , \u0_desIn_r_reg[19]/NET0131  , \u0_desIn_r_reg[1]/NET0131  , \u0_desIn_r_reg[20]/NET0131  , \u0_desIn_r_reg[21]/NET0131  , \u0_desIn_r_reg[22]/NET0131  , \u0_desIn_r_reg[23]/NET0131  , \u0_desIn_r_reg[24]/NET0131  , \u0_desIn_r_reg[25]/NET0131  , \u0_desIn_r_reg[26]/NET0131  , \u0_desIn_r_reg[27]/NET0131  , \u0_desIn_r_reg[28]/NET0131  , \u0_desIn_r_reg[29]/NET0131  , \u0_desIn_r_reg[2]/NET0131  , \u0_desIn_r_reg[30]/NET0131  , \u0_desIn_r_reg[31]/NET0131  , \u0_desIn_r_reg[32]/NET0131  , \u0_desIn_r_reg[33]/NET0131  , \u0_desIn_r_reg[34]/NET0131  , \u0_desIn_r_reg[35]/NET0131  , \u0_desIn_r_reg[36]/NET0131  , \u0_desIn_r_reg[37]/NET0131  , \u0_desIn_r_reg[38]/NET0131  , \u0_desIn_r_reg[39]/NET0131  , \u0_desIn_r_reg[3]/NET0131  , \u0_desIn_r_reg[40]/NET0131  , \u0_desIn_r_reg[41]/NET0131  , \u0_desIn_r_reg[42]/NET0131  , \u0_desIn_r_reg[43]/NET0131  , \u0_desIn_r_reg[44]/NET0131  , \u0_desIn_r_reg[45]/NET0131  , \u0_desIn_r_reg[46]/NET0131  , \u0_desIn_r_reg[47]/NET0131  , \u0_desIn_r_reg[48]/NET0131  , \u0_desIn_r_reg[49]/NET0131  , \u0_desIn_r_reg[4]/NET0131  , \u0_desIn_r_reg[50]/NET0131  , \u0_desIn_r_reg[51]/NET0131  , \u0_desIn_r_reg[52]/NET0131  , \u0_desIn_r_reg[53]/NET0131  , \u0_desIn_r_reg[54]/NET0131  , \u0_desIn_r_reg[55]/NET0131  , \u0_desIn_r_reg[56]/NET0131  , \u0_desIn_r_reg[57]/NET0131  , \u0_desIn_r_reg[58]/NET0131  , \u0_desIn_r_reg[59]/NET0131  , \u0_desIn_r_reg[5]/NET0131  , \u0_desIn_r_reg[60]/NET0131  , \u0_desIn_r_reg[61]/NET0131  , \u0_desIn_r_reg[62]/NET0131  , \u0_desIn_r_reg[63]/NET0131  , \u0_desIn_r_reg[6]/NET0131  , \u0_desIn_r_reg[7]/NET0131  , \u0_desIn_r_reg[8]/NET0131  , \u0_desIn_r_reg[9]/NET0131  , \u0_key_r_reg[0]/NET0131  , \u0_key_r_reg[10]/P0001  , \u0_key_r_reg[11]/NET0131  , \u0_key_r_reg[12]/NET0131  , \u0_key_r_reg[13]/NET0131  , \u0_key_r_reg[14]/NET0131  , \u0_key_r_reg[15]/NET0131  , \u0_key_r_reg[16]/NET0131  , \u0_key_r_reg[17]/NET0131  , \u0_key_r_reg[18]/NET0131  , \u0_key_r_reg[19]/NET0131  , \u0_key_r_reg[1]/NET0131  , \u0_key_r_reg[20]/NET0131  , \u0_key_r_reg[21]/NET0131  , \u0_key_r_reg[22]/NET0131  , \u0_key_r_reg[23]/NET0131  , \u0_key_r_reg[24]/NET0131  , \u0_key_r_reg[25]/NET0131  , \u0_key_r_reg[26]/NET0131  , \u0_key_r_reg[27]/NET0131  , \u0_key_r_reg[28]/NET0131  , \u0_key_r_reg[29]/NET0131  , \u0_key_r_reg[2]/NET0131  , \u0_key_r_reg[30]/NET0131  , \u0_key_r_reg[31]/NET0131  , \u0_key_r_reg[32]/NET0131  , \u0_key_r_reg[33]/NET0131  , \u0_key_r_reg[34]/NET0131  , \u0_key_r_reg[35]/P0001  , \u0_key_r_reg[36]/NET0131  , \u0_key_r_reg[37]/NET0131  , \u0_key_r_reg[38]/NET0131  , \u0_key_r_reg[39]/P0001  , \u0_key_r_reg[3]/NET0131  , \u0_key_r_reg[40]/NET0131  , \u0_key_r_reg[41]/NET0131  , \u0_key_r_reg[42]/P0001  , \u0_key_r_reg[43]/NET0131  , \u0_key_r_reg[44]/NET0131  , \u0_key_r_reg[45]/NET0131  , \u0_key_r_reg[46]/NET0131  , \u0_key_r_reg[47]/NET0131  , \u0_key_r_reg[48]/NET0131  , \u0_key_r_reg[49]/NET0131  , \u0_key_r_reg[4]/NET0131  , \u0_key_r_reg[50]/NET0131  , \u0_key_r_reg[51]/NET0131  , \u0_key_r_reg[52]/NET0131  , \u0_key_r_reg[53]/NET0131  , \u0_key_r_reg[54]/NET0131  , \u0_key_r_reg[55]/NET0131  , \u0_key_r_reg[5]/NET0131  , \u0_key_r_reg[6]/NET0131  , \u0_key_r_reg[7]/NET0131  , \u0_key_r_reg[8]/NET0131  , \u0_key_r_reg[9]/NET0131  , \u0_uk_K_r0_reg[0]/NET0131  , \u0_uk_K_r0_reg[10]/NET0131  , \u0_uk_K_r0_reg[11]/NET0131  , \u0_uk_K_r0_reg[12]/NET0131  , \u0_uk_K_r0_reg[13]/NET0131  , \u0_uk_K_r0_reg[14]/NET0131  , \u0_uk_K_r0_reg[15]/NET0131  , \u0_uk_K_r0_reg[16]/NET0131  , \u0_uk_K_r0_reg[17]/NET0131  , \u0_uk_K_r0_reg[18]/NET0131  , \u0_uk_K_r0_reg[19]/NET0131  , \u0_uk_K_r0_reg[20]/NET0131  , \u0_uk_K_r0_reg[21]/NET0131  , \u0_uk_K_r0_reg[22]/NET0131  , \u0_uk_K_r0_reg[23]/NET0131  , \u0_uk_K_r0_reg[24]/P0001  , \u0_uk_K_r0_reg[25]/P0001  , \u0_uk_K_r0_reg[26]/NET0131  , \u0_uk_K_r0_reg[27]/NET0131  , \u0_uk_K_r0_reg[28]/NET0131  , \u0_uk_K_r0_reg[29]/NET0131  , \u0_uk_K_r0_reg[2]/NET0131  , \u0_uk_K_r0_reg[30]/NET0131  , \u0_uk_K_r0_reg[31]/NET0131  , \u0_uk_K_r0_reg[32]/NET0131  , \u0_uk_K_r0_reg[33]/NET0131  , \u0_uk_K_r0_reg[34]/NET0131  , \u0_uk_K_r0_reg[35]/NET0131  , \u0_uk_K_r0_reg[36]/NET0131  , \u0_uk_K_r0_reg[37]/NET0131  , \u0_uk_K_r0_reg[38]/NET0131  , \u0_uk_K_r0_reg[39]/NET0131  , \u0_uk_K_r0_reg[3]/NET0131  , \u0_uk_K_r0_reg[40]/NET0131  , \u0_uk_K_r0_reg[41]/NET0131  , \u0_uk_K_r0_reg[42]/NET0131  , \u0_uk_K_r0_reg[43]/NET0131  , \u0_uk_K_r0_reg[44]/NET0131  , \u0_uk_K_r0_reg[45]/NET0131  , \u0_uk_K_r0_reg[46]/NET0131  , \u0_uk_K_r0_reg[47]/NET0131  , \u0_uk_K_r0_reg[48]/NET0131  , \u0_uk_K_r0_reg[49]/NET0131  , \u0_uk_K_r0_reg[4]/NET0131  , \u0_uk_K_r0_reg[50]/NET0131  , \u0_uk_K_r0_reg[51]/NET0131  , \u0_uk_K_r0_reg[52]/NET0131  , \u0_uk_K_r0_reg[54]/NET0131  , \u0_uk_K_r0_reg[55]/NET0131  , \u0_uk_K_r0_reg[5]/NET0131  , \u0_uk_K_r0_reg[6]/NET0131  , \u0_uk_K_r0_reg[7]/NET0131  , \u0_uk_K_r0_reg[8]/NET0131  , \u0_uk_K_r0_reg[9]/NET0131  , \u0_uk_K_r10_reg[0]/NET0131  , \u0_uk_K_r10_reg[10]/NET0131  , \u0_uk_K_r10_reg[11]/NET0131  , \u0_uk_K_r10_reg[12]/NET0131  , \u0_uk_K_r10_reg[14]/NET0131  , \u0_uk_K_r10_reg[15]/NET0131  , \u0_uk_K_r10_reg[16]/NET0131  , \u0_uk_K_r10_reg[17]/NET0131  , \u0_uk_K_r10_reg[18]/NET0131  , \u0_uk_K_r10_reg[19]/NET0131  , \u0_uk_K_r10_reg[1]/NET0131  , \u0_uk_K_r10_reg[20]/NET0131  , \u0_uk_K_r10_reg[21]/NET0131  , \u0_uk_K_r10_reg[22]/NET0131  , \u0_uk_K_r10_reg[23]/NET0131  , \u0_uk_K_r10_reg[24]/NET0131  , \u0_uk_K_r10_reg[25]/NET0131  , \u0_uk_K_r10_reg[26]/NET0131  , \u0_uk_K_r10_reg[27]/NET0131  , \u0_uk_K_r10_reg[28]/NET0131  , \u0_uk_K_r10_reg[29]/NET0131  , \u0_uk_K_r10_reg[2]/NET0131  , \u0_uk_K_r10_reg[30]/NET0131  , \u0_uk_K_r10_reg[31]/NET0131  , \u0_uk_K_r10_reg[32]/NET0131  , \u0_uk_K_r10_reg[33]/NET0131  , \u0_uk_K_r10_reg[34]/NET0131  , \u0_uk_K_r10_reg[35]/NET0131  , \u0_uk_K_r10_reg[36]/NET0131  , \u0_uk_K_r10_reg[37]/NET0131  , \u0_uk_K_r10_reg[38]/NET0131  , \u0_uk_K_r10_reg[39]/NET0131  , \u0_uk_K_r10_reg[3]/NET0131  , \u0_uk_K_r10_reg[40]/NET0131  , \u0_uk_K_r10_reg[41]/P0001  , \u0_uk_K_r10_reg[42]/NET0131  , \u0_uk_K_r10_reg[43]/NET0131  , \u0_uk_K_r10_reg[44]/NET0131  , \u0_uk_K_r10_reg[45]/P0001  , \u0_uk_K_r10_reg[46]/NET0131  , \u0_uk_K_r10_reg[47]/NET0131  , \u0_uk_K_r10_reg[48]/NET0131  , \u0_uk_K_r10_reg[49]/NET0131  , \u0_uk_K_r10_reg[4]/NET0131  , \u0_uk_K_r10_reg[50]/NET0131  , \u0_uk_K_r10_reg[51]/NET0131  , \u0_uk_K_r10_reg[52]/NET0131  , \u0_uk_K_r10_reg[53]/NET0131  , \u0_uk_K_r10_reg[54]/NET0131  , \u0_uk_K_r10_reg[55]/NET0131  , \u0_uk_K_r10_reg[5]/NET0131  , \u0_uk_K_r10_reg[6]/NET0131  , \u0_uk_K_r10_reg[7]/NET0131  , \u0_uk_K_r10_reg[8]/NET0131  , \u0_uk_K_r10_reg[9]/NET0131  , \u0_uk_K_r11_reg[0]/NET0131  , \u0_uk_K_r11_reg[10]/NET0131  , \u0_uk_K_r11_reg[11]/NET0131  , \u0_uk_K_r11_reg[12]/NET0131  , \u0_uk_K_r11_reg[13]/NET0131  , \u0_uk_K_r11_reg[14]/NET0131  , \u0_uk_K_r11_reg[15]/NET0131  , \u0_uk_K_r11_reg[16]/NET0131  , \u0_uk_K_r11_reg[17]/NET0131  , \u0_uk_K_r11_reg[18]/NET0131  , \u0_uk_K_r11_reg[19]/NET0131  , \u0_uk_K_r11_reg[1]/NET0131  , \u0_uk_K_r11_reg[20]/NET0131  , \u0_uk_K_r11_reg[21]/NET0131  , \u0_uk_K_r11_reg[22]/NET0131  , \u0_uk_K_r11_reg[23]/NET0131  , \u0_uk_K_r11_reg[24]/NET0131  , \u0_uk_K_r11_reg[25]/NET0131  , \u0_uk_K_r11_reg[26]/NET0131  , \u0_uk_K_r11_reg[27]/P0001  , \u0_uk_K_r11_reg[28]/NET0131  , \u0_uk_K_r11_reg[29]/NET0131  , \u0_uk_K_r11_reg[2]/NET0131  , \u0_uk_K_r11_reg[31]/NET0131  , \u0_uk_K_r11_reg[32]/NET0131  , \u0_uk_K_r11_reg[33]/NET0131  , \u0_uk_K_r11_reg[34]/NET0131  , \u0_uk_K_r11_reg[35]/NET0131  , \u0_uk_K_r11_reg[36]/NET0131  , \u0_uk_K_r11_reg[37]/NET0131  , \u0_uk_K_r11_reg[38]/NET0131  , \u0_uk_K_r11_reg[39]/NET0131  , \u0_uk_K_r11_reg[3]/NET0131  , \u0_uk_K_r11_reg[40]/NET0131  , \u0_uk_K_r11_reg[41]/NET0131  , \u0_uk_K_r11_reg[42]/NET0131  , \u0_uk_K_r11_reg[43]/NET0131  , \u0_uk_K_r11_reg[44]/NET0131  , \u0_uk_K_r11_reg[45]/NET0131  , \u0_uk_K_r11_reg[46]/NET0131  , \u0_uk_K_r11_reg[47]/NET0131  , \u0_uk_K_r11_reg[48]/NET0131  , \u0_uk_K_r11_reg[49]/NET0131  , \u0_uk_K_r11_reg[4]/NET0131  , \u0_uk_K_r11_reg[50]/NET0131  , \u0_uk_K_r11_reg[51]/NET0131  , \u0_uk_K_r11_reg[52]/NET0131  , \u0_uk_K_r11_reg[53]/P0001  , \u0_uk_K_r11_reg[54]/NET0131  , \u0_uk_K_r11_reg[55]/NET0131  , \u0_uk_K_r11_reg[5]/NET0131  , \u0_uk_K_r11_reg[6]/NET0131  , \u0_uk_K_r11_reg[7]/NET0131  , \u0_uk_K_r11_reg[8]/NET0131  , \u0_uk_K_r11_reg[9]/NET0131  , \u0_uk_K_r12_reg[0]/NET0131  , \u0_uk_K_r12_reg[10]/P0001  , \u0_uk_K_r12_reg[11]/NET0131  , \u0_uk_K_r12_reg[12]/NET0131  , \u0_uk_K_r12_reg[13]/NET0131  , \u0_uk_K_r12_reg[14]/NET0131  , \u0_uk_K_r12_reg[15]/NET0131  , \u0_uk_K_r12_reg[16]/NET0131  , \u0_uk_K_r12_reg[17]/NET0131  , \u0_uk_K_r12_reg[18]/NET0131  , \u0_uk_K_r12_reg[19]/NET0131  , \u0_uk_K_r12_reg[1]/NET0131  , \u0_uk_K_r12_reg[20]/NET0131  , \u0_uk_K_r12_reg[21]/NET0131  , \u0_uk_K_r12_reg[22]/NET0131  , \u0_uk_K_r12_reg[23]/NET0131  , \u0_uk_K_r12_reg[24]/NET0131  , \u0_uk_K_r12_reg[25]/NET0131  , \u0_uk_K_r12_reg[26]/NET0131  , \u0_uk_K_r12_reg[27]/NET0131  , \u0_uk_K_r12_reg[28]/NET0131  , \u0_uk_K_r12_reg[29]/NET0131  , \u0_uk_K_r12_reg[2]/NET0131  , \u0_uk_K_r12_reg[30]/NET0131  , \u0_uk_K_r12_reg[31]/NET0131  , \u0_uk_K_r12_reg[32]/NET0131  , \u0_uk_K_r12_reg[33]/NET0131  , \u0_uk_K_r12_reg[34]/NET0131  , \u0_uk_K_r12_reg[35]/NET0131  , \u0_uk_K_r12_reg[36]/NET0131  , \u0_uk_K_r12_reg[37]/NET0131  , \u0_uk_K_r12_reg[38]/NET0131  , \u0_uk_K_r12_reg[3]/NET0131  , \u0_uk_K_r12_reg[40]/NET0131  , \u0_uk_K_r12_reg[41]/NET0131  , \u0_uk_K_r12_reg[42]/NET0131  , \u0_uk_K_r12_reg[43]/NET0131  , \u0_uk_K_r12_reg[44]/P0001  , \u0_uk_K_r12_reg[45]/NET0131  , \u0_uk_K_r12_reg[46]/NET0131  , \u0_uk_K_r12_reg[47]/NET0131  , \u0_uk_K_r12_reg[48]/NET0131  , \u0_uk_K_r12_reg[49]/NET0131  , \u0_uk_K_r12_reg[4]/NET0131  , \u0_uk_K_r12_reg[50]/NET0131  , \u0_uk_K_r12_reg[51]/NET0131  , \u0_uk_K_r12_reg[52]/NET0131  , \u0_uk_K_r12_reg[53]/NET0131  , \u0_uk_K_r12_reg[54]/NET0131  , \u0_uk_K_r12_reg[55]/NET0131  , \u0_uk_K_r12_reg[5]/NET0131  , \u0_uk_K_r12_reg[6]/NET0131  , \u0_uk_K_r12_reg[7]/P0001  , \u0_uk_K_r12_reg[8]/NET0131  , \u0_uk_K_r12_reg[9]/NET0131  , \u0_uk_K_r13_reg[0]/NET0131  , \u0_uk_K_r13_reg[10]/NET0131  , \u0_uk_K_r13_reg[11]/NET0131  , \u0_uk_K_r13_reg[12]/NET0131  , \u0_uk_K_r13_reg[13]/NET0131  , \u0_uk_K_r13_reg[14]/NET0131  , \u0_uk_K_r13_reg[15]/NET0131  , \u0_uk_K_r13_reg[16]/NET0131  , \u0_uk_K_r13_reg[17]/NET0131  , \u0_uk_K_r13_reg[18]/NET0131  , \u0_uk_K_r13_reg[19]/NET0131  , \u0_uk_K_r13_reg[20]/NET0131  , \u0_uk_K_r13_reg[21]/NET0131  , \u0_uk_K_r13_reg[22]/NET0131  , \u0_uk_K_r13_reg[23]/NET0131  , \u0_uk_K_r13_reg[24]/NET0131  , \u0_uk_K_r13_reg[25]/P0001  , \u0_uk_K_r13_reg[26]/NET0131  , \u0_uk_K_r13_reg[27]/NET0131  , \u0_uk_K_r13_reg[28]/NET0131  , \u0_uk_K_r13_reg[29]/NET0131  , \u0_uk_K_r13_reg[2]/NET0131  , \u0_uk_K_r13_reg[30]/NET0131  , \u0_uk_K_r13_reg[31]/NET0131  , \u0_uk_K_r13_reg[32]/NET0131  , \u0_uk_K_r13_reg[33]/NET0131  , \u0_uk_K_r13_reg[34]/NET0131  , \u0_uk_K_r13_reg[35]/NET0131  , \u0_uk_K_r13_reg[36]/NET0131  , \u0_uk_K_r13_reg[37]/NET0131  , \u0_uk_K_r13_reg[38]/NET0131  , \u0_uk_K_r13_reg[39]/NET0131  , \u0_uk_K_r13_reg[3]/NET0131  , \u0_uk_K_r13_reg[40]/NET0131  , \u0_uk_K_r13_reg[41]/NET0131  , \u0_uk_K_r13_reg[42]/NET0131  , \u0_uk_K_r13_reg[43]/NET0131  , \u0_uk_K_r13_reg[44]/NET0131  , \u0_uk_K_r13_reg[45]/NET0131  , \u0_uk_K_r13_reg[46]/NET0131  , \u0_uk_K_r13_reg[47]/NET0131  , \u0_uk_K_r13_reg[48]/NET0131  , \u0_uk_K_r13_reg[49]/NET0131  , \u0_uk_K_r13_reg[4]/NET0131  , \u0_uk_K_r13_reg[50]/NET0131  , \u0_uk_K_r13_reg[51]/NET0131  , \u0_uk_K_r13_reg[52]/P0001  , \u0_uk_K_r13_reg[54]/NET0131  , \u0_uk_K_r13_reg[55]/NET0131  , \u0_uk_K_r13_reg[5]/NET0131  , \u0_uk_K_r13_reg[6]/NET0131  , \u0_uk_K_r13_reg[7]/NET0131  , \u0_uk_K_r13_reg[8]/NET0131  , \u0_uk_K_r13_reg[9]/NET0131  , \u0_uk_K_r14_reg[0]/NET0131  , \u0_uk_K_r14_reg[10]/P0001  , \u0_uk_K_r14_reg[11]/NET0131  , \u0_uk_K_r14_reg[12]/NET0131  , \u0_uk_K_r14_reg[13]/NET0131  , \u0_uk_K_r14_reg[14]/NET0131  , \u0_uk_K_r14_reg[15]/NET0131  , \u0_uk_K_r14_reg[16]/NET0131  , \u0_uk_K_r14_reg[17]/NET0131  , \u0_uk_K_r14_reg[18]/NET0131  , \u0_uk_K_r14_reg[19]/NET0131  , \u0_uk_K_r14_reg[1]/NET0131  , \u0_uk_K_r14_reg[20]/NET0131  , \u0_uk_K_r14_reg[21]/NET0131  , \u0_uk_K_r14_reg[22]/NET0131  , \u0_uk_K_r14_reg[23]/NET0131  , \u0_uk_K_r14_reg[24]/NET0131  , \u0_uk_K_r14_reg[25]/NET0131  , \u0_uk_K_r14_reg[26]/NET0131  , \u0_uk_K_r14_reg[27]/NET0131  , \u0_uk_K_r14_reg[28]/NET0131  , \u0_uk_K_r14_reg[29]/NET0131  , \u0_uk_K_r14_reg[2]/NET0131  , \u0_uk_K_r14_reg[30]/NET0131  , \u0_uk_K_r14_reg[31]/NET0131  , \u0_uk_K_r14_reg[32]/NET0131  , \u0_uk_K_r14_reg[33]/NET0131  , \u0_uk_K_r14_reg[34]/NET0131  , \u0_uk_K_r14_reg[35]/P0001  , \u0_uk_K_r14_reg[36]/NET0131  , \u0_uk_K_r14_reg[37]/NET0131  , \u0_uk_K_r14_reg[38]/NET0131  , \u0_uk_K_r14_reg[39]/P0001  , \u0_uk_K_r14_reg[3]/NET0131  , \u0_uk_K_r14_reg[40]/NET0131  , \u0_uk_K_r14_reg[41]/NET0131  , \u0_uk_K_r14_reg[42]/P0001  , \u0_uk_K_r14_reg[43]/NET0131  , \u0_uk_K_r14_reg[44]/NET0131  , \u0_uk_K_r14_reg[45]/NET0131  , \u0_uk_K_r14_reg[46]/NET0131  , \u0_uk_K_r14_reg[47]/NET0131  , \u0_uk_K_r14_reg[48]/NET0131  , \u0_uk_K_r14_reg[49]/NET0131  , \u0_uk_K_r14_reg[4]/NET0131  , \u0_uk_K_r14_reg[50]/NET0131  , \u0_uk_K_r14_reg[51]/NET0131  , \u0_uk_K_r14_reg[52]/NET0131  , \u0_uk_K_r14_reg[53]/NET0131  , \u0_uk_K_r14_reg[54]/NET0131  , \u0_uk_K_r14_reg[55]/NET0131  , \u0_uk_K_r14_reg[5]/NET0131  , \u0_uk_K_r14_reg[6]/NET0131  , \u0_uk_K_r14_reg[7]/NET0131  , \u0_uk_K_r14_reg[8]/NET0131  , \u0_uk_K_r14_reg[9]/NET0131  , \u0_uk_K_r1_reg[0]/NET0131  , \u0_uk_K_r1_reg[10]/P0001  , \u0_uk_K_r1_reg[11]/NET0131  , \u0_uk_K_r1_reg[12]/NET0131  , \u0_uk_K_r1_reg[13]/NET0131  , \u0_uk_K_r1_reg[14]/NET0131  , \u0_uk_K_r1_reg[15]/NET0131  , \u0_uk_K_r1_reg[16]/NET0131  , \u0_uk_K_r1_reg[17]/NET0131  , \u0_uk_K_r1_reg[18]/NET0131  , \u0_uk_K_r1_reg[19]/NET0131  , \u0_uk_K_r1_reg[1]/NET0131  , \u0_uk_K_r1_reg[20]/NET0131  , \u0_uk_K_r1_reg[21]/NET0131  , \u0_uk_K_r1_reg[22]/NET0131  , \u0_uk_K_r1_reg[23]/NET0131  , \u0_uk_K_r1_reg[24]/NET0131  , \u0_uk_K_r1_reg[25]/NET0131  , \u0_uk_K_r1_reg[26]/NET0131  , \u0_uk_K_r1_reg[27]/NET0131  , \u0_uk_K_r1_reg[28]/NET0131  , \u0_uk_K_r1_reg[29]/NET0131  , \u0_uk_K_r1_reg[2]/NET0131  , \u0_uk_K_r1_reg[30]/NET0131  , \u0_uk_K_r1_reg[31]/NET0131  , \u0_uk_K_r1_reg[32]/NET0131  , \u0_uk_K_r1_reg[33]/NET0131  , \u0_uk_K_r1_reg[34]/NET0131  , \u0_uk_K_r1_reg[35]/NET0131  , \u0_uk_K_r1_reg[36]/NET0131  , \u0_uk_K_r1_reg[37]/NET0131  , \u0_uk_K_r1_reg[38]/NET0131  , \u0_uk_K_r1_reg[3]/NET0131  , \u0_uk_K_r1_reg[40]/NET0131  , \u0_uk_K_r1_reg[41]/NET0131  , \u0_uk_K_r1_reg[42]/NET0131  , \u0_uk_K_r1_reg[43]/NET0131  , \u0_uk_K_r1_reg[44]/P0001  , \u0_uk_K_r1_reg[45]/NET0131  , \u0_uk_K_r1_reg[46]/NET0131  , \u0_uk_K_r1_reg[47]/NET0131  , \u0_uk_K_r1_reg[48]/NET0131  , \u0_uk_K_r1_reg[49]/NET0131  , \u0_uk_K_r1_reg[4]/NET0131  , \u0_uk_K_r1_reg[50]/NET0131  , \u0_uk_K_r1_reg[51]/NET0131  , \u0_uk_K_r1_reg[52]/NET0131  , \u0_uk_K_r1_reg[53]/NET0131  , \u0_uk_K_r1_reg[54]/NET0131  , \u0_uk_K_r1_reg[55]/NET0131  , \u0_uk_K_r1_reg[5]/NET0131  , \u0_uk_K_r1_reg[6]/NET0131  , \u0_uk_K_r1_reg[7]/P0001  , \u0_uk_K_r1_reg[8]/NET0131  , \u0_uk_K_r1_reg[9]/NET0131  , \u0_uk_K_r2_reg[0]/NET0131  , \u0_uk_K_r2_reg[10]/NET0131  , \u0_uk_K_r2_reg[11]/NET0131  , \u0_uk_K_r2_reg[12]/NET0131  , \u0_uk_K_r2_reg[13]/NET0131  , \u0_uk_K_r2_reg[14]/NET0131  , \u0_uk_K_r2_reg[15]/NET0131  , \u0_uk_K_r2_reg[16]/NET0131  , \u0_uk_K_r2_reg[17]/NET0131  , \u0_uk_K_r2_reg[18]/NET0131  , \u0_uk_K_r2_reg[19]/NET0131  , \u0_uk_K_r2_reg[1]/NET0131  , \u0_uk_K_r2_reg[20]/NET0131  , \u0_uk_K_r2_reg[21]/NET0131  , \u0_uk_K_r2_reg[22]/NET0131  , \u0_uk_K_r2_reg[23]/NET0131  , \u0_uk_K_r2_reg[24]/NET0131  , \u0_uk_K_r2_reg[25]/NET0131  , \u0_uk_K_r2_reg[26]/NET0131  , \u0_uk_K_r2_reg[27]/P0001  , \u0_uk_K_r2_reg[28]/NET0131  , \u0_uk_K_r2_reg[29]/NET0131  , \u0_uk_K_r2_reg[2]/NET0131  , \u0_uk_K_r2_reg[31]/NET0131  , \u0_uk_K_r2_reg[32]/NET0131  , \u0_uk_K_r2_reg[33]/NET0131  , \u0_uk_K_r2_reg[34]/NET0131  , \u0_uk_K_r2_reg[35]/NET0131  , \u0_uk_K_r2_reg[36]/NET0131  , \u0_uk_K_r2_reg[37]/NET0131  , \u0_uk_K_r2_reg[38]/NET0131  , \u0_uk_K_r2_reg[39]/NET0131  , \u0_uk_K_r2_reg[3]/NET0131  , \u0_uk_K_r2_reg[40]/NET0131  , \u0_uk_K_r2_reg[41]/NET0131  , \u0_uk_K_r2_reg[42]/NET0131  , \u0_uk_K_r2_reg[43]/NET0131  , \u0_uk_K_r2_reg[44]/NET0131  , \u0_uk_K_r2_reg[45]/NET0131  , \u0_uk_K_r2_reg[46]/NET0131  , \u0_uk_K_r2_reg[47]/NET0131  , \u0_uk_K_r2_reg[48]/NET0131  , \u0_uk_K_r2_reg[49]/NET0131  , \u0_uk_K_r2_reg[4]/NET0131  , \u0_uk_K_r2_reg[50]/NET0131  , \u0_uk_K_r2_reg[51]/NET0131  , \u0_uk_K_r2_reg[52]/NET0131  , \u0_uk_K_r2_reg[53]/P0001  , \u0_uk_K_r2_reg[54]/NET0131  , \u0_uk_K_r2_reg[55]/NET0131  , \u0_uk_K_r2_reg[5]/NET0131  , \u0_uk_K_r2_reg[6]/NET0131  , \u0_uk_K_r2_reg[7]/NET0131  , \u0_uk_K_r2_reg[8]/NET0131  , \u0_uk_K_r2_reg[9]/NET0131  , \u0_uk_K_r3_reg[0]/NET0131  , \u0_uk_K_r3_reg[10]/NET0131  , \u0_uk_K_r3_reg[11]/NET0131  , \u0_uk_K_r3_reg[12]/NET0131  , \u0_uk_K_r3_reg[14]/NET0131  , \u0_uk_K_r3_reg[15]/NET0131  , \u0_uk_K_r3_reg[16]/NET0131  , \u0_uk_K_r3_reg[17]/NET0131  , \u0_uk_K_r3_reg[18]/NET0131  , \u0_uk_K_r3_reg[19]/NET0131  , \u0_uk_K_r3_reg[1]/NET0131  , \u0_uk_K_r3_reg[20]/NET0131  , \u0_uk_K_r3_reg[21]/NET0131  , \u0_uk_K_r3_reg[22]/NET0131  , \u0_uk_K_r3_reg[23]/NET0131  , \u0_uk_K_r3_reg[24]/NET0131  , \u0_uk_K_r3_reg[25]/NET0131  , \u0_uk_K_r3_reg[26]/NET0131  , \u0_uk_K_r3_reg[27]/NET0131  , \u0_uk_K_r3_reg[28]/NET0131  , \u0_uk_K_r3_reg[29]/NET0131  , \u0_uk_K_r3_reg[2]/NET0131  , \u0_uk_K_r3_reg[30]/NET0131  , \u0_uk_K_r3_reg[31]/NET0131  , \u0_uk_K_r3_reg[32]/NET0131  , \u0_uk_K_r3_reg[33]/NET0131  , \u0_uk_K_r3_reg[34]/NET0131  , \u0_uk_K_r3_reg[35]/NET0131  , \u0_uk_K_r3_reg[36]/NET0131  , \u0_uk_K_r3_reg[37]/NET0131  , \u0_uk_K_r3_reg[38]/NET0131  , \u0_uk_K_r3_reg[39]/NET0131  , \u0_uk_K_r3_reg[3]/NET0131  , \u0_uk_K_r3_reg[40]/NET0131  , \u0_uk_K_r3_reg[41]/NET0131  , \u0_uk_K_r3_reg[42]/NET0131  , \u0_uk_K_r3_reg[43]/NET0131  , \u0_uk_K_r3_reg[44]/NET0131  , \u0_uk_K_r3_reg[45]/P0001  , \u0_uk_K_r3_reg[46]/NET0131  , \u0_uk_K_r3_reg[47]/NET0131  , \u0_uk_K_r3_reg[48]/NET0131  , \u0_uk_K_r3_reg[49]/NET0131  , \u0_uk_K_r3_reg[4]/NET0131  , \u0_uk_K_r3_reg[50]/NET0131  , \u0_uk_K_r3_reg[51]/NET0131  , \u0_uk_K_r3_reg[52]/NET0131  , \u0_uk_K_r3_reg[53]/NET0131  , \u0_uk_K_r3_reg[54]/NET0131  , \u0_uk_K_r3_reg[55]/NET0131  , \u0_uk_K_r3_reg[5]/NET0131  , \u0_uk_K_r3_reg[6]/NET0131  , \u0_uk_K_r3_reg[7]/NET0131  , \u0_uk_K_r3_reg[8]/NET0131  , \u0_uk_K_r3_reg[9]/NET0131  , \u0_uk_K_r4_reg[0]/P0001  , \u0_uk_K_r4_reg[10]/NET0131  , \u0_uk_K_r4_reg[11]/NET0131  , \u0_uk_K_r4_reg[12]/NET0131  , \u0_uk_K_r4_reg[13]/NET0131  , \u0_uk_K_r4_reg[14]/NET0131  , \u0_uk_K_r4_reg[15]/NET0131  , \u0_uk_K_r4_reg[16]/NET0131  , \u0_uk_K_r4_reg[17]/NET0131  , \u0_uk_K_r4_reg[18]/NET0131  , \u0_uk_K_r4_reg[19]/NET0131  , \u0_uk_K_r4_reg[1]/NET0131  , \u0_uk_K_r4_reg[20]/NET0131  , \u0_uk_K_r4_reg[21]/NET0131  , \u0_uk_K_r4_reg[22]/NET0131  , \u0_uk_K_r4_reg[23]/P0001  , \u0_uk_K_r4_reg[25]/NET0131  , \u0_uk_K_r4_reg[26]/NET0131  , \u0_uk_K_r4_reg[27]/P0001  , \u0_uk_K_r4_reg[28]/NET0131  , \u0_uk_K_r4_reg[29]/NET0131  , \u0_uk_K_r4_reg[30]/NET0131  , \u0_uk_K_r4_reg[31]/P0001  , \u0_uk_K_r4_reg[32]/NET0131  , \u0_uk_K_r4_reg[33]/NET0131  , \u0_uk_K_r4_reg[34]/NET0131  , \u0_uk_K_r4_reg[35]/NET0131  , \u0_uk_K_r4_reg[36]/NET0131  , \u0_uk_K_r4_reg[37]/NET0131  , \u0_uk_K_r4_reg[38]/NET0131  , \u0_uk_K_r4_reg[39]/NET0131  , \u0_uk_K_r4_reg[3]/NET0131  , \u0_uk_K_r4_reg[40]/NET0131  , \u0_uk_K_r4_reg[41]/NET0131  , \u0_uk_K_r4_reg[42]/NET0131  , \u0_uk_K_r4_reg[43]/NET0131  , \u0_uk_K_r4_reg[44]/NET0131  , \u0_uk_K_r4_reg[45]/NET0131  , \u0_uk_K_r4_reg[46]/NET0131  , \u0_uk_K_r4_reg[47]/NET0131  , \u0_uk_K_r4_reg[48]/NET0131  , \u0_uk_K_r4_reg[49]/NET0131  , \u0_uk_K_r4_reg[4]/NET0131  , \u0_uk_K_r4_reg[50]/NET0131  , \u0_uk_K_r4_reg[51]/NET0131  , \u0_uk_K_r4_reg[52]/NET0131  , \u0_uk_K_r4_reg[53]/NET0131  , \u0_uk_K_r4_reg[54]/NET0131  , \u0_uk_K_r4_reg[55]/NET0131  , \u0_uk_K_r4_reg[5]/NET0131  , \u0_uk_K_r4_reg[6]/NET0131  , \u0_uk_K_r4_reg[7]/NET0131  , \u0_uk_K_r4_reg[8]/NET0131  , \u0_uk_K_r4_reg[9]/NET0131  , \u0_uk_K_r5_reg[0]/NET0131  , \u0_uk_K_r5_reg[10]/NET0131  , \u0_uk_K_r5_reg[11]/NET0131  , \u0_uk_K_r5_reg[12]/NET0131  , \u0_uk_K_r5_reg[13]/P0001  , \u0_uk_K_r5_reg[14]/NET0131  , \u0_uk_K_r5_reg[15]/NET0131  , \u0_uk_K_r5_reg[16]/NET0131  , \u0_uk_K_r5_reg[17]/NET0131  , \u0_uk_K_r5_reg[18]/NET0131  , \u0_uk_K_r5_reg[19]/NET0131  , \u0_uk_K_r5_reg[1]/NET0131  , \u0_uk_K_r5_reg[20]/NET0131  , \u0_uk_K_r5_reg[21]/NET0131  , \u0_uk_K_r5_reg[22]/NET0131  , \u0_uk_K_r5_reg[23]/NET0131  , \u0_uk_K_r5_reg[24]/NET0131  , \u0_uk_K_r5_reg[25]/NET0131  , \u0_uk_K_r5_reg[26]/NET0131  , \u0_uk_K_r5_reg[27]/NET0131  , \u0_uk_K_r5_reg[28]/NET0131  , \u0_uk_K_r5_reg[29]/NET0131  , \u0_uk_K_r5_reg[2]/NET0131  , \u0_uk_K_r5_reg[30]/NET0131  , \u0_uk_K_r5_reg[31]/NET0131  , \u0_uk_K_r5_reg[32]/NET0131  , \u0_uk_K_r5_reg[33]/NET0131  , \u0_uk_K_r5_reg[34]/NET0131  , \u0_uk_K_r5_reg[35]/NET0131  , \u0_uk_K_r5_reg[36]/NET0131  , \u0_uk_K_r5_reg[37]/P0001  , \u0_uk_K_r5_reg[38]/NET0131  , \u0_uk_K_r5_reg[39]/NET0131  , \u0_uk_K_r5_reg[3]/NET0131  , \u0_uk_K_r5_reg[40]/NET0131  , \u0_uk_K_r5_reg[41]/NET0131  , \u0_uk_K_r5_reg[42]/NET0131  , \u0_uk_K_r5_reg[43]/NET0131  , \u0_uk_K_r5_reg[44]/NET0131  , \u0_uk_K_r5_reg[46]/NET0131  , \u0_uk_K_r5_reg[47]/NET0131  , \u0_uk_K_r5_reg[48]/NET0131  , \u0_uk_K_r5_reg[49]/NET0131  , \u0_uk_K_r5_reg[4]/NET0131  , \u0_uk_K_r5_reg[50]/NET0131  , \u0_uk_K_r5_reg[51]/NET0131  , \u0_uk_K_r5_reg[52]/NET0131  , \u0_uk_K_r5_reg[53]/NET0131  , \u0_uk_K_r5_reg[54]/NET0131  , \u0_uk_K_r5_reg[55]/NET0131  , \u0_uk_K_r5_reg[5]/NET0131  , \u0_uk_K_r5_reg[6]/NET0131  , \u0_uk_K_r5_reg[7]/NET0131  , \u0_uk_K_r5_reg[8]/NET0131  , \u0_uk_K_r5_reg[9]/NET0131  , \u0_uk_K_r6_reg[0]/NET0131  , \u0_uk_K_r6_reg[10]/NET0131  , \u0_uk_K_r6_reg[11]/NET0131  , \u0_uk_K_r6_reg[12]/NET0131  , \u0_uk_K_r6_reg[13]/NET0131  , \u0_uk_K_r6_reg[14]/NET0131  , \u0_uk_K_r6_reg[15]/NET0131  , \u0_uk_K_r6_reg[16]/NET0131  , \u0_uk_K_r6_reg[17]/NET0131  , \u0_uk_K_r6_reg[18]/NET0131  , \u0_uk_K_r6_reg[19]/NET0131  , \u0_uk_K_r6_reg[1]/NET0131  , \u0_uk_K_r6_reg[20]/NET0131  , \u0_uk_K_r6_reg[21]/NET0131  , \u0_uk_K_r6_reg[22]/NET0131  , \u0_uk_K_r6_reg[23]/P0001  , \u0_uk_K_r6_reg[24]/NET0131  , \u0_uk_K_r6_reg[25]/NET0131  , \u0_uk_K_r6_reg[26]/P0001  , \u0_uk_K_r6_reg[27]/NET0131  , \u0_uk_K_r6_reg[28]/NET0131  , \u0_uk_K_r6_reg[29]/NET0131  , \u0_uk_K_r6_reg[2]/NET0131  , \u0_uk_K_r6_reg[30]/P0001  , \u0_uk_K_r6_reg[31]/NET0131  , \u0_uk_K_r6_reg[32]/NET0131  , \u0_uk_K_r6_reg[33]/NET0131  , \u0_uk_K_r6_reg[34]/NET0131  , \u0_uk_K_r6_reg[35]/NET0131  , \u0_uk_K_r6_reg[36]/NET0131  , \u0_uk_K_r6_reg[37]/NET0131  , \u0_uk_K_r6_reg[38]/NET0131  , \u0_uk_K_r6_reg[39]/NET0131  , \u0_uk_K_r6_reg[3]/NET0131  , \u0_uk_K_r6_reg[40]/NET0131  , \u0_uk_K_r6_reg[41]/NET0131  , \u0_uk_K_r6_reg[42]/NET0131  , \u0_uk_K_r6_reg[43]/NET0131  , \u0_uk_K_r6_reg[44]/NET0131  , \u0_uk_K_r6_reg[45]/NET0131  , \u0_uk_K_r6_reg[46]/NET0131  , \u0_uk_K_r6_reg[47]/NET0131  , \u0_uk_K_r6_reg[48]/NET0131  , \u0_uk_K_r6_reg[49]/NET0131  , \u0_uk_K_r6_reg[4]/NET0131  , \u0_uk_K_r6_reg[50]/NET0131  , \u0_uk_K_r6_reg[51]/NET0131  , \u0_uk_K_r6_reg[52]/NET0131  , \u0_uk_K_r6_reg[53]/NET0131  , \u0_uk_K_r6_reg[54]/NET0131  , \u0_uk_K_r6_reg[55]/P0001  , \u0_uk_K_r6_reg[5]/NET0131  , \u0_uk_K_r6_reg[6]/NET0131  , \u0_uk_K_r6_reg[7]/NET0131  , \u0_uk_K_r6_reg[8]/NET0131  , \u0_uk_K_r6_reg[9]/NET0131  , \u0_uk_K_r7_reg[0]/NET0131  , \u0_uk_K_r7_reg[10]/NET0131  , \u0_uk_K_r7_reg[11]/NET0131  , \u0_uk_K_r7_reg[12]/NET0131  , \u0_uk_K_r7_reg[13]/NET0131  , \u0_uk_K_r7_reg[14]/NET0131  , \u0_uk_K_r7_reg[15]/NET0131  , \u0_uk_K_r7_reg[16]/NET0131  , \u0_uk_K_r7_reg[17]/NET0131  , \u0_uk_K_r7_reg[18]/NET0131  , \u0_uk_K_r7_reg[19]/NET0131  , \u0_uk_K_r7_reg[1]/NET0131  , \u0_uk_K_r7_reg[20]/NET0131  , \u0_uk_K_r7_reg[21]/NET0131  , \u0_uk_K_r7_reg[22]/NET0131  , \u0_uk_K_r7_reg[23]/P0001  , \u0_uk_K_r7_reg[24]/NET0131  , \u0_uk_K_r7_reg[25]/NET0131  , \u0_uk_K_r7_reg[26]/P0001  , \u0_uk_K_r7_reg[27]/NET0131  , \u0_uk_K_r7_reg[28]/NET0131  , \u0_uk_K_r7_reg[29]/NET0131  , \u0_uk_K_r7_reg[2]/NET0131  , \u0_uk_K_r7_reg[30]/P0001  , \u0_uk_K_r7_reg[31]/NET0131  , \u0_uk_K_r7_reg[32]/NET0131  , \u0_uk_K_r7_reg[33]/NET0131  , \u0_uk_K_r7_reg[34]/NET0131  , \u0_uk_K_r7_reg[35]/NET0131  , \u0_uk_K_r7_reg[36]/NET0131  , \u0_uk_K_r7_reg[37]/NET0131  , \u0_uk_K_r7_reg[38]/NET0131  , \u0_uk_K_r7_reg[39]/NET0131  , \u0_uk_K_r7_reg[3]/NET0131  , \u0_uk_K_r7_reg[40]/NET0131  , \u0_uk_K_r7_reg[41]/NET0131  , \u0_uk_K_r7_reg[42]/NET0131  , \u0_uk_K_r7_reg[43]/NET0131  , \u0_uk_K_r7_reg[44]/NET0131  , \u0_uk_K_r7_reg[45]/NET0131  , \u0_uk_K_r7_reg[46]/NET0131  , \u0_uk_K_r7_reg[47]/NET0131  , \u0_uk_K_r7_reg[48]/NET0131  , \u0_uk_K_r7_reg[49]/NET0131  , \u0_uk_K_r7_reg[4]/NET0131  , \u0_uk_K_r7_reg[50]/NET0131  , \u0_uk_K_r7_reg[51]/NET0131  , \u0_uk_K_r7_reg[52]/NET0131  , \u0_uk_K_r7_reg[53]/NET0131  , \u0_uk_K_r7_reg[54]/NET0131  , \u0_uk_K_r7_reg[55]/P0001  , \u0_uk_K_r7_reg[5]/NET0131  , \u0_uk_K_r7_reg[6]/NET0131  , \u0_uk_K_r7_reg[7]/NET0131  , \u0_uk_K_r7_reg[8]/NET0131  , \u0_uk_K_r7_reg[9]/NET0131  , \u0_uk_K_r8_reg[0]/NET0131  , \u0_uk_K_r8_reg[10]/NET0131  , \u0_uk_K_r8_reg[11]/NET0131  , \u0_uk_K_r8_reg[12]/NET0131  , \u0_uk_K_r8_reg[13]/P0001  , \u0_uk_K_r8_reg[14]/NET0131  , \u0_uk_K_r8_reg[15]/NET0131  , \u0_uk_K_r8_reg[16]/NET0131  , \u0_uk_K_r8_reg[17]/NET0131  , \u0_uk_K_r8_reg[18]/NET0131  , \u0_uk_K_r8_reg[19]/NET0131  , \u0_uk_K_r8_reg[1]/NET0131  , \u0_uk_K_r8_reg[20]/NET0131  , \u0_uk_K_r8_reg[21]/NET0131  , \u0_uk_K_r8_reg[22]/NET0131  , \u0_uk_K_r8_reg[23]/NET0131  , \u0_uk_K_r8_reg[24]/NET0131  , \u0_uk_K_r8_reg[25]/NET0131  , \u0_uk_K_r8_reg[26]/NET0131  , \u0_uk_K_r8_reg[27]/NET0131  , \u0_uk_K_r8_reg[28]/NET0131  , \u0_uk_K_r8_reg[29]/NET0131  , \u0_uk_K_r8_reg[2]/NET0131  , \u0_uk_K_r8_reg[30]/NET0131  , \u0_uk_K_r8_reg[31]/NET0131  , \u0_uk_K_r8_reg[32]/NET0131  , \u0_uk_K_r8_reg[33]/NET0131  , \u0_uk_K_r8_reg[34]/NET0131  , \u0_uk_K_r8_reg[35]/NET0131  , \u0_uk_K_r8_reg[36]/NET0131  , \u0_uk_K_r8_reg[37]/P0001  , \u0_uk_K_r8_reg[38]/NET0131  , \u0_uk_K_r8_reg[39]/NET0131  , \u0_uk_K_r8_reg[3]/NET0131  , \u0_uk_K_r8_reg[40]/NET0131  , \u0_uk_K_r8_reg[41]/NET0131  , \u0_uk_K_r8_reg[42]/NET0131  , \u0_uk_K_r8_reg[43]/NET0131  , \u0_uk_K_r8_reg[44]/NET0131  , \u0_uk_K_r8_reg[46]/NET0131  , \u0_uk_K_r8_reg[47]/NET0131  , \u0_uk_K_r8_reg[48]/NET0131  , \u0_uk_K_r8_reg[49]/NET0131  , \u0_uk_K_r8_reg[4]/NET0131  , \u0_uk_K_r8_reg[50]/NET0131  , \u0_uk_K_r8_reg[51]/NET0131  , \u0_uk_K_r8_reg[52]/NET0131  , \u0_uk_K_r8_reg[53]/NET0131  , \u0_uk_K_r8_reg[54]/NET0131  , \u0_uk_K_r8_reg[55]/NET0131  , \u0_uk_K_r8_reg[5]/NET0131  , \u0_uk_K_r8_reg[6]/NET0131  , \u0_uk_K_r8_reg[7]/NET0131  , \u0_uk_K_r8_reg[8]/NET0131  , \u0_uk_K_r8_reg[9]/P0001  , \u0_uk_K_r9_reg[0]/P0001  , \u0_uk_K_r9_reg[10]/NET0131  , \u0_uk_K_r9_reg[11]/NET0131  , \u0_uk_K_r9_reg[12]/NET0131  , \u0_uk_K_r9_reg[13]/NET0131  , \u0_uk_K_r9_reg[14]/NET0131  , \u0_uk_K_r9_reg[15]/NET0131  , \u0_uk_K_r9_reg[16]/NET0131  , \u0_uk_K_r9_reg[17]/NET0131  , \u0_uk_K_r9_reg[18]/NET0131  , \u0_uk_K_r9_reg[19]/NET0131  , \u0_uk_K_r9_reg[1]/NET0131  , \u0_uk_K_r9_reg[20]/NET0131  , \u0_uk_K_r9_reg[21]/NET0131  , \u0_uk_K_r9_reg[22]/NET0131  , \u0_uk_K_r9_reg[23]/P0001  , \u0_uk_K_r9_reg[25]/NET0131  , \u0_uk_K_r9_reg[26]/NET0131  , \u0_uk_K_r9_reg[27]/P0001  , \u0_uk_K_r9_reg[28]/NET0131  , \u0_uk_K_r9_reg[29]/NET0131  , \u0_uk_K_r9_reg[30]/NET0131  , \u0_uk_K_r9_reg[31]/P0001  , \u0_uk_K_r9_reg[32]/NET0131  , \u0_uk_K_r9_reg[33]/NET0131  , \u0_uk_K_r9_reg[34]/NET0131  , \u0_uk_K_r9_reg[35]/NET0131  , \u0_uk_K_r9_reg[36]/NET0131  , \u0_uk_K_r9_reg[37]/NET0131  , \u0_uk_K_r9_reg[38]/NET0131  , \u0_uk_K_r9_reg[39]/NET0131  , \u0_uk_K_r9_reg[3]/NET0131  , \u0_uk_K_r9_reg[40]/NET0131  , \u0_uk_K_r9_reg[41]/NET0131  , \u0_uk_K_r9_reg[42]/NET0131  , \u0_uk_K_r9_reg[43]/NET0131  , \u0_uk_K_r9_reg[44]/NET0131  , \u0_uk_K_r9_reg[45]/NET0131  , \u0_uk_K_r9_reg[46]/NET0131  , \u0_uk_K_r9_reg[47]/NET0131  , \u0_uk_K_r9_reg[48]/NET0131  , \u0_uk_K_r9_reg[49]/NET0131  , \u0_uk_K_r9_reg[4]/NET0131  , \u0_uk_K_r9_reg[50]/NET0131  , \u0_uk_K_r9_reg[51]/NET0131  , \u0_uk_K_r9_reg[52]/NET0131  , \u0_uk_K_r9_reg[53]/NET0131  , \u0_uk_K_r9_reg[54]/NET0131  , \u0_uk_K_r9_reg[55]/NET0131  , \u0_uk_K_r9_reg[5]/NET0131  , \u0_uk_K_r9_reg[6]/NET0131  , \u0_uk_K_r9_reg[7]/NET0131  , \u0_uk_K_r9_reg[8]/NET0131  , \u0_uk_K_r9_reg[9]/NET0131  , \u1_L0_reg[10]/NET0131  , \u1_L0_reg[11]/NET0131  , \u1_L0_reg[12]/NET0131  , \u1_L0_reg[13]/NET0131  , \u1_L0_reg[14]/NET0131  , \u1_L0_reg[15]/P0001  , \u1_L0_reg[16]/NET0131  , \u1_L0_reg[17]/NET0131  , \u1_L0_reg[18]/NET0131  , \u1_L0_reg[19]/NET0131  , \u1_L0_reg[1]/NET0131  , \u1_L0_reg[20]/NET0131  , \u1_L0_reg[21]/NET0131  , \u1_L0_reg[22]/NET0131  , \u1_L0_reg[23]/NET0131  , \u1_L0_reg[24]/NET0131  , \u1_L0_reg[25]/NET0131  , \u1_L0_reg[26]/NET0131  , \u1_L0_reg[27]/NET0131  , \u1_L0_reg[28]/NET0131  , \u1_L0_reg[29]/NET0131  , \u1_L0_reg[2]/NET0131  , \u1_L0_reg[30]/NET0131  , \u1_L0_reg[31]/NET0131  , \u1_L0_reg[32]/NET0131  , \u1_L0_reg[3]/NET0131  , \u1_L0_reg[4]/NET0131  , \u1_L0_reg[5]/NET0131  , \u1_L0_reg[6]/NET0131  , \u1_L0_reg[7]/NET0131  , \u1_L0_reg[8]/NET0131  , \u1_L0_reg[9]/NET0131  , \u1_L10_reg[10]/NET0131  , \u1_L10_reg[11]/NET0131  , \u1_L10_reg[12]/NET0131  , \u1_L10_reg[13]/NET0131  , \u1_L10_reg[14]/NET0131  , \u1_L10_reg[15]/P0001  , \u1_L10_reg[16]/NET0131  , \u1_L10_reg[17]/NET0131  , \u1_L10_reg[18]/P0001  , \u1_L10_reg[19]/P0001  , \u1_L10_reg[1]/NET0131  , \u1_L10_reg[20]/NET0131  , \u1_L10_reg[21]/NET0131  , \u1_L10_reg[22]/NET0131  , \u1_L10_reg[23]/NET0131  , \u1_L10_reg[24]/NET0131  , \u1_L10_reg[25]/NET0131  , \u1_L10_reg[26]/NET0131  , \u1_L10_reg[27]/NET0131  , \u1_L10_reg[28]/NET0131  , \u1_L10_reg[29]/NET0131  , \u1_L10_reg[2]/NET0131  , \u1_L10_reg[30]/NET0131  , \u1_L10_reg[31]/NET0131  , \u1_L10_reg[32]/NET0131  , \u1_L10_reg[3]/NET0131  , \u1_L10_reg[4]/NET0131  , \u1_L10_reg[5]/NET0131  , \u1_L10_reg[6]/NET0131  , \u1_L10_reg[7]/NET0131  , \u1_L10_reg[8]/NET0131  , \u1_L10_reg[9]/NET0131  , \u1_L11_reg[10]/NET0131  , \u1_L11_reg[11]/NET0131  , \u1_L11_reg[12]/NET0131  , \u1_L11_reg[13]/NET0131  , \u1_L11_reg[14]/NET0131  , \u1_L11_reg[15]/P0001  , \u1_L11_reg[16]/NET0131  , \u1_L11_reg[17]/NET0131  , \u1_L11_reg[18]/P0001  , \u1_L11_reg[19]/P0001  , \u1_L11_reg[1]/NET0131  , \u1_L11_reg[20]/NET0131  , \u1_L11_reg[21]/NET0131  , \u1_L11_reg[22]/NET0131  , \u1_L11_reg[23]/NET0131  , \u1_L11_reg[24]/NET0131  , \u1_L11_reg[25]/NET0131  , \u1_L11_reg[26]/NET0131  , \u1_L11_reg[27]/NET0131  , \u1_L11_reg[28]/NET0131  , \u1_L11_reg[29]/NET0131  , \u1_L11_reg[2]/NET0131  , \u1_L11_reg[30]/NET0131  , \u1_L11_reg[31]/NET0131  , \u1_L11_reg[32]/NET0131  , \u1_L11_reg[3]/NET0131  , \u1_L11_reg[4]/NET0131  , \u1_L11_reg[5]/NET0131  , \u1_L11_reg[6]/NET0131  , \u1_L11_reg[7]/NET0131  , \u1_L11_reg[8]/NET0131  , \u1_L11_reg[9]/NET0131  , \u1_L12_reg[10]/NET0131  , \u1_L12_reg[11]/NET0131  , \u1_L12_reg[12]/NET0131  , \u1_L12_reg[13]/NET0131  , \u1_L12_reg[14]/NET0131  , \u1_L12_reg[15]/P0001  , \u1_L12_reg[16]/NET0131  , \u1_L12_reg[17]/NET0131  , \u1_L12_reg[18]/P0001  , \u1_L12_reg[19]/NET0131  , \u1_L12_reg[1]/NET0131  , \u1_L12_reg[20]/NET0131  , \u1_L12_reg[21]/NET0131  , \u1_L12_reg[22]/NET0131  , \u1_L12_reg[23]/P0001  , \u1_L12_reg[24]/NET0131  , \u1_L12_reg[25]/NET0131  , \u1_L12_reg[26]/NET0131  , \u1_L12_reg[27]/NET0131  , \u1_L12_reg[28]/NET0131  , \u1_L12_reg[29]/NET0131  , \u1_L12_reg[2]/NET0131  , \u1_L12_reg[30]/NET0131  , \u1_L12_reg[31]/NET0131  , \u1_L12_reg[32]/NET0131  , \u1_L12_reg[3]/NET0131  , \u1_L12_reg[4]/NET0131  , \u1_L12_reg[5]/NET0131  , \u1_L12_reg[6]/NET0131  , \u1_L12_reg[7]/NET0131  , \u1_L12_reg[8]/NET0131  , \u1_L12_reg[9]/NET0131  , \u1_L13_reg[10]/NET0131  , \u1_L13_reg[11]/NET0131  , \u1_L13_reg[12]/NET0131  , \u1_L13_reg[13]/NET0131  , \u1_L13_reg[14]/NET0131  , \u1_L13_reg[15]/P0001  , \u1_L13_reg[16]/NET0131  , \u1_L13_reg[17]/NET0131  , \u1_L13_reg[18]/P0001  , \u1_L13_reg[19]/P0001  , \u1_L13_reg[1]/NET0131  , \u1_L13_reg[20]/NET0131  , \u1_L13_reg[21]/NET0131  , \u1_L13_reg[22]/NET0131  , \u1_L13_reg[23]/P0001  , \u1_L13_reg[24]/NET0131  , \u1_L13_reg[25]/NET0131  , \u1_L13_reg[26]/NET0131  , \u1_L13_reg[27]/NET0131  , \u1_L13_reg[28]/NET0131  , \u1_L13_reg[29]/NET0131  , \u1_L13_reg[2]/NET0131  , \u1_L13_reg[30]/NET0131  , \u1_L13_reg[31]/NET0131  , \u1_L13_reg[32]/NET0131  , \u1_L13_reg[3]/NET0131  , \u1_L13_reg[4]/NET0131  , \u1_L13_reg[5]/NET0131  , \u1_L13_reg[6]/NET0131  , \u1_L13_reg[7]/NET0131  , \u1_L13_reg[8]/NET0131  , \u1_L13_reg[9]/NET0131  , \u1_L14_reg[10]/P0001  , \u1_L14_reg[11]/P0001  , \u1_L14_reg[12]/P0001  , \u1_L14_reg[13]/P0001  , \u1_L14_reg[14]/P0001  , \u1_L14_reg[15]/P0001  , \u1_L14_reg[16]/P0001  , \u1_L14_reg[17]/P0001  , \u1_L14_reg[18]/P0001  , \u1_L14_reg[19]/P0001  , \u1_L14_reg[1]/P0001  , \u1_L14_reg[20]/P0001  , \u1_L14_reg[21]/P0001  , \u1_L14_reg[22]/P0001  , \u1_L14_reg[23]/P0001  , \u1_L14_reg[24]/P0001  , \u1_L14_reg[25]/P0001  , \u1_L14_reg[26]/P0001  , \u1_L14_reg[27]/P0001  , \u1_L14_reg[28]/P0001  , \u1_L14_reg[29]/P0001  , \u1_L14_reg[2]/P0001  , \u1_L14_reg[30]/P0001  , \u1_L14_reg[31]/P0001  , \u1_L14_reg[32]/P0001  , \u1_L14_reg[3]/P0001  , \u1_L14_reg[4]/P0001  , \u1_L14_reg[5]/P0001  , \u1_L14_reg[6]/P0001  , \u1_L14_reg[7]/P0001  , \u1_L14_reg[8]/P0001  , \u1_L14_reg[9]/P0001  , \u1_L1_reg[10]/NET0131  , \u1_L1_reg[11]/NET0131  , \u1_L1_reg[12]/NET0131  , \u1_L1_reg[13]/NET0131  , \u1_L1_reg[14]/NET0131  , \u1_L1_reg[15]/P0001  , \u1_L1_reg[16]/NET0131  , \u1_L1_reg[17]/NET0131  , \u1_L1_reg[18]/NET0131  , \u1_L1_reg[19]/P0001  , \u1_L1_reg[1]/NET0131  , \u1_L1_reg[20]/NET0131  , \u1_L1_reg[21]/NET0131  , \u1_L1_reg[22]/NET0131  , \u1_L1_reg[23]/NET0131  , \u1_L1_reg[24]/NET0131  , \u1_L1_reg[25]/NET0131  , \u1_L1_reg[26]/NET0131  , \u1_L1_reg[27]/NET0131  , \u1_L1_reg[28]/NET0131  , \u1_L1_reg[29]/NET0131  , \u1_L1_reg[2]/NET0131  , \u1_L1_reg[30]/NET0131  , \u1_L1_reg[31]/NET0131  , \u1_L1_reg[32]/NET0131  , \u1_L1_reg[3]/NET0131  , \u1_L1_reg[4]/NET0131  , \u1_L1_reg[5]/NET0131  , \u1_L1_reg[6]/NET0131  , \u1_L1_reg[7]/NET0131  , \u1_L1_reg[8]/NET0131  , \u1_L1_reg[9]/NET0131  , \u1_L2_reg[10]/NET0131  , \u1_L2_reg[11]/NET0131  , \u1_L2_reg[12]/NET0131  , \u1_L2_reg[13]/NET0131  , \u1_L2_reg[14]/NET0131  , \u1_L2_reg[15]/P0001  , \u1_L2_reg[16]/NET0131  , \u1_L2_reg[17]/NET0131  , \u1_L2_reg[18]/NET0131  , \u1_L2_reg[19]/NET0131  , \u1_L2_reg[1]/NET0131  , \u1_L2_reg[20]/NET0131  , \u1_L2_reg[21]/NET0131  , \u1_L2_reg[22]/NET0131  , \u1_L2_reg[23]/NET0131  , \u1_L2_reg[24]/NET0131  , \u1_L2_reg[25]/NET0131  , \u1_L2_reg[26]/NET0131  , \u1_L2_reg[27]/NET0131  , \u1_L2_reg[28]/NET0131  , \u1_L2_reg[29]/NET0131  , \u1_L2_reg[2]/NET0131  , \u1_L2_reg[30]/NET0131  , \u1_L2_reg[31]/NET0131  , \u1_L2_reg[32]/NET0131  , \u1_L2_reg[3]/NET0131  , \u1_L2_reg[4]/NET0131  , \u1_L2_reg[5]/NET0131  , \u1_L2_reg[6]/NET0131  , \u1_L2_reg[7]/NET0131  , \u1_L2_reg[8]/NET0131  , \u1_L2_reg[9]/NET0131  , \u1_L3_reg[10]/NET0131  , \u1_L3_reg[11]/NET0131  , \u1_L3_reg[12]/NET0131  , \u1_L3_reg[13]/NET0131  , \u1_L3_reg[14]/NET0131  , \u1_L3_reg[15]/P0001  , \u1_L3_reg[16]/NET0131  , \u1_L3_reg[17]/NET0131  , \u1_L3_reg[18]/NET0131  , \u1_L3_reg[19]/NET0131  , \u1_L3_reg[1]/NET0131  , \u1_L3_reg[20]/NET0131  , \u1_L3_reg[21]/NET0131  , \u1_L3_reg[22]/NET0131  , \u1_L3_reg[23]/NET0131  , \u1_L3_reg[24]/NET0131  , \u1_L3_reg[25]/NET0131  , \u1_L3_reg[26]/NET0131  , \u1_L3_reg[27]/NET0131  , \u1_L3_reg[28]/NET0131  , \u1_L3_reg[29]/NET0131  , \u1_L3_reg[2]/NET0131  , \u1_L3_reg[30]/NET0131  , \u1_L3_reg[31]/NET0131  , \u1_L3_reg[32]/NET0131  , \u1_L3_reg[3]/NET0131  , \u1_L3_reg[4]/NET0131  , \u1_L3_reg[5]/NET0131  , \u1_L3_reg[6]/NET0131  , \u1_L3_reg[7]/NET0131  , \u1_L3_reg[8]/NET0131  , \u1_L3_reg[9]/NET0131  , \u1_L4_reg[10]/NET0131  , \u1_L4_reg[11]/P0001  , \u1_L4_reg[12]/NET0131  , \u1_L4_reg[13]/NET0131  , \u1_L4_reg[14]/NET0131  , \u1_L4_reg[15]/P0001  , \u1_L4_reg[16]/NET0131  , \u1_L4_reg[17]/NET0131  , \u1_L4_reg[18]/NET0131  , \u1_L4_reg[19]/P0001  , \u1_L4_reg[1]/NET0131  , \u1_L4_reg[20]/NET0131  , \u1_L4_reg[21]/NET0131  , \u1_L4_reg[22]/NET0131  , \u1_L4_reg[23]/NET0131  , \u1_L4_reg[24]/NET0131  , \u1_L4_reg[25]/NET0131  , \u1_L4_reg[26]/NET0131  , \u1_L4_reg[27]/NET0131  , \u1_L4_reg[28]/NET0131  , \u1_L4_reg[29]/NET0131  , \u1_L4_reg[2]/NET0131  , \u1_L4_reg[30]/NET0131  , \u1_L4_reg[31]/NET0131  , \u1_L4_reg[32]/NET0131  , \u1_L4_reg[3]/NET0131  , \u1_L4_reg[4]/NET0131  , \u1_L4_reg[5]/NET0131  , \u1_L4_reg[6]/NET0131  , \u1_L4_reg[7]/NET0131  , \u1_L4_reg[8]/NET0131  , \u1_L4_reg[9]/NET0131  , \u1_L5_reg[10]/NET0131  , \u1_L5_reg[11]/NET0131  , \u1_L5_reg[12]/NET0131  , \u1_L5_reg[13]/NET0131  , \u1_L5_reg[14]/NET0131  , \u1_L5_reg[15]/P0001  , \u1_L5_reg[16]/NET0131  , \u1_L5_reg[17]/NET0131  , \u1_L5_reg[18]/NET0131  , \u1_L5_reg[19]/NET0131  , \u1_L5_reg[1]/NET0131  , \u1_L5_reg[20]/NET0131  , \u1_L5_reg[21]/NET0131  , \u1_L5_reg[22]/NET0131  , \u1_L5_reg[23]/NET0131  , \u1_L5_reg[24]/NET0131  , \u1_L5_reg[25]/NET0131  , \u1_L5_reg[26]/NET0131  , \u1_L5_reg[27]/NET0131  , \u1_L5_reg[28]/NET0131  , \u1_L5_reg[29]/NET0131  , \u1_L5_reg[2]/NET0131  , \u1_L5_reg[30]/NET0131  , \u1_L5_reg[31]/NET0131  , \u1_L5_reg[32]/NET0131  , \u1_L5_reg[3]/NET0131  , \u1_L5_reg[4]/NET0131  , \u1_L5_reg[5]/NET0131  , \u1_L5_reg[6]/NET0131  , \u1_L5_reg[7]/NET0131  , \u1_L5_reg[8]/NET0131  , \u1_L5_reg[9]/NET0131  , \u1_L6_reg[10]/NET0131  , \u1_L6_reg[11]/NET0131  , \u1_L6_reg[12]/NET0131  , \u1_L6_reg[13]/NET0131  , \u1_L6_reg[14]/NET0131  , \u1_L6_reg[15]/P0001  , \u1_L6_reg[16]/NET0131  , \u1_L6_reg[17]/NET0131  , \u1_L6_reg[18]/NET0131  , \u1_L6_reg[19]/NET0131  , \u1_L6_reg[1]/NET0131  , \u1_L6_reg[20]/NET0131  , \u1_L6_reg[21]/NET0131  , \u1_L6_reg[22]/NET0131  , \u1_L6_reg[23]/NET0131  , \u1_L6_reg[24]/NET0131  , \u1_L6_reg[25]/NET0131  , \u1_L6_reg[26]/NET0131  , \u1_L6_reg[27]/NET0131  , \u1_L6_reg[28]/NET0131  , \u1_L6_reg[29]/NET0131  , \u1_L6_reg[2]/NET0131  , \u1_L6_reg[30]/NET0131  , \u1_L6_reg[31]/NET0131  , \u1_L6_reg[32]/NET0131  , \u1_L6_reg[3]/NET0131  , \u1_L6_reg[4]/NET0131  , \u1_L6_reg[5]/NET0131  , \u1_L6_reg[6]/NET0131  , \u1_L6_reg[7]/NET0131  , \u1_L6_reg[8]/NET0131  , \u1_L6_reg[9]/NET0131  , \u1_L7_reg[10]/NET0131  , \u1_L7_reg[11]/NET0131  , \u1_L7_reg[12]/NET0131  , \u1_L7_reg[13]/NET0131  , \u1_L7_reg[14]/NET0131  , \u1_L7_reg[15]/P0001  , \u1_L7_reg[16]/NET0131  , \u1_L7_reg[17]/NET0131  , \u1_L7_reg[18]/NET0131  , \u1_L7_reg[19]/P0001  , \u1_L7_reg[1]/NET0131  , \u1_L7_reg[20]/NET0131  , \u1_L7_reg[21]/NET0131  , \u1_L7_reg[22]/NET0131  , \u1_L7_reg[23]/NET0131  , \u1_L7_reg[24]/NET0131  , \u1_L7_reg[25]/NET0131  , \u1_L7_reg[26]/NET0131  , \u1_L7_reg[27]/NET0131  , \u1_L7_reg[28]/NET0131  , \u1_L7_reg[29]/NET0131  , \u1_L7_reg[2]/NET0131  , \u1_L7_reg[30]/NET0131  , \u1_L7_reg[31]/NET0131  , \u1_L7_reg[32]/NET0131  , \u1_L7_reg[3]/NET0131  , \u1_L7_reg[4]/NET0131  , \u1_L7_reg[5]/NET0131  , \u1_L7_reg[6]/NET0131  , \u1_L7_reg[7]/NET0131  , \u1_L7_reg[8]/NET0131  , \u1_L7_reg[9]/NET0131  , \u1_L8_reg[10]/NET0131  , \u1_L8_reg[11]/NET0131  , \u1_L8_reg[12]/NET0131  , \u1_L8_reg[13]/NET0131  , \u1_L8_reg[14]/NET0131  , \u1_L8_reg[15]/P0001  , \u1_L8_reg[16]/NET0131  , \u1_L8_reg[17]/NET0131  , \u1_L8_reg[18]/NET0131  , \u1_L8_reg[19]/P0001  , \u1_L8_reg[1]/NET0131  , \u1_L8_reg[20]/NET0131  , \u1_L8_reg[21]/NET0131  , \u1_L8_reg[22]/NET0131  , \u1_L8_reg[23]/NET0131  , \u1_L8_reg[24]/NET0131  , \u1_L8_reg[25]/NET0131  , \u1_L8_reg[26]/NET0131  , \u1_L8_reg[27]/NET0131  , \u1_L8_reg[28]/NET0131  , \u1_L8_reg[29]/NET0131  , \u1_L8_reg[2]/NET0131  , \u1_L8_reg[30]/NET0131  , \u1_L8_reg[31]/NET0131  , \u1_L8_reg[32]/NET0131  , \u1_L8_reg[3]/NET0131  , \u1_L8_reg[4]/NET0131  , \u1_L8_reg[5]/NET0131  , \u1_L8_reg[6]/NET0131  , \u1_L8_reg[7]/NET0131  , \u1_L8_reg[8]/NET0131  , \u1_L8_reg[9]/NET0131  , \u1_L9_reg[10]/NET0131  , \u1_L9_reg[11]/NET0131  , \u1_L9_reg[12]/NET0131  , \u1_L9_reg[13]/NET0131  , \u1_L9_reg[14]/NET0131  , \u1_L9_reg[15]/P0001  , \u1_L9_reg[16]/NET0131  , \u1_L9_reg[17]/NET0131  , \u1_L9_reg[18]/P0001  , \u1_L9_reg[19]/NET0131  , \u1_L9_reg[1]/NET0131  , \u1_L9_reg[20]/NET0131  , \u1_L9_reg[21]/NET0131  , \u1_L9_reg[22]/NET0131  , \u1_L9_reg[23]/NET0131  , \u1_L9_reg[24]/NET0131  , \u1_L9_reg[25]/NET0131  , \u1_L9_reg[26]/NET0131  , \u1_L9_reg[27]/NET0131  , \u1_L9_reg[28]/NET0131  , \u1_L9_reg[29]/NET0131  , \u1_L9_reg[2]/NET0131  , \u1_L9_reg[30]/NET0131  , \u1_L9_reg[31]/NET0131  , \u1_L9_reg[32]/NET0131  , \u1_L9_reg[3]/NET0131  , \u1_L9_reg[4]/NET0131  , \u1_L9_reg[5]/NET0131  , \u1_L9_reg[6]/NET0131  , \u1_L9_reg[7]/NET0131  , \u1_L9_reg[8]/NET0131  , \u1_L9_reg[9]/NET0131  , \u1_R0_reg[10]/NET0131  , \u1_R0_reg[11]/NET0131  , \u1_R0_reg[12]/NET0131  , \u1_R0_reg[13]/NET0131  , \u1_R0_reg[14]/NET0131  , \u1_R0_reg[15]/NET0131  , \u1_R0_reg[16]/NET0131  , \u1_R0_reg[17]/NET0131  , \u1_R0_reg[18]/NET0131  , \u1_R0_reg[19]/NET0131  , \u1_R0_reg[1]/NET0131  , \u1_R0_reg[20]/NET0131  , \u1_R0_reg[21]/NET0131  , \u1_R0_reg[22]/NET0131  , \u1_R0_reg[23]/NET0131  , \u1_R0_reg[24]/NET0131  , \u1_R0_reg[25]/NET0131  , \u1_R0_reg[26]/NET0131  , \u1_R0_reg[27]/NET0131  , \u1_R0_reg[28]/NET0131  , \u1_R0_reg[29]/NET0131  , \u1_R0_reg[2]/NET0131  , \u1_R0_reg[30]/NET0131  , \u1_R0_reg[31]/P0001  , \u1_R0_reg[32]/NET0131  , \u1_R0_reg[3]/NET0131  , \u1_R0_reg[4]/NET0131  , \u1_R0_reg[5]/NET0131  , \u1_R0_reg[6]/NET0131  , \u1_R0_reg[7]/NET0131  , \u1_R0_reg[8]/NET0131  , \u1_R0_reg[9]/NET0131  , \u1_R10_reg[10]/NET0131  , \u1_R10_reg[11]/NET0131  , \u1_R10_reg[12]/NET0131  , \u1_R10_reg[13]/NET0131  , \u1_R10_reg[14]/NET0131  , \u1_R10_reg[15]/NET0131  , \u1_R10_reg[16]/NET0131  , \u1_R10_reg[17]/NET0131  , \u1_R10_reg[18]/NET0131  , \u1_R10_reg[19]/NET0131  , \u1_R10_reg[1]/NET0131  , \u1_R10_reg[20]/NET0131  , \u1_R10_reg[21]/NET0131  , \u1_R10_reg[22]/NET0131  , \u1_R10_reg[23]/NET0131  , \u1_R10_reg[24]/NET0131  , \u1_R10_reg[25]/NET0131  , \u1_R10_reg[26]/NET0131  , \u1_R10_reg[27]/NET0131  , \u1_R10_reg[28]/NET0131  , \u1_R10_reg[29]/NET0131  , \u1_R10_reg[2]/NET0131  , \u1_R10_reg[30]/NET0131  , \u1_R10_reg[31]/P0001  , \u1_R10_reg[32]/NET0131  , \u1_R10_reg[3]/NET0131  , \u1_R10_reg[4]/NET0131  , \u1_R10_reg[5]/NET0131  , \u1_R10_reg[6]/NET0131  , \u1_R10_reg[7]/NET0131  , \u1_R10_reg[8]/NET0131  , \u1_R10_reg[9]/NET0131  , \u1_R11_reg[10]/NET0131  , \u1_R11_reg[11]/NET0131  , \u1_R11_reg[12]/NET0131  , \u1_R11_reg[13]/NET0131  , \u1_R11_reg[14]/NET0131  , \u1_R11_reg[15]/NET0131  , \u1_R11_reg[16]/NET0131  , \u1_R11_reg[17]/NET0131  , \u1_R11_reg[18]/NET0131  , \u1_R11_reg[19]/NET0131  , \u1_R11_reg[1]/NET0131  , \u1_R11_reg[20]/NET0131  , \u1_R11_reg[21]/NET0131  , \u1_R11_reg[22]/NET0131  , \u1_R11_reg[23]/NET0131  , \u1_R11_reg[24]/NET0131  , \u1_R11_reg[25]/NET0131  , \u1_R11_reg[26]/NET0131  , \u1_R11_reg[27]/NET0131  , \u1_R11_reg[28]/NET0131  , \u1_R11_reg[29]/NET0131  , \u1_R11_reg[2]/NET0131  , \u1_R11_reg[30]/NET0131  , \u1_R11_reg[31]/NET0131  , \u1_R11_reg[32]/NET0131  , \u1_R11_reg[3]/NET0131  , \u1_R11_reg[4]/NET0131  , \u1_R11_reg[5]/NET0131  , \u1_R11_reg[6]/NET0131  , \u1_R11_reg[7]/NET0131  , \u1_R11_reg[8]/NET0131  , \u1_R11_reg[9]/NET0131  , \u1_R12_reg[10]/NET0131  , \u1_R12_reg[11]/NET0131  , \u1_R12_reg[12]/NET0131  , \u1_R12_reg[13]/NET0131  , \u1_R12_reg[14]/NET0131  , \u1_R12_reg[15]/NET0131  , \u1_R12_reg[16]/NET0131  , \u1_R12_reg[17]/NET0131  , \u1_R12_reg[18]/NET0131  , \u1_R12_reg[19]/NET0131  , \u1_R12_reg[1]/NET0131  , \u1_R12_reg[20]/NET0131  , \u1_R12_reg[21]/NET0131  , \u1_R12_reg[22]/NET0131  , \u1_R12_reg[23]/NET0131  , \u1_R12_reg[24]/NET0131  , \u1_R12_reg[25]/NET0131  , \u1_R12_reg[26]/NET0131  , \u1_R12_reg[27]/NET0131  , \u1_R12_reg[28]/NET0131  , \u1_R12_reg[29]/NET0131  , \u1_R12_reg[2]/NET0131  , \u1_R12_reg[30]/NET0131  , \u1_R12_reg[31]/NET0131  , \u1_R12_reg[32]/NET0131  , \u1_R12_reg[3]/NET0131  , \u1_R12_reg[4]/NET0131  , \u1_R12_reg[5]/NET0131  , \u1_R12_reg[6]/NET0131  , \u1_R12_reg[7]/NET0131  , \u1_R12_reg[8]/NET0131  , \u1_R12_reg[9]/NET0131  , \u1_R13_reg[10]/NET0131  , \u1_R13_reg[11]/P0001  , \u1_R13_reg[12]/NET0131  , \u1_R13_reg[13]/NET0131  , \u1_R13_reg[14]/NET0131  , \u1_R13_reg[15]/NET0131  , \u1_R13_reg[16]/NET0131  , \u1_R13_reg[17]/NET0131  , \u1_R13_reg[18]/NET0131  , \u1_R13_reg[19]/NET0131  , \u1_R13_reg[1]/NET0131  , \u1_R13_reg[20]/NET0131  , \u1_R13_reg[21]/NET0131  , \u1_R13_reg[22]/NET0131  , \u1_R13_reg[23]/P0001  , \u1_R13_reg[24]/NET0131  , \u1_R13_reg[25]/NET0131  , \u1_R13_reg[26]/NET0131  , \u1_R13_reg[27]/P0001  , \u1_R13_reg[28]/NET0131  , \u1_R13_reg[29]/NET0131  , \u1_R13_reg[2]/NET0131  , \u1_R13_reg[30]/NET0131  , \u1_R13_reg[31]/P0001  , \u1_R13_reg[32]/NET0131  , \u1_R13_reg[3]/NET0131  , \u1_R13_reg[4]/NET0131  , \u1_R13_reg[5]/NET0131  , \u1_R13_reg[6]/NET0131  , \u1_R13_reg[7]/NET0131  , \u1_R13_reg[8]/NET0131  , \u1_R13_reg[9]/NET0131  , \u1_R14_reg[10]/P0001  , \u1_R14_reg[11]/P0001  , \u1_R14_reg[12]/NET0131  , \u1_R14_reg[13]/NET0131  , \u1_R14_reg[14]/NET0131  , \u1_R14_reg[15]/NET0131  , \u1_R14_reg[16]/NET0131  , \u1_R14_reg[17]/NET0131  , \u1_R14_reg[18]/NET0131  , \u1_R14_reg[19]/P0001  , \u1_R14_reg[1]/NET0131  , \u1_R14_reg[20]/NET0131  , \u1_R14_reg[21]/NET0131  , \u1_R14_reg[22]/P0001  , \u1_R14_reg[23]/P0001  , \u1_R14_reg[24]/NET0131  , \u1_R14_reg[25]/NET0131  , \u1_R14_reg[26]/NET0131  , \u1_R14_reg[27]/P0001  , \u1_R14_reg[28]/NET0131  , \u1_R14_reg[29]/NET0131  , \u1_R14_reg[2]/NET0131  , \u1_R14_reg[30]/NET0131  , \u1_R14_reg[31]/P0001  , \u1_R14_reg[32]/NET0131  , \u1_R14_reg[3]/NET0131  , \u1_R14_reg[4]/NET0131  , \u1_R14_reg[5]/NET0131  , \u1_R14_reg[6]/NET0131  , \u1_R14_reg[7]/P0001  , \u1_R14_reg[8]/NET0131  , \u1_R14_reg[9]/NET0131  , \u1_R1_reg[10]/NET0131  , \u1_R1_reg[11]/NET0131  , \u1_R1_reg[12]/NET0131  , \u1_R1_reg[13]/NET0131  , \u1_R1_reg[14]/NET0131  , \u1_R1_reg[15]/NET0131  , \u1_R1_reg[16]/NET0131  , \u1_R1_reg[17]/NET0131  , \u1_R1_reg[18]/NET0131  , \u1_R1_reg[19]/NET0131  , \u1_R1_reg[1]/NET0131  , \u1_R1_reg[20]/NET0131  , \u1_R1_reg[21]/NET0131  , \u1_R1_reg[22]/NET0131  , \u1_R1_reg[23]/NET0131  , \u1_R1_reg[24]/NET0131  , \u1_R1_reg[25]/NET0131  , \u1_R1_reg[26]/NET0131  , \u1_R1_reg[27]/NET0131  , \u1_R1_reg[28]/NET0131  , \u1_R1_reg[29]/NET0131  , \u1_R1_reg[2]/NET0131  , \u1_R1_reg[30]/NET0131  , \u1_R1_reg[31]/P0001  , \u1_R1_reg[32]/NET0131  , \u1_R1_reg[3]/NET0131  , \u1_R1_reg[4]/NET0131  , \u1_R1_reg[5]/NET0131  , \u1_R1_reg[6]/NET0131  , \u1_R1_reg[7]/NET0131  , \u1_R1_reg[8]/NET0131  , \u1_R1_reg[9]/NET0131  , \u1_R2_reg[10]/NET0131  , \u1_R2_reg[11]/NET0131  , \u1_R2_reg[12]/NET0131  , \u1_R2_reg[13]/NET0131  , \u1_R2_reg[14]/NET0131  , \u1_R2_reg[15]/NET0131  , \u1_R2_reg[16]/NET0131  , \u1_R2_reg[17]/NET0131  , \u1_R2_reg[18]/NET0131  , \u1_R2_reg[19]/NET0131  , \u1_R2_reg[1]/NET0131  , \u1_R2_reg[20]/NET0131  , \u1_R2_reg[21]/NET0131  , \u1_R2_reg[22]/NET0131  , \u1_R2_reg[23]/NET0131  , \u1_R2_reg[24]/NET0131  , \u1_R2_reg[25]/NET0131  , \u1_R2_reg[26]/NET0131  , \u1_R2_reg[27]/NET0131  , \u1_R2_reg[28]/NET0131  , \u1_R2_reg[29]/NET0131  , \u1_R2_reg[2]/NET0131  , \u1_R2_reg[30]/NET0131  , \u1_R2_reg[31]/P0001  , \u1_R2_reg[32]/NET0131  , \u1_R2_reg[3]/NET0131  , \u1_R2_reg[4]/NET0131  , \u1_R2_reg[5]/NET0131  , \u1_R2_reg[6]/NET0131  , \u1_R2_reg[7]/NET0131  , \u1_R2_reg[8]/NET0131  , \u1_R2_reg[9]/NET0131  , \u1_R3_reg[10]/NET0131  , \u1_R3_reg[11]/NET0131  , \u1_R3_reg[12]/NET0131  , \u1_R3_reg[13]/NET0131  , \u1_R3_reg[14]/NET0131  , \u1_R3_reg[15]/NET0131  , \u1_R3_reg[16]/NET0131  , \u1_R3_reg[17]/NET0131  , \u1_R3_reg[18]/NET0131  , \u1_R3_reg[19]/NET0131  , \u1_R3_reg[1]/NET0131  , \u1_R3_reg[20]/NET0131  , \u1_R3_reg[21]/NET0131  , \u1_R3_reg[22]/NET0131  , \u1_R3_reg[23]/NET0131  , \u1_R3_reg[24]/NET0131  , \u1_R3_reg[25]/NET0131  , \u1_R3_reg[26]/NET0131  , \u1_R3_reg[27]/NET0131  , \u1_R3_reg[28]/NET0131  , \u1_R3_reg[29]/NET0131  , \u1_R3_reg[2]/NET0131  , \u1_R3_reg[30]/NET0131  , \u1_R3_reg[31]/P0001  , \u1_R3_reg[32]/NET0131  , \u1_R3_reg[3]/NET0131  , \u1_R3_reg[4]/NET0131  , \u1_R3_reg[5]/NET0131  , \u1_R3_reg[6]/NET0131  , \u1_R3_reg[7]/NET0131  , \u1_R3_reg[8]/NET0131  , \u1_R3_reg[9]/NET0131  , \u1_R4_reg[10]/NET0131  , \u1_R4_reg[11]/P0001  , \u1_R4_reg[12]/NET0131  , \u1_R4_reg[13]/NET0131  , \u1_R4_reg[14]/NET0131  , \u1_R4_reg[15]/NET0131  , \u1_R4_reg[16]/NET0131  , \u1_R4_reg[17]/NET0131  , \u1_R4_reg[18]/NET0131  , \u1_R4_reg[19]/NET0131  , \u1_R4_reg[1]/NET0131  , \u1_R4_reg[20]/NET0131  , \u1_R4_reg[21]/NET0131  , \u1_R4_reg[22]/NET0131  , \u1_R4_reg[23]/NET0131  , \u1_R4_reg[24]/NET0131  , \u1_R4_reg[25]/NET0131  , \u1_R4_reg[26]/NET0131  , \u1_R4_reg[27]/NET0131  , \u1_R4_reg[28]/NET0131  , \u1_R4_reg[29]/NET0131  , \u1_R4_reg[2]/NET0131  , \u1_R4_reg[30]/NET0131  , \u1_R4_reg[31]/P0001  , \u1_R4_reg[32]/NET0131  , \u1_R4_reg[3]/NET0131  , \u1_R4_reg[4]/NET0131  , \u1_R4_reg[5]/NET0131  , \u1_R4_reg[6]/NET0131  , \u1_R4_reg[7]/NET0131  , \u1_R4_reg[8]/NET0131  , \u1_R4_reg[9]/NET0131  , \u1_R5_reg[10]/NET0131  , \u1_R5_reg[11]/NET0131  , \u1_R5_reg[12]/NET0131  , \u1_R5_reg[13]/NET0131  , \u1_R5_reg[14]/NET0131  , \u1_R5_reg[15]/NET0131  , \u1_R5_reg[16]/NET0131  , \u1_R5_reg[17]/NET0131  , \u1_R5_reg[18]/NET0131  , \u1_R5_reg[19]/NET0131  , \u1_R5_reg[1]/NET0131  , \u1_R5_reg[20]/NET0131  , \u1_R5_reg[21]/NET0131  , \u1_R5_reg[22]/NET0131  , \u1_R5_reg[23]/NET0131  , \u1_R5_reg[24]/NET0131  , \u1_R5_reg[25]/NET0131  , \u1_R5_reg[26]/NET0131  , \u1_R5_reg[27]/NET0131  , \u1_R5_reg[28]/NET0131  , \u1_R5_reg[29]/NET0131  , \u1_R5_reg[2]/NET0131  , \u1_R5_reg[30]/NET0131  , \u1_R5_reg[31]/P0001  , \u1_R5_reg[32]/NET0131  , \u1_R5_reg[3]/NET0131  , \u1_R5_reg[4]/NET0131  , \u1_R5_reg[5]/NET0131  , \u1_R5_reg[6]/NET0131  , \u1_R5_reg[7]/NET0131  , \u1_R5_reg[8]/NET0131  , \u1_R5_reg[9]/NET0131  , \u1_R6_reg[10]/NET0131  , \u1_R6_reg[11]/NET0131  , \u1_R6_reg[12]/NET0131  , \u1_R6_reg[13]/NET0131  , \u1_R6_reg[14]/NET0131  , \u1_R6_reg[15]/NET0131  , \u1_R6_reg[16]/NET0131  , \u1_R6_reg[17]/NET0131  , \u1_R6_reg[18]/NET0131  , \u1_R6_reg[19]/NET0131  , \u1_R6_reg[1]/NET0131  , \u1_R6_reg[20]/NET0131  , \u1_R6_reg[21]/NET0131  , \u1_R6_reg[22]/NET0131  , \u1_R6_reg[23]/NET0131  , \u1_R6_reg[24]/NET0131  , \u1_R6_reg[25]/NET0131  , \u1_R6_reg[26]/NET0131  , \u1_R6_reg[27]/NET0131  , \u1_R6_reg[28]/NET0131  , \u1_R6_reg[29]/NET0131  , \u1_R6_reg[2]/NET0131  , \u1_R6_reg[30]/NET0131  , \u1_R6_reg[31]/P0001  , \u1_R6_reg[32]/NET0131  , \u1_R6_reg[3]/NET0131  , \u1_R6_reg[4]/NET0131  , \u1_R6_reg[5]/NET0131  , \u1_R6_reg[6]/NET0131  , \u1_R6_reg[7]/NET0131  , \u1_R6_reg[8]/NET0131  , \u1_R6_reg[9]/NET0131  , \u1_R7_reg[10]/NET0131  , \u1_R7_reg[11]/NET0131  , \u1_R7_reg[12]/NET0131  , \u1_R7_reg[13]/NET0131  , \u1_R7_reg[14]/NET0131  , \u1_R7_reg[15]/NET0131  , \u1_R7_reg[16]/NET0131  , \u1_R7_reg[17]/NET0131  , \u1_R7_reg[18]/NET0131  , \u1_R7_reg[19]/NET0131  , \u1_R7_reg[1]/NET0131  , \u1_R7_reg[20]/NET0131  , \u1_R7_reg[21]/NET0131  , \u1_R7_reg[22]/NET0131  , \u1_R7_reg[23]/NET0131  , \u1_R7_reg[24]/NET0131  , \u1_R7_reg[25]/NET0131  , \u1_R7_reg[26]/NET0131  , \u1_R7_reg[27]/NET0131  , \u1_R7_reg[28]/NET0131  , \u1_R7_reg[29]/NET0131  , \u1_R7_reg[2]/NET0131  , \u1_R7_reg[30]/NET0131  , \u1_R7_reg[31]/P0001  , \u1_R7_reg[32]/NET0131  , \u1_R7_reg[3]/NET0131  , \u1_R7_reg[4]/NET0131  , \u1_R7_reg[5]/NET0131  , \u1_R7_reg[6]/NET0131  , \u1_R7_reg[7]/NET0131  , \u1_R7_reg[8]/NET0131  , \u1_R7_reg[9]/NET0131  , \u1_R8_reg[10]/NET0131  , \u1_R8_reg[11]/NET0131  , \u1_R8_reg[12]/NET0131  , \u1_R8_reg[13]/NET0131  , \u1_R8_reg[14]/NET0131  , \u1_R8_reg[15]/NET0131  , \u1_R8_reg[16]/NET0131  , \u1_R8_reg[17]/NET0131  , \u1_R8_reg[18]/NET0131  , \u1_R8_reg[19]/NET0131  , \u1_R8_reg[1]/NET0131  , \u1_R8_reg[20]/NET0131  , \u1_R8_reg[21]/NET0131  , \u1_R8_reg[22]/NET0131  , \u1_R8_reg[23]/NET0131  , \u1_R8_reg[24]/NET0131  , \u1_R8_reg[25]/NET0131  , \u1_R8_reg[26]/NET0131  , \u1_R8_reg[27]/NET0131  , \u1_R8_reg[28]/NET0131  , \u1_R8_reg[29]/NET0131  , \u1_R8_reg[2]/NET0131  , \u1_R8_reg[30]/NET0131  , \u1_R8_reg[31]/P0001  , \u1_R8_reg[32]/NET0131  , \u1_R8_reg[3]/NET0131  , \u1_R8_reg[4]/NET0131  , \u1_R8_reg[5]/NET0131  , \u1_R8_reg[6]/NET0131  , \u1_R8_reg[7]/NET0131  , \u1_R8_reg[8]/NET0131  , \u1_R8_reg[9]/NET0131  , \u1_R9_reg[10]/NET0131  , \u1_R9_reg[11]/NET0131  , \u1_R9_reg[12]/NET0131  , \u1_R9_reg[13]/NET0131  , \u1_R9_reg[14]/NET0131  , \u1_R9_reg[15]/NET0131  , \u1_R9_reg[16]/NET0131  , \u1_R9_reg[17]/NET0131  , \u1_R9_reg[18]/NET0131  , \u1_R9_reg[19]/NET0131  , \u1_R9_reg[1]/NET0131  , \u1_R9_reg[20]/NET0131  , \u1_R9_reg[21]/NET0131  , \u1_R9_reg[22]/NET0131  , \u1_R9_reg[23]/NET0131  , \u1_R9_reg[24]/NET0131  , \u1_R9_reg[25]/NET0131  , \u1_R9_reg[26]/NET0131  , \u1_R9_reg[27]/NET0131  , \u1_R9_reg[28]/NET0131  , \u1_R9_reg[29]/NET0131  , \u1_R9_reg[2]/NET0131  , \u1_R9_reg[30]/NET0131  , \u1_R9_reg[31]/NET0131  , \u1_R9_reg[32]/NET0131  , \u1_R9_reg[3]/NET0131  , \u1_R9_reg[4]/NET0131  , \u1_R9_reg[5]/NET0131  , \u1_R9_reg[6]/NET0131  , \u1_R9_reg[7]/NET0131  , \u1_R9_reg[8]/NET0131  , \u1_R9_reg[9]/NET0131  , \u1_desIn_r_reg[0]/NET0131  , \u1_desIn_r_reg[10]/NET0131  , \u1_desIn_r_reg[11]/NET0131  , \u1_desIn_r_reg[12]/NET0131  , \u1_desIn_r_reg[13]/NET0131  , \u1_desIn_r_reg[14]/NET0131  , \u1_desIn_r_reg[15]/NET0131  , \u1_desIn_r_reg[16]/NET0131  , \u1_desIn_r_reg[17]/NET0131  , \u1_desIn_r_reg[18]/P0001  , \u1_desIn_r_reg[19]/NET0131  , \u1_desIn_r_reg[1]/NET0131  , \u1_desIn_r_reg[20]/NET0131  , \u1_desIn_r_reg[21]/NET0131  , \u1_desIn_r_reg[22]/NET0131  , \u1_desIn_r_reg[23]/NET0131  , \u1_desIn_r_reg[24]/NET0131  , \u1_desIn_r_reg[25]/NET0131  , \u1_desIn_r_reg[26]/NET0131  , \u1_desIn_r_reg[27]/NET0131  , \u1_desIn_r_reg[28]/NET0131  , \u1_desIn_r_reg[29]/NET0131  , \u1_desIn_r_reg[2]/NET0131  , \u1_desIn_r_reg[30]/NET0131  , \u1_desIn_r_reg[31]/NET0131  , \u1_desIn_r_reg[32]/NET0131  , \u1_desIn_r_reg[33]/NET0131  , \u1_desIn_r_reg[34]/NET0131  , \u1_desIn_r_reg[35]/NET0131  , \u1_desIn_r_reg[36]/NET0131  , \u1_desIn_r_reg[37]/NET0131  , \u1_desIn_r_reg[38]/NET0131  , \u1_desIn_r_reg[39]/NET0131  , \u1_desIn_r_reg[3]/NET0131  , \u1_desIn_r_reg[40]/NET0131  , \u1_desIn_r_reg[41]/NET0131  , \u1_desIn_r_reg[42]/NET0131  , \u1_desIn_r_reg[43]/NET0131  , \u1_desIn_r_reg[44]/NET0131  , \u1_desIn_r_reg[45]/NET0131  , \u1_desIn_r_reg[46]/NET0131  , \u1_desIn_r_reg[47]/NET0131  , \u1_desIn_r_reg[48]/NET0131  , \u1_desIn_r_reg[49]/NET0131  , \u1_desIn_r_reg[4]/NET0131  , \u1_desIn_r_reg[50]/NET0131  , \u1_desIn_r_reg[51]/NET0131  , \u1_desIn_r_reg[52]/P0001  , \u1_desIn_r_reg[53]/NET0131  , \u1_desIn_r_reg[54]/NET0131  , \u1_desIn_r_reg[55]/NET0131  , \u1_desIn_r_reg[56]/NET0131  , \u1_desIn_r_reg[57]/NET0131  , \u1_desIn_r_reg[58]/NET0131  , \u1_desIn_r_reg[59]/NET0131  , \u1_desIn_r_reg[5]/NET0131  , \u1_desIn_r_reg[60]/NET0131  , \u1_desIn_r_reg[61]/NET0131  , \u1_desIn_r_reg[62]/NET0131  , \u1_desIn_r_reg[63]/NET0131  , \u1_desIn_r_reg[6]/NET0131  , \u1_desIn_r_reg[7]/NET0131  , \u1_desIn_r_reg[8]/NET0131  , \u1_desIn_r_reg[9]/NET0131  , \u1_key_r_reg[0]/NET0131  , \u1_key_r_reg[10]/NET0131  , \u1_key_r_reg[11]/NET0131  , \u1_key_r_reg[12]/NET0131  , \u1_key_r_reg[13]/NET0131  , \u1_key_r_reg[14]/NET0131  , \u1_key_r_reg[15]/NET0131  , \u1_key_r_reg[16]/NET0131  , \u1_key_r_reg[17]/NET0131  , \u1_key_r_reg[18]/NET0131  , \u1_key_r_reg[19]/NET0131  , \u1_key_r_reg[1]/NET0131  , \u1_key_r_reg[20]/NET0131  , \u1_key_r_reg[21]/NET0131  , \u1_key_r_reg[22]/NET0131  , \u1_key_r_reg[23]/NET0131  , \u1_key_r_reg[24]/NET0131  , \u1_key_r_reg[25]/NET0131  , \u1_key_r_reg[26]/NET0131  , \u1_key_r_reg[27]/NET0131  , \u1_key_r_reg[28]/NET0131  , \u1_key_r_reg[29]/NET0131  , \u1_key_r_reg[2]/NET0131  , \u1_key_r_reg[30]/NET0131  , \u1_key_r_reg[31]/NET0131  , \u1_key_r_reg[32]/NET0131  , \u1_key_r_reg[33]/NET0131  , \u1_key_r_reg[34]/NET0131  , \u1_key_r_reg[35]/P0001  , \u1_key_r_reg[36]/NET0131  , \u1_key_r_reg[37]/NET0131  , \u1_key_r_reg[38]/NET0131  , \u1_key_r_reg[39]/P0001  , \u1_key_r_reg[3]/NET0131  , \u1_key_r_reg[40]/NET0131  , \u1_key_r_reg[41]/NET0131  , \u1_key_r_reg[42]/P0001  , \u1_key_r_reg[43]/NET0131  , \u1_key_r_reg[44]/NET0131  , \u1_key_r_reg[45]/NET0131  , \u1_key_r_reg[46]/NET0131  , \u1_key_r_reg[47]/NET0131  , \u1_key_r_reg[48]/NET0131  , \u1_key_r_reg[49]/NET0131  , \u1_key_r_reg[4]/NET0131  , \u1_key_r_reg[50]/NET0131  , \u1_key_r_reg[51]/NET0131  , \u1_key_r_reg[52]/NET0131  , \u1_key_r_reg[53]/NET0131  , \u1_key_r_reg[54]/NET0131  , \u1_key_r_reg[55]/NET0131  , \u1_key_r_reg[5]/NET0131  , \u1_key_r_reg[6]/NET0131  , \u1_key_r_reg[7]/NET0131  , \u1_key_r_reg[8]/NET0131  , \u1_key_r_reg[9]/NET0131  , \u1_uk_K_r0_reg[0]/NET0131  , \u1_uk_K_r0_reg[10]/NET0131  , \u1_uk_K_r0_reg[11]/NET0131  , \u1_uk_K_r0_reg[12]/NET0131  , \u1_uk_K_r0_reg[13]/NET0131  , \u1_uk_K_r0_reg[14]/NET0131  , \u1_uk_K_r0_reg[15]/NET0131  , \u1_uk_K_r0_reg[16]/NET0131  , \u1_uk_K_r0_reg[17]/NET0131  , \u1_uk_K_r0_reg[18]/NET0131  , \u1_uk_K_r0_reg[19]/NET0131  , \u1_uk_K_r0_reg[20]/NET0131  , \u1_uk_K_r0_reg[21]/NET0131  , \u1_uk_K_r0_reg[22]/NET0131  , \u1_uk_K_r0_reg[23]/NET0131  , \u1_uk_K_r0_reg[24]/NET0131  , \u1_uk_K_r0_reg[25]/P0001  , \u1_uk_K_r0_reg[26]/NET0131  , \u1_uk_K_r0_reg[27]/NET0131  , \u1_uk_K_r0_reg[28]/NET0131  , \u1_uk_K_r0_reg[29]/NET0131  , \u1_uk_K_r0_reg[2]/NET0131  , \u1_uk_K_r0_reg[30]/NET0131  , \u1_uk_K_r0_reg[31]/NET0131  , \u1_uk_K_r0_reg[32]/NET0131  , \u1_uk_K_r0_reg[33]/NET0131  , \u1_uk_K_r0_reg[34]/NET0131  , \u1_uk_K_r0_reg[35]/NET0131  , \u1_uk_K_r0_reg[36]/NET0131  , \u1_uk_K_r0_reg[37]/NET0131  , \u1_uk_K_r0_reg[38]/NET0131  , \u1_uk_K_r0_reg[39]/NET0131  , \u1_uk_K_r0_reg[3]/NET0131  , \u1_uk_K_r0_reg[40]/NET0131  , \u1_uk_K_r0_reg[41]/NET0131  , \u1_uk_K_r0_reg[42]/NET0131  , \u1_uk_K_r0_reg[43]/NET0131  , \u1_uk_K_r0_reg[44]/NET0131  , \u1_uk_K_r0_reg[45]/NET0131  , \u1_uk_K_r0_reg[46]/NET0131  , \u1_uk_K_r0_reg[47]/NET0131  , \u1_uk_K_r0_reg[48]/NET0131  , \u1_uk_K_r0_reg[49]/NET0131  , \u1_uk_K_r0_reg[4]/NET0131  , \u1_uk_K_r0_reg[50]/NET0131  , \u1_uk_K_r0_reg[51]/NET0131  , \u1_uk_K_r0_reg[52]/P0001  , \u1_uk_K_r0_reg[54]/NET0131  , \u1_uk_K_r0_reg[55]/NET0131  , \u1_uk_K_r0_reg[5]/NET0131  , \u1_uk_K_r0_reg[6]/NET0131  , \u1_uk_K_r0_reg[7]/NET0131  , \u1_uk_K_r0_reg[8]/NET0131  , \u1_uk_K_r0_reg[9]/NET0131  , \u1_uk_K_r10_reg[0]/NET0131  , \u1_uk_K_r10_reg[10]/NET0131  , \u1_uk_K_r10_reg[11]/NET0131  , \u1_uk_K_r10_reg[12]/NET0131  , \u1_uk_K_r10_reg[14]/NET0131  , \u1_uk_K_r10_reg[15]/NET0131  , \u1_uk_K_r10_reg[16]/NET0131  , \u1_uk_K_r10_reg[17]/NET0131  , \u1_uk_K_r10_reg[18]/NET0131  , \u1_uk_K_r10_reg[19]/NET0131  , \u1_uk_K_r10_reg[1]/NET0131  , \u1_uk_K_r10_reg[20]/NET0131  , \u1_uk_K_r10_reg[21]/NET0131  , \u1_uk_K_r10_reg[22]/NET0131  , \u1_uk_K_r10_reg[23]/NET0131  , \u1_uk_K_r10_reg[24]/NET0131  , \u1_uk_K_r10_reg[25]/NET0131  , \u1_uk_K_r10_reg[26]/NET0131  , \u1_uk_K_r10_reg[27]/NET0131  , \u1_uk_K_r10_reg[28]/NET0131  , \u1_uk_K_r10_reg[29]/NET0131  , \u1_uk_K_r10_reg[2]/NET0131  , \u1_uk_K_r10_reg[30]/NET0131  , \u1_uk_K_r10_reg[31]/NET0131  , \u1_uk_K_r10_reg[32]/NET0131  , \u1_uk_K_r10_reg[33]/NET0131  , \u1_uk_K_r10_reg[34]/NET0131  , \u1_uk_K_r10_reg[35]/NET0131  , \u1_uk_K_r10_reg[36]/NET0131  , \u1_uk_K_r10_reg[37]/NET0131  , \u1_uk_K_r10_reg[38]/NET0131  , \u1_uk_K_r10_reg[39]/NET0131  , \u1_uk_K_r10_reg[3]/NET0131  , \u1_uk_K_r10_reg[40]/NET0131  , \u1_uk_K_r10_reg[41]/P0001  , \u1_uk_K_r10_reg[42]/NET0131  , \u1_uk_K_r10_reg[43]/NET0131  , \u1_uk_K_r10_reg[44]/NET0131  , \u1_uk_K_r10_reg[45]/P0001  , \u1_uk_K_r10_reg[46]/NET0131  , \u1_uk_K_r10_reg[47]/NET0131  , \u1_uk_K_r10_reg[48]/NET0131  , \u1_uk_K_r10_reg[49]/NET0131  , \u1_uk_K_r10_reg[4]/NET0131  , \u1_uk_K_r10_reg[50]/NET0131  , \u1_uk_K_r10_reg[51]/NET0131  , \u1_uk_K_r10_reg[52]/NET0131  , \u1_uk_K_r10_reg[53]/NET0131  , \u1_uk_K_r10_reg[54]/NET0131  , \u1_uk_K_r10_reg[55]/NET0131  , \u1_uk_K_r10_reg[5]/NET0131  , \u1_uk_K_r10_reg[6]/NET0131  , \u1_uk_K_r10_reg[7]/NET0131  , \u1_uk_K_r10_reg[8]/NET0131  , \u1_uk_K_r10_reg[9]/NET0131  , \u1_uk_K_r11_reg[0]/NET0131  , \u1_uk_K_r11_reg[10]/NET0131  , \u1_uk_K_r11_reg[11]/NET0131  , \u1_uk_K_r11_reg[12]/NET0131  , \u1_uk_K_r11_reg[13]/NET0131  , \u1_uk_K_r11_reg[14]/NET0131  , \u1_uk_K_r11_reg[15]/NET0131  , \u1_uk_K_r11_reg[16]/NET0131  , \u1_uk_K_r11_reg[17]/NET0131  , \u1_uk_K_r11_reg[18]/NET0131  , \u1_uk_K_r11_reg[19]/NET0131  , \u1_uk_K_r11_reg[1]/NET0131  , \u1_uk_K_r11_reg[20]/NET0131  , \u1_uk_K_r11_reg[21]/NET0131  , \u1_uk_K_r11_reg[22]/NET0131  , \u1_uk_K_r11_reg[23]/NET0131  , \u1_uk_K_r11_reg[24]/NET0131  , \u1_uk_K_r11_reg[25]/NET0131  , \u1_uk_K_r11_reg[26]/NET0131  , \u1_uk_K_r11_reg[27]/P0001  , \u1_uk_K_r11_reg[28]/NET0131  , \u1_uk_K_r11_reg[29]/NET0131  , \u1_uk_K_r11_reg[2]/NET0131  , \u1_uk_K_r11_reg[31]/NET0131  , \u1_uk_K_r11_reg[32]/NET0131  , \u1_uk_K_r11_reg[33]/NET0131  , \u1_uk_K_r11_reg[34]/NET0131  , \u1_uk_K_r11_reg[35]/NET0131  , \u1_uk_K_r11_reg[36]/NET0131  , \u1_uk_K_r11_reg[37]/NET0131  , \u1_uk_K_r11_reg[38]/NET0131  , \u1_uk_K_r11_reg[39]/NET0131  , \u1_uk_K_r11_reg[3]/NET0131  , \u1_uk_K_r11_reg[40]/NET0131  , \u1_uk_K_r11_reg[41]/NET0131  , \u1_uk_K_r11_reg[42]/NET0131  , \u1_uk_K_r11_reg[43]/NET0131  , \u1_uk_K_r11_reg[44]/NET0131  , \u1_uk_K_r11_reg[45]/NET0131  , \u1_uk_K_r11_reg[46]/NET0131  , \u1_uk_K_r11_reg[47]/NET0131  , \u1_uk_K_r11_reg[48]/NET0131  , \u1_uk_K_r11_reg[49]/NET0131  , \u1_uk_K_r11_reg[4]/NET0131  , \u1_uk_K_r11_reg[50]/NET0131  , \u1_uk_K_r11_reg[51]/NET0131  , \u1_uk_K_r11_reg[52]/NET0131  , \u1_uk_K_r11_reg[53]/P0001  , \u1_uk_K_r11_reg[54]/NET0131  , \u1_uk_K_r11_reg[55]/NET0131  , \u1_uk_K_r11_reg[5]/NET0131  , \u1_uk_K_r11_reg[6]/NET0131  , \u1_uk_K_r11_reg[7]/NET0131  , \u1_uk_K_r11_reg[8]/NET0131  , \u1_uk_K_r11_reg[9]/NET0131  , \u1_uk_K_r12_reg[0]/NET0131  , \u1_uk_K_r12_reg[10]/P0001  , \u1_uk_K_r12_reg[11]/NET0131  , \u1_uk_K_r12_reg[12]/NET0131  , \u1_uk_K_r12_reg[13]/NET0131  , \u1_uk_K_r12_reg[14]/NET0131  , \u1_uk_K_r12_reg[15]/NET0131  , \u1_uk_K_r12_reg[16]/NET0131  , \u1_uk_K_r12_reg[17]/NET0131  , \u1_uk_K_r12_reg[18]/NET0131  , \u1_uk_K_r12_reg[19]/NET0131  , \u1_uk_K_r12_reg[1]/NET0131  , \u1_uk_K_r12_reg[20]/NET0131  , \u1_uk_K_r12_reg[21]/NET0131  , \u1_uk_K_r12_reg[22]/NET0131  , \u1_uk_K_r12_reg[23]/NET0131  , \u1_uk_K_r12_reg[24]/NET0131  , \u1_uk_K_r12_reg[25]/NET0131  , \u1_uk_K_r12_reg[26]/NET0131  , \u1_uk_K_r12_reg[27]/NET0131  , \u1_uk_K_r12_reg[28]/NET0131  , \u1_uk_K_r12_reg[29]/NET0131  , \u1_uk_K_r12_reg[2]/NET0131  , \u1_uk_K_r12_reg[30]/NET0131  , \u1_uk_K_r12_reg[31]/NET0131  , \u1_uk_K_r12_reg[32]/NET0131  , \u1_uk_K_r12_reg[33]/NET0131  , \u1_uk_K_r12_reg[34]/NET0131  , \u1_uk_K_r12_reg[35]/NET0131  , \u1_uk_K_r12_reg[36]/NET0131  , \u1_uk_K_r12_reg[37]/NET0131  , \u1_uk_K_r12_reg[38]/NET0131  , \u1_uk_K_r12_reg[3]/NET0131  , \u1_uk_K_r12_reg[40]/NET0131  , \u1_uk_K_r12_reg[41]/NET0131  , \u1_uk_K_r12_reg[42]/NET0131  , \u1_uk_K_r12_reg[43]/NET0131  , \u1_uk_K_r12_reg[44]/P0001  , \u1_uk_K_r12_reg[45]/NET0131  , \u1_uk_K_r12_reg[46]/NET0131  , \u1_uk_K_r12_reg[47]/NET0131  , \u1_uk_K_r12_reg[48]/NET0131  , \u1_uk_K_r12_reg[49]/NET0131  , \u1_uk_K_r12_reg[4]/NET0131  , \u1_uk_K_r12_reg[50]/NET0131  , \u1_uk_K_r12_reg[51]/NET0131  , \u1_uk_K_r12_reg[52]/NET0131  , \u1_uk_K_r12_reg[53]/NET0131  , \u1_uk_K_r12_reg[54]/NET0131  , \u1_uk_K_r12_reg[55]/NET0131  , \u1_uk_K_r12_reg[5]/NET0131  , \u1_uk_K_r12_reg[6]/NET0131  , \u1_uk_K_r12_reg[7]/P0001  , \u1_uk_K_r12_reg[8]/NET0131  , \u1_uk_K_r12_reg[9]/NET0131  , \u1_uk_K_r13_reg[0]/NET0131  , \u1_uk_K_r13_reg[10]/NET0131  , \u1_uk_K_r13_reg[11]/NET0131  , \u1_uk_K_r13_reg[12]/NET0131  , \u1_uk_K_r13_reg[13]/NET0131  , \u1_uk_K_r13_reg[14]/NET0131  , \u1_uk_K_r13_reg[15]/NET0131  , \u1_uk_K_r13_reg[16]/NET0131  , \u1_uk_K_r13_reg[17]/NET0131  , \u1_uk_K_r13_reg[18]/NET0131  , \u1_uk_K_r13_reg[19]/NET0131  , \u1_uk_K_r13_reg[20]/NET0131  , \u1_uk_K_r13_reg[21]/NET0131  , \u1_uk_K_r13_reg[22]/NET0131  , \u1_uk_K_r13_reg[23]/NET0131  , \u1_uk_K_r13_reg[24]/NET0131  , \u1_uk_K_r13_reg[25]/P0001  , \u1_uk_K_r13_reg[26]/NET0131  , \u1_uk_K_r13_reg[27]/NET0131  , \u1_uk_K_r13_reg[28]/NET0131  , \u1_uk_K_r13_reg[29]/NET0131  , \u1_uk_K_r13_reg[2]/NET0131  , \u1_uk_K_r13_reg[30]/NET0131  , \u1_uk_K_r13_reg[31]/NET0131  , \u1_uk_K_r13_reg[32]/NET0131  , \u1_uk_K_r13_reg[33]/NET0131  , \u1_uk_K_r13_reg[34]/NET0131  , \u1_uk_K_r13_reg[35]/NET0131  , \u1_uk_K_r13_reg[36]/NET0131  , \u1_uk_K_r13_reg[37]/NET0131  , \u1_uk_K_r13_reg[38]/NET0131  , \u1_uk_K_r13_reg[39]/NET0131  , \u1_uk_K_r13_reg[3]/NET0131  , \u1_uk_K_r13_reg[40]/NET0131  , \u1_uk_K_r13_reg[41]/NET0131  , \u1_uk_K_r13_reg[42]/NET0131  , \u1_uk_K_r13_reg[43]/NET0131  , \u1_uk_K_r13_reg[44]/NET0131  , \u1_uk_K_r13_reg[45]/NET0131  , \u1_uk_K_r13_reg[46]/NET0131  , \u1_uk_K_r13_reg[47]/NET0131  , \u1_uk_K_r13_reg[48]/NET0131  , \u1_uk_K_r13_reg[49]/NET0131  , \u1_uk_K_r13_reg[4]/NET0131  , \u1_uk_K_r13_reg[50]/NET0131  , \u1_uk_K_r13_reg[51]/NET0131  , \u1_uk_K_r13_reg[52]/P0001  , \u1_uk_K_r13_reg[54]/NET0131  , \u1_uk_K_r13_reg[55]/NET0131  , \u1_uk_K_r13_reg[5]/NET0131  , \u1_uk_K_r13_reg[6]/NET0131  , \u1_uk_K_r13_reg[7]/NET0131  , \u1_uk_K_r13_reg[8]/NET0131  , \u1_uk_K_r13_reg[9]/NET0131  , \u1_uk_K_r14_reg[0]/P0001  , \u1_uk_K_r14_reg[10]/P0001  , \u1_uk_K_r14_reg[11]/NET0131  , \u1_uk_K_r14_reg[12]/NET0131  , \u1_uk_K_r14_reg[13]/NET0131  , \u1_uk_K_r14_reg[14]/NET0131  , \u1_uk_K_r14_reg[15]/NET0131  , \u1_uk_K_r14_reg[16]/NET0131  , \u1_uk_K_r14_reg[17]/NET0131  , \u1_uk_K_r14_reg[18]/NET0131  , \u1_uk_K_r14_reg[19]/NET0131  , \u1_uk_K_r14_reg[1]/NET0131  , \u1_uk_K_r14_reg[20]/NET0131  , \u1_uk_K_r14_reg[21]/NET0131  , \u1_uk_K_r14_reg[22]/NET0131  , \u1_uk_K_r14_reg[23]/NET0131  , \u1_uk_K_r14_reg[24]/NET0131  , \u1_uk_K_r14_reg[25]/NET0131  , \u1_uk_K_r14_reg[26]/NET0131  , \u1_uk_K_r14_reg[27]/NET0131  , \u1_uk_K_r14_reg[28]/NET0131  , \u1_uk_K_r14_reg[29]/NET0131  , \u1_uk_K_r14_reg[2]/NET0131  , \u1_uk_K_r14_reg[30]/NET0131  , \u1_uk_K_r14_reg[31]/NET0131  , \u1_uk_K_r14_reg[32]/NET0131  , \u1_uk_K_r14_reg[33]/NET0131  , \u1_uk_K_r14_reg[34]/NET0131  , \u1_uk_K_r14_reg[35]/P0001  , \u1_uk_K_r14_reg[36]/NET0131  , \u1_uk_K_r14_reg[37]/NET0131  , \u1_uk_K_r14_reg[38]/NET0131  , \u1_uk_K_r14_reg[39]/P0001  , \u1_uk_K_r14_reg[3]/NET0131  , \u1_uk_K_r14_reg[40]/NET0131  , \u1_uk_K_r14_reg[41]/NET0131  , \u1_uk_K_r14_reg[42]/P0001  , \u1_uk_K_r14_reg[43]/NET0131  , \u1_uk_K_r14_reg[44]/NET0131  , \u1_uk_K_r14_reg[45]/NET0131  , \u1_uk_K_r14_reg[46]/NET0131  , \u1_uk_K_r14_reg[47]/NET0131  , \u1_uk_K_r14_reg[48]/NET0131  , \u1_uk_K_r14_reg[49]/NET0131  , \u1_uk_K_r14_reg[4]/NET0131  , \u1_uk_K_r14_reg[50]/NET0131  , \u1_uk_K_r14_reg[51]/NET0131  , \u1_uk_K_r14_reg[52]/NET0131  , \u1_uk_K_r14_reg[53]/NET0131  , \u1_uk_K_r14_reg[54]/NET0131  , \u1_uk_K_r14_reg[55]/NET0131  , \u1_uk_K_r14_reg[5]/NET0131  , \u1_uk_K_r14_reg[6]/NET0131  , \u1_uk_K_r14_reg[7]/NET0131  , \u1_uk_K_r14_reg[8]/P0001  , \u1_uk_K_r14_reg[9]/NET0131  , \u1_uk_K_r1_reg[0]/NET0131  , \u1_uk_K_r1_reg[10]/P0001  , \u1_uk_K_r1_reg[11]/NET0131  , \u1_uk_K_r1_reg[12]/NET0131  , \u1_uk_K_r1_reg[13]/NET0131  , \u1_uk_K_r1_reg[14]/NET0131  , \u1_uk_K_r1_reg[15]/NET0131  , \u1_uk_K_r1_reg[16]/NET0131  , \u1_uk_K_r1_reg[17]/NET0131  , \u1_uk_K_r1_reg[18]/NET0131  , \u1_uk_K_r1_reg[19]/NET0131  , \u1_uk_K_r1_reg[1]/NET0131  , \u1_uk_K_r1_reg[20]/NET0131  , \u1_uk_K_r1_reg[21]/NET0131  , \u1_uk_K_r1_reg[22]/NET0131  , \u1_uk_K_r1_reg[23]/NET0131  , \u1_uk_K_r1_reg[24]/NET0131  , \u1_uk_K_r1_reg[25]/NET0131  , \u1_uk_K_r1_reg[26]/NET0131  , \u1_uk_K_r1_reg[27]/NET0131  , \u1_uk_K_r1_reg[28]/NET0131  , \u1_uk_K_r1_reg[29]/NET0131  , \u1_uk_K_r1_reg[2]/NET0131  , \u1_uk_K_r1_reg[30]/NET0131  , \u1_uk_K_r1_reg[31]/NET0131  , \u1_uk_K_r1_reg[32]/NET0131  , \u1_uk_K_r1_reg[33]/NET0131  , \u1_uk_K_r1_reg[34]/NET0131  , \u1_uk_K_r1_reg[35]/NET0131  , \u1_uk_K_r1_reg[36]/NET0131  , \u1_uk_K_r1_reg[37]/NET0131  , \u1_uk_K_r1_reg[38]/NET0131  , \u1_uk_K_r1_reg[3]/NET0131  , \u1_uk_K_r1_reg[40]/NET0131  , \u1_uk_K_r1_reg[41]/NET0131  , \u1_uk_K_r1_reg[42]/NET0131  , \u1_uk_K_r1_reg[43]/NET0131  , \u1_uk_K_r1_reg[44]/P0001  , \u1_uk_K_r1_reg[45]/NET0131  , \u1_uk_K_r1_reg[46]/NET0131  , \u1_uk_K_r1_reg[47]/NET0131  , \u1_uk_K_r1_reg[48]/NET0131  , \u1_uk_K_r1_reg[49]/NET0131  , \u1_uk_K_r1_reg[4]/NET0131  , \u1_uk_K_r1_reg[50]/NET0131  , \u1_uk_K_r1_reg[51]/NET0131  , \u1_uk_K_r1_reg[52]/NET0131  , \u1_uk_K_r1_reg[53]/NET0131  , \u1_uk_K_r1_reg[54]/NET0131  , \u1_uk_K_r1_reg[55]/NET0131  , \u1_uk_K_r1_reg[5]/NET0131  , \u1_uk_K_r1_reg[6]/NET0131  , \u1_uk_K_r1_reg[7]/P0001  , \u1_uk_K_r1_reg[8]/NET0131  , \u1_uk_K_r1_reg[9]/NET0131  , \u1_uk_K_r2_reg[0]/NET0131  , \u1_uk_K_r2_reg[10]/NET0131  , \u1_uk_K_r2_reg[11]/NET0131  , \u1_uk_K_r2_reg[12]/NET0131  , \u1_uk_K_r2_reg[13]/NET0131  , \u1_uk_K_r2_reg[14]/NET0131  , \u1_uk_K_r2_reg[15]/NET0131  , \u1_uk_K_r2_reg[16]/NET0131  , \u1_uk_K_r2_reg[17]/NET0131  , \u1_uk_K_r2_reg[18]/NET0131  , \u1_uk_K_r2_reg[19]/NET0131  , \u1_uk_K_r2_reg[1]/NET0131  , \u1_uk_K_r2_reg[20]/NET0131  , \u1_uk_K_r2_reg[21]/NET0131  , \u1_uk_K_r2_reg[22]/NET0131  , \u1_uk_K_r2_reg[23]/NET0131  , \u1_uk_K_r2_reg[24]/NET0131  , \u1_uk_K_r2_reg[25]/NET0131  , \u1_uk_K_r2_reg[26]/NET0131  , \u1_uk_K_r2_reg[27]/NET0131  , \u1_uk_K_r2_reg[28]/NET0131  , \u1_uk_K_r2_reg[29]/NET0131  , \u1_uk_K_r2_reg[2]/NET0131  , \u1_uk_K_r2_reg[31]/NET0131  , \u1_uk_K_r2_reg[32]/NET0131  , \u1_uk_K_r2_reg[33]/NET0131  , \u1_uk_K_r2_reg[34]/NET0131  , \u1_uk_K_r2_reg[35]/NET0131  , \u1_uk_K_r2_reg[36]/NET0131  , \u1_uk_K_r2_reg[37]/NET0131  , \u1_uk_K_r2_reg[38]/NET0131  , \u1_uk_K_r2_reg[39]/NET0131  , \u1_uk_K_r2_reg[3]/NET0131  , \u1_uk_K_r2_reg[40]/NET0131  , \u1_uk_K_r2_reg[41]/NET0131  , \u1_uk_K_r2_reg[42]/NET0131  , \u1_uk_K_r2_reg[43]/NET0131  , \u1_uk_K_r2_reg[44]/NET0131  , \u1_uk_K_r2_reg[45]/NET0131  , \u1_uk_K_r2_reg[46]/NET0131  , \u1_uk_K_r2_reg[47]/NET0131  , \u1_uk_K_r2_reg[48]/NET0131  , \u1_uk_K_r2_reg[49]/NET0131  , \u1_uk_K_r2_reg[4]/NET0131  , \u1_uk_K_r2_reg[50]/NET0131  , \u1_uk_K_r2_reg[51]/NET0131  , \u1_uk_K_r2_reg[52]/NET0131  , \u1_uk_K_r2_reg[53]/P0001  , \u1_uk_K_r2_reg[54]/NET0131  , \u1_uk_K_r2_reg[55]/NET0131  , \u1_uk_K_r2_reg[5]/NET0131  , \u1_uk_K_r2_reg[6]/NET0131  , \u1_uk_K_r2_reg[7]/NET0131  , \u1_uk_K_r2_reg[8]/NET0131  , \u1_uk_K_r2_reg[9]/NET0131  , \u1_uk_K_r3_reg[0]/NET0131  , \u1_uk_K_r3_reg[10]/NET0131  , \u1_uk_K_r3_reg[11]/NET0131  , \u1_uk_K_r3_reg[12]/NET0131  , \u1_uk_K_r3_reg[14]/NET0131  , \u1_uk_K_r3_reg[15]/NET0131  , \u1_uk_K_r3_reg[16]/NET0131  , \u1_uk_K_r3_reg[17]/NET0131  , \u1_uk_K_r3_reg[18]/NET0131  , \u1_uk_K_r3_reg[19]/NET0131  , \u1_uk_K_r3_reg[1]/NET0131  , \u1_uk_K_r3_reg[20]/NET0131  , \u1_uk_K_r3_reg[21]/NET0131  , \u1_uk_K_r3_reg[22]/NET0131  , \u1_uk_K_r3_reg[23]/NET0131  , \u1_uk_K_r3_reg[24]/NET0131  , \u1_uk_K_r3_reg[25]/NET0131  , \u1_uk_K_r3_reg[26]/NET0131  , \u1_uk_K_r3_reg[27]/NET0131  , \u1_uk_K_r3_reg[28]/NET0131  , \u1_uk_K_r3_reg[29]/NET0131  , \u1_uk_K_r3_reg[2]/NET0131  , \u1_uk_K_r3_reg[30]/NET0131  , \u1_uk_K_r3_reg[31]/NET0131  , \u1_uk_K_r3_reg[32]/NET0131  , \u1_uk_K_r3_reg[33]/NET0131  , \u1_uk_K_r3_reg[34]/NET0131  , \u1_uk_K_r3_reg[35]/NET0131  , \u1_uk_K_r3_reg[36]/NET0131  , \u1_uk_K_r3_reg[37]/NET0131  , \u1_uk_K_r3_reg[38]/NET0131  , \u1_uk_K_r3_reg[39]/NET0131  , \u1_uk_K_r3_reg[3]/NET0131  , \u1_uk_K_r3_reg[40]/NET0131  , \u1_uk_K_r3_reg[41]/NET0131  , \u1_uk_K_r3_reg[42]/NET0131  , \u1_uk_K_r3_reg[43]/NET0131  , \u1_uk_K_r3_reg[44]/NET0131  , \u1_uk_K_r3_reg[45]/NET0131  , \u1_uk_K_r3_reg[46]/NET0131  , \u1_uk_K_r3_reg[47]/NET0131  , \u1_uk_K_r3_reg[48]/NET0131  , \u1_uk_K_r3_reg[49]/NET0131  , \u1_uk_K_r3_reg[4]/NET0131  , \u1_uk_K_r3_reg[50]/NET0131  , \u1_uk_K_r3_reg[51]/NET0131  , \u1_uk_K_r3_reg[52]/NET0131  , \u1_uk_K_r3_reg[53]/NET0131  , \u1_uk_K_r3_reg[54]/NET0131  , \u1_uk_K_r3_reg[55]/NET0131  , \u1_uk_K_r3_reg[5]/NET0131  , \u1_uk_K_r3_reg[6]/NET0131  , \u1_uk_K_r3_reg[7]/NET0131  , \u1_uk_K_r3_reg[8]/NET0131  , \u1_uk_K_r3_reg[9]/NET0131  , \u1_uk_K_r4_reg[0]/P0001  , \u1_uk_K_r4_reg[10]/NET0131  , \u1_uk_K_r4_reg[11]/NET0131  , \u1_uk_K_r4_reg[12]/NET0131  , \u1_uk_K_r4_reg[13]/NET0131  , \u1_uk_K_r4_reg[14]/NET0131  , \u1_uk_K_r4_reg[15]/NET0131  , \u1_uk_K_r4_reg[16]/NET0131  , \u1_uk_K_r4_reg[17]/NET0131  , \u1_uk_K_r4_reg[18]/NET0131  , \u1_uk_K_r4_reg[19]/NET0131  , \u1_uk_K_r4_reg[1]/NET0131  , \u1_uk_K_r4_reg[20]/NET0131  , \u1_uk_K_r4_reg[21]/NET0131  , \u1_uk_K_r4_reg[22]/NET0131  , \u1_uk_K_r4_reg[23]/P0001  , \u1_uk_K_r4_reg[25]/NET0131  , \u1_uk_K_r4_reg[26]/NET0131  , \u1_uk_K_r4_reg[27]/P0001  , \u1_uk_K_r4_reg[28]/NET0131  , \u1_uk_K_r4_reg[29]/NET0131  , \u1_uk_K_r4_reg[30]/NET0131  , \u1_uk_K_r4_reg[31]/P0001  , \u1_uk_K_r4_reg[32]/NET0131  , \u1_uk_K_r4_reg[33]/NET0131  , \u1_uk_K_r4_reg[34]/NET0131  , \u1_uk_K_r4_reg[35]/NET0131  , \u1_uk_K_r4_reg[36]/NET0131  , \u1_uk_K_r4_reg[37]/NET0131  , \u1_uk_K_r4_reg[38]/NET0131  , \u1_uk_K_r4_reg[39]/NET0131  , \u1_uk_K_r4_reg[3]/NET0131  , \u1_uk_K_r4_reg[40]/NET0131  , \u1_uk_K_r4_reg[41]/NET0131  , \u1_uk_K_r4_reg[42]/NET0131  , \u1_uk_K_r4_reg[43]/NET0131  , \u1_uk_K_r4_reg[44]/NET0131  , \u1_uk_K_r4_reg[45]/NET0131  , \u1_uk_K_r4_reg[46]/NET0131  , \u1_uk_K_r4_reg[47]/NET0131  , \u1_uk_K_r4_reg[48]/NET0131  , \u1_uk_K_r4_reg[49]/NET0131  , \u1_uk_K_r4_reg[4]/NET0131  , \u1_uk_K_r4_reg[50]/NET0131  , \u1_uk_K_r4_reg[51]/NET0131  , \u1_uk_K_r4_reg[52]/NET0131  , \u1_uk_K_r4_reg[53]/NET0131  , \u1_uk_K_r4_reg[54]/NET0131  , \u1_uk_K_r4_reg[55]/NET0131  , \u1_uk_K_r4_reg[5]/NET0131  , \u1_uk_K_r4_reg[6]/NET0131  , \u1_uk_K_r4_reg[7]/NET0131  , \u1_uk_K_r4_reg[8]/NET0131  , \u1_uk_K_r4_reg[9]/NET0131  , \u1_uk_K_r5_reg[0]/NET0131  , \u1_uk_K_r5_reg[10]/NET0131  , \u1_uk_K_r5_reg[11]/NET0131  , \u1_uk_K_r5_reg[12]/P0001  , \u1_uk_K_r5_reg[13]/P0001  , \u1_uk_K_r5_reg[14]/NET0131  , \u1_uk_K_r5_reg[15]/NET0131  , \u1_uk_K_r5_reg[16]/NET0131  , \u1_uk_K_r5_reg[17]/NET0131  , \u1_uk_K_r5_reg[18]/NET0131  , \u1_uk_K_r5_reg[19]/NET0131  , \u1_uk_K_r5_reg[1]/NET0131  , \u1_uk_K_r5_reg[20]/NET0131  , \u1_uk_K_r5_reg[21]/NET0131  , \u1_uk_K_r5_reg[22]/NET0131  , \u1_uk_K_r5_reg[23]/NET0131  , \u1_uk_K_r5_reg[24]/NET0131  , \u1_uk_K_r5_reg[25]/NET0131  , \u1_uk_K_r5_reg[26]/NET0131  , \u1_uk_K_r5_reg[27]/NET0131  , \u1_uk_K_r5_reg[28]/NET0131  , \u1_uk_K_r5_reg[29]/NET0131  , \u1_uk_K_r5_reg[2]/NET0131  , \u1_uk_K_r5_reg[30]/NET0131  , \u1_uk_K_r5_reg[31]/NET0131  , \u1_uk_K_r5_reg[32]/NET0131  , \u1_uk_K_r5_reg[33]/NET0131  , \u1_uk_K_r5_reg[34]/NET0131  , \u1_uk_K_r5_reg[35]/NET0131  , \u1_uk_K_r5_reg[36]/NET0131  , \u1_uk_K_r5_reg[37]/P0001  , \u1_uk_K_r5_reg[38]/NET0131  , \u1_uk_K_r5_reg[39]/NET0131  , \u1_uk_K_r5_reg[3]/NET0131  , \u1_uk_K_r5_reg[40]/NET0131  , \u1_uk_K_r5_reg[41]/NET0131  , \u1_uk_K_r5_reg[42]/NET0131  , \u1_uk_K_r5_reg[43]/NET0131  , \u1_uk_K_r5_reg[44]/NET0131  , \u1_uk_K_r5_reg[46]/NET0131  , \u1_uk_K_r5_reg[47]/NET0131  , \u1_uk_K_r5_reg[48]/NET0131  , \u1_uk_K_r5_reg[49]/NET0131  , \u1_uk_K_r5_reg[4]/NET0131  , \u1_uk_K_r5_reg[50]/NET0131  , \u1_uk_K_r5_reg[51]/NET0131  , \u1_uk_K_r5_reg[52]/NET0131  , \u1_uk_K_r5_reg[53]/NET0131  , \u1_uk_K_r5_reg[54]/NET0131  , \u1_uk_K_r5_reg[55]/NET0131  , \u1_uk_K_r5_reg[5]/NET0131  , \u1_uk_K_r5_reg[6]/NET0131  , \u1_uk_K_r5_reg[7]/NET0131  , \u1_uk_K_r5_reg[8]/NET0131  , \u1_uk_K_r5_reg[9]/NET0131  , \u1_uk_K_r6_reg[0]/NET0131  , \u1_uk_K_r6_reg[10]/NET0131  , \u1_uk_K_r6_reg[11]/NET0131  , \u1_uk_K_r6_reg[12]/NET0131  , \u1_uk_K_r6_reg[13]/NET0131  , \u1_uk_K_r6_reg[14]/NET0131  , \u1_uk_K_r6_reg[15]/NET0131  , \u1_uk_K_r6_reg[16]/NET0131  , \u1_uk_K_r6_reg[17]/NET0131  , \u1_uk_K_r6_reg[18]/NET0131  , \u1_uk_K_r6_reg[19]/NET0131  , \u1_uk_K_r6_reg[1]/NET0131  , \u1_uk_K_r6_reg[20]/NET0131  , \u1_uk_K_r6_reg[21]/NET0131  , \u1_uk_K_r6_reg[22]/NET0131  , \u1_uk_K_r6_reg[23]/P0001  , \u1_uk_K_r6_reg[24]/NET0131  , \u1_uk_K_r6_reg[25]/NET0131  , \u1_uk_K_r6_reg[26]/NET0131  , \u1_uk_K_r6_reg[27]/NET0131  , \u1_uk_K_r6_reg[28]/NET0131  , \u1_uk_K_r6_reg[29]/NET0131  , \u1_uk_K_r6_reg[2]/NET0131  , \u1_uk_K_r6_reg[30]/P0001  , \u1_uk_K_r6_reg[31]/NET0131  , \u1_uk_K_r6_reg[32]/NET0131  , \u1_uk_K_r6_reg[33]/NET0131  , \u1_uk_K_r6_reg[34]/NET0131  , \u1_uk_K_r6_reg[35]/NET0131  , \u1_uk_K_r6_reg[36]/NET0131  , \u1_uk_K_r6_reg[37]/NET0131  , \u1_uk_K_r6_reg[38]/NET0131  , \u1_uk_K_r6_reg[39]/NET0131  , \u1_uk_K_r6_reg[3]/NET0131  , \u1_uk_K_r6_reg[40]/NET0131  , \u1_uk_K_r6_reg[41]/NET0131  , \u1_uk_K_r6_reg[42]/NET0131  , \u1_uk_K_r6_reg[43]/NET0131  , \u1_uk_K_r6_reg[44]/NET0131  , \u1_uk_K_r6_reg[45]/NET0131  , \u1_uk_K_r6_reg[46]/NET0131  , \u1_uk_K_r6_reg[47]/NET0131  , \u1_uk_K_r6_reg[48]/NET0131  , \u1_uk_K_r6_reg[49]/NET0131  , \u1_uk_K_r6_reg[4]/NET0131  , \u1_uk_K_r6_reg[50]/NET0131  , \u1_uk_K_r6_reg[51]/NET0131  , \u1_uk_K_r6_reg[52]/NET0131  , \u1_uk_K_r6_reg[53]/NET0131  , \u1_uk_K_r6_reg[54]/NET0131  , \u1_uk_K_r6_reg[55]/P0001  , \u1_uk_K_r6_reg[5]/NET0131  , \u1_uk_K_r6_reg[6]/NET0131  , \u1_uk_K_r6_reg[7]/NET0131  , \u1_uk_K_r6_reg[8]/NET0131  , \u1_uk_K_r6_reg[9]/NET0131  , \u1_uk_K_r7_reg[0]/NET0131  , \u1_uk_K_r7_reg[10]/NET0131  , \u1_uk_K_r7_reg[11]/NET0131  , \u1_uk_K_r7_reg[12]/NET0131  , \u1_uk_K_r7_reg[13]/NET0131  , \u1_uk_K_r7_reg[14]/NET0131  , \u1_uk_K_r7_reg[15]/NET0131  , \u1_uk_K_r7_reg[16]/NET0131  , \u1_uk_K_r7_reg[17]/NET0131  , \u1_uk_K_r7_reg[18]/NET0131  , \u1_uk_K_r7_reg[19]/NET0131  , \u1_uk_K_r7_reg[1]/NET0131  , \u1_uk_K_r7_reg[20]/NET0131  , \u1_uk_K_r7_reg[21]/NET0131  , \u1_uk_K_r7_reg[22]/NET0131  , \u1_uk_K_r7_reg[23]/P0001  , \u1_uk_K_r7_reg[24]/NET0131  , \u1_uk_K_r7_reg[25]/NET0131  , \u1_uk_K_r7_reg[26]/P0001  , \u1_uk_K_r7_reg[27]/NET0131  , \u1_uk_K_r7_reg[28]/NET0131  , \u1_uk_K_r7_reg[29]/NET0131  , \u1_uk_K_r7_reg[2]/NET0131  , \u1_uk_K_r7_reg[30]/P0001  , \u1_uk_K_r7_reg[31]/NET0131  , \u1_uk_K_r7_reg[32]/NET0131  , \u1_uk_K_r7_reg[33]/NET0131  , \u1_uk_K_r7_reg[34]/NET0131  , \u1_uk_K_r7_reg[35]/NET0131  , \u1_uk_K_r7_reg[36]/NET0131  , \u1_uk_K_r7_reg[37]/NET0131  , \u1_uk_K_r7_reg[38]/NET0131  , \u1_uk_K_r7_reg[39]/NET0131  , \u1_uk_K_r7_reg[3]/NET0131  , \u1_uk_K_r7_reg[40]/NET0131  , \u1_uk_K_r7_reg[41]/NET0131  , \u1_uk_K_r7_reg[42]/NET0131  , \u1_uk_K_r7_reg[43]/NET0131  , \u1_uk_K_r7_reg[44]/NET0131  , \u1_uk_K_r7_reg[45]/NET0131  , \u1_uk_K_r7_reg[46]/NET0131  , \u1_uk_K_r7_reg[47]/NET0131  , \u1_uk_K_r7_reg[48]/NET0131  , \u1_uk_K_r7_reg[49]/NET0131  , \u1_uk_K_r7_reg[4]/NET0131  , \u1_uk_K_r7_reg[50]/NET0131  , \u1_uk_K_r7_reg[51]/NET0131  , \u1_uk_K_r7_reg[52]/NET0131  , \u1_uk_K_r7_reg[53]/NET0131  , \u1_uk_K_r7_reg[54]/NET0131  , \u1_uk_K_r7_reg[55]/P0001  , \u1_uk_K_r7_reg[5]/NET0131  , \u1_uk_K_r7_reg[6]/NET0131  , \u1_uk_K_r7_reg[7]/NET0131  , \u1_uk_K_r7_reg[8]/NET0131  , \u1_uk_K_r7_reg[9]/NET0131  , \u1_uk_K_r8_reg[0]/NET0131  , \u1_uk_K_r8_reg[10]/NET0131  , \u1_uk_K_r8_reg[11]/NET0131  , \u1_uk_K_r8_reg[12]/NET0131  , \u1_uk_K_r8_reg[13]/P0001  , \u1_uk_K_r8_reg[14]/NET0131  , \u1_uk_K_r8_reg[15]/NET0131  , \u1_uk_K_r8_reg[16]/NET0131  , \u1_uk_K_r8_reg[17]/NET0131  , \u1_uk_K_r8_reg[18]/NET0131  , \u1_uk_K_r8_reg[19]/NET0131  , \u1_uk_K_r8_reg[1]/NET0131  , \u1_uk_K_r8_reg[20]/NET0131  , \u1_uk_K_r8_reg[21]/NET0131  , \u1_uk_K_r8_reg[22]/NET0131  , \u1_uk_K_r8_reg[23]/NET0131  , \u1_uk_K_r8_reg[24]/NET0131  , \u1_uk_K_r8_reg[25]/NET0131  , \u1_uk_K_r8_reg[26]/NET0131  , \u1_uk_K_r8_reg[27]/NET0131  , \u1_uk_K_r8_reg[28]/NET0131  , \u1_uk_K_r8_reg[29]/NET0131  , \u1_uk_K_r8_reg[2]/NET0131  , \u1_uk_K_r8_reg[30]/NET0131  , \u1_uk_K_r8_reg[31]/NET0131  , \u1_uk_K_r8_reg[32]/NET0131  , \u1_uk_K_r8_reg[33]/NET0131  , \u1_uk_K_r8_reg[34]/NET0131  , \u1_uk_K_r8_reg[35]/NET0131  , \u1_uk_K_r8_reg[36]/NET0131  , \u1_uk_K_r8_reg[37]/P0001  , \u1_uk_K_r8_reg[38]/NET0131  , \u1_uk_K_r8_reg[39]/NET0131  , \u1_uk_K_r8_reg[3]/NET0131  , \u1_uk_K_r8_reg[40]/NET0131  , \u1_uk_K_r8_reg[41]/NET0131  , \u1_uk_K_r8_reg[42]/NET0131  , \u1_uk_K_r8_reg[43]/NET0131  , \u1_uk_K_r8_reg[44]/NET0131  , \u1_uk_K_r8_reg[46]/NET0131  , \u1_uk_K_r8_reg[47]/NET0131  , \u1_uk_K_r8_reg[48]/NET0131  , \u1_uk_K_r8_reg[49]/NET0131  , \u1_uk_K_r8_reg[4]/NET0131  , \u1_uk_K_r8_reg[50]/NET0131  , \u1_uk_K_r8_reg[51]/NET0131  , \u1_uk_K_r8_reg[52]/NET0131  , \u1_uk_K_r8_reg[53]/NET0131  , \u1_uk_K_r8_reg[54]/NET0131  , \u1_uk_K_r8_reg[55]/NET0131  , \u1_uk_K_r8_reg[5]/NET0131  , \u1_uk_K_r8_reg[6]/NET0131  , \u1_uk_K_r8_reg[7]/NET0131  , \u1_uk_K_r8_reg[8]/NET0131  , \u1_uk_K_r8_reg[9]/NET0131  , \u1_uk_K_r9_reg[0]/P0001  , \u1_uk_K_r9_reg[10]/NET0131  , \u1_uk_K_r9_reg[11]/NET0131  , \u1_uk_K_r9_reg[12]/NET0131  , \u1_uk_K_r9_reg[13]/NET0131  , \u1_uk_K_r9_reg[14]/NET0131  , \u1_uk_K_r9_reg[15]/NET0131  , \u1_uk_K_r9_reg[16]/NET0131  , \u1_uk_K_r9_reg[17]/NET0131  , \u1_uk_K_r9_reg[18]/NET0131  , \u1_uk_K_r9_reg[19]/NET0131  , \u1_uk_K_r9_reg[1]/NET0131  , \u1_uk_K_r9_reg[20]/NET0131  , \u1_uk_K_r9_reg[21]/NET0131  , \u1_uk_K_r9_reg[22]/NET0131  , \u1_uk_K_r9_reg[23]/NET0131  , \u1_uk_K_r9_reg[25]/NET0131  , \u1_uk_K_r9_reg[26]/NET0131  , \u1_uk_K_r9_reg[27]/P0001  , \u1_uk_K_r9_reg[28]/NET0131  , \u1_uk_K_r9_reg[29]/NET0131  , \u1_uk_K_r9_reg[30]/NET0131  , \u1_uk_K_r9_reg[31]/P0001  , \u1_uk_K_r9_reg[32]/NET0131  , \u1_uk_K_r9_reg[33]/NET0131  , \u1_uk_K_r9_reg[34]/NET0131  , \u1_uk_K_r9_reg[35]/NET0131  , \u1_uk_K_r9_reg[36]/NET0131  , \u1_uk_K_r9_reg[37]/NET0131  , \u1_uk_K_r9_reg[38]/NET0131  , \u1_uk_K_r9_reg[39]/NET0131  , \u1_uk_K_r9_reg[3]/NET0131  , \u1_uk_K_r9_reg[40]/NET0131  , \u1_uk_K_r9_reg[41]/NET0131  , \u1_uk_K_r9_reg[42]/NET0131  , \u1_uk_K_r9_reg[43]/NET0131  , \u1_uk_K_r9_reg[44]/NET0131  , \u1_uk_K_r9_reg[45]/NET0131  , \u1_uk_K_r9_reg[46]/NET0131  , \u1_uk_K_r9_reg[47]/NET0131  , \u1_uk_K_r9_reg[48]/NET0131  , \u1_uk_K_r9_reg[49]/NET0131  , \u1_uk_K_r9_reg[4]/NET0131  , \u1_uk_K_r9_reg[50]/NET0131  , \u1_uk_K_r9_reg[51]/NET0131  , \u1_uk_K_r9_reg[52]/NET0131  , \u1_uk_K_r9_reg[53]/NET0131  , \u1_uk_K_r9_reg[54]/NET0131  , \u1_uk_K_r9_reg[55]/NET0131  , \u1_uk_K_r9_reg[5]/NET0131  , \u1_uk_K_r9_reg[6]/NET0131  , \u1_uk_K_r9_reg[7]/NET0131  , \u1_uk_K_r9_reg[8]/NET0131  , \u1_uk_K_r9_reg[9]/NET0131  , \u2_L0_reg[10]/NET0131  , \u2_L0_reg[11]/NET0131  , \u2_L0_reg[12]/NET0131  , \u2_L0_reg[13]/NET0131  , \u2_L0_reg[14]/NET0131  , \u2_L0_reg[15]/NET0131  , \u2_L0_reg[16]/NET0131  , \u2_L0_reg[17]/NET0131  , \u2_L0_reg[18]/P0001  , \u2_L0_reg[19]/NET0131  , \u2_L0_reg[1]/NET0131  , \u2_L0_reg[20]/NET0131  , \u2_L0_reg[21]/NET0131  , \u2_L0_reg[22]/NET0131  , \u2_L0_reg[23]/NET0131  , \u2_L0_reg[24]/NET0131  , \u2_L0_reg[25]/NET0131  , \u2_L0_reg[26]/NET0131  , \u2_L0_reg[27]/NET0131  , \u2_L0_reg[28]/NET0131  , \u2_L0_reg[29]/NET0131  , \u2_L0_reg[2]/NET0131  , \u2_L0_reg[30]/NET0131  , \u2_L0_reg[31]/NET0131  , \u2_L0_reg[32]/NET0131  , \u2_L0_reg[3]/NET0131  , \u2_L0_reg[4]/NET0131  , \u2_L0_reg[5]/NET0131  , \u2_L0_reg[6]/NET0131  , \u2_L0_reg[7]/NET0131  , \u2_L0_reg[8]/NET0131  , \u2_L0_reg[9]/NET0131  , \u2_L10_reg[10]/NET0131  , \u2_L10_reg[11]/NET0131  , \u2_L10_reg[12]/NET0131  , \u2_L10_reg[13]/NET0131  , \u2_L10_reg[14]/NET0131  , \u2_L10_reg[15]/NET0131  , \u2_L10_reg[16]/NET0131  , \u2_L10_reg[17]/NET0131  , \u2_L10_reg[18]/P0001  , \u2_L10_reg[19]/NET0131  , \u2_L10_reg[1]/NET0131  , \u2_L10_reg[20]/NET0131  , \u2_L10_reg[21]/NET0131  , \u2_L10_reg[22]/NET0131  , \u2_L10_reg[23]/NET0131  , \u2_L10_reg[24]/NET0131  , \u2_L10_reg[25]/NET0131  , \u2_L10_reg[26]/NET0131  , \u2_L10_reg[27]/NET0131  , \u2_L10_reg[28]/NET0131  , \u2_L10_reg[29]/NET0131  , \u2_L10_reg[2]/NET0131  , \u2_L10_reg[30]/NET0131  , \u2_L10_reg[31]/NET0131  , \u2_L10_reg[32]/NET0131  , \u2_L10_reg[3]/NET0131  , \u2_L10_reg[4]/NET0131  , \u2_L10_reg[5]/NET0131  , \u2_L10_reg[6]/NET0131  , \u2_L10_reg[7]/NET0131  , \u2_L10_reg[8]/NET0131  , \u2_L10_reg[9]/NET0131  , \u2_L11_reg[10]/NET0131  , \u2_L11_reg[11]/NET0131  , \u2_L11_reg[12]/NET0131  , \u2_L11_reg[13]/NET0131  , \u2_L11_reg[14]/NET0131  , \u2_L11_reg[15]/NET0131  , \u2_L11_reg[16]/NET0131  , \u2_L11_reg[17]/NET0131  , \u2_L11_reg[18]/P0001  , \u2_L11_reg[19]/NET0131  , \u2_L11_reg[1]/NET0131  , \u2_L11_reg[20]/NET0131  , \u2_L11_reg[21]/NET0131  , \u2_L11_reg[22]/NET0131  , \u2_L11_reg[23]/NET0131  , \u2_L11_reg[24]/NET0131  , \u2_L11_reg[25]/NET0131  , \u2_L11_reg[26]/NET0131  , \u2_L11_reg[27]/NET0131  , \u2_L11_reg[28]/NET0131  , \u2_L11_reg[29]/NET0131  , \u2_L11_reg[2]/NET0131  , \u2_L11_reg[30]/NET0131  , \u2_L11_reg[31]/NET0131  , \u2_L11_reg[32]/NET0131  , \u2_L11_reg[3]/NET0131  , \u2_L11_reg[4]/NET0131  , \u2_L11_reg[5]/NET0131  , \u2_L11_reg[6]/NET0131  , \u2_L11_reg[7]/NET0131  , \u2_L11_reg[8]/NET0131  , \u2_L11_reg[9]/NET0131  , \u2_L12_reg[10]/NET0131  , \u2_L12_reg[11]/NET0131  , \u2_L12_reg[12]/NET0131  , \u2_L12_reg[13]/NET0131  , \u2_L12_reg[14]/NET0131  , \u2_L12_reg[15]/NET0131  , \u2_L12_reg[16]/NET0131  , \u2_L12_reg[17]/NET0131  , \u2_L12_reg[18]/P0001  , \u2_L12_reg[19]/NET0131  , \u2_L12_reg[1]/NET0131  , \u2_L12_reg[20]/NET0131  , \u2_L12_reg[21]/NET0131  , \u2_L12_reg[22]/NET0131  , \u2_L12_reg[23]/NET0131  , \u2_L12_reg[24]/NET0131  , \u2_L12_reg[25]/NET0131  , \u2_L12_reg[26]/NET0131  , \u2_L12_reg[27]/NET0131  , \u2_L12_reg[28]/NET0131  , \u2_L12_reg[29]/NET0131  , \u2_L12_reg[2]/NET0131  , \u2_L12_reg[30]/NET0131  , \u2_L12_reg[31]/NET0131  , \u2_L12_reg[32]/NET0131  , \u2_L12_reg[3]/NET0131  , \u2_L12_reg[4]/NET0131  , \u2_L12_reg[5]/NET0131  , \u2_L12_reg[6]/NET0131  , \u2_L12_reg[7]/NET0131  , \u2_L12_reg[8]/NET0131  , \u2_L12_reg[9]/NET0131  , \u2_L13_reg[10]/NET0131  , \u2_L13_reg[11]/NET0131  , \u2_L13_reg[12]/NET0131  , \u2_L13_reg[13]/NET0131  , \u2_L13_reg[14]/NET0131  , \u2_L13_reg[15]/NET0131  , \u2_L13_reg[16]/NET0131  , \u2_L13_reg[17]/NET0131  , \u2_L13_reg[18]/P0001  , \u2_L13_reg[19]/P0001  , \u2_L13_reg[1]/NET0131  , \u2_L13_reg[20]/NET0131  , \u2_L13_reg[21]/NET0131  , \u2_L13_reg[22]/NET0131  , \u2_L13_reg[23]/P0001  , \u2_L13_reg[24]/NET0131  , \u2_L13_reg[25]/NET0131  , \u2_L13_reg[26]/NET0131  , \u2_L13_reg[27]/NET0131  , \u2_L13_reg[28]/NET0131  , \u2_L13_reg[29]/NET0131  , \u2_L13_reg[2]/NET0131  , \u2_L13_reg[30]/NET0131  , \u2_L13_reg[31]/NET0131  , \u2_L13_reg[32]/NET0131  , \u2_L13_reg[3]/NET0131  , \u2_L13_reg[4]/NET0131  , \u2_L13_reg[5]/NET0131  , \u2_L13_reg[6]/NET0131  , \u2_L13_reg[7]/NET0131  , \u2_L13_reg[8]/NET0131  , \u2_L13_reg[9]/NET0131  , \u2_L14_reg[10]/P0001  , \u2_L14_reg[11]/P0001  , \u2_L14_reg[12]/P0001  , \u2_L14_reg[13]/P0001  , \u2_L14_reg[14]/P0001  , \u2_L14_reg[15]/P0001  , \u2_L14_reg[16]/P0001  , \u2_L14_reg[17]/P0001  , \u2_L14_reg[18]/P0001  , \u2_L14_reg[19]/P0001  , \u2_L14_reg[1]/P0001  , \u2_L14_reg[20]/P0001  , \u2_L14_reg[21]/P0001  , \u2_L14_reg[22]/P0001  , \u2_L14_reg[23]/P0001  , \u2_L14_reg[24]/P0001  , \u2_L14_reg[25]/P0001  , \u2_L14_reg[26]/P0001  , \u2_L14_reg[27]/P0001  , \u2_L14_reg[28]/P0001  , \u2_L14_reg[29]/P0001  , \u2_L14_reg[2]/P0001  , \u2_L14_reg[30]/P0001  , \u2_L14_reg[31]/P0001  , \u2_L14_reg[32]/P0001  , \u2_L14_reg[3]/P0001  , \u2_L14_reg[4]/P0001  , \u2_L14_reg[5]/P0001  , \u2_L14_reg[6]/P0001  , \u2_L14_reg[7]/P0001  , \u2_L14_reg[8]/P0001  , \u2_L14_reg[9]/P0001  , \u2_L1_reg[10]/NET0131  , \u2_L1_reg[11]/NET0131  , \u2_L1_reg[12]/NET0131  , \u2_L1_reg[13]/NET0131  , \u2_L1_reg[14]/NET0131  , \u2_L1_reg[15]/NET0131  , \u2_L1_reg[16]/NET0131  , \u2_L1_reg[17]/NET0131  , \u2_L1_reg[18]/P0001  , \u2_L1_reg[19]/NET0131  , \u2_L1_reg[1]/NET0131  , \u2_L1_reg[20]/NET0131  , \u2_L1_reg[21]/NET0131  , \u2_L1_reg[22]/NET0131  , \u2_L1_reg[23]/NET0131  , \u2_L1_reg[24]/NET0131  , \u2_L1_reg[25]/NET0131  , \u2_L1_reg[26]/NET0131  , \u2_L1_reg[27]/NET0131  , \u2_L1_reg[28]/NET0131  , \u2_L1_reg[29]/NET0131  , \u2_L1_reg[2]/NET0131  , \u2_L1_reg[30]/NET0131  , \u2_L1_reg[31]/NET0131  , \u2_L1_reg[32]/NET0131  , \u2_L1_reg[3]/NET0131  , \u2_L1_reg[4]/NET0131  , \u2_L1_reg[5]/NET0131  , \u2_L1_reg[6]/NET0131  , \u2_L1_reg[7]/NET0131  , \u2_L1_reg[8]/NET0131  , \u2_L1_reg[9]/NET0131  , \u2_L2_reg[10]/NET0131  , \u2_L2_reg[11]/NET0131  , \u2_L2_reg[12]/NET0131  , \u2_L2_reg[13]/NET0131  , \u2_L2_reg[14]/NET0131  , \u2_L2_reg[15]/NET0131  , \u2_L2_reg[16]/NET0131  , \u2_L2_reg[17]/NET0131  , \u2_L2_reg[18]/P0001  , \u2_L2_reg[19]/NET0131  , \u2_L2_reg[1]/NET0131  , \u2_L2_reg[20]/NET0131  , \u2_L2_reg[21]/NET0131  , \u2_L2_reg[22]/NET0131  , \u2_L2_reg[23]/NET0131  , \u2_L2_reg[24]/NET0131  , \u2_L2_reg[25]/NET0131  , \u2_L2_reg[26]/NET0131  , \u2_L2_reg[27]/NET0131  , \u2_L2_reg[28]/NET0131  , \u2_L2_reg[29]/NET0131  , \u2_L2_reg[2]/NET0131  , \u2_L2_reg[30]/NET0131  , \u2_L2_reg[31]/NET0131  , \u2_L2_reg[32]/NET0131  , \u2_L2_reg[3]/NET0131  , \u2_L2_reg[4]/NET0131  , \u2_L2_reg[5]/NET0131  , \u2_L2_reg[6]/NET0131  , \u2_L2_reg[7]/NET0131  , \u2_L2_reg[8]/NET0131  , \u2_L2_reg[9]/NET0131  , \u2_L3_reg[10]/NET0131  , \u2_L3_reg[11]/NET0131  , \u2_L3_reg[12]/NET0131  , \u2_L3_reg[13]/NET0131  , \u2_L3_reg[14]/NET0131  , \u2_L3_reg[15]/NET0131  , \u2_L3_reg[16]/NET0131  , \u2_L3_reg[17]/NET0131  , \u2_L3_reg[18]/P0001  , \u2_L3_reg[19]/NET0131  , \u2_L3_reg[1]/NET0131  , \u2_L3_reg[20]/NET0131  , \u2_L3_reg[21]/NET0131  , \u2_L3_reg[22]/NET0131  , \u2_L3_reg[23]/NET0131  , \u2_L3_reg[24]/NET0131  , \u2_L3_reg[25]/NET0131  , \u2_L3_reg[26]/NET0131  , \u2_L3_reg[27]/NET0131  , \u2_L3_reg[28]/NET0131  , \u2_L3_reg[29]/NET0131  , \u2_L3_reg[2]/NET0131  , \u2_L3_reg[30]/NET0131  , \u2_L3_reg[31]/NET0131  , \u2_L3_reg[32]/NET0131  , \u2_L3_reg[3]/NET0131  , \u2_L3_reg[4]/NET0131  , \u2_L3_reg[5]/NET0131  , \u2_L3_reg[6]/NET0131  , \u2_L3_reg[7]/NET0131  , \u2_L3_reg[8]/NET0131  , \u2_L3_reg[9]/NET0131  , \u2_L4_reg[10]/NET0131  , \u2_L4_reg[11]/NET0131  , \u2_L4_reg[12]/NET0131  , \u2_L4_reg[13]/NET0131  , \u2_L4_reg[14]/NET0131  , \u2_L4_reg[15]/NET0131  , \u2_L4_reg[16]/NET0131  , \u2_L4_reg[17]/NET0131  , \u2_L4_reg[18]/P0001  , \u2_L4_reg[19]/NET0131  , \u2_L4_reg[1]/NET0131  , \u2_L4_reg[20]/NET0131  , \u2_L4_reg[21]/NET0131  , \u2_L4_reg[22]/NET0131  , \u2_L4_reg[23]/NET0131  , \u2_L4_reg[24]/NET0131  , \u2_L4_reg[25]/NET0131  , \u2_L4_reg[26]/NET0131  , \u2_L4_reg[27]/NET0131  , \u2_L4_reg[28]/NET0131  , \u2_L4_reg[29]/NET0131  , \u2_L4_reg[2]/NET0131  , \u2_L4_reg[30]/NET0131  , \u2_L4_reg[31]/NET0131  , \u2_L4_reg[32]/NET0131  , \u2_L4_reg[3]/NET0131  , \u2_L4_reg[4]/NET0131  , \u2_L4_reg[5]/NET0131  , \u2_L4_reg[6]/NET0131  , \u2_L4_reg[7]/NET0131  , \u2_L4_reg[8]/NET0131  , \u2_L4_reg[9]/NET0131  , \u2_L5_reg[10]/NET0131  , \u2_L5_reg[11]/NET0131  , \u2_L5_reg[12]/NET0131  , \u2_L5_reg[13]/NET0131  , \u2_L5_reg[14]/NET0131  , \u2_L5_reg[15]/NET0131  , \u2_L5_reg[16]/NET0131  , \u2_L5_reg[17]/NET0131  , \u2_L5_reg[18]/NET0131  , \u2_L5_reg[19]/NET0131  , \u2_L5_reg[1]/NET0131  , \u2_L5_reg[20]/NET0131  , \u2_L5_reg[21]/NET0131  , \u2_L5_reg[22]/NET0131  , \u2_L5_reg[23]/NET0131  , \u2_L5_reg[24]/NET0131  , \u2_L5_reg[25]/NET0131  , \u2_L5_reg[26]/NET0131  , \u2_L5_reg[27]/NET0131  , \u2_L5_reg[28]/NET0131  , \u2_L5_reg[29]/NET0131  , \u2_L5_reg[2]/NET0131  , \u2_L5_reg[30]/NET0131  , \u2_L5_reg[31]/NET0131  , \u2_L5_reg[32]/NET0131  , \u2_L5_reg[3]/NET0131  , \u2_L5_reg[4]/NET0131  , \u2_L5_reg[5]/NET0131  , \u2_L5_reg[6]/NET0131  , \u2_L5_reg[7]/NET0131  , \u2_L5_reg[8]/NET0131  , \u2_L5_reg[9]/NET0131  , \u2_L6_reg[10]/NET0131  , \u2_L6_reg[11]/NET0131  , \u2_L6_reg[12]/NET0131  , \u2_L6_reg[13]/NET0131  , \u2_L6_reg[14]/NET0131  , \u2_L6_reg[15]/NET0131  , \u2_L6_reg[16]/NET0131  , \u2_L6_reg[17]/NET0131  , \u2_L6_reg[18]/P0001  , \u2_L6_reg[19]/NET0131  , \u2_L6_reg[1]/NET0131  , \u2_L6_reg[20]/NET0131  , \u2_L6_reg[21]/NET0131  , \u2_L6_reg[22]/NET0131  , \u2_L6_reg[23]/NET0131  , \u2_L6_reg[24]/NET0131  , \u2_L6_reg[25]/NET0131  , \u2_L6_reg[26]/NET0131  , \u2_L6_reg[27]/NET0131  , \u2_L6_reg[28]/NET0131  , \u2_L6_reg[29]/NET0131  , \u2_L6_reg[2]/NET0131  , \u2_L6_reg[30]/NET0131  , \u2_L6_reg[31]/NET0131  , \u2_L6_reg[32]/NET0131  , \u2_L6_reg[3]/NET0131  , \u2_L6_reg[4]/NET0131  , \u2_L6_reg[5]/NET0131  , \u2_L6_reg[6]/NET0131  , \u2_L6_reg[7]/NET0131  , \u2_L6_reg[8]/NET0131  , \u2_L6_reg[9]/NET0131  , \u2_L7_reg[10]/NET0131  , \u2_L7_reg[11]/NET0131  , \u2_L7_reg[12]/NET0131  , \u2_L7_reg[13]/NET0131  , \u2_L7_reg[14]/NET0131  , \u2_L7_reg[15]/NET0131  , \u2_L7_reg[16]/NET0131  , \u2_L7_reg[17]/NET0131  , \u2_L7_reg[18]/P0001  , \u2_L7_reg[19]/NET0131  , \u2_L7_reg[1]/NET0131  , \u2_L7_reg[20]/NET0131  , \u2_L7_reg[21]/NET0131  , \u2_L7_reg[22]/NET0131  , \u2_L7_reg[23]/NET0131  , \u2_L7_reg[24]/NET0131  , \u2_L7_reg[25]/NET0131  , \u2_L7_reg[26]/NET0131  , \u2_L7_reg[27]/NET0131  , \u2_L7_reg[28]/NET0131  , \u2_L7_reg[29]/NET0131  , \u2_L7_reg[2]/NET0131  , \u2_L7_reg[30]/NET0131  , \u2_L7_reg[31]/NET0131  , \u2_L7_reg[32]/NET0131  , \u2_L7_reg[3]/NET0131  , \u2_L7_reg[4]/NET0131  , \u2_L7_reg[5]/NET0131  , \u2_L7_reg[6]/NET0131  , \u2_L7_reg[7]/NET0131  , \u2_L7_reg[8]/NET0131  , \u2_L7_reg[9]/NET0131  , \u2_L8_reg[10]/NET0131  , \u2_L8_reg[11]/NET0131  , \u2_L8_reg[12]/NET0131  , \u2_L8_reg[13]/NET0131  , \u2_L8_reg[14]/NET0131  , \u2_L8_reg[15]/NET0131  , \u2_L8_reg[16]/NET0131  , \u2_L8_reg[17]/NET0131  , \u2_L8_reg[18]/P0001  , \u2_L8_reg[19]/NET0131  , \u2_L8_reg[1]/NET0131  , \u2_L8_reg[20]/NET0131  , \u2_L8_reg[21]/NET0131  , \u2_L8_reg[22]/NET0131  , \u2_L8_reg[23]/NET0131  , \u2_L8_reg[24]/NET0131  , \u2_L8_reg[25]/NET0131  , \u2_L8_reg[26]/NET0131  , \u2_L8_reg[27]/NET0131  , \u2_L8_reg[28]/NET0131  , \u2_L8_reg[29]/NET0131  , \u2_L8_reg[2]/NET0131  , \u2_L8_reg[30]/NET0131  , \u2_L8_reg[31]/NET0131  , \u2_L8_reg[32]/NET0131  , \u2_L8_reg[3]/NET0131  , \u2_L8_reg[4]/NET0131  , \u2_L8_reg[5]/NET0131  , \u2_L8_reg[6]/NET0131  , \u2_L8_reg[7]/NET0131  , \u2_L8_reg[8]/NET0131  , \u2_L8_reg[9]/NET0131  , \u2_L9_reg[10]/NET0131  , \u2_L9_reg[11]/NET0131  , \u2_L9_reg[12]/NET0131  , \u2_L9_reg[13]/NET0131  , \u2_L9_reg[14]/NET0131  , \u2_L9_reg[15]/NET0131  , \u2_L9_reg[16]/NET0131  , \u2_L9_reg[17]/NET0131  , \u2_L9_reg[18]/P0001  , \u2_L9_reg[19]/NET0131  , \u2_L9_reg[1]/NET0131  , \u2_L9_reg[20]/NET0131  , \u2_L9_reg[21]/NET0131  , \u2_L9_reg[22]/NET0131  , \u2_L9_reg[23]/NET0131  , \u2_L9_reg[24]/NET0131  , \u2_L9_reg[25]/NET0131  , \u2_L9_reg[26]/NET0131  , \u2_L9_reg[27]/NET0131  , \u2_L9_reg[28]/NET0131  , \u2_L9_reg[29]/NET0131  , \u2_L9_reg[2]/NET0131  , \u2_L9_reg[30]/NET0131  , \u2_L9_reg[31]/NET0131  , \u2_L9_reg[32]/NET0131  , \u2_L9_reg[3]/NET0131  , \u2_L9_reg[4]/NET0131  , \u2_L9_reg[5]/NET0131  , \u2_L9_reg[6]/NET0131  , \u2_L9_reg[7]/NET0131  , \u2_L9_reg[8]/NET0131  , \u2_L9_reg[9]/NET0131  , \u2_R0_reg[10]/NET0131  , \u2_R0_reg[11]/P0001  , \u2_R0_reg[12]/NET0131  , \u2_R0_reg[13]/NET0131  , \u2_R0_reg[14]/NET0131  , \u2_R0_reg[15]/NET0131  , \u2_R0_reg[16]/NET0131  , \u2_R0_reg[17]/NET0131  , \u2_R0_reg[18]/NET0131  , \u2_R0_reg[19]/NET0131  , \u2_R0_reg[1]/NET0131  , \u2_R0_reg[20]/NET0131  , \u2_R0_reg[21]/NET0131  , \u2_R0_reg[22]/NET0131  , \u2_R0_reg[23]/NET0131  , \u2_R0_reg[24]/NET0131  , \u2_R0_reg[25]/NET0131  , \u2_R0_reg[26]/NET0131  , \u2_R0_reg[27]/NET0131  , \u2_R0_reg[28]/NET0131  , \u2_R0_reg[29]/NET0131  , \u2_R0_reg[2]/NET0131  , \u2_R0_reg[30]/NET0131  , \u2_R0_reg[31]/P0001  , \u2_R0_reg[32]/NET0131  , \u2_R0_reg[3]/NET0131  , \u2_R0_reg[4]/NET0131  , \u2_R0_reg[5]/NET0131  , \u2_R0_reg[6]/NET0131  , \u2_R0_reg[7]/NET0131  , \u2_R0_reg[8]/NET0131  , \u2_R0_reg[9]/NET0131  , \u2_R10_reg[10]/NET0131  , \u2_R10_reg[11]/NET0131  , \u2_R10_reg[12]/NET0131  , \u2_R10_reg[13]/NET0131  , \u2_R10_reg[14]/NET0131  , \u2_R10_reg[15]/NET0131  , \u2_R10_reg[16]/NET0131  , \u2_R10_reg[17]/NET0131  , \u2_R10_reg[18]/NET0131  , \u2_R10_reg[19]/NET0131  , \u2_R10_reg[1]/NET0131  , \u2_R10_reg[20]/NET0131  , \u2_R10_reg[21]/NET0131  , \u2_R10_reg[22]/NET0131  , \u2_R10_reg[23]/NET0131  , \u2_R10_reg[24]/NET0131  , \u2_R10_reg[25]/NET0131  , \u2_R10_reg[26]/NET0131  , \u2_R10_reg[27]/NET0131  , \u2_R10_reg[28]/NET0131  , \u2_R10_reg[29]/NET0131  , \u2_R10_reg[2]/NET0131  , \u2_R10_reg[30]/NET0131  , \u2_R10_reg[31]/P0001  , \u2_R10_reg[32]/NET0131  , \u2_R10_reg[3]/NET0131  , \u2_R10_reg[4]/NET0131  , \u2_R10_reg[5]/NET0131  , \u2_R10_reg[6]/NET0131  , \u2_R10_reg[7]/NET0131  , \u2_R10_reg[8]/NET0131  , \u2_R10_reg[9]/NET0131  , \u2_R11_reg[10]/NET0131  , \u2_R11_reg[11]/NET0131  , \u2_R11_reg[12]/NET0131  , \u2_R11_reg[13]/NET0131  , \u2_R11_reg[14]/NET0131  , \u2_R11_reg[15]/NET0131  , \u2_R11_reg[16]/NET0131  , \u2_R11_reg[17]/NET0131  , \u2_R11_reg[18]/NET0131  , \u2_R11_reg[19]/NET0131  , \u2_R11_reg[1]/NET0131  , \u2_R11_reg[20]/NET0131  , \u2_R11_reg[21]/NET0131  , \u2_R11_reg[22]/NET0131  , \u2_R11_reg[23]/NET0131  , \u2_R11_reg[24]/NET0131  , \u2_R11_reg[25]/NET0131  , \u2_R11_reg[26]/NET0131  , \u2_R11_reg[27]/NET0131  , \u2_R11_reg[28]/NET0131  , \u2_R11_reg[29]/NET0131  , \u2_R11_reg[2]/NET0131  , \u2_R11_reg[30]/NET0131  , \u2_R11_reg[31]/P0001  , \u2_R11_reg[32]/NET0131  , \u2_R11_reg[3]/NET0131  , \u2_R11_reg[4]/NET0131  , \u2_R11_reg[5]/NET0131  , \u2_R11_reg[6]/NET0131  , \u2_R11_reg[7]/NET0131  , \u2_R11_reg[8]/NET0131  , \u2_R11_reg[9]/NET0131  , \u2_R12_reg[10]/NET0131  , \u2_R12_reg[11]/NET0131  , \u2_R12_reg[12]/NET0131  , \u2_R12_reg[13]/NET0131  , \u2_R12_reg[14]/NET0131  , \u2_R12_reg[15]/NET0131  , \u2_R12_reg[16]/NET0131  , \u2_R12_reg[17]/NET0131  , \u2_R12_reg[18]/NET0131  , \u2_R12_reg[19]/NET0131  , \u2_R12_reg[1]/NET0131  , \u2_R12_reg[20]/NET0131  , \u2_R12_reg[21]/NET0131  , \u2_R12_reg[22]/NET0131  , \u2_R12_reg[23]/NET0131  , \u2_R12_reg[24]/NET0131  , \u2_R12_reg[25]/NET0131  , \u2_R12_reg[26]/NET0131  , \u2_R12_reg[27]/NET0131  , \u2_R12_reg[28]/NET0131  , \u2_R12_reg[29]/NET0131  , \u2_R12_reg[2]/NET0131  , \u2_R12_reg[30]/NET0131  , \u2_R12_reg[31]/P0001  , \u2_R12_reg[32]/NET0131  , \u2_R12_reg[3]/NET0131  , \u2_R12_reg[4]/NET0131  , \u2_R12_reg[5]/NET0131  , \u2_R12_reg[6]/NET0131  , \u2_R12_reg[7]/NET0131  , \u2_R12_reg[8]/NET0131  , \u2_R12_reg[9]/NET0131  , \u2_R13_reg[10]/NET0131  , \u2_R13_reg[11]/NET0131  , \u2_R13_reg[12]/NET0131  , \u2_R13_reg[13]/NET0131  , \u2_R13_reg[14]/NET0131  , \u2_R13_reg[15]/NET0131  , \u2_R13_reg[16]/NET0131  , \u2_R13_reg[17]/NET0131  , \u2_R13_reg[18]/NET0131  , \u2_R13_reg[19]/NET0131  , \u2_R13_reg[1]/NET0131  , \u2_R13_reg[20]/NET0131  , \u2_R13_reg[21]/NET0131  , \u2_R13_reg[22]/NET0131  , \u2_R13_reg[23]/NET0131  , \u2_R13_reg[24]/NET0131  , \u2_R13_reg[25]/NET0131  , \u2_R13_reg[26]/NET0131  , \u2_R13_reg[27]/P0001  , \u2_R13_reg[28]/NET0131  , \u2_R13_reg[29]/NET0131  , \u2_R13_reg[2]/NET0131  , \u2_R13_reg[30]/NET0131  , \u2_R13_reg[31]/P0001  , \u2_R13_reg[32]/NET0131  , \u2_R13_reg[3]/NET0131  , \u2_R13_reg[4]/NET0131  , \u2_R13_reg[5]/NET0131  , \u2_R13_reg[6]/NET0131  , \u2_R13_reg[7]/NET0131  , \u2_R13_reg[8]/NET0131  , \u2_R13_reg[9]/NET0131  , \u2_R14_reg[10]/P0001  , \u2_R14_reg[11]/P0001  , \u2_R14_reg[12]/NET0131  , \u2_R14_reg[13]/NET0131  , \u2_R14_reg[14]/NET0131  , \u2_R14_reg[15]/NET0131  , \u2_R14_reg[16]/NET0131  , \u2_R14_reg[17]/NET0131  , \u2_R14_reg[18]/NET0131  , \u2_R14_reg[19]/P0001  , \u2_R14_reg[1]/NET0131  , \u2_R14_reg[20]/NET0131  , \u2_R14_reg[21]/NET0131  , \u2_R14_reg[22]/P0001  , \u2_R14_reg[23]/P0001  , \u2_R14_reg[24]/NET0131  , \u2_R14_reg[25]/NET0131  , \u2_R14_reg[26]/P0001  , \u2_R14_reg[27]/P0001  , \u2_R14_reg[28]/NET0131  , \u2_R14_reg[29]/NET0131  , \u2_R14_reg[2]/NET0131  , \u2_R14_reg[30]/NET0131  , \u2_R14_reg[31]/P0001  , \u2_R14_reg[32]/NET0131  , \u2_R14_reg[3]/NET0131  , \u2_R14_reg[4]/NET0131  , \u2_R14_reg[5]/NET0131  , \u2_R14_reg[6]/NET0131  , \u2_R14_reg[7]/P0001  , \u2_R14_reg[8]/NET0131  , \u2_R14_reg[9]/NET0131  , \u2_R1_reg[10]/NET0131  , \u2_R1_reg[11]/P0001  , \u2_R1_reg[12]/NET0131  , \u2_R1_reg[13]/NET0131  , \u2_R1_reg[14]/NET0131  , \u2_R1_reg[15]/NET0131  , \u2_R1_reg[16]/NET0131  , \u2_R1_reg[17]/NET0131  , \u2_R1_reg[18]/NET0131  , \u2_R1_reg[19]/NET0131  , \u2_R1_reg[1]/NET0131  , \u2_R1_reg[20]/NET0131  , \u2_R1_reg[21]/NET0131  , \u2_R1_reg[22]/NET0131  , \u2_R1_reg[23]/NET0131  , \u2_R1_reg[24]/NET0131  , \u2_R1_reg[25]/NET0131  , \u2_R1_reg[26]/NET0131  , \u2_R1_reg[27]/NET0131  , \u2_R1_reg[28]/NET0131  , \u2_R1_reg[29]/NET0131  , \u2_R1_reg[2]/NET0131  , \u2_R1_reg[30]/NET0131  , \u2_R1_reg[31]/P0001  , \u2_R1_reg[32]/NET0131  , \u2_R1_reg[3]/NET0131  , \u2_R1_reg[4]/NET0131  , \u2_R1_reg[5]/NET0131  , \u2_R1_reg[6]/NET0131  , \u2_R1_reg[7]/NET0131  , \u2_R1_reg[8]/NET0131  , \u2_R1_reg[9]/NET0131  , \u2_R2_reg[10]/NET0131  , \u2_R2_reg[11]/NET0131  , \u2_R2_reg[12]/NET0131  , \u2_R2_reg[13]/NET0131  , \u2_R2_reg[14]/NET0131  , \u2_R2_reg[15]/NET0131  , \u2_R2_reg[16]/NET0131  , \u2_R2_reg[17]/NET0131  , \u2_R2_reg[18]/NET0131  , \u2_R2_reg[19]/NET0131  , \u2_R2_reg[1]/NET0131  , \u2_R2_reg[20]/NET0131  , \u2_R2_reg[21]/NET0131  , \u2_R2_reg[22]/NET0131  , \u2_R2_reg[23]/NET0131  , \u2_R2_reg[24]/NET0131  , \u2_R2_reg[25]/NET0131  , \u2_R2_reg[26]/NET0131  , \u2_R2_reg[27]/NET0131  , \u2_R2_reg[28]/NET0131  , \u2_R2_reg[29]/NET0131  , \u2_R2_reg[2]/NET0131  , \u2_R2_reg[30]/NET0131  , \u2_R2_reg[31]/P0001  , \u2_R2_reg[32]/NET0131  , \u2_R2_reg[3]/NET0131  , \u2_R2_reg[4]/NET0131  , \u2_R2_reg[5]/NET0131  , \u2_R2_reg[6]/NET0131  , \u2_R2_reg[7]/NET0131  , \u2_R2_reg[8]/NET0131  , \u2_R2_reg[9]/NET0131  , \u2_R3_reg[10]/NET0131  , \u2_R3_reg[11]/P0001  , \u2_R3_reg[12]/NET0131  , \u2_R3_reg[13]/NET0131  , \u2_R3_reg[14]/NET0131  , \u2_R3_reg[15]/NET0131  , \u2_R3_reg[16]/NET0131  , \u2_R3_reg[17]/NET0131  , \u2_R3_reg[18]/NET0131  , \u2_R3_reg[19]/NET0131  , \u2_R3_reg[1]/NET0131  , \u2_R3_reg[20]/NET0131  , \u2_R3_reg[21]/NET0131  , \u2_R3_reg[22]/NET0131  , \u2_R3_reg[23]/NET0131  , \u2_R3_reg[24]/NET0131  , \u2_R3_reg[25]/NET0131  , \u2_R3_reg[26]/NET0131  , \u2_R3_reg[27]/NET0131  , \u2_R3_reg[28]/NET0131  , \u2_R3_reg[29]/NET0131  , \u2_R3_reg[2]/NET0131  , \u2_R3_reg[30]/NET0131  , \u2_R3_reg[31]/P0001  , \u2_R3_reg[32]/NET0131  , \u2_R3_reg[3]/NET0131  , \u2_R3_reg[4]/NET0131  , \u2_R3_reg[5]/NET0131  , \u2_R3_reg[6]/NET0131  , \u2_R3_reg[7]/NET0131  , \u2_R3_reg[8]/NET0131  , \u2_R3_reg[9]/NET0131  , \u2_R4_reg[10]/NET0131  , \u2_R4_reg[11]/NET0131  , \u2_R4_reg[12]/NET0131  , \u2_R4_reg[13]/NET0131  , \u2_R4_reg[14]/NET0131  , \u2_R4_reg[15]/NET0131  , \u2_R4_reg[16]/NET0131  , \u2_R4_reg[17]/NET0131  , \u2_R4_reg[18]/NET0131  , \u2_R4_reg[19]/NET0131  , \u2_R4_reg[1]/NET0131  , \u2_R4_reg[20]/NET0131  , \u2_R4_reg[21]/NET0131  , \u2_R4_reg[22]/NET0131  , \u2_R4_reg[23]/NET0131  , \u2_R4_reg[24]/NET0131  , \u2_R4_reg[25]/NET0131  , \u2_R4_reg[26]/NET0131  , \u2_R4_reg[27]/NET0131  , \u2_R4_reg[28]/NET0131  , \u2_R4_reg[29]/NET0131  , \u2_R4_reg[2]/NET0131  , \u2_R4_reg[30]/NET0131  , \u2_R4_reg[31]/P0001  , \u2_R4_reg[32]/NET0131  , \u2_R4_reg[3]/NET0131  , \u2_R4_reg[4]/NET0131  , \u2_R4_reg[5]/NET0131  , \u2_R4_reg[6]/NET0131  , \u2_R4_reg[7]/NET0131  , \u2_R4_reg[8]/NET0131  , \u2_R4_reg[9]/NET0131  , \u2_R5_reg[10]/NET0131  , \u2_R5_reg[11]/NET0131  , \u2_R5_reg[12]/NET0131  , \u2_R5_reg[13]/NET0131  , \u2_R5_reg[14]/NET0131  , \u2_R5_reg[15]/NET0131  , \u2_R5_reg[16]/NET0131  , \u2_R5_reg[17]/NET0131  , \u2_R5_reg[18]/NET0131  , \u2_R5_reg[19]/NET0131  , \u2_R5_reg[1]/NET0131  , \u2_R5_reg[20]/NET0131  , \u2_R5_reg[21]/NET0131  , \u2_R5_reg[22]/NET0131  , \u2_R5_reg[23]/NET0131  , \u2_R5_reg[24]/NET0131  , \u2_R5_reg[25]/NET0131  , \u2_R5_reg[26]/NET0131  , \u2_R5_reg[27]/NET0131  , \u2_R5_reg[28]/NET0131  , \u2_R5_reg[29]/NET0131  , \u2_R5_reg[2]/NET0131  , \u2_R5_reg[30]/NET0131  , \u2_R5_reg[31]/P0001  , \u2_R5_reg[32]/NET0131  , \u2_R5_reg[3]/NET0131  , \u2_R5_reg[4]/NET0131  , \u2_R5_reg[5]/NET0131  , \u2_R5_reg[6]/NET0131  , \u2_R5_reg[7]/NET0131  , \u2_R5_reg[8]/NET0131  , \u2_R5_reg[9]/NET0131  , \u2_R6_reg[10]/NET0131  , \u2_R6_reg[11]/NET0131  , \u2_R6_reg[12]/NET0131  , \u2_R6_reg[13]/NET0131  , \u2_R6_reg[14]/NET0131  , \u2_R6_reg[15]/NET0131  , \u2_R6_reg[16]/NET0131  , \u2_R6_reg[17]/NET0131  , \u2_R6_reg[18]/NET0131  , \u2_R6_reg[19]/NET0131  , \u2_R6_reg[1]/NET0131  , \u2_R6_reg[20]/NET0131  , \u2_R6_reg[21]/NET0131  , \u2_R6_reg[22]/NET0131  , \u2_R6_reg[23]/NET0131  , \u2_R6_reg[24]/NET0131  , \u2_R6_reg[25]/NET0131  , \u2_R6_reg[26]/NET0131  , \u2_R6_reg[27]/NET0131  , \u2_R6_reg[28]/NET0131  , \u2_R6_reg[29]/NET0131  , \u2_R6_reg[2]/NET0131  , \u2_R6_reg[30]/NET0131  , \u2_R6_reg[31]/P0001  , \u2_R6_reg[32]/NET0131  , \u2_R6_reg[3]/NET0131  , \u2_R6_reg[4]/NET0131  , \u2_R6_reg[5]/NET0131  , \u2_R6_reg[6]/NET0131  , \u2_R6_reg[7]/NET0131  , \u2_R6_reg[8]/NET0131  , \u2_R6_reg[9]/NET0131  , \u2_R7_reg[10]/NET0131  , \u2_R7_reg[11]/NET0131  , \u2_R7_reg[12]/NET0131  , \u2_R7_reg[13]/NET0131  , \u2_R7_reg[14]/NET0131  , \u2_R7_reg[15]/NET0131  , \u2_R7_reg[16]/NET0131  , \u2_R7_reg[17]/NET0131  , \u2_R7_reg[18]/NET0131  , \u2_R7_reg[19]/NET0131  , \u2_R7_reg[1]/NET0131  , \u2_R7_reg[20]/NET0131  , \u2_R7_reg[21]/NET0131  , \u2_R7_reg[22]/NET0131  , \u2_R7_reg[23]/NET0131  , \u2_R7_reg[24]/NET0131  , \u2_R7_reg[25]/NET0131  , \u2_R7_reg[26]/NET0131  , \u2_R7_reg[27]/NET0131  , \u2_R7_reg[28]/NET0131  , \u2_R7_reg[29]/NET0131  , \u2_R7_reg[2]/NET0131  , \u2_R7_reg[30]/NET0131  , \u2_R7_reg[31]/P0001  , \u2_R7_reg[32]/NET0131  , \u2_R7_reg[3]/NET0131  , \u2_R7_reg[4]/NET0131  , \u2_R7_reg[5]/NET0131  , \u2_R7_reg[6]/NET0131  , \u2_R7_reg[7]/NET0131  , \u2_R7_reg[8]/NET0131  , \u2_R7_reg[9]/NET0131  , \u2_R8_reg[10]/NET0131  , \u2_R8_reg[11]/NET0131  , \u2_R8_reg[12]/NET0131  , \u2_R8_reg[13]/NET0131  , \u2_R8_reg[14]/NET0131  , \u2_R8_reg[15]/NET0131  , \u2_R8_reg[16]/NET0131  , \u2_R8_reg[17]/NET0131  , \u2_R8_reg[18]/NET0131  , \u2_R8_reg[19]/NET0131  , \u2_R8_reg[1]/NET0131  , \u2_R8_reg[20]/NET0131  , \u2_R8_reg[21]/NET0131  , \u2_R8_reg[22]/NET0131  , \u2_R8_reg[23]/NET0131  , \u2_R8_reg[24]/NET0131  , \u2_R8_reg[25]/NET0131  , \u2_R8_reg[26]/NET0131  , \u2_R8_reg[27]/NET0131  , \u2_R8_reg[28]/NET0131  , \u2_R8_reg[29]/NET0131  , \u2_R8_reg[2]/NET0131  , \u2_R8_reg[30]/NET0131  , \u2_R8_reg[31]/P0001  , \u2_R8_reg[32]/NET0131  , \u2_R8_reg[3]/NET0131  , \u2_R8_reg[4]/NET0131  , \u2_R8_reg[5]/NET0131  , \u2_R8_reg[6]/NET0131  , \u2_R8_reg[7]/NET0131  , \u2_R8_reg[8]/NET0131  , \u2_R8_reg[9]/NET0131  , \u2_R9_reg[10]/NET0131  , \u2_R9_reg[11]/NET0131  , \u2_R9_reg[12]/NET0131  , \u2_R9_reg[13]/NET0131  , \u2_R9_reg[14]/NET0131  , \u2_R9_reg[15]/NET0131  , \u2_R9_reg[16]/NET0131  , \u2_R9_reg[17]/NET0131  , \u2_R9_reg[18]/NET0131  , \u2_R9_reg[19]/NET0131  , \u2_R9_reg[1]/NET0131  , \u2_R9_reg[20]/NET0131  , \u2_R9_reg[21]/NET0131  , \u2_R9_reg[22]/NET0131  , \u2_R9_reg[23]/NET0131  , \u2_R9_reg[24]/NET0131  , \u2_R9_reg[25]/NET0131  , \u2_R9_reg[26]/NET0131  , \u2_R9_reg[27]/NET0131  , \u2_R9_reg[28]/NET0131  , \u2_R9_reg[29]/NET0131  , \u2_R9_reg[2]/NET0131  , \u2_R9_reg[30]/NET0131  , \u2_R9_reg[31]/P0001  , \u2_R9_reg[32]/NET0131  , \u2_R9_reg[3]/NET0131  , \u2_R9_reg[4]/NET0131  , \u2_R9_reg[5]/NET0131  , \u2_R9_reg[6]/NET0131  , \u2_R9_reg[7]/NET0131  , \u2_R9_reg[8]/NET0131  , \u2_R9_reg[9]/NET0131  , \u2_desIn_r_reg[0]/NET0131  , \u2_desIn_r_reg[10]/P0001  , \u2_desIn_r_reg[11]/NET0131  , \u2_desIn_r_reg[12]/NET0131  , \u2_desIn_r_reg[13]/NET0131  , \u2_desIn_r_reg[14]/NET0131  , \u2_desIn_r_reg[15]/NET0131  , \u2_desIn_r_reg[16]/NET0131  , \u2_desIn_r_reg[17]/NET0131  , \u2_desIn_r_reg[18]/NET0131  , \u2_desIn_r_reg[19]/NET0131  , \u2_desIn_r_reg[1]/NET0131  , \u2_desIn_r_reg[20]/NET0131  , \u2_desIn_r_reg[21]/NET0131  , \u2_desIn_r_reg[22]/NET0131  , \u2_desIn_r_reg[23]/NET0131  , \u2_desIn_r_reg[24]/NET0131  , \u2_desIn_r_reg[25]/NET0131  , \u2_desIn_r_reg[26]/NET0131  , \u2_desIn_r_reg[27]/NET0131  , \u2_desIn_r_reg[28]/NET0131  , \u2_desIn_r_reg[29]/NET0131  , \u2_desIn_r_reg[2]/NET0131  , \u2_desIn_r_reg[30]/NET0131  , \u2_desIn_r_reg[31]/NET0131  , \u2_desIn_r_reg[32]/NET0131  , \u2_desIn_r_reg[33]/NET0131  , \u2_desIn_r_reg[34]/NET0131  , \u2_desIn_r_reg[35]/NET0131  , \u2_desIn_r_reg[36]/NET0131  , \u2_desIn_r_reg[37]/NET0131  , \u2_desIn_r_reg[38]/NET0131  , \u2_desIn_r_reg[39]/NET0131  , \u2_desIn_r_reg[3]/NET0131  , \u2_desIn_r_reg[40]/NET0131  , \u2_desIn_r_reg[41]/NET0131  , \u2_desIn_r_reg[42]/NET0131  , \u2_desIn_r_reg[43]/NET0131  , \u2_desIn_r_reg[44]/NET0131  , \u2_desIn_r_reg[45]/NET0131  , \u2_desIn_r_reg[46]/NET0131  , \u2_desIn_r_reg[47]/NET0131  , \u2_desIn_r_reg[48]/NET0131  , \u2_desIn_r_reg[49]/NET0131  , \u2_desIn_r_reg[4]/NET0131  , \u2_desIn_r_reg[50]/NET0131  , \u2_desIn_r_reg[51]/NET0131  , \u2_desIn_r_reg[52]/NET0131  , \u2_desIn_r_reg[53]/NET0131  , \u2_desIn_r_reg[54]/NET0131  , \u2_desIn_r_reg[55]/NET0131  , \u2_desIn_r_reg[56]/NET0131  , \u2_desIn_r_reg[57]/NET0131  , \u2_desIn_r_reg[58]/NET0131  , \u2_desIn_r_reg[59]/NET0131  , \u2_desIn_r_reg[5]/NET0131  , \u2_desIn_r_reg[60]/NET0131  , \u2_desIn_r_reg[61]/NET0131  , \u2_desIn_r_reg[62]/NET0131  , \u2_desIn_r_reg[63]/NET0131  , \u2_desIn_r_reg[6]/NET0131  , \u2_desIn_r_reg[7]/NET0131  , \u2_desIn_r_reg[8]/NET0131  , \u2_desIn_r_reg[9]/NET0131  , \u2_key_r_reg[0]/NET0131  , \u2_key_r_reg[10]/NET0131  , \u2_key_r_reg[11]/NET0131  , \u2_key_r_reg[12]/NET0131  , \u2_key_r_reg[13]/NET0131  , \u2_key_r_reg[14]/NET0131  , \u2_key_r_reg[15]/NET0131  , \u2_key_r_reg[16]/NET0131  , \u2_key_r_reg[17]/NET0131  , \u2_key_r_reg[18]/NET0131  , \u2_key_r_reg[19]/NET0131  , \u2_key_r_reg[1]/NET0131  , \u2_key_r_reg[20]/NET0131  , \u2_key_r_reg[21]/NET0131  , \u2_key_r_reg[22]/NET0131  , \u2_key_r_reg[23]/NET0131  , \u2_key_r_reg[24]/NET0131  , \u2_key_r_reg[25]/NET0131  , \u2_key_r_reg[26]/NET0131  , \u2_key_r_reg[27]/NET0131  , \u2_key_r_reg[28]/NET0131  , \u2_key_r_reg[29]/NET0131  , \u2_key_r_reg[2]/NET0131  , \u2_key_r_reg[30]/NET0131  , \u2_key_r_reg[31]/NET0131  , \u2_key_r_reg[32]/NET0131  , \u2_key_r_reg[33]/NET0131  , \u2_key_r_reg[34]/NET0131  , \u2_key_r_reg[35]/P0001  , \u2_key_r_reg[36]/NET0131  , \u2_key_r_reg[37]/NET0131  , \u2_key_r_reg[38]/NET0131  , \u2_key_r_reg[39]/P0001  , \u2_key_r_reg[3]/NET0131  , \u2_key_r_reg[40]/NET0131  , \u2_key_r_reg[41]/NET0131  , \u2_key_r_reg[42]/P0001  , \u2_key_r_reg[43]/NET0131  , \u2_key_r_reg[44]/NET0131  , \u2_key_r_reg[45]/NET0131  , \u2_key_r_reg[46]/NET0131  , \u2_key_r_reg[47]/NET0131  , \u2_key_r_reg[48]/NET0131  , \u2_key_r_reg[49]/NET0131  , \u2_key_r_reg[4]/NET0131  , \u2_key_r_reg[50]/NET0131  , \u2_key_r_reg[51]/NET0131  , \u2_key_r_reg[52]/NET0131  , \u2_key_r_reg[53]/NET0131  , \u2_key_r_reg[54]/NET0131  , \u2_key_r_reg[55]/NET0131  , \u2_key_r_reg[5]/NET0131  , \u2_key_r_reg[6]/NET0131  , \u2_key_r_reg[7]/NET0131  , \u2_key_r_reg[8]/NET0131  , \u2_key_r_reg[9]/NET0131  , \u2_uk_K_r0_reg[0]/NET0131  , \u2_uk_K_r0_reg[10]/NET0131  , \u2_uk_K_r0_reg[11]/NET0131  , \u2_uk_K_r0_reg[12]/NET0131  , \u2_uk_K_r0_reg[13]/NET0131  , \u2_uk_K_r0_reg[14]/NET0131  , \u2_uk_K_r0_reg[15]/NET0131  , \u2_uk_K_r0_reg[16]/NET0131  , \u2_uk_K_r0_reg[17]/NET0131  , \u2_uk_K_r0_reg[18]/NET0131  , \u2_uk_K_r0_reg[19]/NET0131  , \u2_uk_K_r0_reg[20]/NET0131  , \u2_uk_K_r0_reg[21]/NET0131  , \u2_uk_K_r0_reg[22]/NET0131  , \u2_uk_K_r0_reg[23]/NET0131  , \u2_uk_K_r0_reg[24]/P0001  , \u2_uk_K_r0_reg[25]/P0001  , \u2_uk_K_r0_reg[26]/NET0131  , \u2_uk_K_r0_reg[27]/NET0131  , \u2_uk_K_r0_reg[28]/NET0131  , \u2_uk_K_r0_reg[29]/NET0131  , \u2_uk_K_r0_reg[2]/NET0131  , \u2_uk_K_r0_reg[30]/NET0131  , \u2_uk_K_r0_reg[31]/NET0131  , \u2_uk_K_r0_reg[32]/NET0131  , \u2_uk_K_r0_reg[33]/NET0131  , \u2_uk_K_r0_reg[34]/NET0131  , \u2_uk_K_r0_reg[35]/NET0131  , \u2_uk_K_r0_reg[36]/NET0131  , \u2_uk_K_r0_reg[37]/NET0131  , \u2_uk_K_r0_reg[38]/NET0131  , \u2_uk_K_r0_reg[39]/NET0131  , \u2_uk_K_r0_reg[3]/NET0131  , \u2_uk_K_r0_reg[40]/NET0131  , \u2_uk_K_r0_reg[41]/NET0131  , \u2_uk_K_r0_reg[42]/NET0131  , \u2_uk_K_r0_reg[43]/NET0131  , \u2_uk_K_r0_reg[44]/NET0131  , \u2_uk_K_r0_reg[45]/NET0131  , \u2_uk_K_r0_reg[46]/NET0131  , \u2_uk_K_r0_reg[47]/NET0131  , \u2_uk_K_r0_reg[48]/NET0131  , \u2_uk_K_r0_reg[49]/NET0131  , \u2_uk_K_r0_reg[4]/NET0131  , \u2_uk_K_r0_reg[50]/NET0131  , \u2_uk_K_r0_reg[51]/NET0131  , \u2_uk_K_r0_reg[52]/P0001  , \u2_uk_K_r0_reg[54]/NET0131  , \u2_uk_K_r0_reg[55]/NET0131  , \u2_uk_K_r0_reg[5]/NET0131  , \u2_uk_K_r0_reg[6]/NET0131  , \u2_uk_K_r0_reg[7]/NET0131  , \u2_uk_K_r0_reg[8]/NET0131  , \u2_uk_K_r0_reg[9]/NET0131  , \u2_uk_K_r10_reg[0]/NET0131  , \u2_uk_K_r10_reg[10]/NET0131  , \u2_uk_K_r10_reg[11]/NET0131  , \u2_uk_K_r10_reg[12]/NET0131  , \u2_uk_K_r10_reg[14]/NET0131  , \u2_uk_K_r10_reg[15]/NET0131  , \u2_uk_K_r10_reg[16]/NET0131  , \u2_uk_K_r10_reg[17]/NET0131  , \u2_uk_K_r10_reg[18]/NET0131  , \u2_uk_K_r10_reg[19]/NET0131  , \u2_uk_K_r10_reg[1]/NET0131  , \u2_uk_K_r10_reg[20]/NET0131  , \u2_uk_K_r10_reg[21]/NET0131  , \u2_uk_K_r10_reg[22]/NET0131  , \u2_uk_K_r10_reg[23]/NET0131  , \u2_uk_K_r10_reg[24]/NET0131  , \u2_uk_K_r10_reg[25]/NET0131  , \u2_uk_K_r10_reg[26]/NET0131  , \u2_uk_K_r10_reg[27]/NET0131  , \u2_uk_K_r10_reg[28]/NET0131  , \u2_uk_K_r10_reg[29]/NET0131  , \u2_uk_K_r10_reg[2]/NET0131  , \u2_uk_K_r10_reg[30]/NET0131  , \u2_uk_K_r10_reg[31]/NET0131  , \u2_uk_K_r10_reg[32]/NET0131  , \u2_uk_K_r10_reg[33]/NET0131  , \u2_uk_K_r10_reg[34]/NET0131  , \u2_uk_K_r10_reg[35]/NET0131  , \u2_uk_K_r10_reg[36]/NET0131  , \u2_uk_K_r10_reg[37]/NET0131  , \u2_uk_K_r10_reg[38]/NET0131  , \u2_uk_K_r10_reg[39]/NET0131  , \u2_uk_K_r10_reg[3]/NET0131  , \u2_uk_K_r10_reg[40]/NET0131  , \u2_uk_K_r10_reg[41]/NET0131  , \u2_uk_K_r10_reg[42]/NET0131  , \u2_uk_K_r10_reg[43]/NET0131  , \u2_uk_K_r10_reg[44]/NET0131  , \u2_uk_K_r10_reg[45]/P0001  , \u2_uk_K_r10_reg[46]/NET0131  , \u2_uk_K_r10_reg[47]/NET0131  , \u2_uk_K_r10_reg[48]/NET0131  , \u2_uk_K_r10_reg[49]/NET0131  , \u2_uk_K_r10_reg[4]/NET0131  , \u2_uk_K_r10_reg[50]/NET0131  , \u2_uk_K_r10_reg[51]/NET0131  , \u2_uk_K_r10_reg[52]/NET0131  , \u2_uk_K_r10_reg[53]/NET0131  , \u2_uk_K_r10_reg[54]/NET0131  , \u2_uk_K_r10_reg[55]/NET0131  , \u2_uk_K_r10_reg[5]/NET0131  , \u2_uk_K_r10_reg[6]/NET0131  , \u2_uk_K_r10_reg[7]/NET0131  , \u2_uk_K_r10_reg[8]/NET0131  , \u2_uk_K_r10_reg[9]/NET0131  , \u2_uk_K_r11_reg[0]/NET0131  , \u2_uk_K_r11_reg[10]/NET0131  , \u2_uk_K_r11_reg[11]/NET0131  , \u2_uk_K_r11_reg[12]/NET0131  , \u2_uk_K_r11_reg[13]/NET0131  , \u2_uk_K_r11_reg[14]/NET0131  , \u2_uk_K_r11_reg[15]/NET0131  , \u2_uk_K_r11_reg[16]/NET0131  , \u2_uk_K_r11_reg[17]/NET0131  , \u2_uk_K_r11_reg[18]/NET0131  , \u2_uk_K_r11_reg[19]/NET0131  , \u2_uk_K_r11_reg[1]/NET0131  , \u2_uk_K_r11_reg[20]/NET0131  , \u2_uk_K_r11_reg[21]/NET0131  , \u2_uk_K_r11_reg[22]/NET0131  , \u2_uk_K_r11_reg[23]/NET0131  , \u2_uk_K_r11_reg[24]/NET0131  , \u2_uk_K_r11_reg[25]/NET0131  , \u2_uk_K_r11_reg[26]/NET0131  , \u2_uk_K_r11_reg[27]/NET0131  , \u2_uk_K_r11_reg[28]/NET0131  , \u2_uk_K_r11_reg[29]/NET0131  , \u2_uk_K_r11_reg[2]/NET0131  , \u2_uk_K_r11_reg[31]/NET0131  , \u2_uk_K_r11_reg[32]/NET0131  , \u2_uk_K_r11_reg[33]/NET0131  , \u2_uk_K_r11_reg[34]/NET0131  , \u2_uk_K_r11_reg[35]/NET0131  , \u2_uk_K_r11_reg[36]/NET0131  , \u2_uk_K_r11_reg[37]/NET0131  , \u2_uk_K_r11_reg[38]/NET0131  , \u2_uk_K_r11_reg[39]/NET0131  , \u2_uk_K_r11_reg[3]/NET0131  , \u2_uk_K_r11_reg[40]/NET0131  , \u2_uk_K_r11_reg[41]/NET0131  , \u2_uk_K_r11_reg[42]/NET0131  , \u2_uk_K_r11_reg[43]/NET0131  , \u2_uk_K_r11_reg[44]/NET0131  , \u2_uk_K_r11_reg[45]/NET0131  , \u2_uk_K_r11_reg[46]/NET0131  , \u2_uk_K_r11_reg[47]/NET0131  , \u2_uk_K_r11_reg[48]/NET0131  , \u2_uk_K_r11_reg[49]/NET0131  , \u2_uk_K_r11_reg[4]/NET0131  , \u2_uk_K_r11_reg[50]/NET0131  , \u2_uk_K_r11_reg[51]/NET0131  , \u2_uk_K_r11_reg[52]/NET0131  , \u2_uk_K_r11_reg[53]/P0001  , \u2_uk_K_r11_reg[54]/NET0131  , \u2_uk_K_r11_reg[55]/NET0131  , \u2_uk_K_r11_reg[5]/NET0131  , \u2_uk_K_r11_reg[6]/NET0131  , \u2_uk_K_r11_reg[7]/NET0131  , \u2_uk_K_r11_reg[8]/NET0131  , \u2_uk_K_r11_reg[9]/NET0131  , \u2_uk_K_r12_reg[0]/NET0131  , \u2_uk_K_r12_reg[10]/P0001  , \u2_uk_K_r12_reg[11]/NET0131  , \u2_uk_K_r12_reg[12]/NET0131  , \u2_uk_K_r12_reg[13]/NET0131  , \u2_uk_K_r12_reg[14]/NET0131  , \u2_uk_K_r12_reg[15]/NET0131  , \u2_uk_K_r12_reg[16]/NET0131  , \u2_uk_K_r12_reg[17]/NET0131  , \u2_uk_K_r12_reg[18]/NET0131  , \u2_uk_K_r12_reg[19]/NET0131  , \u2_uk_K_r12_reg[1]/NET0131  , \u2_uk_K_r12_reg[20]/NET0131  , \u2_uk_K_r12_reg[21]/NET0131  , \u2_uk_K_r12_reg[22]/NET0131  , \u2_uk_K_r12_reg[23]/NET0131  , \u2_uk_K_r12_reg[24]/NET0131  , \u2_uk_K_r12_reg[25]/NET0131  , \u2_uk_K_r12_reg[26]/NET0131  , \u2_uk_K_r12_reg[27]/NET0131  , \u2_uk_K_r12_reg[28]/NET0131  , \u2_uk_K_r12_reg[29]/NET0131  , \u2_uk_K_r12_reg[2]/NET0131  , \u2_uk_K_r12_reg[30]/NET0131  , \u2_uk_K_r12_reg[31]/NET0131  , \u2_uk_K_r12_reg[32]/NET0131  , \u2_uk_K_r12_reg[33]/NET0131  , \u2_uk_K_r12_reg[34]/NET0131  , \u2_uk_K_r12_reg[35]/NET0131  , \u2_uk_K_r12_reg[36]/NET0131  , \u2_uk_K_r12_reg[37]/NET0131  , \u2_uk_K_r12_reg[38]/NET0131  , \u2_uk_K_r12_reg[3]/NET0131  , \u2_uk_K_r12_reg[40]/NET0131  , \u2_uk_K_r12_reg[41]/NET0131  , \u2_uk_K_r12_reg[42]/NET0131  , \u2_uk_K_r12_reg[43]/NET0131  , \u2_uk_K_r12_reg[44]/P0001  , \u2_uk_K_r12_reg[45]/NET0131  , \u2_uk_K_r12_reg[46]/NET0131  , \u2_uk_K_r12_reg[47]/NET0131  , \u2_uk_K_r12_reg[48]/NET0131  , \u2_uk_K_r12_reg[49]/NET0131  , \u2_uk_K_r12_reg[4]/NET0131  , \u2_uk_K_r12_reg[50]/NET0131  , \u2_uk_K_r12_reg[51]/NET0131  , \u2_uk_K_r12_reg[52]/NET0131  , \u2_uk_K_r12_reg[53]/NET0131  , \u2_uk_K_r12_reg[54]/NET0131  , \u2_uk_K_r12_reg[55]/NET0131  , \u2_uk_K_r12_reg[5]/NET0131  , \u2_uk_K_r12_reg[6]/NET0131  , \u2_uk_K_r12_reg[7]/P0001  , \u2_uk_K_r12_reg[8]/NET0131  , \u2_uk_K_r12_reg[9]/NET0131  , \u2_uk_K_r13_reg[0]/NET0131  , \u2_uk_K_r13_reg[10]/NET0131  , \u2_uk_K_r13_reg[11]/NET0131  , \u2_uk_K_r13_reg[12]/NET0131  , \u2_uk_K_r13_reg[13]/NET0131  , \u2_uk_K_r13_reg[14]/NET0131  , \u2_uk_K_r13_reg[15]/NET0131  , \u2_uk_K_r13_reg[16]/NET0131  , \u2_uk_K_r13_reg[17]/NET0131  , \u2_uk_K_r13_reg[18]/NET0131  , \u2_uk_K_r13_reg[19]/NET0131  , \u2_uk_K_r13_reg[20]/NET0131  , \u2_uk_K_r13_reg[21]/NET0131  , \u2_uk_K_r13_reg[22]/NET0131  , \u2_uk_K_r13_reg[23]/NET0131  , \u2_uk_K_r13_reg[24]/NET0131  , \u2_uk_K_r13_reg[25]/P0001  , \u2_uk_K_r13_reg[26]/NET0131  , \u2_uk_K_r13_reg[27]/NET0131  , \u2_uk_K_r13_reg[28]/NET0131  , \u2_uk_K_r13_reg[29]/NET0131  , \u2_uk_K_r13_reg[2]/NET0131  , \u2_uk_K_r13_reg[30]/NET0131  , \u2_uk_K_r13_reg[31]/NET0131  , \u2_uk_K_r13_reg[32]/NET0131  , \u2_uk_K_r13_reg[33]/NET0131  , \u2_uk_K_r13_reg[34]/NET0131  , \u2_uk_K_r13_reg[35]/NET0131  , \u2_uk_K_r13_reg[36]/NET0131  , \u2_uk_K_r13_reg[37]/NET0131  , \u2_uk_K_r13_reg[38]/NET0131  , \u2_uk_K_r13_reg[39]/NET0131  , \u2_uk_K_r13_reg[3]/NET0131  , \u2_uk_K_r13_reg[40]/NET0131  , \u2_uk_K_r13_reg[41]/NET0131  , \u2_uk_K_r13_reg[42]/NET0131  , \u2_uk_K_r13_reg[43]/NET0131  , \u2_uk_K_r13_reg[44]/NET0131  , \u2_uk_K_r13_reg[45]/NET0131  , \u2_uk_K_r13_reg[46]/NET0131  , \u2_uk_K_r13_reg[47]/NET0131  , \u2_uk_K_r13_reg[48]/NET0131  , \u2_uk_K_r13_reg[49]/NET0131  , \u2_uk_K_r13_reg[4]/NET0131  , \u2_uk_K_r13_reg[50]/NET0131  , \u2_uk_K_r13_reg[51]/NET0131  , \u2_uk_K_r13_reg[52]/NET0131  , \u2_uk_K_r13_reg[54]/NET0131  , \u2_uk_K_r13_reg[55]/NET0131  , \u2_uk_K_r13_reg[5]/NET0131  , \u2_uk_K_r13_reg[6]/NET0131  , \u2_uk_K_r13_reg[7]/NET0131  , \u2_uk_K_r13_reg[8]/NET0131  , \u2_uk_K_r13_reg[9]/NET0131  , \u2_uk_K_r14_reg[0]/NET0131  , \u2_uk_K_r14_reg[10]/P0001  , \u2_uk_K_r14_reg[11]/NET0131  , \u2_uk_K_r14_reg[12]/NET0131  , \u2_uk_K_r14_reg[13]/NET0131  , \u2_uk_K_r14_reg[14]/NET0131  , \u2_uk_K_r14_reg[15]/NET0131  , \u2_uk_K_r14_reg[16]/NET0131  , \u2_uk_K_r14_reg[17]/NET0131  , \u2_uk_K_r14_reg[18]/NET0131  , \u2_uk_K_r14_reg[19]/NET0131  , \u2_uk_K_r14_reg[1]/NET0131  , \u2_uk_K_r14_reg[20]/NET0131  , \u2_uk_K_r14_reg[21]/NET0131  , \u2_uk_K_r14_reg[22]/NET0131  , \u2_uk_K_r14_reg[23]/NET0131  , \u2_uk_K_r14_reg[24]/NET0131  , \u2_uk_K_r14_reg[25]/NET0131  , \u2_uk_K_r14_reg[26]/NET0131  , \u2_uk_K_r14_reg[27]/NET0131  , \u2_uk_K_r14_reg[28]/NET0131  , \u2_uk_K_r14_reg[29]/NET0131  , \u2_uk_K_r14_reg[2]/NET0131  , \u2_uk_K_r14_reg[30]/NET0131  , \u2_uk_K_r14_reg[31]/NET0131  , \u2_uk_K_r14_reg[32]/NET0131  , \u2_uk_K_r14_reg[33]/NET0131  , \u2_uk_K_r14_reg[34]/NET0131  , \u2_uk_K_r14_reg[35]/P0001  , \u2_uk_K_r14_reg[36]/NET0131  , \u2_uk_K_r14_reg[37]/NET0131  , \u2_uk_K_r14_reg[38]/NET0131  , \u2_uk_K_r14_reg[39]/P0001  , \u2_uk_K_r14_reg[3]/NET0131  , \u2_uk_K_r14_reg[40]/NET0131  , \u2_uk_K_r14_reg[41]/NET0131  , \u2_uk_K_r14_reg[42]/P0001  , \u2_uk_K_r14_reg[43]/NET0131  , \u2_uk_K_r14_reg[44]/NET0131  , \u2_uk_K_r14_reg[45]/NET0131  , \u2_uk_K_r14_reg[46]/NET0131  , \u2_uk_K_r14_reg[47]/NET0131  , \u2_uk_K_r14_reg[48]/NET0131  , \u2_uk_K_r14_reg[49]/P0001  , \u2_uk_K_r14_reg[4]/NET0131  , \u2_uk_K_r14_reg[50]/NET0131  , \u2_uk_K_r14_reg[51]/NET0131  , \u2_uk_K_r14_reg[52]/NET0131  , \u2_uk_K_r14_reg[53]/NET0131  , \u2_uk_K_r14_reg[54]/NET0131  , \u2_uk_K_r14_reg[55]/NET0131  , \u2_uk_K_r14_reg[5]/NET0131  , \u2_uk_K_r14_reg[6]/NET0131  , \u2_uk_K_r14_reg[7]/NET0131  , \u2_uk_K_r14_reg[8]/NET0131  , \u2_uk_K_r14_reg[9]/NET0131  , \u2_uk_K_r1_reg[0]/NET0131  , \u2_uk_K_r1_reg[10]/P0001  , \u2_uk_K_r1_reg[11]/NET0131  , \u2_uk_K_r1_reg[12]/NET0131  , \u2_uk_K_r1_reg[13]/NET0131  , \u2_uk_K_r1_reg[14]/NET0131  , \u2_uk_K_r1_reg[15]/NET0131  , \u2_uk_K_r1_reg[16]/NET0131  , \u2_uk_K_r1_reg[17]/NET0131  , \u2_uk_K_r1_reg[18]/NET0131  , \u2_uk_K_r1_reg[19]/NET0131  , \u2_uk_K_r1_reg[1]/NET0131  , \u2_uk_K_r1_reg[20]/NET0131  , \u2_uk_K_r1_reg[21]/NET0131  , \u2_uk_K_r1_reg[22]/NET0131  , \u2_uk_K_r1_reg[23]/NET0131  , \u2_uk_K_r1_reg[24]/NET0131  , \u2_uk_K_r1_reg[25]/NET0131  , \u2_uk_K_r1_reg[26]/NET0131  , \u2_uk_K_r1_reg[27]/NET0131  , \u2_uk_K_r1_reg[28]/NET0131  , \u2_uk_K_r1_reg[29]/NET0131  , \u2_uk_K_r1_reg[2]/NET0131  , \u2_uk_K_r1_reg[30]/NET0131  , \u2_uk_K_r1_reg[31]/NET0131  , \u2_uk_K_r1_reg[32]/NET0131  , \u2_uk_K_r1_reg[33]/NET0131  , \u2_uk_K_r1_reg[34]/NET0131  , \u2_uk_K_r1_reg[35]/NET0131  , \u2_uk_K_r1_reg[36]/NET0131  , \u2_uk_K_r1_reg[37]/NET0131  , \u2_uk_K_r1_reg[38]/NET0131  , \u2_uk_K_r1_reg[3]/NET0131  , \u2_uk_K_r1_reg[40]/NET0131  , \u2_uk_K_r1_reg[41]/NET0131  , \u2_uk_K_r1_reg[42]/NET0131  , \u2_uk_K_r1_reg[43]/NET0131  , \u2_uk_K_r1_reg[44]/P0001  , \u2_uk_K_r1_reg[45]/NET0131  , \u2_uk_K_r1_reg[46]/NET0131  , \u2_uk_K_r1_reg[47]/NET0131  , \u2_uk_K_r1_reg[48]/NET0131  , \u2_uk_K_r1_reg[49]/NET0131  , \u2_uk_K_r1_reg[4]/NET0131  , \u2_uk_K_r1_reg[50]/NET0131  , \u2_uk_K_r1_reg[51]/NET0131  , \u2_uk_K_r1_reg[52]/NET0131  , \u2_uk_K_r1_reg[53]/NET0131  , \u2_uk_K_r1_reg[54]/NET0131  , \u2_uk_K_r1_reg[55]/NET0131  , \u2_uk_K_r1_reg[5]/NET0131  , \u2_uk_K_r1_reg[6]/NET0131  , \u2_uk_K_r1_reg[7]/P0001  , \u2_uk_K_r1_reg[8]/NET0131  , \u2_uk_K_r1_reg[9]/NET0131  , \u2_uk_K_r2_reg[0]/NET0131  , \u2_uk_K_r2_reg[10]/NET0131  , \u2_uk_K_r2_reg[11]/NET0131  , \u2_uk_K_r2_reg[12]/NET0131  , \u2_uk_K_r2_reg[13]/NET0131  , \u2_uk_K_r2_reg[14]/NET0131  , \u2_uk_K_r2_reg[15]/NET0131  , \u2_uk_K_r2_reg[16]/NET0131  , \u2_uk_K_r2_reg[17]/NET0131  , \u2_uk_K_r2_reg[18]/NET0131  , \u2_uk_K_r2_reg[19]/NET0131  , \u2_uk_K_r2_reg[1]/NET0131  , \u2_uk_K_r2_reg[20]/NET0131  , \u2_uk_K_r2_reg[21]/NET0131  , \u2_uk_K_r2_reg[22]/NET0131  , \u2_uk_K_r2_reg[23]/NET0131  , \u2_uk_K_r2_reg[24]/NET0131  , \u2_uk_K_r2_reg[25]/NET0131  , \u2_uk_K_r2_reg[26]/NET0131  , \u2_uk_K_r2_reg[27]/NET0131  , \u2_uk_K_r2_reg[28]/NET0131  , \u2_uk_K_r2_reg[29]/NET0131  , \u2_uk_K_r2_reg[2]/NET0131  , \u2_uk_K_r2_reg[31]/NET0131  , \u2_uk_K_r2_reg[32]/NET0131  , \u2_uk_K_r2_reg[33]/NET0131  , \u2_uk_K_r2_reg[34]/NET0131  , \u2_uk_K_r2_reg[35]/NET0131  , \u2_uk_K_r2_reg[36]/NET0131  , \u2_uk_K_r2_reg[37]/NET0131  , \u2_uk_K_r2_reg[38]/NET0131  , \u2_uk_K_r2_reg[39]/NET0131  , \u2_uk_K_r2_reg[3]/NET0131  , \u2_uk_K_r2_reg[40]/NET0131  , \u2_uk_K_r2_reg[41]/NET0131  , \u2_uk_K_r2_reg[42]/NET0131  , \u2_uk_K_r2_reg[43]/NET0131  , \u2_uk_K_r2_reg[44]/NET0131  , \u2_uk_K_r2_reg[45]/NET0131  , \u2_uk_K_r2_reg[46]/NET0131  , \u2_uk_K_r2_reg[47]/NET0131  , \u2_uk_K_r2_reg[48]/NET0131  , \u2_uk_K_r2_reg[49]/NET0131  , \u2_uk_K_r2_reg[4]/NET0131  , \u2_uk_K_r2_reg[50]/NET0131  , \u2_uk_K_r2_reg[51]/NET0131  , \u2_uk_K_r2_reg[52]/NET0131  , \u2_uk_K_r2_reg[53]/P0001  , \u2_uk_K_r2_reg[54]/NET0131  , \u2_uk_K_r2_reg[55]/NET0131  , \u2_uk_K_r2_reg[5]/NET0131  , \u2_uk_K_r2_reg[6]/NET0131  , \u2_uk_K_r2_reg[7]/NET0131  , \u2_uk_K_r2_reg[8]/NET0131  , \u2_uk_K_r2_reg[9]/NET0131  , \u2_uk_K_r3_reg[0]/NET0131  , \u2_uk_K_r3_reg[10]/NET0131  , \u2_uk_K_r3_reg[11]/NET0131  , \u2_uk_K_r3_reg[12]/NET0131  , \u2_uk_K_r3_reg[14]/NET0131  , \u2_uk_K_r3_reg[15]/NET0131  , \u2_uk_K_r3_reg[16]/NET0131  , \u2_uk_K_r3_reg[17]/NET0131  , \u2_uk_K_r3_reg[18]/NET0131  , \u2_uk_K_r3_reg[19]/NET0131  , \u2_uk_K_r3_reg[1]/NET0131  , \u2_uk_K_r3_reg[20]/NET0131  , \u2_uk_K_r3_reg[21]/NET0131  , \u2_uk_K_r3_reg[22]/NET0131  , \u2_uk_K_r3_reg[23]/NET0131  , \u2_uk_K_r3_reg[24]/NET0131  , \u2_uk_K_r3_reg[25]/NET0131  , \u2_uk_K_r3_reg[26]/NET0131  , \u2_uk_K_r3_reg[27]/NET0131  , \u2_uk_K_r3_reg[28]/NET0131  , \u2_uk_K_r3_reg[29]/NET0131  , \u2_uk_K_r3_reg[2]/NET0131  , \u2_uk_K_r3_reg[30]/NET0131  , \u2_uk_K_r3_reg[31]/NET0131  , \u2_uk_K_r3_reg[32]/NET0131  , \u2_uk_K_r3_reg[33]/NET0131  , \u2_uk_K_r3_reg[34]/NET0131  , \u2_uk_K_r3_reg[35]/NET0131  , \u2_uk_K_r3_reg[36]/NET0131  , \u2_uk_K_r3_reg[37]/NET0131  , \u2_uk_K_r3_reg[38]/NET0131  , \u2_uk_K_r3_reg[39]/NET0131  , \u2_uk_K_r3_reg[3]/NET0131  , \u2_uk_K_r3_reg[40]/NET0131  , \u2_uk_K_r3_reg[41]/NET0131  , \u2_uk_K_r3_reg[42]/NET0131  , \u2_uk_K_r3_reg[43]/NET0131  , \u2_uk_K_r3_reg[44]/NET0131  , \u2_uk_K_r3_reg[45]/P0001  , \u2_uk_K_r3_reg[46]/NET0131  , \u2_uk_K_r3_reg[47]/NET0131  , \u2_uk_K_r3_reg[48]/NET0131  , \u2_uk_K_r3_reg[49]/NET0131  , \u2_uk_K_r3_reg[4]/NET0131  , \u2_uk_K_r3_reg[50]/NET0131  , \u2_uk_K_r3_reg[51]/NET0131  , \u2_uk_K_r3_reg[52]/NET0131  , \u2_uk_K_r3_reg[53]/NET0131  , \u2_uk_K_r3_reg[54]/NET0131  , \u2_uk_K_r3_reg[55]/NET0131  , \u2_uk_K_r3_reg[5]/NET0131  , \u2_uk_K_r3_reg[6]/NET0131  , \u2_uk_K_r3_reg[7]/NET0131  , \u2_uk_K_r3_reg[8]/NET0131  , \u2_uk_K_r3_reg[9]/NET0131  , \u2_uk_K_r4_reg[0]/P0001  , \u2_uk_K_r4_reg[10]/NET0131  , \u2_uk_K_r4_reg[11]/NET0131  , \u2_uk_K_r4_reg[12]/NET0131  , \u2_uk_K_r4_reg[13]/NET0131  , \u2_uk_K_r4_reg[14]/NET0131  , \u2_uk_K_r4_reg[15]/NET0131  , \u2_uk_K_r4_reg[16]/NET0131  , \u2_uk_K_r4_reg[17]/NET0131  , \u2_uk_K_r4_reg[18]/NET0131  , \u2_uk_K_r4_reg[19]/NET0131  , \u2_uk_K_r4_reg[1]/NET0131  , \u2_uk_K_r4_reg[20]/NET0131  , \u2_uk_K_r4_reg[21]/NET0131  , \u2_uk_K_r4_reg[22]/NET0131  , \u2_uk_K_r4_reg[23]/NET0131  , \u2_uk_K_r4_reg[25]/NET0131  , \u2_uk_K_r4_reg[26]/NET0131  , \u2_uk_K_r4_reg[27]/P0001  , \u2_uk_K_r4_reg[28]/NET0131  , \u2_uk_K_r4_reg[29]/NET0131  , \u2_uk_K_r4_reg[30]/NET0131  , \u2_uk_K_r4_reg[31]/P0001  , \u2_uk_K_r4_reg[32]/NET0131  , \u2_uk_K_r4_reg[33]/NET0131  , \u2_uk_K_r4_reg[34]/NET0131  , \u2_uk_K_r4_reg[35]/NET0131  , \u2_uk_K_r4_reg[36]/NET0131  , \u2_uk_K_r4_reg[37]/NET0131  , \u2_uk_K_r4_reg[38]/NET0131  , \u2_uk_K_r4_reg[39]/NET0131  , \u2_uk_K_r4_reg[3]/NET0131  , \u2_uk_K_r4_reg[40]/NET0131  , \u2_uk_K_r4_reg[41]/NET0131  , \u2_uk_K_r4_reg[42]/NET0131  , \u2_uk_K_r4_reg[43]/NET0131  , \u2_uk_K_r4_reg[44]/NET0131  , \u2_uk_K_r4_reg[45]/NET0131  , \u2_uk_K_r4_reg[46]/NET0131  , \u2_uk_K_r4_reg[47]/NET0131  , \u2_uk_K_r4_reg[48]/NET0131  , \u2_uk_K_r4_reg[49]/NET0131  , \u2_uk_K_r4_reg[4]/NET0131  , \u2_uk_K_r4_reg[50]/NET0131  , \u2_uk_K_r4_reg[51]/NET0131  , \u2_uk_K_r4_reg[52]/NET0131  , \u2_uk_K_r4_reg[53]/NET0131  , \u2_uk_K_r4_reg[54]/NET0131  , \u2_uk_K_r4_reg[55]/NET0131  , \u2_uk_K_r4_reg[5]/NET0131  , \u2_uk_K_r4_reg[6]/NET0131  , \u2_uk_K_r4_reg[7]/NET0131  , \u2_uk_K_r4_reg[8]/NET0131  , \u2_uk_K_r4_reg[9]/NET0131  , \u2_uk_K_r5_reg[0]/NET0131  , \u2_uk_K_r5_reg[10]/NET0131  , \u2_uk_K_r5_reg[11]/NET0131  , \u2_uk_K_r5_reg[12]/NET0131  , \u2_uk_K_r5_reg[13]/P0001  , \u2_uk_K_r5_reg[14]/NET0131  , \u2_uk_K_r5_reg[15]/NET0131  , \u2_uk_K_r5_reg[16]/NET0131  , \u2_uk_K_r5_reg[17]/NET0131  , \u2_uk_K_r5_reg[18]/NET0131  , \u2_uk_K_r5_reg[19]/NET0131  , \u2_uk_K_r5_reg[1]/NET0131  , \u2_uk_K_r5_reg[20]/NET0131  , \u2_uk_K_r5_reg[21]/NET0131  , \u2_uk_K_r5_reg[22]/NET0131  , \u2_uk_K_r5_reg[23]/NET0131  , \u2_uk_K_r5_reg[24]/NET0131  , \u2_uk_K_r5_reg[25]/NET0131  , \u2_uk_K_r5_reg[26]/NET0131  , \u2_uk_K_r5_reg[27]/NET0131  , \u2_uk_K_r5_reg[28]/NET0131  , \u2_uk_K_r5_reg[29]/NET0131  , \u2_uk_K_r5_reg[2]/NET0131  , \u2_uk_K_r5_reg[30]/NET0131  , \u2_uk_K_r5_reg[31]/NET0131  , \u2_uk_K_r5_reg[32]/NET0131  , \u2_uk_K_r5_reg[33]/NET0131  , \u2_uk_K_r5_reg[34]/NET0131  , \u2_uk_K_r5_reg[35]/NET0131  , \u2_uk_K_r5_reg[36]/NET0131  , \u2_uk_K_r5_reg[37]/P0001  , \u2_uk_K_r5_reg[38]/NET0131  , \u2_uk_K_r5_reg[39]/NET0131  , \u2_uk_K_r5_reg[3]/NET0131  , \u2_uk_K_r5_reg[40]/NET0131  , \u2_uk_K_r5_reg[41]/NET0131  , \u2_uk_K_r5_reg[42]/NET0131  , \u2_uk_K_r5_reg[43]/NET0131  , \u2_uk_K_r5_reg[44]/NET0131  , \u2_uk_K_r5_reg[46]/NET0131  , \u2_uk_K_r5_reg[47]/NET0131  , \u2_uk_K_r5_reg[48]/NET0131  , \u2_uk_K_r5_reg[49]/NET0131  , \u2_uk_K_r5_reg[4]/NET0131  , \u2_uk_K_r5_reg[50]/NET0131  , \u2_uk_K_r5_reg[51]/NET0131  , \u2_uk_K_r5_reg[52]/NET0131  , \u2_uk_K_r5_reg[53]/NET0131  , \u2_uk_K_r5_reg[54]/NET0131  , \u2_uk_K_r5_reg[55]/NET0131  , \u2_uk_K_r5_reg[5]/NET0131  , \u2_uk_K_r5_reg[6]/NET0131  , \u2_uk_K_r5_reg[7]/NET0131  , \u2_uk_K_r5_reg[8]/NET0131  , \u2_uk_K_r5_reg[9]/P0001  , \u2_uk_K_r6_reg[0]/NET0131  , \u2_uk_K_r6_reg[10]/NET0131  , \u2_uk_K_r6_reg[11]/NET0131  , \u2_uk_K_r6_reg[12]/NET0131  , \u2_uk_K_r6_reg[13]/NET0131  , \u2_uk_K_r6_reg[14]/NET0131  , \u2_uk_K_r6_reg[15]/NET0131  , \u2_uk_K_r6_reg[16]/NET0131  , \u2_uk_K_r6_reg[17]/NET0131  , \u2_uk_K_r6_reg[18]/NET0131  , \u2_uk_K_r6_reg[19]/NET0131  , \u2_uk_K_r6_reg[1]/NET0131  , \u2_uk_K_r6_reg[20]/NET0131  , \u2_uk_K_r6_reg[21]/NET0131  , \u2_uk_K_r6_reg[22]/NET0131  , \u2_uk_K_r6_reg[23]/P0001  , \u2_uk_K_r6_reg[24]/NET0131  , \u2_uk_K_r6_reg[25]/NET0131  , \u2_uk_K_r6_reg[26]/NET0131  , \u2_uk_K_r6_reg[27]/NET0131  , \u2_uk_K_r6_reg[28]/NET0131  , \u2_uk_K_r6_reg[29]/NET0131  , \u2_uk_K_r6_reg[2]/NET0131  , \u2_uk_K_r6_reg[30]/P0001  , \u2_uk_K_r6_reg[31]/NET0131  , \u2_uk_K_r6_reg[32]/NET0131  , \u2_uk_K_r6_reg[33]/NET0131  , \u2_uk_K_r6_reg[34]/NET0131  , \u2_uk_K_r6_reg[35]/NET0131  , \u2_uk_K_r6_reg[36]/NET0131  , \u2_uk_K_r6_reg[37]/NET0131  , \u2_uk_K_r6_reg[38]/NET0131  , \u2_uk_K_r6_reg[39]/NET0131  , \u2_uk_K_r6_reg[3]/NET0131  , \u2_uk_K_r6_reg[40]/NET0131  , \u2_uk_K_r6_reg[41]/NET0131  , \u2_uk_K_r6_reg[42]/NET0131  , \u2_uk_K_r6_reg[43]/NET0131  , \u2_uk_K_r6_reg[44]/NET0131  , \u2_uk_K_r6_reg[45]/NET0131  , \u2_uk_K_r6_reg[46]/NET0131  , \u2_uk_K_r6_reg[47]/NET0131  , \u2_uk_K_r6_reg[48]/NET0131  , \u2_uk_K_r6_reg[49]/NET0131  , \u2_uk_K_r6_reg[4]/NET0131  , \u2_uk_K_r6_reg[50]/NET0131  , \u2_uk_K_r6_reg[51]/NET0131  , \u2_uk_K_r6_reg[52]/NET0131  , \u2_uk_K_r6_reg[53]/NET0131  , \u2_uk_K_r6_reg[54]/NET0131  , \u2_uk_K_r6_reg[55]/P0001  , \u2_uk_K_r6_reg[5]/NET0131  , \u2_uk_K_r6_reg[6]/NET0131  , \u2_uk_K_r6_reg[7]/NET0131  , \u2_uk_K_r6_reg[8]/NET0131  , \u2_uk_K_r6_reg[9]/NET0131  , \u2_uk_K_r7_reg[0]/NET0131  , \u2_uk_K_r7_reg[10]/NET0131  , \u2_uk_K_r7_reg[11]/NET0131  , \u2_uk_K_r7_reg[12]/NET0131  , \u2_uk_K_r7_reg[13]/NET0131  , \u2_uk_K_r7_reg[14]/NET0131  , \u2_uk_K_r7_reg[15]/NET0131  , \u2_uk_K_r7_reg[16]/NET0131  , \u2_uk_K_r7_reg[17]/NET0131  , \u2_uk_K_r7_reg[18]/NET0131  , \u2_uk_K_r7_reg[19]/NET0131  , \u2_uk_K_r7_reg[1]/NET0131  , \u2_uk_K_r7_reg[20]/NET0131  , \u2_uk_K_r7_reg[21]/NET0131  , \u2_uk_K_r7_reg[22]/NET0131  , \u2_uk_K_r7_reg[23]/P0001  , \u2_uk_K_r7_reg[24]/NET0131  , \u2_uk_K_r7_reg[25]/NET0131  , \u2_uk_K_r7_reg[26]/NET0131  , \u2_uk_K_r7_reg[27]/NET0131  , \u2_uk_K_r7_reg[28]/NET0131  , \u2_uk_K_r7_reg[29]/NET0131  , \u2_uk_K_r7_reg[2]/NET0131  , \u2_uk_K_r7_reg[30]/P0001  , \u2_uk_K_r7_reg[31]/NET0131  , \u2_uk_K_r7_reg[32]/NET0131  , \u2_uk_K_r7_reg[33]/NET0131  , \u2_uk_K_r7_reg[34]/NET0131  , \u2_uk_K_r7_reg[35]/NET0131  , \u2_uk_K_r7_reg[36]/NET0131  , \u2_uk_K_r7_reg[37]/NET0131  , \u2_uk_K_r7_reg[38]/NET0131  , \u2_uk_K_r7_reg[39]/NET0131  , \u2_uk_K_r7_reg[3]/NET0131  , \u2_uk_K_r7_reg[40]/NET0131  , \u2_uk_K_r7_reg[41]/NET0131  , \u2_uk_K_r7_reg[42]/NET0131  , \u2_uk_K_r7_reg[43]/NET0131  , \u2_uk_K_r7_reg[44]/NET0131  , \u2_uk_K_r7_reg[45]/NET0131  , \u2_uk_K_r7_reg[46]/NET0131  , \u2_uk_K_r7_reg[47]/NET0131  , \u2_uk_K_r7_reg[48]/NET0131  , \u2_uk_K_r7_reg[49]/NET0131  , \u2_uk_K_r7_reg[4]/NET0131  , \u2_uk_K_r7_reg[50]/NET0131  , \u2_uk_K_r7_reg[51]/NET0131  , \u2_uk_K_r7_reg[52]/NET0131  , \u2_uk_K_r7_reg[53]/NET0131  , \u2_uk_K_r7_reg[54]/NET0131  , \u2_uk_K_r7_reg[55]/P0001  , \u2_uk_K_r7_reg[5]/NET0131  , \u2_uk_K_r7_reg[6]/NET0131  , \u2_uk_K_r7_reg[7]/NET0131  , \u2_uk_K_r7_reg[8]/NET0131  , \u2_uk_K_r7_reg[9]/NET0131  , \u2_uk_K_r8_reg[0]/NET0131  , \u2_uk_K_r8_reg[10]/NET0131  , \u2_uk_K_r8_reg[11]/NET0131  , \u2_uk_K_r8_reg[12]/NET0131  , \u2_uk_K_r8_reg[13]/P0001  , \u2_uk_K_r8_reg[14]/NET0131  , \u2_uk_K_r8_reg[15]/NET0131  , \u2_uk_K_r8_reg[16]/NET0131  , \u2_uk_K_r8_reg[17]/NET0131  , \u2_uk_K_r8_reg[18]/NET0131  , \u2_uk_K_r8_reg[19]/NET0131  , \u2_uk_K_r8_reg[1]/NET0131  , \u2_uk_K_r8_reg[20]/NET0131  , \u2_uk_K_r8_reg[21]/NET0131  , \u2_uk_K_r8_reg[22]/NET0131  , \u2_uk_K_r8_reg[23]/NET0131  , \u2_uk_K_r8_reg[24]/NET0131  , \u2_uk_K_r8_reg[25]/NET0131  , \u2_uk_K_r8_reg[26]/NET0131  , \u2_uk_K_r8_reg[27]/NET0131  , \u2_uk_K_r8_reg[28]/NET0131  , \u2_uk_K_r8_reg[29]/NET0131  , \u2_uk_K_r8_reg[2]/NET0131  , \u2_uk_K_r8_reg[30]/NET0131  , \u2_uk_K_r8_reg[31]/NET0131  , \u2_uk_K_r8_reg[32]/NET0131  , \u2_uk_K_r8_reg[33]/NET0131  , \u2_uk_K_r8_reg[34]/NET0131  , \u2_uk_K_r8_reg[35]/NET0131  , \u2_uk_K_r8_reg[36]/NET0131  , \u2_uk_K_r8_reg[37]/P0001  , \u2_uk_K_r8_reg[38]/NET0131  , \u2_uk_K_r8_reg[39]/NET0131  , \u2_uk_K_r8_reg[3]/NET0131  , \u2_uk_K_r8_reg[40]/NET0131  , \u2_uk_K_r8_reg[41]/NET0131  , \u2_uk_K_r8_reg[42]/NET0131  , \u2_uk_K_r8_reg[43]/NET0131  , \u2_uk_K_r8_reg[44]/NET0131  , \u2_uk_K_r8_reg[46]/NET0131  , \u2_uk_K_r8_reg[47]/NET0131  , \u2_uk_K_r8_reg[48]/NET0131  , \u2_uk_K_r8_reg[49]/NET0131  , \u2_uk_K_r8_reg[4]/NET0131  , \u2_uk_K_r8_reg[50]/NET0131  , \u2_uk_K_r8_reg[51]/NET0131  , \u2_uk_K_r8_reg[52]/NET0131  , \u2_uk_K_r8_reg[53]/NET0131  , \u2_uk_K_r8_reg[54]/NET0131  , \u2_uk_K_r8_reg[55]/NET0131  , \u2_uk_K_r8_reg[5]/NET0131  , \u2_uk_K_r8_reg[6]/NET0131  , \u2_uk_K_r8_reg[7]/NET0131  , \u2_uk_K_r8_reg[8]/NET0131  , \u2_uk_K_r8_reg[9]/NET0131  , \u2_uk_K_r9_reg[0]/P0001  , \u2_uk_K_r9_reg[10]/NET0131  , \u2_uk_K_r9_reg[11]/NET0131  , \u2_uk_K_r9_reg[12]/NET0131  , \u2_uk_K_r9_reg[13]/NET0131  , \u2_uk_K_r9_reg[14]/NET0131  , \u2_uk_K_r9_reg[15]/NET0131  , \u2_uk_K_r9_reg[16]/NET0131  , \u2_uk_K_r9_reg[17]/NET0131  , \u2_uk_K_r9_reg[18]/NET0131  , \u2_uk_K_r9_reg[19]/NET0131  , \u2_uk_K_r9_reg[1]/NET0131  , \u2_uk_K_r9_reg[20]/NET0131  , \u2_uk_K_r9_reg[21]/NET0131  , \u2_uk_K_r9_reg[22]/NET0131  , \u2_uk_K_r9_reg[23]/NET0131  , \u2_uk_K_r9_reg[25]/NET0131  , \u2_uk_K_r9_reg[26]/NET0131  , \u2_uk_K_r9_reg[27]/NET0131  , \u2_uk_K_r9_reg[28]/NET0131  , \u2_uk_K_r9_reg[29]/NET0131  , \u2_uk_K_r9_reg[30]/NET0131  , \u2_uk_K_r9_reg[31]/P0001  , \u2_uk_K_r9_reg[32]/NET0131  , \u2_uk_K_r9_reg[33]/NET0131  , \u2_uk_K_r9_reg[34]/NET0131  , \u2_uk_K_r9_reg[35]/NET0131  , \u2_uk_K_r9_reg[36]/NET0131  , \u2_uk_K_r9_reg[37]/NET0131  , \u2_uk_K_r9_reg[38]/NET0131  , \u2_uk_K_r9_reg[39]/NET0131  , \u2_uk_K_r9_reg[3]/NET0131  , \u2_uk_K_r9_reg[40]/NET0131  , \u2_uk_K_r9_reg[41]/NET0131  , \u2_uk_K_r9_reg[42]/NET0131  , \u2_uk_K_r9_reg[43]/NET0131  , \u2_uk_K_r9_reg[44]/NET0131  , \u2_uk_K_r9_reg[45]/NET0131  , \u2_uk_K_r9_reg[46]/NET0131  , \u2_uk_K_r9_reg[47]/NET0131  , \u2_uk_K_r9_reg[48]/NET0131  , \u2_uk_K_r9_reg[49]/NET0131  , \u2_uk_K_r9_reg[4]/NET0131  , \u2_uk_K_r9_reg[50]/NET0131  , \u2_uk_K_r9_reg[51]/NET0131  , \u2_uk_K_r9_reg[52]/NET0131  , \u2_uk_K_r9_reg[53]/NET0131  , \u2_uk_K_r9_reg[54]/NET0131  , \u2_uk_K_r9_reg[55]/NET0131  , \u2_uk_K_r9_reg[5]/NET0131  , \u2_uk_K_r9_reg[6]/NET0131  , \u2_uk_K_r9_reg[7]/NET0131  , \u2_uk_K_r9_reg[8]/NET0131  , \u2_uk_K_r9_reg[9]/NET0131  , \_al_n0  , \_al_n1  , \g16/_0_  , \g191647/_3_  , \g191648/_3_  , \g191819/_3_  , \g191821/_0_  , \g191940/_3_  , \g191941/_0_  , \g191942/_0_  , \g191944/_0_  , \g191945/_0_  , \g191946/_0_  , \g191947/_3_  , \g191948/_0_  , \g191949/_0_  , \g191950/_0_  , \g191951/_3_  , \g191952/_0_  , \g192015/_3_  , \g192016/_3_  , \g192017/_3_  , \g192018/_3_  , \g192019/_3_  , \g192020/_0_  , \g192021/_3_  , \g192022/_0_  , \g192047/_0_  , \g192048/_0_  , \g192049/_0_  , \g192050/_0_  , \g192051/_0_  , \g192081/_0_  , \g193428/_3_  , \g193720/_0_  , \g193721/_0_  , \g193877/_0_  , \g193878/_0_  , \g193879/_0_  , \g193880/_3_  , \g193881/_0_  , \g193882/_0_  , \g193998/_0_  , \g193999/_0_  , \g194000/_3_  , \g194001/_0_  , \g194002/_0_  , \g194003/_0_  , \g194004/_0_  , \g194005/_0_  , \g194006/_0_  , \g194007/_0_  , \g194008/_0_  , \g194009/_0_  , \g194010/_0_  , \g194055/_3_  , \g194056/_3_  , \g194057/_0_  , \g194058/_0_  , \g194059/_0_  , \g194060/_0_  , \g194090/_0_  , \g194091/_0_  , \g194092/_0_  , \g194093/_0_  , \g195671/_0_  , \g195672/_3_  , \g195868/_0_  , \g195869/_0_  , \g195870/_0_  , \g196010/_0_  , \g196011/_0_  , \g196012/_0_  , \g196013/_0_  , \g196014/_0_  , \g196015/_0_  , \g196016/_0_  , \g196017/_0_  , \g196018/_0_  , \g196019/_3_  , \g196020/_0_  , \g196021/_0_  , \g196022/_0_  , \g196096/_3_  , \g196097/_0_  , \g196098/_0_  , \g196099/_0_  , \g196100/_3_  , \g196101/_0_  , \g196102/_0_  , \g196103/_0_  , \g196136/_0_  , \g196137/_0_  , \g196138/_0_  , \g196139/_0_  , \g196140/_0_  , \g196170/_0_  , \g197520/_3_  , \g197821/_0_  , \g197923/_0_  , \g197996/_0_  , \g197997/_3_  , \g197998/_0_  , \g197999/_0_  , \g198000/_0_  , \g198071/_0_  , \g198123/_0_  , \g198124/_0_  , \g198125/_0_  , \g198126/_0_  , \g198127/_0_  , \g198128/_0_  , \g198129/_0_  , \g198130/_0_  , \g198131/_0_  , \g198132/_0_  , \g198133/_0_  , \g198134/_3_  , \g198135/_0_  , \g198182/_0_  , \g198183/_3_  , \g198184/_0_  , \g198185/_0_  , \g198186/_0_  , \g198187/_0_  , \g198219/_0_  , \g198220/_0_  , \g198221/_0_  , \g198222/_0_  , \g199794/_0_  , \g199795/_3_  , \g200006/_0_  , \g200007/_0_  , \g200008/_0_  , \g200139/_0_  , \g200140/_0_  , \g200141/_0_  , \g200142/_0_  , \g200143/_0_  , \g200144/_0_  , \g200145/_0_  , \g200146/_0_  , \g200147/_0_  , \g200148/_0_  , \g200149/_0_  , \g200150/_3_  , \g200151/_0_  , \g200228/_3_  , \g200229/_0_  , \g200230/_0_  , \g200231/_0_  , \g200232/_3_  , \g200233/_0_  , \g200234/_0_  , \g200235/_0_  , \g200268/_0_  , \g200269/_0_  , \g200270/_0_  , \g200271/_0_  , \g200272/_0_  , \g200299/_0_  , \g201655/_3_  , \g201960/_0_  , \g201961/_0_  , \g202131/_0_  , \g202132/_0_  , \g202133/_3_  , \g202134/_0_  , \g202135/_0_  , \g202136/_0_  , \g202257/_0_  , \g202258/_0_  , \g202259/_3_  , \g202260/_0_  , \g202261/_0_  , \g202262/_0_  , \g202263/_0_  , \g202264/_0_  , \g202265/_0_  , \g202266/_0_  , \g202267/_0_  , \g202268/_0_  , \g202269/_0_  , \g202317/_0_  , \g202318/_3_  , \g202319/_0_  , \g202320/_0_  , \g202321/_0_  , \g202322/_0_  , \g202354/_0_  , \g202355/_0_  , \g202356/_0_  , \g202357/_0_  , \g203927/_0_  , \g203928/_3_  , \g204142/_0_  , \g204143/_0_  , \g204144/_0_  , \g204275/_0_  , \g204276/_0_  , \g204277/_0_  , \g204278/_0_  , \g204279/_0_  , \g204280/_0_  , \g204281/_0_  , \g204282/_0_  , \g204283/_0_  , \g204284/_0_  , \g204285/_0_  , \g204286/_3_  , \g204287/_0_  , \g204363/_3_  , \g204364/_0_  , \g204365/_0_  , \g204366/_0_  , \g204367/_3_  , \g204368/_0_  , \g204369/_0_  , \g204370/_0_  , \g204403/_0_  , \g204404/_0_  , \g204405/_0_  , \g204406/_0_  , \g204407/_0_  , \g204434/_0_  , \g205833/_3_  , \g206103/_0_  , \g206104/_0_  , \g206266/_0_  , \g206267/_0_  , \g206268/_0_  , \g206269/_3_  , \g206270/_0_  , \g206271/_0_  , \g206387/_0_  , \g206388/_0_  , \g206389/_3_  , \g206390/_0_  , \g206391/_0_  , \g206392/_0_  , \g206393/_0_  , \g206394/_0_  , \g206395/_0_  , \g206396/_0_  , \g206397/_0_  , \g206398/_0_  , \g206399/_0_  , \g206446/_0_  , \g206447/_3_  , \g206448/_0_  , \g206449/_0_  , \g206450/_0_  , \g206451/_0_  , \g206483/_0_  , \g206484/_0_  , \g206485/_0_  , \g206486/_0_  , \g208069/_0_  , \g208070/_3_  , \g208253/_0_  , \g208254/_0_  , \g208255/_0_  , \g208406/_0_  , \g208407/_0_  , \g208408/_0_  , \g208409/_0_  , \g208410/_0_  , \g208411/_0_  , \g208412/_0_  , \g208413/_0_  , \g208414/_0_  , \g208415/_3_  , \g208416/_0_  , \g208417/_0_  , \g208418/_0_  , \g208493/_3_  , \g208494/_0_  , \g208495/_0_  , \g208496/_0_  , \g208497/_3_  , \g208498/_0_  , \g208499/_0_  , \g208500/_0_  , \g208533/_0_  , \g208534/_0_  , \g208535/_0_  , \g208536/_0_  , \g208537/_0_  , \g208564/_0_  , \g209938/_3_  , \g210205/_0_  , \g210206/_0_  , \g210380/_0_  , \g210381/_0_  , \g210382/_0_  , \g210383/_3_  , \g210384/_0_  , \g210385/_0_  , \g210499/_0_  , \g210500/_0_  , \g210501/_3_  , \g210502/_0_  , \g210503/_0_  , \g210504/_0_  , \g210505/_0_  , \g210506/_0_  , \g210507/_0_  , \g210508/_0_  , \g210509/_0_  , \g210510/_0_  , \g210511/_0_  , \g210558/_0_  , \g210559/_3_  , \g210560/_0_  , \g210561/_0_  , \g210562/_0_  , \g210563/_0_  , \g210595/_0_  , \g210596/_0_  , \g210597/_0_  , \g210598/_0_  , \g212159/_0_  , \g212160/_3_  , \g212384/_0_  , \g212385/_0_  , \g212386/_0_  , \g212536/_0_  , \g212537/_0_  , \g212538/_0_  , \g212539/_0_  , \g212540/_0_  , \g212541/_0_  , \g212542/_0_  , \g212543/_0_  , \g212544/_0_  , \g212545/_0_  , \g212546/_3_  , \g212547/_0_  , \g212623/_3_  , \g212624/_0_  , \g212625/_0_  , \g212626/_0_  , \g212627/_0_  , \g212628/_3_  , \g212629/_0_  , \g212630/_0_  , \g212631/_0_  , \g212667/_0_  , \g212668/_0_  , \g212669/_0_  , \g212670/_0_  , \g212671/_0_  , \g212699/_0_  , \g214033/_3_  , \g214309/_3_  , \g214310/_0_  , \g214494/_0_  , \g214495/_0_  , \g214496/_0_  , \g214497/_3_  , \g214632/_0_  , \g214633/_0_  , \g214634/_3_  , \g214635/_0_  , \g214636/_0_  , \g214637/_0_  , \g214638/_0_  , \g214639/_0_  , \g214640/_0_  , \g214641/_0_  , \g214642/_0_  , \g214643/_0_  , \g214691/_0_  , \g214692/_0_  , \g214693/_3_  , \g214694/_0_  , \g214695/_0_  , \g214696/_0_  , \g214697/_0_  , \g214729/_0_  , \g214730/_0_  , \g214731/_0_  , \g214732/_0_  , \g214733/_0_  , \g216157/_0_  , \g216158/_3_  , \g216492/_0_  , \g216493/_0_  , \g216671/_0_  , \g216672/_0_  , \g216673/_0_  , \g216674/_0_  , \g216675/_0_  , \g216676/_3_  , \g216677/_0_  , \g216735/_0_  , \g216736/_3_  , \g216737/_0_  , \g216738/_0_  , \g216739/_0_  , \g216740/_0_  , \g216741/_0_  , \g216742/_0_  , \g216743/_0_  , \g216744/_0_  , \g216745/_0_  , \g216746/_3_  , \g216747/_0_  , \g216748/_0_  , \g216749/_0_  , \g216788/_0_  , \g216789/_0_  , \g216790/_0_  , \g216791/_0_  , \g216792/_0_  , \g216829/_0_  , \g218407/_3_  , \g218408/_0_  , \g218423/_3_  , \g218601/_0_  , \g218602/_0_  , \g218603/_0_  , \g218604/_0_  , \g218724/_0_  , \g218725/_0_  , \g218726/_0_  , \g218727/_0_  , \g218728/_0_  , \g218729/_0_  , \g218730/_0_  , \g218731/_0_  , \g218732/_0_  , \g218733/_0_  , \g218734/_0_  , \g218735/_3_  , \g218736/_0_  , \g218808/_3_  , \g218809/_0_  , \g218810/_0_  , \g218811/_3_  , \g218812/_0_  , \g218813/_0_  , \g218814/_0_  , \g218846/_0_  , \g218847/_0_  , \g218848/_0_  , \g218849/_0_  , \g218877/_0_  , \g22/_0_  , \g220545/_0_  , \g220546/_3_  , \g220725/_3_  , \g220726/_0_  , \g220793/_0_  , \g220794/_0_  , \g220795/_0_  , \g220796/_0_  , \g220797/_0_  , \g220798/_0_  , \g220799/_0_  , \g220800/_0_  , \g220801/_0_  , \g220802/_0_  , \g220803/_0_  , \g220804/_3_  , \g220805/_0_  , \g220806/_0_  , \g220807/_0_  , \g220872/_3_  , \g220873/_0_  , \g220874/_3_  , \g220875/_0_  , \g220876/_0_  , \g220877/_0_  , \g220921/_0_  , \g220922/_0_  , \g220923/_0_  , \g220924/_0_  , \g220925/_0_  , \g220926/_0_  , \g220969/_0_  , \g221011/_3_  , \g221039/_3_  , \g221086/_3_  , \g221131/_0_  , \g224010/_3_  , \g224368/_3_  , \g224369/_3_  , \g224532/_0_  , \g224533/_0_  , \g224534/_0_  , \g224535/_3_  , \g224536/_0_  , \g224537/_0_  , \g224640/_3_  , \g224641/_0_  , \g224642/_0_  , \g224643/_3_  , \g224644/_0_  , \g224645/_0_  , \g224646/_3_  , \g224647/_0_  , \g224648/_3_  , \g224649/_0_  , \g224650/_0_  , \g224651/_0_  , \g224652/_0_  , \g224690/_0_  , \g224691/_3_  , \g224692/_3_  , \g224693/_0_  , \g224694/_0_  , \g224695/_3_  , \g224723/_0_  , \g224724/_0_  , \g224725/_0_  , \g224726/_0_  , \g226372/_0_  , \g226373/_3_  , \g226549/_3_  , \g226550/_0_  , \g226616/_0_  , \g226635/_0_  , \g226636/_0_  , \g226637/_0_  , \g226638/_0_  , \g226639/_0_  , \g226640/_0_  , \g226641/_3_  , \g226642/_0_  , \g226643/_0_  , \g226644/_0_  , \g226645/_0_  , \g226646/_0_  , \g226692/_3_  , \g226693/_0_  , \g226694/_3_  , \g226695/_3_  , \g226696/_3_  , \g226697/_0_  , \g226698/_0_  , \g226699/_0_  , \g226728/_0_  , \g226729/_0_  , \g226730/_0_  , \g226731/_0_  , \g226732/_0_  , \g226759/_0_  , \g228250/_0_  , \g228396/_0_  , \g228397/_0_  , \g228566/_0_  , \g228567/_0_  , \g228568/_0_  , \g228609/_0_  , \g228610/_3_  , \g228688/_0_  , \g228689/_0_  , \g228690/_3_  , \g228691/_0_  , \g228692/_0_  , \g228693/_0_  , \g228694/_0_  , \g228695/_0_  , \g228696/_0_  , \g228697/_0_  , \g228698/_0_  , \g228699/_0_  , \g228700/_0_  , \g228748/_0_  , \g228749/_3_  , \g228750/_0_  , \g228751/_0_  , \g228752/_0_  , \g228753/_0_  , \g228784/_0_  , \g228785/_0_  , \g228786/_0_  , \g228787/_3_  , \g230339/_0_  , \g230340/_0_  , \g230546/_0_  , \g230580/_0_  , \g230679/_0_  , \g230680/_0_  , \g230681/_0_  , \g230682/_0_  , \g230683/_0_  , \g230684/_0_  , \g230685/_0_  , \g230686/_0_  , \g230687/_0_  , \g230688/_0_  , \g230689/_3_  , \g230690/_0_  , \g230710/_0_  , \g230766/_0_  , \g230767/_0_  , \g230768/_0_  , \g230769/_3_  , \g230770/_0_  , \g230771/_0_  , \g230772/_0_  , \g230773/_3_  , \g230810/_0_  , \g230811/_0_  , \g230812/_0_  , \g230813/_0_  , \g230814/_0_  , \g230840/_3_  , \g232196/_3_  , \g232469/_0_  , \g232470/_0_  , \g232633/_0_  , \g232635/_3_  , \g232636/_0_  , \g232637/_0_  , \g232691/_0_  , \g232747/_0_  , \g232748/_0_  , \g232749/_3_  , \g232750/_0_  , \g232751/_0_  , \g232752/_0_  , \g232753/_0_  , \g232754/_0_  , \g232755/_0_  , \g232756/_0_  , \g232757/_0_  , \g232758/_0_  , \g232759/_0_  , \g232804/_0_  , \g232805/_0_  , \g232806/_0_  , \g232807/_0_  , \g232808/_3_  , \g232809/_0_  , \g232841/_0_  , \g232842/_3_  , \g232843/_0_  , \g232844/_0_  , \g234520/_0_  , \g234687/_0_  , \g234688/_0_  , \g234689/_0_  , \g234764/_0_  , \g234765/_0_  , \g234766/_0_  , \g234767/_3_  , \g234768/_0_  , \g234769/_0_  , \g234770/_0_  , \g234771/_0_  , \g234772/_0_  , \g234773/_0_  , \g234774/_3_  , \g234775/_0_  , \g234776/_0_  , \g234824/_3_  , \g234825/_0_  , \g234826/_0_  , \g234827/_0_  , \g234828/_3_  , \g234829/_0_  , \g234830/_0_  , \g234831/_0_  , \g234867/_0_  , \g234868/_0_  , \g234869/_0_  , \g234870/_0_  , \g234896/_0_  , \g236294/_3_  , \g236541/_0_  , \g236542/_0_  , \g236724/_0_  , \g236725/_0_  , \g236726/_0_  , \g236727/_3_  , \g236728/_0_  , \g236729/_0_  , \g236821/_0_  , \g236822/_3_  , \g236823/_0_  , \g236824/_3_  , \g236825/_0_  , \g236826/_0_  , \g236827/_0_  , \g236828/_0_  , \g236829/_0_  , \g236830/_0_  , \g236831/_0_  , \g236832/_0_  , \g236877/_0_  , \g236878/_3_  , \g236879/_0_  , \g236880/_0_  , \g236881/_0_  , \g236882/_0_  , \g236914/_0_  , \g236915/_0_  , \g236916/_0_  , \g236917/_0_  , \g238530/_0_  , \g238531/_3_  , \g238723/_0_  , \g238724/_0_  , \g238725/_0_  , \g238840/_0_  , \g238841/_0_  , \g238842/_0_  , \g238843/_3_  , \g238844/_0_  , \g238845/_0_  , \g238846/_0_  , \g238847/_0_  , \g238848/_0_  , \g238849/_0_  , \g238850/_0_  , \g238851/_3_  , \g238852/_0_  , \g238924/_0_  , \g238925/_0_  , \g238926/_0_  , \g238927/_3_  , \g238928/_0_  , \g238929/_0_  , \g238930/_0_  , \g238965/_0_  , \g238966/_0_  , \g238967/_0_  , \g238968/_0_  , \g238969/_0_  , \g238996/_0_  , \g240353/_3_  , \g240640/_0_  , \g240641/_0_  , \g240813/_0_  , \g240814/_0_  , \g240815/_3_  , \g240816/_0_  , \g240817/_0_  , \g240818/_0_  , \g240925/_0_  , \g240926/_0_  , \g240927/_3_  , \g240928/_0_  , \g240929/_3_  , \g240930/_0_  , \g240931/_0_  , \g240932/_0_  , \g240933/_0_  , \g240934/_0_  , \g240935/_0_  , \g240936/_0_  , \g240937/_0_  , \g240984/_0_  , \g240985/_3_  , \g240986/_0_  , \g240987/_0_  , \g240988/_0_  , \g240989/_0_  , \g241021/_0_  , \g241022/_0_  , \g241023/_0_  , \g241024/_0_  , \g242616/_0_  , \g242617/_3_  , \g242815/_0_  , \g242816/_0_  , \g242817/_0_  , \g242955/_0_  , \g242956/_0_  , \g242957/_0_  , \g242958/_3_  , \g242959/_0_  , \g242960/_0_  , \g242961/_0_  , \g242962/_0_  , \g242963/_3_  , \g242964/_0_  , \g242965/_0_  , \g242966/_0_  , \g242967/_0_  , \g243037/_3_  , \g243038/_0_  , \g243039/_0_  , \g243040/_0_  , \g243041/_3_  , \g243042/_0_  , \g243043/_0_  , \g243044/_0_  , \g243078/_0_  , \g243079/_0_  , \g243080/_0_  , \g243081/_0_  , \g243082/_0_  , \g243109/_0_  , \g244465/_3_  , \g244753/_3_  , \g244754/_0_  , \g244924/_0_  , \g244925/_0_  , \g244926/_3_  , \g244927/_0_  , \g244928/_0_  , \g245035/_0_  , \g245036/_0_  , \g245037/_0_  , \g245038/_3_  , \g245039/_3_  , \g245040/_0_  , \g245041/_0_  , \g245043/_0_  , \g245045/_0_  , \g245046/_0_  , \g245047/_0_  , \g245092/_0_  , \g245093/_3_  , \g245094/_0_  , \g245095/_0_  , \g245096/_0_  , \g245097/_0_  , \g245129/_0_  , \g245130/_0_  , \g245131/_0_  , \g245132/_0_  , \g246715/_0_  , \g246716/_3_  , \g246911/_0_  , \g246912/_0_  , \g246913/_0_  , \g247057/_0_  , \g247058/_0_  , \g247059/_0_  , \g247060/_0_  , \g247061/_0_  , \g247062/_3_  , \g247063/_0_  , \g247064/_0_  , \g247065/_0_  , \g247066/_0_  , \g247067/_3_  , \g247068/_0_  , \g247069/_0_  , \g247137/_3_  , \g247138/_0_  , \g247139/_0_  , \g247140/_0_  , \g247141/_3_  , \g247142/_0_  , \g247143/_0_  , \g247144/_0_  , \g247179/_0_  , \g247180/_0_  , \g247181/_0_  , \g247182/_0_  , \g247183/_0_  , \g247210/_0_  , \g248581/_3_  , \g248828/_0_  , \g248829/_0_  , \g249033/_0_  , \g249035/_0_  , \g249036/_3_  , \g249037/_0_  , \g249038/_0_  , \g249147/_0_  , \g249148/_0_  , \g249149/_3_  , \g249150/_0_  , \g249152/_0_  , \g249153/_0_  , \g249155/_0_  , \g249156/_0_  , \g249157/_0_  , \g249200/_3_  , \g249201/_0_  , \g249202/_0_  , \g249203/_3_  , \g249204/_0_  , \g249205/_0_  , \g249206/_0_  , \g249207/_0_  , \g249239/_0_  , \g249240/_0_  , \g249241/_0_  , \g249242/_0_  , \g250815/_0_  , \g251006/_0_  , \g251007/_0_  , \g251008/_0_  , \g251009/_3_  , \g251160/_0_  , \g251161/_0_  , \g251162/_0_  , \g251163/_3_  , \g251164/_0_  , \g251165/_0_  , \g251166/_0_  , \g251167/_0_  , \g251168/_0_  , \g251169/_0_  , \g251170/_3_  , \g251171/_0_  , \g251245/_3_  , \g251246/_0_  , \g251247/_0_  , \g251248/_0_  , \g251249/_3_  , \g251250/_0_  , \g251251/_0_  , \g251252/_0_  , \g251286/_0_  , \g251287/_0_  , \g251288/_0_  , \g251289/_0_  , \g251290/_0_  , \g251291/_0_  , \g251318/_0_  , \g252698/_3_  , \g252942/_0_  , \g252943/_0_  , \g253118/_0_  , \g253119/_0_  , \g253120/_0_  , \g253121/_0_  , \g253122/_3_  , \g253123/_0_  , \g253236/_0_  , \g253237/_3_  , \g253238/_3_  , \g253239/_0_  , \g253240/_0_  , \g253241/_0_  , \g253242/_0_  , \g253243/_0_  , \g253244/_0_  , \g253245/_0_  , \g253246/_0_  , \g253247/_0_  , \g253248/_0_  , \g253306/_0_  , \g253307/_3_  , \g253308/_0_  , \g253309/_0_  , \g253310/_0_  , \g253311/_0_  , \g253356/_0_  , \g253357/_0_  , \g253358/_0_  , \g253359/_0_  , \g253436/_3_  , \g253437/_0_  , \g253438/_0_  , \g253469/_3_  , \g253470/_3_  , \g253471/_3_  , \g253521/_0_  , \g253522/_0_  , \g253523/_0_  , \g253524/_3_  , \g256730/_3_  , \g256731/_3_  , \g256927/_0_  , \g256928/_0_  , \g256929/_3_  , \g257049/_0_  , \g257050/_0_  , \g257051/_3_  , \g257052/_0_  , \g257053/_0_  , \g257054/_0_  , \g257055/_3_  , \g257056/_0_  , \g257057/_0_  , \g257058/_3_  , \g257059/_0_  , \g257060/_0_  , \g257082/_0_  , \g257125/_3_  , \g257126/_0_  , \g257127/_0_  , \g257128/_3_  , \g257129/_3_  , \g257130/_0_  , \g257131/_0_  , \g257132/_0_  , \g257163/_0_  , \g257164/_0_  , \g257165/_0_  , \g257166/_0_  , \g257167/_0_  , \g257194/_0_  , \g258552/_0_  , \g258850/_0_  , \g258851/_3_  , \g258993/_0_  , \g258994/_0_  , \g258995/_0_  , \g258996/_0_  , \g259026/_3_  , \g259027/_0_  , \g259105/_0_  , \g259106/_0_  , \g259107/_3_  , \g259108/_0_  , \g259109/_3_  , \g259110/_0_  , \g259111/_0_  , \g259112/_0_  , \g259113/_0_  , \g259114/_0_  , \g259115/_0_  , \g259116/_0_  , \g259117/_0_  , \g259163/_3_  , \g259164/_3_  , \g259165/_0_  , \g259166/_0_  , \g259167/_0_  , \g259168/_0_  , \g259197/_0_  , \g259198/_0_  , \g259199/_0_  , \g259200/_0_  , \g260774/_0_  , \g260792/_3_  , \g260991/_0_  , \g261013/_0_  , \g261070/_0_  , \g261125/_0_  , \g261126/_0_  , \g261128/_0_  , \g261129/_0_  , \g261130/_0_  , \g261131/_0_  , \g261132/_0_  , \g261133/_0_  , \g261134/_3_  , \g261135/_0_  , \g261136/_0_  , \g261158/_3_  , \g261206/_0_  , \g261207/_0_  , \g261208/_0_  , \g261209/_0_  , \g261210/_3_  , \g261211/_0_  , \g261212/_3_  , \g261213/_0_  , \g261248/_0_  , \g261249/_0_  , \g261250/_0_  , \g261251/_0_  , \g261252/_0_  , \g261279/_0_  , \g262658/_3_  , \g262949/_0_  , \g263008/_3_  , \g263092/_0_  , \g263093/_0_  , \g263099/_0_  , \g263100/_0_  , \g263101/_0_  , \g263159/_3_  , \g263204/_3_  , \g263205/_0_  , \g263206/_0_  , \g263208/_0_  , \g263209/_0_  , \g263210/_0_  , \g263211/_0_  , \g263212/_0_  , \g263213/_0_  , \g263214/_0_  , \g263215/_3_  , \g263216/_0_  , \g263260/_0_  , \g263261/_0_  , \g263262/_3_  , \g263263/_0_  , \g263264/_0_  , \g263265/_0_  , \g263297/_0_  , \g263298/_0_  , \g263299/_0_  , \g263300/_0_  , \g264930/_0_  , \g264946/_3_  , \g265143/_0_  , \g265144/_0_  , \g265152/_0_  , \g265222/_0_  , \g265223/_0_  , \g265224/_0_  , \g265225/_0_  , \g265226/_0_  , \g265227/_3_  , \g265228/_0_  , \g265229/_0_  , \g265230/_0_  , \g265231/_0_  , \g265232/_0_  , \g265233/_3_  , \g265234/_0_  , \g265306/_0_  , \g265307/_0_  , \g265308/_3_  , \g265309/_3_  , \g265310/_0_  , \g265311/_0_  , \g265312/_0_  , \g265313/_0_  , \g265348/_0_  , \g265349/_0_  , \g265350/_0_  , \g265351/_0_  , \g265379/_0_  , \g266965/_3_  , \g267049/_3_  , \g267050/_0_  , \g267215/_0_  , \g267216/_0_  , \g267263/_0_  , \g267264/_3_  , \g267265/_0_  , \g267266/_0_  , \g267314/_3_  , \g267315/_0_  , \g267316/_0_  , \g267317/_0_  , \g267318/_0_  , \g267319/_0_  , \g267320/_3_  , \g267321/_0_  , \g267322/_0_  , \g267324/_0_  , \g267325/_0_  , \g267326/_0_  , \g267372/_0_  , \g267373/_3_  , \g267374/_0_  , \g267375/_0_  , \g267376/_0_  , \g267377/_0_  , \g267409/_0_  , \g267410/_0_  , \g267411/_0_  , \g267412/_0_  , \g269004/_0_  , \g269099/_3_  , \g269202/_0_  , \g269226/_0_  , \g269333/_3_  , \g269334/_0_  , \g269335/_0_  , \g269355/_0_  , \g269356/_0_  , \g269357/_3_  , \g269358/_0_  , \g269359/_0_  , \g269360/_0_  , \g269361/_0_  , \g269362/_0_  , \g269363/_0_  , \g269364/_0_  , \g269414/_0_  , \g269415/_0_  , \g269416/_0_  , \g269417/_0_  , \g269418/_3_  , \g269419/_0_  , \g269420/_3_  , \g269421/_0_  , \g269456/_0_  , \g269457/_0_  , \g269458/_0_  , \g269459/_0_  , \g269460/_0_  , \g269487/_0_  , \g271006/_3_  , \g271186/_3_  , \g271187/_0_  , \g271299/_0_  , \g271300/_0_  , \g271301/_3_  , \g271302/_0_  , \g271303/_0_  , \g271352/_0_  , \g271410/_0_  , \g271411/_0_  , \g271412/_0_  , \g271413/_0_  , \g271414/_0_  , \g271415/_0_  , \g271416/_0_  , \g271417/_3_  , \g271418/_3_  , \g271419/_0_  , \g271420/_0_  , \g271421/_0_  , \g271422/_0_  , \g271468/_3_  , \g271469/_0_  , \g271470/_0_  , \g271471/_0_  , \g271472/_0_  , \g271473/_0_  , \g271505/_0_  , \g271506/_0_  , \g271507/_0_  , \g271508/_0_  , \g273135/_0_  , \g273136/_3_  , \g273362/_0_  , \g273373/_0_  , \g273374/_0_  , \g273431/_0_  , \g273432/_0_  , \g273433/_3_  , \g273434/_0_  , \g273435/_0_  , \g273436/_0_  , \g273437/_3_  , \g273438/_0_  , \g273439/_0_  , \g273441/_0_  , \g273442/_0_  , \g273443/_0_  , \g273515/_3_  , \g273516/_0_  , \g273517/_0_  , \g273518/_3_  , \g273519/_0_  , \g273520/_0_  , \g273521/_0_  , \g273522/_0_  , \g273557/_0_  , \g273558/_0_  , \g273559/_0_  , \g273560/_0_  , \g273561/_0_  , \g273588/_0_  , \g274960/_3_  , \g275266/_3_  , \g275327/_0_  , \g275396/_0_  , \g275397/_3_  , \g275398/_0_  , \g275455/_0_  , \g275456/_0_  , \g275463/_0_  , \g275510/_3_  , \g275511/_0_  , \g275512/_0_  , \g275513/_0_  , \g275514/_3_  , \g275515/_0_  , \g275516/_0_  , \g275517/_0_  , \g275518/_0_  , \g275519/_0_  , \g275520/_0_  , \g275521/_0_  , \g275522/_0_  , \g275568/_0_  , \g275569/_0_  , \g275570/_0_  , \g275571/_0_  , \g275572/_3_  , \g275573/_0_  , \g275605/_0_  , \g275606/_0_  , \g275607/_0_  , \g275608/_0_  , \g277189/_0_  , \g277294/_3_  , \g277367/_0_  , \g277456/_0_  , \g277457/_0_  , \g277512/_0_  , \g277513/_0_  , \g277514/_3_  , \g277515/_0_  , \g277516/_0_  , \g277517/_3_  , \g277518/_0_  , \g277519/_0_  , \g277520/_0_  , \g277521/_0_  , \g277594/_0_  , \g277595/_0_  , \g277596/_3_  , \g277597/_0_  , \g277598/_0_  , \g277599/_0_  , \g277600/_0_  , \g277601/_3_  , \g277635/_0_  , \g277636/_0_  , \g277637/_0_  , \g277638/_0_  , \g277639/_0_  , \g277666/_0_  , \g279090/_3_  , \g279330/_0_  , \g279331/_0_  , \g279493/_3_  , \g279494/_0_  , \g279495/_0_  , \g279502/_0_  , \g279503/_0_  , \g279504/_0_  , \g279590/_0_  , \g279591/_0_  , \g279592/_0_  , \g279593/_0_  , \g279594/_3_  , \g279595/_3_  , \g279596/_0_  , \g279597/_0_  , \g279598/_0_  , \g279599/_0_  , \g279600/_0_  , \g279601/_0_  , \g279602/_0_  , \g279649/_0_  , \g279650/_0_  , \g279651/_0_  , \g279652/_0_  , \g279653/_0_  , \g279654/_3_  , \g279686/_0_  , \g279687/_0_  , \g279688/_0_  , \g279689/_0_  , \g281329/_0_  , \g281394/_0_  , \g281483/_0_  , \g281498/_0_  , \g281532/_0_  , \g281616/_0_  , \g281617/_0_  , \g281618/_0_  , \g281619/_0_  , \g281620/_0_  , \g281621/_0_  , \g281622/_0_  , \g281623/_3_  , \g281624/_0_  , \g281642/_0_  , \g281643/_0_  , \g281644/_3_  , \g281645/_0_  , \g281696/_0_  , \g281697/_3_  , \g281698/_0_  , \g281699/_0_  , \g281700/_0_  , \g281701/_0_  , \g281702/_3_  , \g281703/_0_  , \g281799/_0_  , \g281800/_0_  , \g281801/_0_  , \g281802/_0_  , \g281803/_0_  , \g281965/_0_  , \g287377/_0_  , \g287867/_0_  , \g287899/_0_  , \g288304/_0_  , \g288334/_0_  , \g288350/_0_  , \g288351/_0_  , \g288352/_3_  , \g288353/_0_  , \g288668/_0_  , \g288669/_0_  , \g288670/_0_  , \g288671/_0_  , \g288673/_0_  , \g288674/_3_  , \g288675/_0_  , \g288676/_0_  , \g288677/_0_  , \g288678/_0_  , \g288679/_0_  , \g288680/_3_  , \g288889/_0_  , \g288890/_0_  , \g288891/_0_  , \g288892/_0_  , \g288893/_3_  , \g288894/_0_  , \g288895/_0_  , \g288984/_0_  , \g288985/_0_  , \g288986/_0_  , \g294974/_0_  , \g295054/_0_  , \g295601/_0_  , \g295607/_0_  , \g296036/_0_  , \g296037/_0_  , \g296038/_0_  , \g296039/_0_  , \g296040/_0_  , \g296041/_0_  , \g296042/_0_  , \g296043/_3_  , \g296044/_0_  , \g296045/_0_  , \g296046/_0_  , \g296047/_0_  , \g296048/_0_  , \g296049/_3_  , \g296522/_3_  , \g296523/_3_  , \g296524/_0_  , \g296525/_0_  , \g296526/_0_  , \g296527/_0_  , \g296528/_3_  , \g296529/_0_  , \g296530/_0_  , \g296531/_0_  , \g297026/_0_  , \g297027/_0_  , \g305620/_3_  , \g305621/_3_  , \g305622/_3_  , \g305623/_3_  , \g305624/_3_  , \g305625/_3_  , \g305626/_3_  , \g305627/_3_  , \g305628/_3_  , \g305629/_3_  , \g305630/_3_  , \g305631/_3_  , \g305632/_3_  , \g305633/_3_  , \g305634/_3_  , \g305635/_3_  , \g305636/_3_  , \g305637/_3_  , \g305638/_3_  , \g305639/_3_  , \g305640/_3_  , \g305641/_3_  , \g305642/_3_  , \g305643/_3_  , \g305644/_3_  , \g305645/_3_  , \g305646/_3_  , \g305647/_3_  , \g305648/_3_  , \g305649/_3_  , \g305650/_3_  , \g305651/_3_  , \g305652/_3_  , \g305653/_3_  , \g305654/_3_  , \g305655/_3_  , \g305656/_3_  , \g305657/_3_  , \g305658/_3_  , \g305659/_3_  , \g305660/_3_  , \g305661/_3_  , \g305662/_3_  , \g305663/_3_  , \g305664/_3_  , \g305665/_3_  , \g305666/_3_  , \g305667/_3_  , \g305668/_3_  , \g305669/_3_  , \g305670/_3_  , \g305671/_3_  , \g305672/_3_  , \g305673/_3_  , \g305674/_3_  , \g305675/_3_  , \g305676/_3_  , \g305677/_3_  , \g305678/_3_  , \g305679/_3_  , \g305680/_3_  , \g305681/_3_  , \g305682/_3_  , \g305683/_3_  , \g305684/_3_  , \g305685/_3_  , \g305686/_3_  , \g305687/_3_  , \g305688/_3_  , \g305689/_3_  , \g305690/_3_  , \g305691/_3_  , \g305692/_3_  , \g305693/_3_  , \g305694/_3_  , \g305695/_3_  , \g305696/_3_  , \g305697/_3_  , \g305698/_3_  , \g305699/_3_  , \g305700/_3_  , \g305701/_3_  , \g305702/_3_  , \g305703/_3_  , \g305704/_3_  , \g305705/_3_  , \g305706/_3_  , \g305707/_3_  , \g305708/_3_  , \g305709/_3_  , \g305710/_3_  , \g305711/_3_  , \g305712/_3_  , \g305713/_3_  , \g305714/_3_  , \g305715/_3_  , \g305716/_3_  , \g305717/_3_  , \g305718/_3_  , \g305719/_3_  , \g305720/_3_  , \g305721/_3_  , \g305722/_3_  , \g305723/_3_  , \g305724/_3_  , \g305725/_3_  , \g305726/_3_  , \g305727/_3_  , \g305728/_3_  , \g305729/_3_  , \g305730/_3_  , \g305731/_3_  , \g321371/_0_  , \g321424/_0_  , \g321474/_3_  , \g321637/_3_  , \g321688/_0_  , \g321712/_0_  , \g321772/_3_  , \g321832/_0_  , \g321999/_0_  , \g322013/_3_  , \g322109/_0_  , \g322184/_0_  , \g322250/_0_  , \g322274/_0_  , \g322293/_3_  , \g322437/_0_  , \g322537/_3_  , \g322584/_0_  , \g322830/_0_  , \g322871/_0_  , \g322882/_0_  , \g322933/_0_  , \g323004/_0_  , \g323104/_0_  , \g323125/_0_  , \g323138/_3_  , \g323273/_0_  , \u0_desOut_reg[0]/_05_  , \u0_desOut_reg[12]/_05_  , \u0_desOut_reg[14]/_05_  , \u0_desOut_reg[18]/_05_  , \u0_desOut_reg[20]/_05_  , \u0_desOut_reg[24]/_05_  , \u0_desOut_reg[26]/_05_  , \u0_desOut_reg[28]/_05_  , \u0_desOut_reg[2]/_05_  , \u0_desOut_reg[30]/_05_  , \u0_desOut_reg[32]/_05_  , \u0_desOut_reg[34]/_05_  , \u0_desOut_reg[36]/_05_  , \u0_desOut_reg[42]/_05_  , \u0_desOut_reg[44]/_05_  , \u0_desOut_reg[46]/_05_  , \u0_desOut_reg[48]/_05_  , \u0_desOut_reg[54]/_05_  , \u0_desOut_reg[56]/_05_  , \u0_desOut_reg[62]/_05_  , \u0_desOut_reg[6]/_05_  , \u0_desOut_reg[8]/_05_  , \u1_desOut_reg[0]/_05_  , \u1_desOut_reg[12]/_05_  , \u1_desOut_reg[14]/_05_  , \u1_desOut_reg[16]/_05_  , \u1_desOut_reg[18]/_05_  , \u1_desOut_reg[20]/_05_  , \u1_desOut_reg[22]/_05_  , \u1_desOut_reg[24]/_05_  , \u1_desOut_reg[26]/_05_  , \u1_desOut_reg[28]/_05_  , \u1_desOut_reg[2]/_05_  , \u1_desOut_reg[30]/_05_  , \u1_desOut_reg[32]/_05_  , \u1_desOut_reg[34]/_05_  , \u1_desOut_reg[36]/_05_  , \u1_desOut_reg[38]/_05_  , \u1_desOut_reg[42]/_05_  , \u1_desOut_reg[44]/_05_  , \u1_desOut_reg[46]/_05_  , \u1_desOut_reg[48]/_05_  , \u1_desOut_reg[4]/_05_  , \u1_desOut_reg[54]/_05_  , \u1_desOut_reg[56]/_05_  , \u1_desOut_reg[58]/_05_  , \u1_desOut_reg[60]/_05_  , \u1_desOut_reg[62]/_05_  , \u1_desOut_reg[6]/_05_  , \u1_desOut_reg[8]/_05_  , \u2_desOut_reg[0]/_05_  , \u2_desOut_reg[10]/_05_  , \u2_desOut_reg[12]/_05_  , \u2_desOut_reg[14]/_05_  , \u2_desOut_reg[16]/_05_  , \u2_desOut_reg[18]/_05_  , \u2_desOut_reg[20]/_05_  , \u2_desOut_reg[22]/_05_  , \u2_desOut_reg[24]/_05_  , \u2_desOut_reg[26]/_05_  , \u2_desOut_reg[28]/_05_  , \u2_desOut_reg[2]/_05_  , \u2_desOut_reg[30]/_05_  , \u2_desOut_reg[32]/_05_  , \u2_desOut_reg[34]/_05_  , \u2_desOut_reg[36]/_05_  , \u2_desOut_reg[38]/_05_  , \u2_desOut_reg[40]/_05_  , \u2_desOut_reg[42]/_05_  , \u2_desOut_reg[44]/_05_  , \u2_desOut_reg[46]/_05_  , \u2_desOut_reg[48]/_05_  , \u2_desOut_reg[4]/_05_  , \u2_desOut_reg[50]/_05_  , \u2_desOut_reg[52]/_05_  , \u2_desOut_reg[54]/_05_  , \u2_desOut_reg[56]/_05_  , \u2_desOut_reg[58]/_05_  , \u2_desOut_reg[60]/_05_  , \u2_desOut_reg[62]/_05_  , \u2_desOut_reg[6]/_05_  , \u2_desOut_reg[8]/_05_  );
  input decrypt_pad ;
  input \key1[0]_pad  ;
  input \key1[10]_pad  ;
  input \key1[11]_pad  ;
  input \key1[12]_pad  ;
  input \key1[13]_pad  ;
  input \key1[14]_pad  ;
  input \key1[15]_pad  ;
  input \key1[16]_pad  ;
  input \key1[17]_pad  ;
  input \key1[18]_pad  ;
  input \key1[19]_pad  ;
  input \key1[1]_pad  ;
  input \key1[20]_pad  ;
  input \key1[21]_pad  ;
  input \key1[22]_pad  ;
  input \key1[23]_pad  ;
  input \key1[24]_pad  ;
  input \key1[25]_pad  ;
  input \key1[26]_pad  ;
  input \key1[27]_pad  ;
  input \key1[28]_pad  ;
  input \key1[29]_pad  ;
  input \key1[2]_pad  ;
  input \key1[30]_pad  ;
  input \key1[31]_pad  ;
  input \key1[32]_pad  ;
  input \key1[33]_pad  ;
  input \key1[34]_pad  ;
  input \key1[35]_pad  ;
  input \key1[36]_pad  ;
  input \key1[37]_pad  ;
  input \key1[38]_pad  ;
  input \key1[39]_pad  ;
  input \key1[3]_pad  ;
  input \key1[40]_pad  ;
  input \key1[41]_pad  ;
  input \key1[42]_pad  ;
  input \key1[43]_pad  ;
  input \key1[44]_pad  ;
  input \key1[45]_pad  ;
  input \key1[46]_pad  ;
  input \key1[47]_pad  ;
  input \key1[48]_pad  ;
  input \key1[49]_pad  ;
  input \key1[4]_pad  ;
  input \key1[50]_pad  ;
  input \key1[51]_pad  ;
  input \key1[52]_pad  ;
  input \key1[53]_pad  ;
  input \key1[54]_pad  ;
  input \key1[55]_pad  ;
  input \key1[5]_pad  ;
  input \key1[6]_pad  ;
  input \key1[7]_pad  ;
  input \key1[8]_pad  ;
  input \key1[9]_pad  ;
  input \key3[0]_pad  ;
  input \key3[10]_pad  ;
  input \key3[11]_pad  ;
  input \key3[12]_pad  ;
  input \key3[13]_pad  ;
  input \key3[14]_pad  ;
  input \key3[15]_pad  ;
  input \key3[16]_pad  ;
  input \key3[17]_pad  ;
  input \key3[18]_pad  ;
  input \key3[19]_pad  ;
  input \key3[1]_pad  ;
  input \key3[20]_pad  ;
  input \key3[21]_pad  ;
  input \key3[22]_pad  ;
  input \key3[23]_pad  ;
  input \key3[24]_pad  ;
  input \key3[25]_pad  ;
  input \key3[26]_pad  ;
  input \key3[27]_pad  ;
  input \key3[28]_pad  ;
  input \key3[29]_pad  ;
  input \key3[2]_pad  ;
  input \key3[30]_pad  ;
  input \key3[31]_pad  ;
  input \key3[32]_pad  ;
  input \key3[33]_pad  ;
  input \key3[34]_pad  ;
  input \key3[35]_pad  ;
  input \key3[36]_pad  ;
  input \key3[37]_pad  ;
  input \key3[38]_pad  ;
  input \key3[39]_pad  ;
  input \key3[3]_pad  ;
  input \key3[40]_pad  ;
  input \key3[41]_pad  ;
  input \key3[42]_pad  ;
  input \key3[43]_pad  ;
  input \key3[44]_pad  ;
  input \key3[45]_pad  ;
  input \key3[46]_pad  ;
  input \key3[47]_pad  ;
  input \key3[48]_pad  ;
  input \key3[49]_pad  ;
  input \key3[4]_pad  ;
  input \key3[50]_pad  ;
  input \key3[51]_pad  ;
  input \key3[52]_pad  ;
  input \key3[53]_pad  ;
  input \key3[54]_pad  ;
  input \key3[55]_pad  ;
  input \key3[5]_pad  ;
  input \key3[6]_pad  ;
  input \key3[7]_pad  ;
  input \key3[8]_pad  ;
  input \key3[9]_pad  ;
  input \u0_L0_reg[10]/NET0131  ;
  input \u0_L0_reg[11]/NET0131  ;
  input \u0_L0_reg[12]/NET0131  ;
  input \u0_L0_reg[13]/NET0131  ;
  input \u0_L0_reg[14]/NET0131  ;
  input \u0_L0_reg[15]/P0001  ;
  input \u0_L0_reg[16]/NET0131  ;
  input \u0_L0_reg[17]/NET0131  ;
  input \u0_L0_reg[18]/NET0131  ;
  input \u0_L0_reg[19]/P0001  ;
  input \u0_L0_reg[1]/NET0131  ;
  input \u0_L0_reg[20]/NET0131  ;
  input \u0_L0_reg[21]/NET0131  ;
  input \u0_L0_reg[22]/NET0131  ;
  input \u0_L0_reg[23]/NET0131  ;
  input \u0_L0_reg[24]/NET0131  ;
  input \u0_L0_reg[25]/NET0131  ;
  input \u0_L0_reg[26]/NET0131  ;
  input \u0_L0_reg[27]/NET0131  ;
  input \u0_L0_reg[28]/NET0131  ;
  input \u0_L0_reg[29]/NET0131  ;
  input \u0_L0_reg[2]/NET0131  ;
  input \u0_L0_reg[30]/P0001  ;
  input \u0_L0_reg[31]/NET0131  ;
  input \u0_L0_reg[32]/NET0131  ;
  input \u0_L0_reg[3]/NET0131  ;
  input \u0_L0_reg[4]/NET0131  ;
  input \u0_L0_reg[5]/NET0131  ;
  input \u0_L0_reg[6]/NET0131  ;
  input \u0_L0_reg[7]/NET0131  ;
  input \u0_L0_reg[8]/NET0131  ;
  input \u0_L0_reg[9]/NET0131  ;
  input \u0_L10_reg[10]/NET0131  ;
  input \u0_L10_reg[11]/NET0131  ;
  input \u0_L10_reg[12]/NET0131  ;
  input \u0_L10_reg[13]/NET0131  ;
  input \u0_L10_reg[14]/NET0131  ;
  input \u0_L10_reg[15]/P0001  ;
  input \u0_L10_reg[16]/NET0131  ;
  input \u0_L10_reg[17]/NET0131  ;
  input \u0_L10_reg[18]/NET0131  ;
  input \u0_L10_reg[19]/NET0131  ;
  input \u0_L10_reg[1]/NET0131  ;
  input \u0_L10_reg[20]/NET0131  ;
  input \u0_L10_reg[21]/NET0131  ;
  input \u0_L10_reg[22]/NET0131  ;
  input \u0_L10_reg[23]/NET0131  ;
  input \u0_L10_reg[24]/NET0131  ;
  input \u0_L10_reg[25]/NET0131  ;
  input \u0_L10_reg[26]/NET0131  ;
  input \u0_L10_reg[27]/NET0131  ;
  input \u0_L10_reg[28]/NET0131  ;
  input \u0_L10_reg[29]/NET0131  ;
  input \u0_L10_reg[2]/NET0131  ;
  input \u0_L10_reg[30]/NET0131  ;
  input \u0_L10_reg[31]/NET0131  ;
  input \u0_L10_reg[32]/NET0131  ;
  input \u0_L10_reg[3]/NET0131  ;
  input \u0_L10_reg[4]/NET0131  ;
  input \u0_L10_reg[5]/NET0131  ;
  input \u0_L10_reg[6]/NET0131  ;
  input \u0_L10_reg[7]/NET0131  ;
  input \u0_L10_reg[8]/NET0131  ;
  input \u0_L10_reg[9]/NET0131  ;
  input \u0_L11_reg[10]/NET0131  ;
  input \u0_L11_reg[11]/P0001  ;
  input \u0_L11_reg[12]/NET0131  ;
  input \u0_L11_reg[13]/NET0131  ;
  input \u0_L11_reg[14]/NET0131  ;
  input \u0_L11_reg[15]/P0001  ;
  input \u0_L11_reg[16]/NET0131  ;
  input \u0_L11_reg[17]/NET0131  ;
  input \u0_L11_reg[18]/NET0131  ;
  input \u0_L11_reg[19]/NET0131  ;
  input \u0_L11_reg[1]/NET0131  ;
  input \u0_L11_reg[20]/NET0131  ;
  input \u0_L11_reg[21]/NET0131  ;
  input \u0_L11_reg[22]/NET0131  ;
  input \u0_L11_reg[23]/NET0131  ;
  input \u0_L11_reg[24]/NET0131  ;
  input \u0_L11_reg[25]/NET0131  ;
  input \u0_L11_reg[26]/NET0131  ;
  input \u0_L11_reg[27]/NET0131  ;
  input \u0_L11_reg[28]/NET0131  ;
  input \u0_L11_reg[29]/NET0131  ;
  input \u0_L11_reg[2]/NET0131  ;
  input \u0_L11_reg[30]/NET0131  ;
  input \u0_L11_reg[31]/NET0131  ;
  input \u0_L11_reg[32]/NET0131  ;
  input \u0_L11_reg[3]/NET0131  ;
  input \u0_L11_reg[4]/NET0131  ;
  input \u0_L11_reg[5]/NET0131  ;
  input \u0_L11_reg[6]/NET0131  ;
  input \u0_L11_reg[7]/NET0131  ;
  input \u0_L11_reg[8]/NET0131  ;
  input \u0_L11_reg[9]/NET0131  ;
  input \u0_L12_reg[10]/NET0131  ;
  input \u0_L12_reg[11]/NET0131  ;
  input \u0_L12_reg[12]/NET0131  ;
  input \u0_L12_reg[13]/NET0131  ;
  input \u0_L12_reg[14]/NET0131  ;
  input \u0_L12_reg[15]/P0001  ;
  input \u0_L12_reg[16]/NET0131  ;
  input \u0_L12_reg[17]/NET0131  ;
  input \u0_L12_reg[18]/NET0131  ;
  input \u0_L12_reg[19]/P0001  ;
  input \u0_L12_reg[1]/NET0131  ;
  input \u0_L12_reg[20]/NET0131  ;
  input \u0_L12_reg[21]/NET0131  ;
  input \u0_L12_reg[22]/NET0131  ;
  input \u0_L12_reg[23]/NET0131  ;
  input \u0_L12_reg[24]/NET0131  ;
  input \u0_L12_reg[25]/NET0131  ;
  input \u0_L12_reg[26]/NET0131  ;
  input \u0_L12_reg[27]/NET0131  ;
  input \u0_L12_reg[28]/NET0131  ;
  input \u0_L12_reg[29]/NET0131  ;
  input \u0_L12_reg[2]/NET0131  ;
  input \u0_L12_reg[30]/NET0131  ;
  input \u0_L12_reg[31]/NET0131  ;
  input \u0_L12_reg[32]/NET0131  ;
  input \u0_L12_reg[3]/NET0131  ;
  input \u0_L12_reg[4]/NET0131  ;
  input \u0_L12_reg[5]/NET0131  ;
  input \u0_L12_reg[6]/NET0131  ;
  input \u0_L12_reg[7]/NET0131  ;
  input \u0_L12_reg[8]/NET0131  ;
  input \u0_L12_reg[9]/NET0131  ;
  input \u0_L13_reg[10]/NET0131  ;
  input \u0_L13_reg[11]/NET0131  ;
  input \u0_L13_reg[12]/NET0131  ;
  input \u0_L13_reg[13]/NET0131  ;
  input \u0_L13_reg[14]/NET0131  ;
  input \u0_L13_reg[15]/P0001  ;
  input \u0_L13_reg[16]/NET0131  ;
  input \u0_L13_reg[17]/NET0131  ;
  input \u0_L13_reg[18]/NET0131  ;
  input \u0_L13_reg[19]/NET0131  ;
  input \u0_L13_reg[1]/NET0131  ;
  input \u0_L13_reg[20]/NET0131  ;
  input \u0_L13_reg[21]/NET0131  ;
  input \u0_L13_reg[22]/NET0131  ;
  input \u0_L13_reg[23]/NET0131  ;
  input \u0_L13_reg[24]/NET0131  ;
  input \u0_L13_reg[25]/NET0131  ;
  input \u0_L13_reg[26]/NET0131  ;
  input \u0_L13_reg[27]/NET0131  ;
  input \u0_L13_reg[28]/NET0131  ;
  input \u0_L13_reg[29]/NET0131  ;
  input \u0_L13_reg[2]/NET0131  ;
  input \u0_L13_reg[30]/NET0131  ;
  input \u0_L13_reg[31]/NET0131  ;
  input \u0_L13_reg[32]/NET0131  ;
  input \u0_L13_reg[3]/NET0131  ;
  input \u0_L13_reg[4]/NET0131  ;
  input \u0_L13_reg[5]/NET0131  ;
  input \u0_L13_reg[6]/NET0131  ;
  input \u0_L13_reg[7]/NET0131  ;
  input \u0_L13_reg[8]/NET0131  ;
  input \u0_L13_reg[9]/NET0131  ;
  input \u0_L14_reg[10]/P0001  ;
  input \u0_L14_reg[11]/P0001  ;
  input \u0_L14_reg[12]/P0001  ;
  input \u0_L14_reg[13]/P0001  ;
  input \u0_L14_reg[14]/P0001  ;
  input \u0_L14_reg[15]/P0001  ;
  input \u0_L14_reg[16]/P0001  ;
  input \u0_L14_reg[17]/P0001  ;
  input \u0_L14_reg[18]/P0001  ;
  input \u0_L14_reg[19]/P0001  ;
  input \u0_L14_reg[1]/P0001  ;
  input \u0_L14_reg[20]/P0001  ;
  input \u0_L14_reg[21]/P0001  ;
  input \u0_L14_reg[22]/P0001  ;
  input \u0_L14_reg[23]/P0001  ;
  input \u0_L14_reg[24]/P0001  ;
  input \u0_L14_reg[25]/P0001  ;
  input \u0_L14_reg[26]/P0001  ;
  input \u0_L14_reg[27]/P0001  ;
  input \u0_L14_reg[28]/P0001  ;
  input \u0_L14_reg[29]/P0001  ;
  input \u0_L14_reg[2]/P0001  ;
  input \u0_L14_reg[30]/P0001  ;
  input \u0_L14_reg[31]/P0001  ;
  input \u0_L14_reg[32]/P0001  ;
  input \u0_L14_reg[3]/P0001  ;
  input \u0_L14_reg[4]/P0001  ;
  input \u0_L14_reg[5]/P0001  ;
  input \u0_L14_reg[6]/P0001  ;
  input \u0_L14_reg[7]/P0001  ;
  input \u0_L14_reg[8]/P0001  ;
  input \u0_L14_reg[9]/P0001  ;
  input \u0_L1_reg[10]/NET0131  ;
  input \u0_L1_reg[11]/NET0131  ;
  input \u0_L1_reg[12]/NET0131  ;
  input \u0_L1_reg[13]/NET0131  ;
  input \u0_L1_reg[14]/NET0131  ;
  input \u0_L1_reg[15]/P0001  ;
  input \u0_L1_reg[16]/NET0131  ;
  input \u0_L1_reg[17]/NET0131  ;
  input \u0_L1_reg[18]/NET0131  ;
  input \u0_L1_reg[19]/NET0131  ;
  input \u0_L1_reg[1]/NET0131  ;
  input \u0_L1_reg[20]/NET0131  ;
  input \u0_L1_reg[21]/NET0131  ;
  input \u0_L1_reg[22]/NET0131  ;
  input \u0_L1_reg[23]/NET0131  ;
  input \u0_L1_reg[24]/NET0131  ;
  input \u0_L1_reg[25]/NET0131  ;
  input \u0_L1_reg[26]/NET0131  ;
  input \u0_L1_reg[27]/NET0131  ;
  input \u0_L1_reg[28]/NET0131  ;
  input \u0_L1_reg[29]/NET0131  ;
  input \u0_L1_reg[2]/NET0131  ;
  input \u0_L1_reg[30]/NET0131  ;
  input \u0_L1_reg[31]/NET0131  ;
  input \u0_L1_reg[32]/NET0131  ;
  input \u0_L1_reg[3]/NET0131  ;
  input \u0_L1_reg[4]/NET0131  ;
  input \u0_L1_reg[5]/NET0131  ;
  input \u0_L1_reg[6]/NET0131  ;
  input \u0_L1_reg[7]/NET0131  ;
  input \u0_L1_reg[8]/NET0131  ;
  input \u0_L1_reg[9]/NET0131  ;
  input \u0_L2_reg[10]/NET0131  ;
  input \u0_L2_reg[11]/NET0131  ;
  input \u0_L2_reg[12]/NET0131  ;
  input \u0_L2_reg[13]/NET0131  ;
  input \u0_L2_reg[14]/NET0131  ;
  input \u0_L2_reg[15]/P0001  ;
  input \u0_L2_reg[16]/NET0131  ;
  input \u0_L2_reg[17]/NET0131  ;
  input \u0_L2_reg[18]/NET0131  ;
  input \u0_L2_reg[19]/P0001  ;
  input \u0_L2_reg[1]/NET0131  ;
  input \u0_L2_reg[20]/NET0131  ;
  input \u0_L2_reg[21]/NET0131  ;
  input \u0_L2_reg[22]/NET0131  ;
  input \u0_L2_reg[23]/NET0131  ;
  input \u0_L2_reg[24]/NET0131  ;
  input \u0_L2_reg[25]/NET0131  ;
  input \u0_L2_reg[26]/NET0131  ;
  input \u0_L2_reg[27]/NET0131  ;
  input \u0_L2_reg[28]/NET0131  ;
  input \u0_L2_reg[29]/NET0131  ;
  input \u0_L2_reg[2]/NET0131  ;
  input \u0_L2_reg[30]/NET0131  ;
  input \u0_L2_reg[31]/NET0131  ;
  input \u0_L2_reg[32]/NET0131  ;
  input \u0_L2_reg[3]/NET0131  ;
  input \u0_L2_reg[4]/NET0131  ;
  input \u0_L2_reg[5]/NET0131  ;
  input \u0_L2_reg[6]/NET0131  ;
  input \u0_L2_reg[7]/NET0131  ;
  input \u0_L2_reg[8]/NET0131  ;
  input \u0_L2_reg[9]/NET0131  ;
  input \u0_L3_reg[10]/NET0131  ;
  input \u0_L3_reg[11]/NET0131  ;
  input \u0_L3_reg[12]/NET0131  ;
  input \u0_L3_reg[13]/NET0131  ;
  input \u0_L3_reg[14]/NET0131  ;
  input \u0_L3_reg[15]/P0001  ;
  input \u0_L3_reg[16]/NET0131  ;
  input \u0_L3_reg[17]/NET0131  ;
  input \u0_L3_reg[18]/NET0131  ;
  input \u0_L3_reg[19]/P0001  ;
  input \u0_L3_reg[1]/NET0131  ;
  input \u0_L3_reg[20]/NET0131  ;
  input \u0_L3_reg[21]/NET0131  ;
  input \u0_L3_reg[22]/NET0131  ;
  input \u0_L3_reg[23]/NET0131  ;
  input \u0_L3_reg[24]/NET0131  ;
  input \u0_L3_reg[25]/NET0131  ;
  input \u0_L3_reg[26]/NET0131  ;
  input \u0_L3_reg[27]/NET0131  ;
  input \u0_L3_reg[28]/NET0131  ;
  input \u0_L3_reg[29]/NET0131  ;
  input \u0_L3_reg[2]/NET0131  ;
  input \u0_L3_reg[30]/NET0131  ;
  input \u0_L3_reg[31]/NET0131  ;
  input \u0_L3_reg[32]/NET0131  ;
  input \u0_L3_reg[3]/NET0131  ;
  input \u0_L3_reg[4]/NET0131  ;
  input \u0_L3_reg[5]/NET0131  ;
  input \u0_L3_reg[6]/NET0131  ;
  input \u0_L3_reg[7]/NET0131  ;
  input \u0_L3_reg[8]/NET0131  ;
  input \u0_L3_reg[9]/NET0131  ;
  input \u0_L4_reg[10]/NET0131  ;
  input \u0_L4_reg[11]/NET0131  ;
  input \u0_L4_reg[12]/NET0131  ;
  input \u0_L4_reg[13]/NET0131  ;
  input \u0_L4_reg[14]/NET0131  ;
  input \u0_L4_reg[15]/P0001  ;
  input \u0_L4_reg[16]/NET0131  ;
  input \u0_L4_reg[17]/NET0131  ;
  input \u0_L4_reg[18]/NET0131  ;
  input \u0_L4_reg[19]/NET0131  ;
  input \u0_L4_reg[1]/NET0131  ;
  input \u0_L4_reg[20]/NET0131  ;
  input \u0_L4_reg[21]/NET0131  ;
  input \u0_L4_reg[22]/NET0131  ;
  input \u0_L4_reg[23]/NET0131  ;
  input \u0_L4_reg[24]/NET0131  ;
  input \u0_L4_reg[25]/NET0131  ;
  input \u0_L4_reg[26]/NET0131  ;
  input \u0_L4_reg[27]/NET0131  ;
  input \u0_L4_reg[28]/NET0131  ;
  input \u0_L4_reg[29]/NET0131  ;
  input \u0_L4_reg[2]/NET0131  ;
  input \u0_L4_reg[30]/NET0131  ;
  input \u0_L4_reg[31]/NET0131  ;
  input \u0_L4_reg[32]/NET0131  ;
  input \u0_L4_reg[3]/NET0131  ;
  input \u0_L4_reg[4]/NET0131  ;
  input \u0_L4_reg[5]/NET0131  ;
  input \u0_L4_reg[6]/NET0131  ;
  input \u0_L4_reg[7]/NET0131  ;
  input \u0_L4_reg[8]/NET0131  ;
  input \u0_L4_reg[9]/NET0131  ;
  input \u0_L5_reg[10]/NET0131  ;
  input \u0_L5_reg[11]/NET0131  ;
  input \u0_L5_reg[12]/NET0131  ;
  input \u0_L5_reg[13]/NET0131  ;
  input \u0_L5_reg[14]/NET0131  ;
  input \u0_L5_reg[15]/P0001  ;
  input \u0_L5_reg[16]/NET0131  ;
  input \u0_L5_reg[17]/NET0131  ;
  input \u0_L5_reg[18]/NET0131  ;
  input \u0_L5_reg[19]/P0001  ;
  input \u0_L5_reg[1]/NET0131  ;
  input \u0_L5_reg[20]/NET0131  ;
  input \u0_L5_reg[21]/NET0131  ;
  input \u0_L5_reg[22]/NET0131  ;
  input \u0_L5_reg[23]/NET0131  ;
  input \u0_L5_reg[24]/NET0131  ;
  input \u0_L5_reg[25]/NET0131  ;
  input \u0_L5_reg[26]/NET0131  ;
  input \u0_L5_reg[27]/NET0131  ;
  input \u0_L5_reg[28]/NET0131  ;
  input \u0_L5_reg[29]/NET0131  ;
  input \u0_L5_reg[2]/NET0131  ;
  input \u0_L5_reg[30]/NET0131  ;
  input \u0_L5_reg[31]/NET0131  ;
  input \u0_L5_reg[32]/NET0131  ;
  input \u0_L5_reg[3]/NET0131  ;
  input \u0_L5_reg[4]/NET0131  ;
  input \u0_L5_reg[5]/NET0131  ;
  input \u0_L5_reg[6]/NET0131  ;
  input \u0_L5_reg[7]/NET0131  ;
  input \u0_L5_reg[8]/NET0131  ;
  input \u0_L5_reg[9]/NET0131  ;
  input \u0_L6_reg[10]/NET0131  ;
  input \u0_L6_reg[11]/NET0131  ;
  input \u0_L6_reg[12]/NET0131  ;
  input \u0_L6_reg[13]/NET0131  ;
  input \u0_L6_reg[14]/NET0131  ;
  input \u0_L6_reg[15]/P0001  ;
  input \u0_L6_reg[16]/NET0131  ;
  input \u0_L6_reg[17]/NET0131  ;
  input \u0_L6_reg[18]/NET0131  ;
  input \u0_L6_reg[19]/P0001  ;
  input \u0_L6_reg[1]/NET0131  ;
  input \u0_L6_reg[20]/NET0131  ;
  input \u0_L6_reg[21]/NET0131  ;
  input \u0_L6_reg[22]/NET0131  ;
  input \u0_L6_reg[23]/NET0131  ;
  input \u0_L6_reg[24]/NET0131  ;
  input \u0_L6_reg[25]/NET0131  ;
  input \u0_L6_reg[26]/NET0131  ;
  input \u0_L6_reg[27]/NET0131  ;
  input \u0_L6_reg[28]/NET0131  ;
  input \u0_L6_reg[29]/NET0131  ;
  input \u0_L6_reg[2]/NET0131  ;
  input \u0_L6_reg[30]/NET0131  ;
  input \u0_L6_reg[31]/NET0131  ;
  input \u0_L6_reg[32]/NET0131  ;
  input \u0_L6_reg[3]/NET0131  ;
  input \u0_L6_reg[4]/NET0131  ;
  input \u0_L6_reg[5]/NET0131  ;
  input \u0_L6_reg[6]/NET0131  ;
  input \u0_L6_reg[7]/NET0131  ;
  input \u0_L6_reg[8]/NET0131  ;
  input \u0_L6_reg[9]/NET0131  ;
  input \u0_L7_reg[10]/NET0131  ;
  input \u0_L7_reg[11]/NET0131  ;
  input \u0_L7_reg[12]/NET0131  ;
  input \u0_L7_reg[13]/NET0131  ;
  input \u0_L7_reg[14]/NET0131  ;
  input \u0_L7_reg[15]/P0001  ;
  input \u0_L7_reg[16]/NET0131  ;
  input \u0_L7_reg[17]/NET0131  ;
  input \u0_L7_reg[18]/NET0131  ;
  input \u0_L7_reg[19]/NET0131  ;
  input \u0_L7_reg[1]/NET0131  ;
  input \u0_L7_reg[20]/NET0131  ;
  input \u0_L7_reg[21]/NET0131  ;
  input \u0_L7_reg[22]/NET0131  ;
  input \u0_L7_reg[23]/NET0131  ;
  input \u0_L7_reg[24]/NET0131  ;
  input \u0_L7_reg[25]/NET0131  ;
  input \u0_L7_reg[26]/NET0131  ;
  input \u0_L7_reg[27]/NET0131  ;
  input \u0_L7_reg[28]/NET0131  ;
  input \u0_L7_reg[29]/NET0131  ;
  input \u0_L7_reg[2]/NET0131  ;
  input \u0_L7_reg[30]/NET0131  ;
  input \u0_L7_reg[31]/NET0131  ;
  input \u0_L7_reg[32]/NET0131  ;
  input \u0_L7_reg[3]/NET0131  ;
  input \u0_L7_reg[4]/NET0131  ;
  input \u0_L7_reg[5]/NET0131  ;
  input \u0_L7_reg[6]/NET0131  ;
  input \u0_L7_reg[7]/NET0131  ;
  input \u0_L7_reg[8]/NET0131  ;
  input \u0_L7_reg[9]/NET0131  ;
  input \u0_L8_reg[10]/NET0131  ;
  input \u0_L8_reg[11]/NET0131  ;
  input \u0_L8_reg[12]/NET0131  ;
  input \u0_L8_reg[13]/NET0131  ;
  input \u0_L8_reg[14]/NET0131  ;
  input \u0_L8_reg[15]/P0001  ;
  input \u0_L8_reg[16]/NET0131  ;
  input \u0_L8_reg[17]/NET0131  ;
  input \u0_L8_reg[18]/NET0131  ;
  input \u0_L8_reg[19]/NET0131  ;
  input \u0_L8_reg[1]/NET0131  ;
  input \u0_L8_reg[20]/NET0131  ;
  input \u0_L8_reg[21]/NET0131  ;
  input \u0_L8_reg[22]/NET0131  ;
  input \u0_L8_reg[23]/NET0131  ;
  input \u0_L8_reg[24]/NET0131  ;
  input \u0_L8_reg[25]/NET0131  ;
  input \u0_L8_reg[26]/NET0131  ;
  input \u0_L8_reg[27]/NET0131  ;
  input \u0_L8_reg[28]/NET0131  ;
  input \u0_L8_reg[29]/NET0131  ;
  input \u0_L8_reg[2]/NET0131  ;
  input \u0_L8_reg[30]/NET0131  ;
  input \u0_L8_reg[31]/NET0131  ;
  input \u0_L8_reg[32]/NET0131  ;
  input \u0_L8_reg[3]/NET0131  ;
  input \u0_L8_reg[4]/NET0131  ;
  input \u0_L8_reg[5]/NET0131  ;
  input \u0_L8_reg[6]/NET0131  ;
  input \u0_L8_reg[7]/NET0131  ;
  input \u0_L8_reg[8]/NET0131  ;
  input \u0_L8_reg[9]/NET0131  ;
  input \u0_L9_reg[10]/NET0131  ;
  input \u0_L9_reg[11]/NET0131  ;
  input \u0_L9_reg[12]/NET0131  ;
  input \u0_L9_reg[13]/NET0131  ;
  input \u0_L9_reg[14]/NET0131  ;
  input \u0_L9_reg[15]/P0001  ;
  input \u0_L9_reg[16]/NET0131  ;
  input \u0_L9_reg[17]/NET0131  ;
  input \u0_L9_reg[18]/NET0131  ;
  input \u0_L9_reg[19]/P0001  ;
  input \u0_L9_reg[1]/NET0131  ;
  input \u0_L9_reg[20]/NET0131  ;
  input \u0_L9_reg[21]/NET0131  ;
  input \u0_L9_reg[22]/NET0131  ;
  input \u0_L9_reg[23]/NET0131  ;
  input \u0_L9_reg[24]/NET0131  ;
  input \u0_L9_reg[25]/NET0131  ;
  input \u0_L9_reg[26]/NET0131  ;
  input \u0_L9_reg[27]/NET0131  ;
  input \u0_L9_reg[28]/NET0131  ;
  input \u0_L9_reg[29]/NET0131  ;
  input \u0_L9_reg[2]/NET0131  ;
  input \u0_L9_reg[30]/NET0131  ;
  input \u0_L9_reg[31]/NET0131  ;
  input \u0_L9_reg[32]/NET0131  ;
  input \u0_L9_reg[3]/NET0131  ;
  input \u0_L9_reg[4]/NET0131  ;
  input \u0_L9_reg[5]/NET0131  ;
  input \u0_L9_reg[6]/NET0131  ;
  input \u0_L9_reg[7]/NET0131  ;
  input \u0_L9_reg[8]/NET0131  ;
  input \u0_L9_reg[9]/NET0131  ;
  input \u0_R0_reg[10]/NET0131  ;
  input \u0_R0_reg[11]/NET0131  ;
  input \u0_R0_reg[12]/NET0131  ;
  input \u0_R0_reg[13]/NET0131  ;
  input \u0_R0_reg[14]/NET0131  ;
  input \u0_R0_reg[15]/NET0131  ;
  input \u0_R0_reg[16]/NET0131  ;
  input \u0_R0_reg[17]/NET0131  ;
  input \u0_R0_reg[18]/NET0131  ;
  input \u0_R0_reg[19]/NET0131  ;
  input \u0_R0_reg[1]/NET0131  ;
  input \u0_R0_reg[20]/NET0131  ;
  input \u0_R0_reg[21]/NET0131  ;
  input \u0_R0_reg[22]/NET0131  ;
  input \u0_R0_reg[23]/NET0131  ;
  input \u0_R0_reg[24]/NET0131  ;
  input \u0_R0_reg[25]/NET0131  ;
  input \u0_R0_reg[26]/NET0131  ;
  input \u0_R0_reg[27]/NET0131  ;
  input \u0_R0_reg[28]/NET0131  ;
  input \u0_R0_reg[29]/NET0131  ;
  input \u0_R0_reg[2]/NET0131  ;
  input \u0_R0_reg[30]/NET0131  ;
  input \u0_R0_reg[31]/NET0131  ;
  input \u0_R0_reg[32]/NET0131  ;
  input \u0_R0_reg[3]/NET0131  ;
  input \u0_R0_reg[4]/NET0131  ;
  input \u0_R0_reg[5]/NET0131  ;
  input \u0_R0_reg[6]/NET0131  ;
  input \u0_R0_reg[7]/NET0131  ;
  input \u0_R0_reg[8]/NET0131  ;
  input \u0_R0_reg[9]/NET0131  ;
  input \u0_R10_reg[10]/NET0131  ;
  input \u0_R10_reg[11]/NET0131  ;
  input \u0_R10_reg[12]/NET0131  ;
  input \u0_R10_reg[13]/NET0131  ;
  input \u0_R10_reg[14]/NET0131  ;
  input \u0_R10_reg[15]/NET0131  ;
  input \u0_R10_reg[16]/NET0131  ;
  input \u0_R10_reg[17]/NET0131  ;
  input \u0_R10_reg[18]/NET0131  ;
  input \u0_R10_reg[19]/NET0131  ;
  input \u0_R10_reg[1]/NET0131  ;
  input \u0_R10_reg[20]/NET0131  ;
  input \u0_R10_reg[21]/NET0131  ;
  input \u0_R10_reg[22]/NET0131  ;
  input \u0_R10_reg[23]/NET0131  ;
  input \u0_R10_reg[24]/NET0131  ;
  input \u0_R10_reg[25]/NET0131  ;
  input \u0_R10_reg[26]/NET0131  ;
  input \u0_R10_reg[27]/NET0131  ;
  input \u0_R10_reg[28]/NET0131  ;
  input \u0_R10_reg[29]/NET0131  ;
  input \u0_R10_reg[2]/NET0131  ;
  input \u0_R10_reg[30]/NET0131  ;
  input \u0_R10_reg[31]/P0001  ;
  input \u0_R10_reg[32]/NET0131  ;
  input \u0_R10_reg[3]/NET0131  ;
  input \u0_R10_reg[4]/NET0131  ;
  input \u0_R10_reg[5]/NET0131  ;
  input \u0_R10_reg[6]/NET0131  ;
  input \u0_R10_reg[7]/NET0131  ;
  input \u0_R10_reg[8]/NET0131  ;
  input \u0_R10_reg[9]/NET0131  ;
  input \u0_R11_reg[10]/NET0131  ;
  input \u0_R11_reg[11]/P0001  ;
  input \u0_R11_reg[12]/NET0131  ;
  input \u0_R11_reg[13]/NET0131  ;
  input \u0_R11_reg[14]/NET0131  ;
  input \u0_R11_reg[15]/NET0131  ;
  input \u0_R11_reg[16]/NET0131  ;
  input \u0_R11_reg[17]/NET0131  ;
  input \u0_R11_reg[18]/NET0131  ;
  input \u0_R11_reg[19]/NET0131  ;
  input \u0_R11_reg[1]/NET0131  ;
  input \u0_R11_reg[20]/NET0131  ;
  input \u0_R11_reg[21]/NET0131  ;
  input \u0_R11_reg[22]/NET0131  ;
  input \u0_R11_reg[23]/NET0131  ;
  input \u0_R11_reg[24]/NET0131  ;
  input \u0_R11_reg[25]/NET0131  ;
  input \u0_R11_reg[26]/NET0131  ;
  input \u0_R11_reg[27]/NET0131  ;
  input \u0_R11_reg[28]/NET0131  ;
  input \u0_R11_reg[29]/NET0131  ;
  input \u0_R11_reg[2]/NET0131  ;
  input \u0_R11_reg[30]/NET0131  ;
  input \u0_R11_reg[31]/P0001  ;
  input \u0_R11_reg[32]/NET0131  ;
  input \u0_R11_reg[3]/NET0131  ;
  input \u0_R11_reg[4]/NET0131  ;
  input \u0_R11_reg[5]/NET0131  ;
  input \u0_R11_reg[6]/NET0131  ;
  input \u0_R11_reg[7]/NET0131  ;
  input \u0_R11_reg[8]/NET0131  ;
  input \u0_R11_reg[9]/NET0131  ;
  input \u0_R12_reg[10]/NET0131  ;
  input \u0_R12_reg[11]/NET0131  ;
  input \u0_R12_reg[12]/NET0131  ;
  input \u0_R12_reg[13]/NET0131  ;
  input \u0_R12_reg[14]/NET0131  ;
  input \u0_R12_reg[15]/NET0131  ;
  input \u0_R12_reg[16]/NET0131  ;
  input \u0_R12_reg[17]/NET0131  ;
  input \u0_R12_reg[18]/NET0131  ;
  input \u0_R12_reg[19]/NET0131  ;
  input \u0_R12_reg[1]/NET0131  ;
  input \u0_R12_reg[20]/NET0131  ;
  input \u0_R12_reg[21]/NET0131  ;
  input \u0_R12_reg[22]/NET0131  ;
  input \u0_R12_reg[23]/NET0131  ;
  input \u0_R12_reg[24]/NET0131  ;
  input \u0_R12_reg[25]/NET0131  ;
  input \u0_R12_reg[26]/NET0131  ;
  input \u0_R12_reg[27]/NET0131  ;
  input \u0_R12_reg[28]/NET0131  ;
  input \u0_R12_reg[29]/NET0131  ;
  input \u0_R12_reg[2]/NET0131  ;
  input \u0_R12_reg[30]/NET0131  ;
  input \u0_R12_reg[31]/P0001  ;
  input \u0_R12_reg[32]/NET0131  ;
  input \u0_R12_reg[3]/NET0131  ;
  input \u0_R12_reg[4]/NET0131  ;
  input \u0_R12_reg[5]/NET0131  ;
  input \u0_R12_reg[6]/NET0131  ;
  input \u0_R12_reg[7]/NET0131  ;
  input \u0_R12_reg[8]/NET0131  ;
  input \u0_R12_reg[9]/NET0131  ;
  input \u0_R13_reg[10]/NET0131  ;
  input \u0_R13_reg[11]/NET0131  ;
  input \u0_R13_reg[12]/NET0131  ;
  input \u0_R13_reg[13]/NET0131  ;
  input \u0_R13_reg[14]/NET0131  ;
  input \u0_R13_reg[15]/NET0131  ;
  input \u0_R13_reg[16]/NET0131  ;
  input \u0_R13_reg[17]/NET0131  ;
  input \u0_R13_reg[18]/NET0131  ;
  input \u0_R13_reg[19]/NET0131  ;
  input \u0_R13_reg[1]/NET0131  ;
  input \u0_R13_reg[20]/NET0131  ;
  input \u0_R13_reg[21]/NET0131  ;
  input \u0_R13_reg[22]/P0001  ;
  input \u0_R13_reg[23]/NET0131  ;
  input \u0_R13_reg[24]/NET0131  ;
  input \u0_R13_reg[25]/NET0131  ;
  input \u0_R13_reg[26]/NET0131  ;
  input \u0_R13_reg[27]/P0001  ;
  input \u0_R13_reg[28]/NET0131  ;
  input \u0_R13_reg[29]/NET0131  ;
  input \u0_R13_reg[2]/NET0131  ;
  input \u0_R13_reg[30]/NET0131  ;
  input \u0_R13_reg[31]/NET0131  ;
  input \u0_R13_reg[32]/NET0131  ;
  input \u0_R13_reg[3]/NET0131  ;
  input \u0_R13_reg[4]/NET0131  ;
  input \u0_R13_reg[5]/NET0131  ;
  input \u0_R13_reg[6]/NET0131  ;
  input \u0_R13_reg[7]/NET0131  ;
  input \u0_R13_reg[8]/NET0131  ;
  input \u0_R13_reg[9]/NET0131  ;
  input \u0_R14_reg[10]/NET0131  ;
  input \u0_R14_reg[11]/P0001  ;
  input \u0_R14_reg[12]/NET0131  ;
  input \u0_R14_reg[13]/NET0131  ;
  input \u0_R14_reg[14]/NET0131  ;
  input \u0_R14_reg[15]/NET0131  ;
  input \u0_R14_reg[16]/NET0131  ;
  input \u0_R14_reg[17]/NET0131  ;
  input \u0_R14_reg[18]/NET0131  ;
  input \u0_R14_reg[19]/NET0131  ;
  input \u0_R14_reg[1]/NET0131  ;
  input \u0_R14_reg[20]/NET0131  ;
  input \u0_R14_reg[21]/NET0131  ;
  input \u0_R14_reg[22]/P0001  ;
  input \u0_R14_reg[23]/NET0131  ;
  input \u0_R14_reg[24]/NET0131  ;
  input \u0_R14_reg[25]/NET0131  ;
  input \u0_R14_reg[26]/P0001  ;
  input \u0_R14_reg[27]/P0001  ;
  input \u0_R14_reg[28]/NET0131  ;
  input \u0_R14_reg[29]/NET0131  ;
  input \u0_R14_reg[2]/NET0131  ;
  input \u0_R14_reg[30]/NET0131  ;
  input \u0_R14_reg[31]/P0001  ;
  input \u0_R14_reg[32]/NET0131  ;
  input \u0_R14_reg[3]/NET0131  ;
  input \u0_R14_reg[4]/NET0131  ;
  input \u0_R14_reg[5]/NET0131  ;
  input \u0_R14_reg[6]/NET0131  ;
  input \u0_R14_reg[7]/NET0131  ;
  input \u0_R14_reg[8]/NET0131  ;
  input \u0_R14_reg[9]/NET0131  ;
  input \u0_R1_reg[10]/NET0131  ;
  input \u0_R1_reg[11]/NET0131  ;
  input \u0_R1_reg[12]/NET0131  ;
  input \u0_R1_reg[13]/NET0131  ;
  input \u0_R1_reg[14]/NET0131  ;
  input \u0_R1_reg[15]/NET0131  ;
  input \u0_R1_reg[16]/NET0131  ;
  input \u0_R1_reg[17]/NET0131  ;
  input \u0_R1_reg[18]/NET0131  ;
  input \u0_R1_reg[19]/NET0131  ;
  input \u0_R1_reg[1]/NET0131  ;
  input \u0_R1_reg[20]/NET0131  ;
  input \u0_R1_reg[21]/NET0131  ;
  input \u0_R1_reg[22]/NET0131  ;
  input \u0_R1_reg[23]/NET0131  ;
  input \u0_R1_reg[24]/NET0131  ;
  input \u0_R1_reg[25]/NET0131  ;
  input \u0_R1_reg[26]/NET0131  ;
  input \u0_R1_reg[27]/NET0131  ;
  input \u0_R1_reg[28]/NET0131  ;
  input \u0_R1_reg[29]/NET0131  ;
  input \u0_R1_reg[2]/NET0131  ;
  input \u0_R1_reg[30]/NET0131  ;
  input \u0_R1_reg[31]/NET0131  ;
  input \u0_R1_reg[32]/NET0131  ;
  input \u0_R1_reg[3]/NET0131  ;
  input \u0_R1_reg[4]/NET0131  ;
  input \u0_R1_reg[5]/NET0131  ;
  input \u0_R1_reg[6]/NET0131  ;
  input \u0_R1_reg[7]/NET0131  ;
  input \u0_R1_reg[8]/NET0131  ;
  input \u0_R1_reg[9]/NET0131  ;
  input \u0_R2_reg[10]/NET0131  ;
  input \u0_R2_reg[11]/NET0131  ;
  input \u0_R2_reg[12]/NET0131  ;
  input \u0_R2_reg[13]/NET0131  ;
  input \u0_R2_reg[14]/NET0131  ;
  input \u0_R2_reg[15]/NET0131  ;
  input \u0_R2_reg[16]/NET0131  ;
  input \u0_R2_reg[17]/NET0131  ;
  input \u0_R2_reg[18]/NET0131  ;
  input \u0_R2_reg[19]/NET0131  ;
  input \u0_R2_reg[1]/NET0131  ;
  input \u0_R2_reg[20]/NET0131  ;
  input \u0_R2_reg[21]/NET0131  ;
  input \u0_R2_reg[22]/NET0131  ;
  input \u0_R2_reg[23]/NET0131  ;
  input \u0_R2_reg[24]/NET0131  ;
  input \u0_R2_reg[25]/NET0131  ;
  input \u0_R2_reg[26]/NET0131  ;
  input \u0_R2_reg[27]/NET0131  ;
  input \u0_R2_reg[28]/NET0131  ;
  input \u0_R2_reg[29]/NET0131  ;
  input \u0_R2_reg[2]/NET0131  ;
  input \u0_R2_reg[30]/NET0131  ;
  input \u0_R2_reg[31]/NET0131  ;
  input \u0_R2_reg[32]/NET0131  ;
  input \u0_R2_reg[3]/NET0131  ;
  input \u0_R2_reg[4]/NET0131  ;
  input \u0_R2_reg[5]/NET0131  ;
  input \u0_R2_reg[6]/NET0131  ;
  input \u0_R2_reg[7]/NET0131  ;
  input \u0_R2_reg[8]/NET0131  ;
  input \u0_R2_reg[9]/NET0131  ;
  input \u0_R3_reg[10]/NET0131  ;
  input \u0_R3_reg[11]/NET0131  ;
  input \u0_R3_reg[12]/NET0131  ;
  input \u0_R3_reg[13]/NET0131  ;
  input \u0_R3_reg[14]/NET0131  ;
  input \u0_R3_reg[15]/NET0131  ;
  input \u0_R3_reg[16]/NET0131  ;
  input \u0_R3_reg[17]/NET0131  ;
  input \u0_R3_reg[18]/NET0131  ;
  input \u0_R3_reg[19]/NET0131  ;
  input \u0_R3_reg[1]/NET0131  ;
  input \u0_R3_reg[20]/NET0131  ;
  input \u0_R3_reg[21]/NET0131  ;
  input \u0_R3_reg[22]/NET0131  ;
  input \u0_R3_reg[23]/NET0131  ;
  input \u0_R3_reg[24]/NET0131  ;
  input \u0_R3_reg[25]/NET0131  ;
  input \u0_R3_reg[26]/NET0131  ;
  input \u0_R3_reg[27]/NET0131  ;
  input \u0_R3_reg[28]/NET0131  ;
  input \u0_R3_reg[29]/NET0131  ;
  input \u0_R3_reg[2]/NET0131  ;
  input \u0_R3_reg[30]/NET0131  ;
  input \u0_R3_reg[31]/P0001  ;
  input \u0_R3_reg[32]/NET0131  ;
  input \u0_R3_reg[3]/NET0131  ;
  input \u0_R3_reg[4]/NET0131  ;
  input \u0_R3_reg[5]/NET0131  ;
  input \u0_R3_reg[6]/NET0131  ;
  input \u0_R3_reg[7]/NET0131  ;
  input \u0_R3_reg[8]/NET0131  ;
  input \u0_R3_reg[9]/NET0131  ;
  input \u0_R4_reg[10]/NET0131  ;
  input \u0_R4_reg[11]/NET0131  ;
  input \u0_R4_reg[12]/NET0131  ;
  input \u0_R4_reg[13]/NET0131  ;
  input \u0_R4_reg[14]/NET0131  ;
  input \u0_R4_reg[15]/NET0131  ;
  input \u0_R4_reg[16]/NET0131  ;
  input \u0_R4_reg[17]/NET0131  ;
  input \u0_R4_reg[18]/NET0131  ;
  input \u0_R4_reg[19]/NET0131  ;
  input \u0_R4_reg[1]/NET0131  ;
  input \u0_R4_reg[20]/NET0131  ;
  input \u0_R4_reg[21]/NET0131  ;
  input \u0_R4_reg[22]/NET0131  ;
  input \u0_R4_reg[23]/NET0131  ;
  input \u0_R4_reg[24]/NET0131  ;
  input \u0_R4_reg[25]/NET0131  ;
  input \u0_R4_reg[26]/NET0131  ;
  input \u0_R4_reg[27]/NET0131  ;
  input \u0_R4_reg[28]/NET0131  ;
  input \u0_R4_reg[29]/NET0131  ;
  input \u0_R4_reg[2]/NET0131  ;
  input \u0_R4_reg[30]/NET0131  ;
  input \u0_R4_reg[31]/P0001  ;
  input \u0_R4_reg[32]/NET0131  ;
  input \u0_R4_reg[3]/NET0131  ;
  input \u0_R4_reg[4]/NET0131  ;
  input \u0_R4_reg[5]/NET0131  ;
  input \u0_R4_reg[6]/NET0131  ;
  input \u0_R4_reg[7]/NET0131  ;
  input \u0_R4_reg[8]/NET0131  ;
  input \u0_R4_reg[9]/NET0131  ;
  input \u0_R5_reg[10]/NET0131  ;
  input \u0_R5_reg[11]/P0001  ;
  input \u0_R5_reg[12]/NET0131  ;
  input \u0_R5_reg[13]/NET0131  ;
  input \u0_R5_reg[14]/NET0131  ;
  input \u0_R5_reg[15]/NET0131  ;
  input \u0_R5_reg[16]/NET0131  ;
  input \u0_R5_reg[17]/NET0131  ;
  input \u0_R5_reg[18]/NET0131  ;
  input \u0_R5_reg[19]/NET0131  ;
  input \u0_R5_reg[1]/NET0131  ;
  input \u0_R5_reg[20]/NET0131  ;
  input \u0_R5_reg[21]/NET0131  ;
  input \u0_R5_reg[22]/NET0131  ;
  input \u0_R5_reg[23]/NET0131  ;
  input \u0_R5_reg[24]/NET0131  ;
  input \u0_R5_reg[25]/NET0131  ;
  input \u0_R5_reg[26]/NET0131  ;
  input \u0_R5_reg[27]/NET0131  ;
  input \u0_R5_reg[28]/NET0131  ;
  input \u0_R5_reg[29]/NET0131  ;
  input \u0_R5_reg[2]/NET0131  ;
  input \u0_R5_reg[30]/NET0131  ;
  input \u0_R5_reg[31]/P0001  ;
  input \u0_R5_reg[32]/NET0131  ;
  input \u0_R5_reg[3]/NET0131  ;
  input \u0_R5_reg[4]/NET0131  ;
  input \u0_R5_reg[5]/NET0131  ;
  input \u0_R5_reg[6]/NET0131  ;
  input \u0_R5_reg[7]/NET0131  ;
  input \u0_R5_reg[8]/NET0131  ;
  input \u0_R5_reg[9]/NET0131  ;
  input \u0_R6_reg[10]/NET0131  ;
  input \u0_R6_reg[11]/NET0131  ;
  input \u0_R6_reg[12]/NET0131  ;
  input \u0_R6_reg[13]/NET0131  ;
  input \u0_R6_reg[14]/NET0131  ;
  input \u0_R6_reg[15]/NET0131  ;
  input \u0_R6_reg[16]/NET0131  ;
  input \u0_R6_reg[17]/NET0131  ;
  input \u0_R6_reg[18]/NET0131  ;
  input \u0_R6_reg[19]/NET0131  ;
  input \u0_R6_reg[1]/NET0131  ;
  input \u0_R6_reg[20]/NET0131  ;
  input \u0_R6_reg[21]/NET0131  ;
  input \u0_R6_reg[22]/NET0131  ;
  input \u0_R6_reg[23]/NET0131  ;
  input \u0_R6_reg[24]/NET0131  ;
  input \u0_R6_reg[25]/NET0131  ;
  input \u0_R6_reg[26]/NET0131  ;
  input \u0_R6_reg[27]/NET0131  ;
  input \u0_R6_reg[28]/NET0131  ;
  input \u0_R6_reg[29]/NET0131  ;
  input \u0_R6_reg[2]/NET0131  ;
  input \u0_R6_reg[30]/NET0131  ;
  input \u0_R6_reg[31]/P0001  ;
  input \u0_R6_reg[32]/NET0131  ;
  input \u0_R6_reg[3]/NET0131  ;
  input \u0_R6_reg[4]/NET0131  ;
  input \u0_R6_reg[5]/NET0131  ;
  input \u0_R6_reg[6]/NET0131  ;
  input \u0_R6_reg[7]/NET0131  ;
  input \u0_R6_reg[8]/NET0131  ;
  input \u0_R6_reg[9]/NET0131  ;
  input \u0_R7_reg[10]/NET0131  ;
  input \u0_R7_reg[11]/P0001  ;
  input \u0_R7_reg[12]/NET0131  ;
  input \u0_R7_reg[13]/NET0131  ;
  input \u0_R7_reg[14]/NET0131  ;
  input \u0_R7_reg[15]/NET0131  ;
  input \u0_R7_reg[16]/NET0131  ;
  input \u0_R7_reg[17]/NET0131  ;
  input \u0_R7_reg[18]/NET0131  ;
  input \u0_R7_reg[19]/NET0131  ;
  input \u0_R7_reg[1]/NET0131  ;
  input \u0_R7_reg[20]/NET0131  ;
  input \u0_R7_reg[21]/NET0131  ;
  input \u0_R7_reg[22]/NET0131  ;
  input \u0_R7_reg[23]/NET0131  ;
  input \u0_R7_reg[24]/NET0131  ;
  input \u0_R7_reg[25]/NET0131  ;
  input \u0_R7_reg[26]/NET0131  ;
  input \u0_R7_reg[27]/NET0131  ;
  input \u0_R7_reg[28]/NET0131  ;
  input \u0_R7_reg[29]/NET0131  ;
  input \u0_R7_reg[2]/NET0131  ;
  input \u0_R7_reg[30]/NET0131  ;
  input \u0_R7_reg[31]/P0001  ;
  input \u0_R7_reg[32]/NET0131  ;
  input \u0_R7_reg[3]/NET0131  ;
  input \u0_R7_reg[4]/NET0131  ;
  input \u0_R7_reg[5]/NET0131  ;
  input \u0_R7_reg[6]/NET0131  ;
  input \u0_R7_reg[7]/NET0131  ;
  input \u0_R7_reg[8]/NET0131  ;
  input \u0_R7_reg[9]/NET0131  ;
  input \u0_R8_reg[10]/NET0131  ;
  input \u0_R8_reg[11]/NET0131  ;
  input \u0_R8_reg[12]/NET0131  ;
  input \u0_R8_reg[13]/NET0131  ;
  input \u0_R8_reg[14]/NET0131  ;
  input \u0_R8_reg[15]/NET0131  ;
  input \u0_R8_reg[16]/NET0131  ;
  input \u0_R8_reg[17]/NET0131  ;
  input \u0_R8_reg[18]/NET0131  ;
  input \u0_R8_reg[19]/NET0131  ;
  input \u0_R8_reg[1]/NET0131  ;
  input \u0_R8_reg[20]/NET0131  ;
  input \u0_R8_reg[21]/NET0131  ;
  input \u0_R8_reg[22]/NET0131  ;
  input \u0_R8_reg[23]/NET0131  ;
  input \u0_R8_reg[24]/NET0131  ;
  input \u0_R8_reg[25]/NET0131  ;
  input \u0_R8_reg[26]/NET0131  ;
  input \u0_R8_reg[27]/NET0131  ;
  input \u0_R8_reg[28]/NET0131  ;
  input \u0_R8_reg[29]/NET0131  ;
  input \u0_R8_reg[2]/NET0131  ;
  input \u0_R8_reg[30]/NET0131  ;
  input \u0_R8_reg[31]/P0001  ;
  input \u0_R8_reg[32]/NET0131  ;
  input \u0_R8_reg[3]/NET0131  ;
  input \u0_R8_reg[4]/NET0131  ;
  input \u0_R8_reg[5]/NET0131  ;
  input \u0_R8_reg[6]/NET0131  ;
  input \u0_R8_reg[7]/NET0131  ;
  input \u0_R8_reg[8]/NET0131  ;
  input \u0_R8_reg[9]/NET0131  ;
  input \u0_R9_reg[10]/NET0131  ;
  input \u0_R9_reg[11]/P0001  ;
  input \u0_R9_reg[12]/NET0131  ;
  input \u0_R9_reg[13]/NET0131  ;
  input \u0_R9_reg[14]/NET0131  ;
  input \u0_R9_reg[15]/NET0131  ;
  input \u0_R9_reg[16]/NET0131  ;
  input \u0_R9_reg[17]/NET0131  ;
  input \u0_R9_reg[18]/NET0131  ;
  input \u0_R9_reg[19]/NET0131  ;
  input \u0_R9_reg[1]/NET0131  ;
  input \u0_R9_reg[20]/NET0131  ;
  input \u0_R9_reg[21]/NET0131  ;
  input \u0_R9_reg[22]/NET0131  ;
  input \u0_R9_reg[23]/NET0131  ;
  input \u0_R9_reg[24]/NET0131  ;
  input \u0_R9_reg[25]/NET0131  ;
  input \u0_R9_reg[26]/NET0131  ;
  input \u0_R9_reg[27]/NET0131  ;
  input \u0_R9_reg[28]/NET0131  ;
  input \u0_R9_reg[29]/NET0131  ;
  input \u0_R9_reg[2]/NET0131  ;
  input \u0_R9_reg[30]/NET0131  ;
  input \u0_R9_reg[31]/P0001  ;
  input \u0_R9_reg[32]/NET0131  ;
  input \u0_R9_reg[3]/NET0131  ;
  input \u0_R9_reg[4]/NET0131  ;
  input \u0_R9_reg[5]/NET0131  ;
  input \u0_R9_reg[6]/NET0131  ;
  input \u0_R9_reg[7]/NET0131  ;
  input \u0_R9_reg[8]/NET0131  ;
  input \u0_R9_reg[9]/NET0131  ;
  input \u0_desIn_r_reg[0]/NET0131  ;
  input \u0_desIn_r_reg[10]/NET0131  ;
  input \u0_desIn_r_reg[11]/NET0131  ;
  input \u0_desIn_r_reg[12]/NET0131  ;
  input \u0_desIn_r_reg[13]/NET0131  ;
  input \u0_desIn_r_reg[14]/NET0131  ;
  input \u0_desIn_r_reg[15]/NET0131  ;
  input \u0_desIn_r_reg[16]/NET0131  ;
  input \u0_desIn_r_reg[17]/NET0131  ;
  input \u0_desIn_r_reg[18]/NET0131  ;
  input \u0_desIn_r_reg[19]/NET0131  ;
  input \u0_desIn_r_reg[1]/NET0131  ;
  input \u0_desIn_r_reg[20]/NET0131  ;
  input \u0_desIn_r_reg[21]/NET0131  ;
  input \u0_desIn_r_reg[22]/NET0131  ;
  input \u0_desIn_r_reg[23]/NET0131  ;
  input \u0_desIn_r_reg[24]/NET0131  ;
  input \u0_desIn_r_reg[25]/NET0131  ;
  input \u0_desIn_r_reg[26]/NET0131  ;
  input \u0_desIn_r_reg[27]/NET0131  ;
  input \u0_desIn_r_reg[28]/NET0131  ;
  input \u0_desIn_r_reg[29]/NET0131  ;
  input \u0_desIn_r_reg[2]/NET0131  ;
  input \u0_desIn_r_reg[30]/NET0131  ;
  input \u0_desIn_r_reg[31]/NET0131  ;
  input \u0_desIn_r_reg[32]/NET0131  ;
  input \u0_desIn_r_reg[33]/NET0131  ;
  input \u0_desIn_r_reg[34]/NET0131  ;
  input \u0_desIn_r_reg[35]/NET0131  ;
  input \u0_desIn_r_reg[36]/NET0131  ;
  input \u0_desIn_r_reg[37]/NET0131  ;
  input \u0_desIn_r_reg[38]/NET0131  ;
  input \u0_desIn_r_reg[39]/NET0131  ;
  input \u0_desIn_r_reg[3]/NET0131  ;
  input \u0_desIn_r_reg[40]/NET0131  ;
  input \u0_desIn_r_reg[41]/NET0131  ;
  input \u0_desIn_r_reg[42]/NET0131  ;
  input \u0_desIn_r_reg[43]/NET0131  ;
  input \u0_desIn_r_reg[44]/NET0131  ;
  input \u0_desIn_r_reg[45]/NET0131  ;
  input \u0_desIn_r_reg[46]/NET0131  ;
  input \u0_desIn_r_reg[47]/NET0131  ;
  input \u0_desIn_r_reg[48]/NET0131  ;
  input \u0_desIn_r_reg[49]/NET0131  ;
  input \u0_desIn_r_reg[4]/NET0131  ;
  input \u0_desIn_r_reg[50]/NET0131  ;
  input \u0_desIn_r_reg[51]/NET0131  ;
  input \u0_desIn_r_reg[52]/NET0131  ;
  input \u0_desIn_r_reg[53]/NET0131  ;
  input \u0_desIn_r_reg[54]/NET0131  ;
  input \u0_desIn_r_reg[55]/NET0131  ;
  input \u0_desIn_r_reg[56]/NET0131  ;
  input \u0_desIn_r_reg[57]/NET0131  ;
  input \u0_desIn_r_reg[58]/NET0131  ;
  input \u0_desIn_r_reg[59]/NET0131  ;
  input \u0_desIn_r_reg[5]/NET0131  ;
  input \u0_desIn_r_reg[60]/NET0131  ;
  input \u0_desIn_r_reg[61]/NET0131  ;
  input \u0_desIn_r_reg[62]/NET0131  ;
  input \u0_desIn_r_reg[63]/NET0131  ;
  input \u0_desIn_r_reg[6]/NET0131  ;
  input \u0_desIn_r_reg[7]/NET0131  ;
  input \u0_desIn_r_reg[8]/NET0131  ;
  input \u0_desIn_r_reg[9]/NET0131  ;
  input \u0_key_r_reg[0]/NET0131  ;
  input \u0_key_r_reg[10]/P0001  ;
  input \u0_key_r_reg[11]/NET0131  ;
  input \u0_key_r_reg[12]/NET0131  ;
  input \u0_key_r_reg[13]/NET0131  ;
  input \u0_key_r_reg[14]/NET0131  ;
  input \u0_key_r_reg[15]/NET0131  ;
  input \u0_key_r_reg[16]/NET0131  ;
  input \u0_key_r_reg[17]/NET0131  ;
  input \u0_key_r_reg[18]/NET0131  ;
  input \u0_key_r_reg[19]/NET0131  ;
  input \u0_key_r_reg[1]/NET0131  ;
  input \u0_key_r_reg[20]/NET0131  ;
  input \u0_key_r_reg[21]/NET0131  ;
  input \u0_key_r_reg[22]/NET0131  ;
  input \u0_key_r_reg[23]/NET0131  ;
  input \u0_key_r_reg[24]/NET0131  ;
  input \u0_key_r_reg[25]/NET0131  ;
  input \u0_key_r_reg[26]/NET0131  ;
  input \u0_key_r_reg[27]/NET0131  ;
  input \u0_key_r_reg[28]/NET0131  ;
  input \u0_key_r_reg[29]/NET0131  ;
  input \u0_key_r_reg[2]/NET0131  ;
  input \u0_key_r_reg[30]/NET0131  ;
  input \u0_key_r_reg[31]/NET0131  ;
  input \u0_key_r_reg[32]/NET0131  ;
  input \u0_key_r_reg[33]/NET0131  ;
  input \u0_key_r_reg[34]/NET0131  ;
  input \u0_key_r_reg[35]/P0001  ;
  input \u0_key_r_reg[36]/NET0131  ;
  input \u0_key_r_reg[37]/NET0131  ;
  input \u0_key_r_reg[38]/NET0131  ;
  input \u0_key_r_reg[39]/P0001  ;
  input \u0_key_r_reg[3]/NET0131  ;
  input \u0_key_r_reg[40]/NET0131  ;
  input \u0_key_r_reg[41]/NET0131  ;
  input \u0_key_r_reg[42]/P0001  ;
  input \u0_key_r_reg[43]/NET0131  ;
  input \u0_key_r_reg[44]/NET0131  ;
  input \u0_key_r_reg[45]/NET0131  ;
  input \u0_key_r_reg[46]/NET0131  ;
  input \u0_key_r_reg[47]/NET0131  ;
  input \u0_key_r_reg[48]/NET0131  ;
  input \u0_key_r_reg[49]/NET0131  ;
  input \u0_key_r_reg[4]/NET0131  ;
  input \u0_key_r_reg[50]/NET0131  ;
  input \u0_key_r_reg[51]/NET0131  ;
  input \u0_key_r_reg[52]/NET0131  ;
  input \u0_key_r_reg[53]/NET0131  ;
  input \u0_key_r_reg[54]/NET0131  ;
  input \u0_key_r_reg[55]/NET0131  ;
  input \u0_key_r_reg[5]/NET0131  ;
  input \u0_key_r_reg[6]/NET0131  ;
  input \u0_key_r_reg[7]/NET0131  ;
  input \u0_key_r_reg[8]/NET0131  ;
  input \u0_key_r_reg[9]/NET0131  ;
  input \u0_uk_K_r0_reg[0]/NET0131  ;
  input \u0_uk_K_r0_reg[10]/NET0131  ;
  input \u0_uk_K_r0_reg[11]/NET0131  ;
  input \u0_uk_K_r0_reg[12]/NET0131  ;
  input \u0_uk_K_r0_reg[13]/NET0131  ;
  input \u0_uk_K_r0_reg[14]/NET0131  ;
  input \u0_uk_K_r0_reg[15]/NET0131  ;
  input \u0_uk_K_r0_reg[16]/NET0131  ;
  input \u0_uk_K_r0_reg[17]/NET0131  ;
  input \u0_uk_K_r0_reg[18]/NET0131  ;
  input \u0_uk_K_r0_reg[19]/NET0131  ;
  input \u0_uk_K_r0_reg[20]/NET0131  ;
  input \u0_uk_K_r0_reg[21]/NET0131  ;
  input \u0_uk_K_r0_reg[22]/NET0131  ;
  input \u0_uk_K_r0_reg[23]/NET0131  ;
  input \u0_uk_K_r0_reg[24]/P0001  ;
  input \u0_uk_K_r0_reg[25]/P0001  ;
  input \u0_uk_K_r0_reg[26]/NET0131  ;
  input \u0_uk_K_r0_reg[27]/NET0131  ;
  input \u0_uk_K_r0_reg[28]/NET0131  ;
  input \u0_uk_K_r0_reg[29]/NET0131  ;
  input \u0_uk_K_r0_reg[2]/NET0131  ;
  input \u0_uk_K_r0_reg[30]/NET0131  ;
  input \u0_uk_K_r0_reg[31]/NET0131  ;
  input \u0_uk_K_r0_reg[32]/NET0131  ;
  input \u0_uk_K_r0_reg[33]/NET0131  ;
  input \u0_uk_K_r0_reg[34]/NET0131  ;
  input \u0_uk_K_r0_reg[35]/NET0131  ;
  input \u0_uk_K_r0_reg[36]/NET0131  ;
  input \u0_uk_K_r0_reg[37]/NET0131  ;
  input \u0_uk_K_r0_reg[38]/NET0131  ;
  input \u0_uk_K_r0_reg[39]/NET0131  ;
  input \u0_uk_K_r0_reg[3]/NET0131  ;
  input \u0_uk_K_r0_reg[40]/NET0131  ;
  input \u0_uk_K_r0_reg[41]/NET0131  ;
  input \u0_uk_K_r0_reg[42]/NET0131  ;
  input \u0_uk_K_r0_reg[43]/NET0131  ;
  input \u0_uk_K_r0_reg[44]/NET0131  ;
  input \u0_uk_K_r0_reg[45]/NET0131  ;
  input \u0_uk_K_r0_reg[46]/NET0131  ;
  input \u0_uk_K_r0_reg[47]/NET0131  ;
  input \u0_uk_K_r0_reg[48]/NET0131  ;
  input \u0_uk_K_r0_reg[49]/NET0131  ;
  input \u0_uk_K_r0_reg[4]/NET0131  ;
  input \u0_uk_K_r0_reg[50]/NET0131  ;
  input \u0_uk_K_r0_reg[51]/NET0131  ;
  input \u0_uk_K_r0_reg[52]/NET0131  ;
  input \u0_uk_K_r0_reg[54]/NET0131  ;
  input \u0_uk_K_r0_reg[55]/NET0131  ;
  input \u0_uk_K_r0_reg[5]/NET0131  ;
  input \u0_uk_K_r0_reg[6]/NET0131  ;
  input \u0_uk_K_r0_reg[7]/NET0131  ;
  input \u0_uk_K_r0_reg[8]/NET0131  ;
  input \u0_uk_K_r0_reg[9]/NET0131  ;
  input \u0_uk_K_r10_reg[0]/NET0131  ;
  input \u0_uk_K_r10_reg[10]/NET0131  ;
  input \u0_uk_K_r10_reg[11]/NET0131  ;
  input \u0_uk_K_r10_reg[12]/NET0131  ;
  input \u0_uk_K_r10_reg[14]/NET0131  ;
  input \u0_uk_K_r10_reg[15]/NET0131  ;
  input \u0_uk_K_r10_reg[16]/NET0131  ;
  input \u0_uk_K_r10_reg[17]/NET0131  ;
  input \u0_uk_K_r10_reg[18]/NET0131  ;
  input \u0_uk_K_r10_reg[19]/NET0131  ;
  input \u0_uk_K_r10_reg[1]/NET0131  ;
  input \u0_uk_K_r10_reg[20]/NET0131  ;
  input \u0_uk_K_r10_reg[21]/NET0131  ;
  input \u0_uk_K_r10_reg[22]/NET0131  ;
  input \u0_uk_K_r10_reg[23]/NET0131  ;
  input \u0_uk_K_r10_reg[24]/NET0131  ;
  input \u0_uk_K_r10_reg[25]/NET0131  ;
  input \u0_uk_K_r10_reg[26]/NET0131  ;
  input \u0_uk_K_r10_reg[27]/NET0131  ;
  input \u0_uk_K_r10_reg[28]/NET0131  ;
  input \u0_uk_K_r10_reg[29]/NET0131  ;
  input \u0_uk_K_r10_reg[2]/NET0131  ;
  input \u0_uk_K_r10_reg[30]/NET0131  ;
  input \u0_uk_K_r10_reg[31]/NET0131  ;
  input \u0_uk_K_r10_reg[32]/NET0131  ;
  input \u0_uk_K_r10_reg[33]/NET0131  ;
  input \u0_uk_K_r10_reg[34]/NET0131  ;
  input \u0_uk_K_r10_reg[35]/NET0131  ;
  input \u0_uk_K_r10_reg[36]/NET0131  ;
  input \u0_uk_K_r10_reg[37]/NET0131  ;
  input \u0_uk_K_r10_reg[38]/NET0131  ;
  input \u0_uk_K_r10_reg[39]/NET0131  ;
  input \u0_uk_K_r10_reg[3]/NET0131  ;
  input \u0_uk_K_r10_reg[40]/NET0131  ;
  input \u0_uk_K_r10_reg[41]/P0001  ;
  input \u0_uk_K_r10_reg[42]/NET0131  ;
  input \u0_uk_K_r10_reg[43]/NET0131  ;
  input \u0_uk_K_r10_reg[44]/NET0131  ;
  input \u0_uk_K_r10_reg[45]/P0001  ;
  input \u0_uk_K_r10_reg[46]/NET0131  ;
  input \u0_uk_K_r10_reg[47]/NET0131  ;
  input \u0_uk_K_r10_reg[48]/NET0131  ;
  input \u0_uk_K_r10_reg[49]/NET0131  ;
  input \u0_uk_K_r10_reg[4]/NET0131  ;
  input \u0_uk_K_r10_reg[50]/NET0131  ;
  input \u0_uk_K_r10_reg[51]/NET0131  ;
  input \u0_uk_K_r10_reg[52]/NET0131  ;
  input \u0_uk_K_r10_reg[53]/NET0131  ;
  input \u0_uk_K_r10_reg[54]/NET0131  ;
  input \u0_uk_K_r10_reg[55]/NET0131  ;
  input \u0_uk_K_r10_reg[5]/NET0131  ;
  input \u0_uk_K_r10_reg[6]/NET0131  ;
  input \u0_uk_K_r10_reg[7]/NET0131  ;
  input \u0_uk_K_r10_reg[8]/NET0131  ;
  input \u0_uk_K_r10_reg[9]/NET0131  ;
  input \u0_uk_K_r11_reg[0]/NET0131  ;
  input \u0_uk_K_r11_reg[10]/NET0131  ;
  input \u0_uk_K_r11_reg[11]/NET0131  ;
  input \u0_uk_K_r11_reg[12]/NET0131  ;
  input \u0_uk_K_r11_reg[13]/NET0131  ;
  input \u0_uk_K_r11_reg[14]/NET0131  ;
  input \u0_uk_K_r11_reg[15]/NET0131  ;
  input \u0_uk_K_r11_reg[16]/NET0131  ;
  input \u0_uk_K_r11_reg[17]/NET0131  ;
  input \u0_uk_K_r11_reg[18]/NET0131  ;
  input \u0_uk_K_r11_reg[19]/NET0131  ;
  input \u0_uk_K_r11_reg[1]/NET0131  ;
  input \u0_uk_K_r11_reg[20]/NET0131  ;
  input \u0_uk_K_r11_reg[21]/NET0131  ;
  input \u0_uk_K_r11_reg[22]/NET0131  ;
  input \u0_uk_K_r11_reg[23]/NET0131  ;
  input \u0_uk_K_r11_reg[24]/NET0131  ;
  input \u0_uk_K_r11_reg[25]/NET0131  ;
  input \u0_uk_K_r11_reg[26]/NET0131  ;
  input \u0_uk_K_r11_reg[27]/P0001  ;
  input \u0_uk_K_r11_reg[28]/NET0131  ;
  input \u0_uk_K_r11_reg[29]/NET0131  ;
  input \u0_uk_K_r11_reg[2]/NET0131  ;
  input \u0_uk_K_r11_reg[31]/NET0131  ;
  input \u0_uk_K_r11_reg[32]/NET0131  ;
  input \u0_uk_K_r11_reg[33]/NET0131  ;
  input \u0_uk_K_r11_reg[34]/NET0131  ;
  input \u0_uk_K_r11_reg[35]/NET0131  ;
  input \u0_uk_K_r11_reg[36]/NET0131  ;
  input \u0_uk_K_r11_reg[37]/NET0131  ;
  input \u0_uk_K_r11_reg[38]/NET0131  ;
  input \u0_uk_K_r11_reg[39]/NET0131  ;
  input \u0_uk_K_r11_reg[3]/NET0131  ;
  input \u0_uk_K_r11_reg[40]/NET0131  ;
  input \u0_uk_K_r11_reg[41]/NET0131  ;
  input \u0_uk_K_r11_reg[42]/NET0131  ;
  input \u0_uk_K_r11_reg[43]/NET0131  ;
  input \u0_uk_K_r11_reg[44]/NET0131  ;
  input \u0_uk_K_r11_reg[45]/NET0131  ;
  input \u0_uk_K_r11_reg[46]/NET0131  ;
  input \u0_uk_K_r11_reg[47]/NET0131  ;
  input \u0_uk_K_r11_reg[48]/NET0131  ;
  input \u0_uk_K_r11_reg[49]/NET0131  ;
  input \u0_uk_K_r11_reg[4]/NET0131  ;
  input \u0_uk_K_r11_reg[50]/NET0131  ;
  input \u0_uk_K_r11_reg[51]/NET0131  ;
  input \u0_uk_K_r11_reg[52]/NET0131  ;
  input \u0_uk_K_r11_reg[53]/P0001  ;
  input \u0_uk_K_r11_reg[54]/NET0131  ;
  input \u0_uk_K_r11_reg[55]/NET0131  ;
  input \u0_uk_K_r11_reg[5]/NET0131  ;
  input \u0_uk_K_r11_reg[6]/NET0131  ;
  input \u0_uk_K_r11_reg[7]/NET0131  ;
  input \u0_uk_K_r11_reg[8]/NET0131  ;
  input \u0_uk_K_r11_reg[9]/NET0131  ;
  input \u0_uk_K_r12_reg[0]/NET0131  ;
  input \u0_uk_K_r12_reg[10]/P0001  ;
  input \u0_uk_K_r12_reg[11]/NET0131  ;
  input \u0_uk_K_r12_reg[12]/NET0131  ;
  input \u0_uk_K_r12_reg[13]/NET0131  ;
  input \u0_uk_K_r12_reg[14]/NET0131  ;
  input \u0_uk_K_r12_reg[15]/NET0131  ;
  input \u0_uk_K_r12_reg[16]/NET0131  ;
  input \u0_uk_K_r12_reg[17]/NET0131  ;
  input \u0_uk_K_r12_reg[18]/NET0131  ;
  input \u0_uk_K_r12_reg[19]/NET0131  ;
  input \u0_uk_K_r12_reg[1]/NET0131  ;
  input \u0_uk_K_r12_reg[20]/NET0131  ;
  input \u0_uk_K_r12_reg[21]/NET0131  ;
  input \u0_uk_K_r12_reg[22]/NET0131  ;
  input \u0_uk_K_r12_reg[23]/NET0131  ;
  input \u0_uk_K_r12_reg[24]/NET0131  ;
  input \u0_uk_K_r12_reg[25]/NET0131  ;
  input \u0_uk_K_r12_reg[26]/NET0131  ;
  input \u0_uk_K_r12_reg[27]/NET0131  ;
  input \u0_uk_K_r12_reg[28]/NET0131  ;
  input \u0_uk_K_r12_reg[29]/NET0131  ;
  input \u0_uk_K_r12_reg[2]/NET0131  ;
  input \u0_uk_K_r12_reg[30]/NET0131  ;
  input \u0_uk_K_r12_reg[31]/NET0131  ;
  input \u0_uk_K_r12_reg[32]/NET0131  ;
  input \u0_uk_K_r12_reg[33]/NET0131  ;
  input \u0_uk_K_r12_reg[34]/NET0131  ;
  input \u0_uk_K_r12_reg[35]/NET0131  ;
  input \u0_uk_K_r12_reg[36]/NET0131  ;
  input \u0_uk_K_r12_reg[37]/NET0131  ;
  input \u0_uk_K_r12_reg[38]/NET0131  ;
  input \u0_uk_K_r12_reg[3]/NET0131  ;
  input \u0_uk_K_r12_reg[40]/NET0131  ;
  input \u0_uk_K_r12_reg[41]/NET0131  ;
  input \u0_uk_K_r12_reg[42]/NET0131  ;
  input \u0_uk_K_r12_reg[43]/NET0131  ;
  input \u0_uk_K_r12_reg[44]/P0001  ;
  input \u0_uk_K_r12_reg[45]/NET0131  ;
  input \u0_uk_K_r12_reg[46]/NET0131  ;
  input \u0_uk_K_r12_reg[47]/NET0131  ;
  input \u0_uk_K_r12_reg[48]/NET0131  ;
  input \u0_uk_K_r12_reg[49]/NET0131  ;
  input \u0_uk_K_r12_reg[4]/NET0131  ;
  input \u0_uk_K_r12_reg[50]/NET0131  ;
  input \u0_uk_K_r12_reg[51]/NET0131  ;
  input \u0_uk_K_r12_reg[52]/NET0131  ;
  input \u0_uk_K_r12_reg[53]/NET0131  ;
  input \u0_uk_K_r12_reg[54]/NET0131  ;
  input \u0_uk_K_r12_reg[55]/NET0131  ;
  input \u0_uk_K_r12_reg[5]/NET0131  ;
  input \u0_uk_K_r12_reg[6]/NET0131  ;
  input \u0_uk_K_r12_reg[7]/P0001  ;
  input \u0_uk_K_r12_reg[8]/NET0131  ;
  input \u0_uk_K_r12_reg[9]/NET0131  ;
  input \u0_uk_K_r13_reg[0]/NET0131  ;
  input \u0_uk_K_r13_reg[10]/NET0131  ;
  input \u0_uk_K_r13_reg[11]/NET0131  ;
  input \u0_uk_K_r13_reg[12]/NET0131  ;
  input \u0_uk_K_r13_reg[13]/NET0131  ;
  input \u0_uk_K_r13_reg[14]/NET0131  ;
  input \u0_uk_K_r13_reg[15]/NET0131  ;
  input \u0_uk_K_r13_reg[16]/NET0131  ;
  input \u0_uk_K_r13_reg[17]/NET0131  ;
  input \u0_uk_K_r13_reg[18]/NET0131  ;
  input \u0_uk_K_r13_reg[19]/NET0131  ;
  input \u0_uk_K_r13_reg[20]/NET0131  ;
  input \u0_uk_K_r13_reg[21]/NET0131  ;
  input \u0_uk_K_r13_reg[22]/NET0131  ;
  input \u0_uk_K_r13_reg[23]/NET0131  ;
  input \u0_uk_K_r13_reg[24]/NET0131  ;
  input \u0_uk_K_r13_reg[25]/P0001  ;
  input \u0_uk_K_r13_reg[26]/NET0131  ;
  input \u0_uk_K_r13_reg[27]/NET0131  ;
  input \u0_uk_K_r13_reg[28]/NET0131  ;
  input \u0_uk_K_r13_reg[29]/NET0131  ;
  input \u0_uk_K_r13_reg[2]/NET0131  ;
  input \u0_uk_K_r13_reg[30]/NET0131  ;
  input \u0_uk_K_r13_reg[31]/NET0131  ;
  input \u0_uk_K_r13_reg[32]/NET0131  ;
  input \u0_uk_K_r13_reg[33]/NET0131  ;
  input \u0_uk_K_r13_reg[34]/NET0131  ;
  input \u0_uk_K_r13_reg[35]/NET0131  ;
  input \u0_uk_K_r13_reg[36]/NET0131  ;
  input \u0_uk_K_r13_reg[37]/NET0131  ;
  input \u0_uk_K_r13_reg[38]/NET0131  ;
  input \u0_uk_K_r13_reg[39]/NET0131  ;
  input \u0_uk_K_r13_reg[3]/NET0131  ;
  input \u0_uk_K_r13_reg[40]/NET0131  ;
  input \u0_uk_K_r13_reg[41]/NET0131  ;
  input \u0_uk_K_r13_reg[42]/NET0131  ;
  input \u0_uk_K_r13_reg[43]/NET0131  ;
  input \u0_uk_K_r13_reg[44]/NET0131  ;
  input \u0_uk_K_r13_reg[45]/NET0131  ;
  input \u0_uk_K_r13_reg[46]/NET0131  ;
  input \u0_uk_K_r13_reg[47]/NET0131  ;
  input \u0_uk_K_r13_reg[48]/NET0131  ;
  input \u0_uk_K_r13_reg[49]/NET0131  ;
  input \u0_uk_K_r13_reg[4]/NET0131  ;
  input \u0_uk_K_r13_reg[50]/NET0131  ;
  input \u0_uk_K_r13_reg[51]/NET0131  ;
  input \u0_uk_K_r13_reg[52]/P0001  ;
  input \u0_uk_K_r13_reg[54]/NET0131  ;
  input \u0_uk_K_r13_reg[55]/NET0131  ;
  input \u0_uk_K_r13_reg[5]/NET0131  ;
  input \u0_uk_K_r13_reg[6]/NET0131  ;
  input \u0_uk_K_r13_reg[7]/NET0131  ;
  input \u0_uk_K_r13_reg[8]/NET0131  ;
  input \u0_uk_K_r13_reg[9]/NET0131  ;
  input \u0_uk_K_r14_reg[0]/NET0131  ;
  input \u0_uk_K_r14_reg[10]/P0001  ;
  input \u0_uk_K_r14_reg[11]/NET0131  ;
  input \u0_uk_K_r14_reg[12]/NET0131  ;
  input \u0_uk_K_r14_reg[13]/NET0131  ;
  input \u0_uk_K_r14_reg[14]/NET0131  ;
  input \u0_uk_K_r14_reg[15]/NET0131  ;
  input \u0_uk_K_r14_reg[16]/NET0131  ;
  input \u0_uk_K_r14_reg[17]/NET0131  ;
  input \u0_uk_K_r14_reg[18]/NET0131  ;
  input \u0_uk_K_r14_reg[19]/NET0131  ;
  input \u0_uk_K_r14_reg[1]/NET0131  ;
  input \u0_uk_K_r14_reg[20]/NET0131  ;
  input \u0_uk_K_r14_reg[21]/NET0131  ;
  input \u0_uk_K_r14_reg[22]/NET0131  ;
  input \u0_uk_K_r14_reg[23]/NET0131  ;
  input \u0_uk_K_r14_reg[24]/NET0131  ;
  input \u0_uk_K_r14_reg[25]/NET0131  ;
  input \u0_uk_K_r14_reg[26]/NET0131  ;
  input \u0_uk_K_r14_reg[27]/NET0131  ;
  input \u0_uk_K_r14_reg[28]/NET0131  ;
  input \u0_uk_K_r14_reg[29]/NET0131  ;
  input \u0_uk_K_r14_reg[2]/NET0131  ;
  input \u0_uk_K_r14_reg[30]/NET0131  ;
  input \u0_uk_K_r14_reg[31]/NET0131  ;
  input \u0_uk_K_r14_reg[32]/NET0131  ;
  input \u0_uk_K_r14_reg[33]/NET0131  ;
  input \u0_uk_K_r14_reg[34]/NET0131  ;
  input \u0_uk_K_r14_reg[35]/P0001  ;
  input \u0_uk_K_r14_reg[36]/NET0131  ;
  input \u0_uk_K_r14_reg[37]/NET0131  ;
  input \u0_uk_K_r14_reg[38]/NET0131  ;
  input \u0_uk_K_r14_reg[39]/P0001  ;
  input \u0_uk_K_r14_reg[3]/NET0131  ;
  input \u0_uk_K_r14_reg[40]/NET0131  ;
  input \u0_uk_K_r14_reg[41]/NET0131  ;
  input \u0_uk_K_r14_reg[42]/P0001  ;
  input \u0_uk_K_r14_reg[43]/NET0131  ;
  input \u0_uk_K_r14_reg[44]/NET0131  ;
  input \u0_uk_K_r14_reg[45]/NET0131  ;
  input \u0_uk_K_r14_reg[46]/NET0131  ;
  input \u0_uk_K_r14_reg[47]/NET0131  ;
  input \u0_uk_K_r14_reg[48]/NET0131  ;
  input \u0_uk_K_r14_reg[49]/NET0131  ;
  input \u0_uk_K_r14_reg[4]/NET0131  ;
  input \u0_uk_K_r14_reg[50]/NET0131  ;
  input \u0_uk_K_r14_reg[51]/NET0131  ;
  input \u0_uk_K_r14_reg[52]/NET0131  ;
  input \u0_uk_K_r14_reg[53]/NET0131  ;
  input \u0_uk_K_r14_reg[54]/NET0131  ;
  input \u0_uk_K_r14_reg[55]/NET0131  ;
  input \u0_uk_K_r14_reg[5]/NET0131  ;
  input \u0_uk_K_r14_reg[6]/NET0131  ;
  input \u0_uk_K_r14_reg[7]/NET0131  ;
  input \u0_uk_K_r14_reg[8]/NET0131  ;
  input \u0_uk_K_r14_reg[9]/NET0131  ;
  input \u0_uk_K_r1_reg[0]/NET0131  ;
  input \u0_uk_K_r1_reg[10]/P0001  ;
  input \u0_uk_K_r1_reg[11]/NET0131  ;
  input \u0_uk_K_r1_reg[12]/NET0131  ;
  input \u0_uk_K_r1_reg[13]/NET0131  ;
  input \u0_uk_K_r1_reg[14]/NET0131  ;
  input \u0_uk_K_r1_reg[15]/NET0131  ;
  input \u0_uk_K_r1_reg[16]/NET0131  ;
  input \u0_uk_K_r1_reg[17]/NET0131  ;
  input \u0_uk_K_r1_reg[18]/NET0131  ;
  input \u0_uk_K_r1_reg[19]/NET0131  ;
  input \u0_uk_K_r1_reg[1]/NET0131  ;
  input \u0_uk_K_r1_reg[20]/NET0131  ;
  input \u0_uk_K_r1_reg[21]/NET0131  ;
  input \u0_uk_K_r1_reg[22]/NET0131  ;
  input \u0_uk_K_r1_reg[23]/NET0131  ;
  input \u0_uk_K_r1_reg[24]/NET0131  ;
  input \u0_uk_K_r1_reg[25]/NET0131  ;
  input \u0_uk_K_r1_reg[26]/NET0131  ;
  input \u0_uk_K_r1_reg[27]/NET0131  ;
  input \u0_uk_K_r1_reg[28]/NET0131  ;
  input \u0_uk_K_r1_reg[29]/NET0131  ;
  input \u0_uk_K_r1_reg[2]/NET0131  ;
  input \u0_uk_K_r1_reg[30]/NET0131  ;
  input \u0_uk_K_r1_reg[31]/NET0131  ;
  input \u0_uk_K_r1_reg[32]/NET0131  ;
  input \u0_uk_K_r1_reg[33]/NET0131  ;
  input \u0_uk_K_r1_reg[34]/NET0131  ;
  input \u0_uk_K_r1_reg[35]/NET0131  ;
  input \u0_uk_K_r1_reg[36]/NET0131  ;
  input \u0_uk_K_r1_reg[37]/NET0131  ;
  input \u0_uk_K_r1_reg[38]/NET0131  ;
  input \u0_uk_K_r1_reg[3]/NET0131  ;
  input \u0_uk_K_r1_reg[40]/NET0131  ;
  input \u0_uk_K_r1_reg[41]/NET0131  ;
  input \u0_uk_K_r1_reg[42]/NET0131  ;
  input \u0_uk_K_r1_reg[43]/NET0131  ;
  input \u0_uk_K_r1_reg[44]/P0001  ;
  input \u0_uk_K_r1_reg[45]/NET0131  ;
  input \u0_uk_K_r1_reg[46]/NET0131  ;
  input \u0_uk_K_r1_reg[47]/NET0131  ;
  input \u0_uk_K_r1_reg[48]/NET0131  ;
  input \u0_uk_K_r1_reg[49]/NET0131  ;
  input \u0_uk_K_r1_reg[4]/NET0131  ;
  input \u0_uk_K_r1_reg[50]/NET0131  ;
  input \u0_uk_K_r1_reg[51]/NET0131  ;
  input \u0_uk_K_r1_reg[52]/NET0131  ;
  input \u0_uk_K_r1_reg[53]/NET0131  ;
  input \u0_uk_K_r1_reg[54]/NET0131  ;
  input \u0_uk_K_r1_reg[55]/NET0131  ;
  input \u0_uk_K_r1_reg[5]/NET0131  ;
  input \u0_uk_K_r1_reg[6]/NET0131  ;
  input \u0_uk_K_r1_reg[7]/P0001  ;
  input \u0_uk_K_r1_reg[8]/NET0131  ;
  input \u0_uk_K_r1_reg[9]/NET0131  ;
  input \u0_uk_K_r2_reg[0]/NET0131  ;
  input \u0_uk_K_r2_reg[10]/NET0131  ;
  input \u0_uk_K_r2_reg[11]/NET0131  ;
  input \u0_uk_K_r2_reg[12]/NET0131  ;
  input \u0_uk_K_r2_reg[13]/NET0131  ;
  input \u0_uk_K_r2_reg[14]/NET0131  ;
  input \u0_uk_K_r2_reg[15]/NET0131  ;
  input \u0_uk_K_r2_reg[16]/NET0131  ;
  input \u0_uk_K_r2_reg[17]/NET0131  ;
  input \u0_uk_K_r2_reg[18]/NET0131  ;
  input \u0_uk_K_r2_reg[19]/NET0131  ;
  input \u0_uk_K_r2_reg[1]/NET0131  ;
  input \u0_uk_K_r2_reg[20]/NET0131  ;
  input \u0_uk_K_r2_reg[21]/NET0131  ;
  input \u0_uk_K_r2_reg[22]/NET0131  ;
  input \u0_uk_K_r2_reg[23]/NET0131  ;
  input \u0_uk_K_r2_reg[24]/NET0131  ;
  input \u0_uk_K_r2_reg[25]/NET0131  ;
  input \u0_uk_K_r2_reg[26]/NET0131  ;
  input \u0_uk_K_r2_reg[27]/P0001  ;
  input \u0_uk_K_r2_reg[28]/NET0131  ;
  input \u0_uk_K_r2_reg[29]/NET0131  ;
  input \u0_uk_K_r2_reg[2]/NET0131  ;
  input \u0_uk_K_r2_reg[31]/NET0131  ;
  input \u0_uk_K_r2_reg[32]/NET0131  ;
  input \u0_uk_K_r2_reg[33]/NET0131  ;
  input \u0_uk_K_r2_reg[34]/NET0131  ;
  input \u0_uk_K_r2_reg[35]/NET0131  ;
  input \u0_uk_K_r2_reg[36]/NET0131  ;
  input \u0_uk_K_r2_reg[37]/NET0131  ;
  input \u0_uk_K_r2_reg[38]/NET0131  ;
  input \u0_uk_K_r2_reg[39]/NET0131  ;
  input \u0_uk_K_r2_reg[3]/NET0131  ;
  input \u0_uk_K_r2_reg[40]/NET0131  ;
  input \u0_uk_K_r2_reg[41]/NET0131  ;
  input \u0_uk_K_r2_reg[42]/NET0131  ;
  input \u0_uk_K_r2_reg[43]/NET0131  ;
  input \u0_uk_K_r2_reg[44]/NET0131  ;
  input \u0_uk_K_r2_reg[45]/NET0131  ;
  input \u0_uk_K_r2_reg[46]/NET0131  ;
  input \u0_uk_K_r2_reg[47]/NET0131  ;
  input \u0_uk_K_r2_reg[48]/NET0131  ;
  input \u0_uk_K_r2_reg[49]/NET0131  ;
  input \u0_uk_K_r2_reg[4]/NET0131  ;
  input \u0_uk_K_r2_reg[50]/NET0131  ;
  input \u0_uk_K_r2_reg[51]/NET0131  ;
  input \u0_uk_K_r2_reg[52]/NET0131  ;
  input \u0_uk_K_r2_reg[53]/P0001  ;
  input \u0_uk_K_r2_reg[54]/NET0131  ;
  input \u0_uk_K_r2_reg[55]/NET0131  ;
  input \u0_uk_K_r2_reg[5]/NET0131  ;
  input \u0_uk_K_r2_reg[6]/NET0131  ;
  input \u0_uk_K_r2_reg[7]/NET0131  ;
  input \u0_uk_K_r2_reg[8]/NET0131  ;
  input \u0_uk_K_r2_reg[9]/NET0131  ;
  input \u0_uk_K_r3_reg[0]/NET0131  ;
  input \u0_uk_K_r3_reg[10]/NET0131  ;
  input \u0_uk_K_r3_reg[11]/NET0131  ;
  input \u0_uk_K_r3_reg[12]/NET0131  ;
  input \u0_uk_K_r3_reg[14]/NET0131  ;
  input \u0_uk_K_r3_reg[15]/NET0131  ;
  input \u0_uk_K_r3_reg[16]/NET0131  ;
  input \u0_uk_K_r3_reg[17]/NET0131  ;
  input \u0_uk_K_r3_reg[18]/NET0131  ;
  input \u0_uk_K_r3_reg[19]/NET0131  ;
  input \u0_uk_K_r3_reg[1]/NET0131  ;
  input \u0_uk_K_r3_reg[20]/NET0131  ;
  input \u0_uk_K_r3_reg[21]/NET0131  ;
  input \u0_uk_K_r3_reg[22]/NET0131  ;
  input \u0_uk_K_r3_reg[23]/NET0131  ;
  input \u0_uk_K_r3_reg[24]/NET0131  ;
  input \u0_uk_K_r3_reg[25]/NET0131  ;
  input \u0_uk_K_r3_reg[26]/NET0131  ;
  input \u0_uk_K_r3_reg[27]/NET0131  ;
  input \u0_uk_K_r3_reg[28]/NET0131  ;
  input \u0_uk_K_r3_reg[29]/NET0131  ;
  input \u0_uk_K_r3_reg[2]/NET0131  ;
  input \u0_uk_K_r3_reg[30]/NET0131  ;
  input \u0_uk_K_r3_reg[31]/NET0131  ;
  input \u0_uk_K_r3_reg[32]/NET0131  ;
  input \u0_uk_K_r3_reg[33]/NET0131  ;
  input \u0_uk_K_r3_reg[34]/NET0131  ;
  input \u0_uk_K_r3_reg[35]/NET0131  ;
  input \u0_uk_K_r3_reg[36]/NET0131  ;
  input \u0_uk_K_r3_reg[37]/NET0131  ;
  input \u0_uk_K_r3_reg[38]/NET0131  ;
  input \u0_uk_K_r3_reg[39]/NET0131  ;
  input \u0_uk_K_r3_reg[3]/NET0131  ;
  input \u0_uk_K_r3_reg[40]/NET0131  ;
  input \u0_uk_K_r3_reg[41]/NET0131  ;
  input \u0_uk_K_r3_reg[42]/NET0131  ;
  input \u0_uk_K_r3_reg[43]/NET0131  ;
  input \u0_uk_K_r3_reg[44]/NET0131  ;
  input \u0_uk_K_r3_reg[45]/P0001  ;
  input \u0_uk_K_r3_reg[46]/NET0131  ;
  input \u0_uk_K_r3_reg[47]/NET0131  ;
  input \u0_uk_K_r3_reg[48]/NET0131  ;
  input \u0_uk_K_r3_reg[49]/NET0131  ;
  input \u0_uk_K_r3_reg[4]/NET0131  ;
  input \u0_uk_K_r3_reg[50]/NET0131  ;
  input \u0_uk_K_r3_reg[51]/NET0131  ;
  input \u0_uk_K_r3_reg[52]/NET0131  ;
  input \u0_uk_K_r3_reg[53]/NET0131  ;
  input \u0_uk_K_r3_reg[54]/NET0131  ;
  input \u0_uk_K_r3_reg[55]/NET0131  ;
  input \u0_uk_K_r3_reg[5]/NET0131  ;
  input \u0_uk_K_r3_reg[6]/NET0131  ;
  input \u0_uk_K_r3_reg[7]/NET0131  ;
  input \u0_uk_K_r3_reg[8]/NET0131  ;
  input \u0_uk_K_r3_reg[9]/NET0131  ;
  input \u0_uk_K_r4_reg[0]/P0001  ;
  input \u0_uk_K_r4_reg[10]/NET0131  ;
  input \u0_uk_K_r4_reg[11]/NET0131  ;
  input \u0_uk_K_r4_reg[12]/NET0131  ;
  input \u0_uk_K_r4_reg[13]/NET0131  ;
  input \u0_uk_K_r4_reg[14]/NET0131  ;
  input \u0_uk_K_r4_reg[15]/NET0131  ;
  input \u0_uk_K_r4_reg[16]/NET0131  ;
  input \u0_uk_K_r4_reg[17]/NET0131  ;
  input \u0_uk_K_r4_reg[18]/NET0131  ;
  input \u0_uk_K_r4_reg[19]/NET0131  ;
  input \u0_uk_K_r4_reg[1]/NET0131  ;
  input \u0_uk_K_r4_reg[20]/NET0131  ;
  input \u0_uk_K_r4_reg[21]/NET0131  ;
  input \u0_uk_K_r4_reg[22]/NET0131  ;
  input \u0_uk_K_r4_reg[23]/P0001  ;
  input \u0_uk_K_r4_reg[25]/NET0131  ;
  input \u0_uk_K_r4_reg[26]/NET0131  ;
  input \u0_uk_K_r4_reg[27]/P0001  ;
  input \u0_uk_K_r4_reg[28]/NET0131  ;
  input \u0_uk_K_r4_reg[29]/NET0131  ;
  input \u0_uk_K_r4_reg[30]/NET0131  ;
  input \u0_uk_K_r4_reg[31]/P0001  ;
  input \u0_uk_K_r4_reg[32]/NET0131  ;
  input \u0_uk_K_r4_reg[33]/NET0131  ;
  input \u0_uk_K_r4_reg[34]/NET0131  ;
  input \u0_uk_K_r4_reg[35]/NET0131  ;
  input \u0_uk_K_r4_reg[36]/NET0131  ;
  input \u0_uk_K_r4_reg[37]/NET0131  ;
  input \u0_uk_K_r4_reg[38]/NET0131  ;
  input \u0_uk_K_r4_reg[39]/NET0131  ;
  input \u0_uk_K_r4_reg[3]/NET0131  ;
  input \u0_uk_K_r4_reg[40]/NET0131  ;
  input \u0_uk_K_r4_reg[41]/NET0131  ;
  input \u0_uk_K_r4_reg[42]/NET0131  ;
  input \u0_uk_K_r4_reg[43]/NET0131  ;
  input \u0_uk_K_r4_reg[44]/NET0131  ;
  input \u0_uk_K_r4_reg[45]/NET0131  ;
  input \u0_uk_K_r4_reg[46]/NET0131  ;
  input \u0_uk_K_r4_reg[47]/NET0131  ;
  input \u0_uk_K_r4_reg[48]/NET0131  ;
  input \u0_uk_K_r4_reg[49]/NET0131  ;
  input \u0_uk_K_r4_reg[4]/NET0131  ;
  input \u0_uk_K_r4_reg[50]/NET0131  ;
  input \u0_uk_K_r4_reg[51]/NET0131  ;
  input \u0_uk_K_r4_reg[52]/NET0131  ;
  input \u0_uk_K_r4_reg[53]/NET0131  ;
  input \u0_uk_K_r4_reg[54]/NET0131  ;
  input \u0_uk_K_r4_reg[55]/NET0131  ;
  input \u0_uk_K_r4_reg[5]/NET0131  ;
  input \u0_uk_K_r4_reg[6]/NET0131  ;
  input \u0_uk_K_r4_reg[7]/NET0131  ;
  input \u0_uk_K_r4_reg[8]/NET0131  ;
  input \u0_uk_K_r4_reg[9]/NET0131  ;
  input \u0_uk_K_r5_reg[0]/NET0131  ;
  input \u0_uk_K_r5_reg[10]/NET0131  ;
  input \u0_uk_K_r5_reg[11]/NET0131  ;
  input \u0_uk_K_r5_reg[12]/NET0131  ;
  input \u0_uk_K_r5_reg[13]/P0001  ;
  input \u0_uk_K_r5_reg[14]/NET0131  ;
  input \u0_uk_K_r5_reg[15]/NET0131  ;
  input \u0_uk_K_r5_reg[16]/NET0131  ;
  input \u0_uk_K_r5_reg[17]/NET0131  ;
  input \u0_uk_K_r5_reg[18]/NET0131  ;
  input \u0_uk_K_r5_reg[19]/NET0131  ;
  input \u0_uk_K_r5_reg[1]/NET0131  ;
  input \u0_uk_K_r5_reg[20]/NET0131  ;
  input \u0_uk_K_r5_reg[21]/NET0131  ;
  input \u0_uk_K_r5_reg[22]/NET0131  ;
  input \u0_uk_K_r5_reg[23]/NET0131  ;
  input \u0_uk_K_r5_reg[24]/NET0131  ;
  input \u0_uk_K_r5_reg[25]/NET0131  ;
  input \u0_uk_K_r5_reg[26]/NET0131  ;
  input \u0_uk_K_r5_reg[27]/NET0131  ;
  input \u0_uk_K_r5_reg[28]/NET0131  ;
  input \u0_uk_K_r5_reg[29]/NET0131  ;
  input \u0_uk_K_r5_reg[2]/NET0131  ;
  input \u0_uk_K_r5_reg[30]/NET0131  ;
  input \u0_uk_K_r5_reg[31]/NET0131  ;
  input \u0_uk_K_r5_reg[32]/NET0131  ;
  input \u0_uk_K_r5_reg[33]/NET0131  ;
  input \u0_uk_K_r5_reg[34]/NET0131  ;
  input \u0_uk_K_r5_reg[35]/NET0131  ;
  input \u0_uk_K_r5_reg[36]/NET0131  ;
  input \u0_uk_K_r5_reg[37]/P0001  ;
  input \u0_uk_K_r5_reg[38]/NET0131  ;
  input \u0_uk_K_r5_reg[39]/NET0131  ;
  input \u0_uk_K_r5_reg[3]/NET0131  ;
  input \u0_uk_K_r5_reg[40]/NET0131  ;
  input \u0_uk_K_r5_reg[41]/NET0131  ;
  input \u0_uk_K_r5_reg[42]/NET0131  ;
  input \u0_uk_K_r5_reg[43]/NET0131  ;
  input \u0_uk_K_r5_reg[44]/NET0131  ;
  input \u0_uk_K_r5_reg[46]/NET0131  ;
  input \u0_uk_K_r5_reg[47]/NET0131  ;
  input \u0_uk_K_r5_reg[48]/NET0131  ;
  input \u0_uk_K_r5_reg[49]/NET0131  ;
  input \u0_uk_K_r5_reg[4]/NET0131  ;
  input \u0_uk_K_r5_reg[50]/NET0131  ;
  input \u0_uk_K_r5_reg[51]/NET0131  ;
  input \u0_uk_K_r5_reg[52]/NET0131  ;
  input \u0_uk_K_r5_reg[53]/NET0131  ;
  input \u0_uk_K_r5_reg[54]/NET0131  ;
  input \u0_uk_K_r5_reg[55]/NET0131  ;
  input \u0_uk_K_r5_reg[5]/NET0131  ;
  input \u0_uk_K_r5_reg[6]/NET0131  ;
  input \u0_uk_K_r5_reg[7]/NET0131  ;
  input \u0_uk_K_r5_reg[8]/NET0131  ;
  input \u0_uk_K_r5_reg[9]/NET0131  ;
  input \u0_uk_K_r6_reg[0]/NET0131  ;
  input \u0_uk_K_r6_reg[10]/NET0131  ;
  input \u0_uk_K_r6_reg[11]/NET0131  ;
  input \u0_uk_K_r6_reg[12]/NET0131  ;
  input \u0_uk_K_r6_reg[13]/NET0131  ;
  input \u0_uk_K_r6_reg[14]/NET0131  ;
  input \u0_uk_K_r6_reg[15]/NET0131  ;
  input \u0_uk_K_r6_reg[16]/NET0131  ;
  input \u0_uk_K_r6_reg[17]/NET0131  ;
  input \u0_uk_K_r6_reg[18]/NET0131  ;
  input \u0_uk_K_r6_reg[19]/NET0131  ;
  input \u0_uk_K_r6_reg[1]/NET0131  ;
  input \u0_uk_K_r6_reg[20]/NET0131  ;
  input \u0_uk_K_r6_reg[21]/NET0131  ;
  input \u0_uk_K_r6_reg[22]/NET0131  ;
  input \u0_uk_K_r6_reg[23]/P0001  ;
  input \u0_uk_K_r6_reg[24]/NET0131  ;
  input \u0_uk_K_r6_reg[25]/NET0131  ;
  input \u0_uk_K_r6_reg[26]/P0001  ;
  input \u0_uk_K_r6_reg[27]/NET0131  ;
  input \u0_uk_K_r6_reg[28]/NET0131  ;
  input \u0_uk_K_r6_reg[29]/NET0131  ;
  input \u0_uk_K_r6_reg[2]/NET0131  ;
  input \u0_uk_K_r6_reg[30]/P0001  ;
  input \u0_uk_K_r6_reg[31]/NET0131  ;
  input \u0_uk_K_r6_reg[32]/NET0131  ;
  input \u0_uk_K_r6_reg[33]/NET0131  ;
  input \u0_uk_K_r6_reg[34]/NET0131  ;
  input \u0_uk_K_r6_reg[35]/NET0131  ;
  input \u0_uk_K_r6_reg[36]/NET0131  ;
  input \u0_uk_K_r6_reg[37]/NET0131  ;
  input \u0_uk_K_r6_reg[38]/NET0131  ;
  input \u0_uk_K_r6_reg[39]/NET0131  ;
  input \u0_uk_K_r6_reg[3]/NET0131  ;
  input \u0_uk_K_r6_reg[40]/NET0131  ;
  input \u0_uk_K_r6_reg[41]/NET0131  ;
  input \u0_uk_K_r6_reg[42]/NET0131  ;
  input \u0_uk_K_r6_reg[43]/NET0131  ;
  input \u0_uk_K_r6_reg[44]/NET0131  ;
  input \u0_uk_K_r6_reg[45]/NET0131  ;
  input \u0_uk_K_r6_reg[46]/NET0131  ;
  input \u0_uk_K_r6_reg[47]/NET0131  ;
  input \u0_uk_K_r6_reg[48]/NET0131  ;
  input \u0_uk_K_r6_reg[49]/NET0131  ;
  input \u0_uk_K_r6_reg[4]/NET0131  ;
  input \u0_uk_K_r6_reg[50]/NET0131  ;
  input \u0_uk_K_r6_reg[51]/NET0131  ;
  input \u0_uk_K_r6_reg[52]/NET0131  ;
  input \u0_uk_K_r6_reg[53]/NET0131  ;
  input \u0_uk_K_r6_reg[54]/NET0131  ;
  input \u0_uk_K_r6_reg[55]/P0001  ;
  input \u0_uk_K_r6_reg[5]/NET0131  ;
  input \u0_uk_K_r6_reg[6]/NET0131  ;
  input \u0_uk_K_r6_reg[7]/NET0131  ;
  input \u0_uk_K_r6_reg[8]/NET0131  ;
  input \u0_uk_K_r6_reg[9]/NET0131  ;
  input \u0_uk_K_r7_reg[0]/NET0131  ;
  input \u0_uk_K_r7_reg[10]/NET0131  ;
  input \u0_uk_K_r7_reg[11]/NET0131  ;
  input \u0_uk_K_r7_reg[12]/NET0131  ;
  input \u0_uk_K_r7_reg[13]/NET0131  ;
  input \u0_uk_K_r7_reg[14]/NET0131  ;
  input \u0_uk_K_r7_reg[15]/NET0131  ;
  input \u0_uk_K_r7_reg[16]/NET0131  ;
  input \u0_uk_K_r7_reg[17]/NET0131  ;
  input \u0_uk_K_r7_reg[18]/NET0131  ;
  input \u0_uk_K_r7_reg[19]/NET0131  ;
  input \u0_uk_K_r7_reg[1]/NET0131  ;
  input \u0_uk_K_r7_reg[20]/NET0131  ;
  input \u0_uk_K_r7_reg[21]/NET0131  ;
  input \u0_uk_K_r7_reg[22]/NET0131  ;
  input \u0_uk_K_r7_reg[23]/P0001  ;
  input \u0_uk_K_r7_reg[24]/NET0131  ;
  input \u0_uk_K_r7_reg[25]/NET0131  ;
  input \u0_uk_K_r7_reg[26]/P0001  ;
  input \u0_uk_K_r7_reg[27]/NET0131  ;
  input \u0_uk_K_r7_reg[28]/NET0131  ;
  input \u0_uk_K_r7_reg[29]/NET0131  ;
  input \u0_uk_K_r7_reg[2]/NET0131  ;
  input \u0_uk_K_r7_reg[30]/P0001  ;
  input \u0_uk_K_r7_reg[31]/NET0131  ;
  input \u0_uk_K_r7_reg[32]/NET0131  ;
  input \u0_uk_K_r7_reg[33]/NET0131  ;
  input \u0_uk_K_r7_reg[34]/NET0131  ;
  input \u0_uk_K_r7_reg[35]/NET0131  ;
  input \u0_uk_K_r7_reg[36]/NET0131  ;
  input \u0_uk_K_r7_reg[37]/NET0131  ;
  input \u0_uk_K_r7_reg[38]/NET0131  ;
  input \u0_uk_K_r7_reg[39]/NET0131  ;
  input \u0_uk_K_r7_reg[3]/NET0131  ;
  input \u0_uk_K_r7_reg[40]/NET0131  ;
  input \u0_uk_K_r7_reg[41]/NET0131  ;
  input \u0_uk_K_r7_reg[42]/NET0131  ;
  input \u0_uk_K_r7_reg[43]/NET0131  ;
  input \u0_uk_K_r7_reg[44]/NET0131  ;
  input \u0_uk_K_r7_reg[45]/NET0131  ;
  input \u0_uk_K_r7_reg[46]/NET0131  ;
  input \u0_uk_K_r7_reg[47]/NET0131  ;
  input \u0_uk_K_r7_reg[48]/NET0131  ;
  input \u0_uk_K_r7_reg[49]/NET0131  ;
  input \u0_uk_K_r7_reg[4]/NET0131  ;
  input \u0_uk_K_r7_reg[50]/NET0131  ;
  input \u0_uk_K_r7_reg[51]/NET0131  ;
  input \u0_uk_K_r7_reg[52]/NET0131  ;
  input \u0_uk_K_r7_reg[53]/NET0131  ;
  input \u0_uk_K_r7_reg[54]/NET0131  ;
  input \u0_uk_K_r7_reg[55]/P0001  ;
  input \u0_uk_K_r7_reg[5]/NET0131  ;
  input \u0_uk_K_r7_reg[6]/NET0131  ;
  input \u0_uk_K_r7_reg[7]/NET0131  ;
  input \u0_uk_K_r7_reg[8]/NET0131  ;
  input \u0_uk_K_r7_reg[9]/NET0131  ;
  input \u0_uk_K_r8_reg[0]/NET0131  ;
  input \u0_uk_K_r8_reg[10]/NET0131  ;
  input \u0_uk_K_r8_reg[11]/NET0131  ;
  input \u0_uk_K_r8_reg[12]/NET0131  ;
  input \u0_uk_K_r8_reg[13]/P0001  ;
  input \u0_uk_K_r8_reg[14]/NET0131  ;
  input \u0_uk_K_r8_reg[15]/NET0131  ;
  input \u0_uk_K_r8_reg[16]/NET0131  ;
  input \u0_uk_K_r8_reg[17]/NET0131  ;
  input \u0_uk_K_r8_reg[18]/NET0131  ;
  input \u0_uk_K_r8_reg[19]/NET0131  ;
  input \u0_uk_K_r8_reg[1]/NET0131  ;
  input \u0_uk_K_r8_reg[20]/NET0131  ;
  input \u0_uk_K_r8_reg[21]/NET0131  ;
  input \u0_uk_K_r8_reg[22]/NET0131  ;
  input \u0_uk_K_r8_reg[23]/NET0131  ;
  input \u0_uk_K_r8_reg[24]/NET0131  ;
  input \u0_uk_K_r8_reg[25]/NET0131  ;
  input \u0_uk_K_r8_reg[26]/NET0131  ;
  input \u0_uk_K_r8_reg[27]/NET0131  ;
  input \u0_uk_K_r8_reg[28]/NET0131  ;
  input \u0_uk_K_r8_reg[29]/NET0131  ;
  input \u0_uk_K_r8_reg[2]/NET0131  ;
  input \u0_uk_K_r8_reg[30]/NET0131  ;
  input \u0_uk_K_r8_reg[31]/NET0131  ;
  input \u0_uk_K_r8_reg[32]/NET0131  ;
  input \u0_uk_K_r8_reg[33]/NET0131  ;
  input \u0_uk_K_r8_reg[34]/NET0131  ;
  input \u0_uk_K_r8_reg[35]/NET0131  ;
  input \u0_uk_K_r8_reg[36]/NET0131  ;
  input \u0_uk_K_r8_reg[37]/P0001  ;
  input \u0_uk_K_r8_reg[38]/NET0131  ;
  input \u0_uk_K_r8_reg[39]/NET0131  ;
  input \u0_uk_K_r8_reg[3]/NET0131  ;
  input \u0_uk_K_r8_reg[40]/NET0131  ;
  input \u0_uk_K_r8_reg[41]/NET0131  ;
  input \u0_uk_K_r8_reg[42]/NET0131  ;
  input \u0_uk_K_r8_reg[43]/NET0131  ;
  input \u0_uk_K_r8_reg[44]/NET0131  ;
  input \u0_uk_K_r8_reg[46]/NET0131  ;
  input \u0_uk_K_r8_reg[47]/NET0131  ;
  input \u0_uk_K_r8_reg[48]/NET0131  ;
  input \u0_uk_K_r8_reg[49]/NET0131  ;
  input \u0_uk_K_r8_reg[4]/NET0131  ;
  input \u0_uk_K_r8_reg[50]/NET0131  ;
  input \u0_uk_K_r8_reg[51]/NET0131  ;
  input \u0_uk_K_r8_reg[52]/NET0131  ;
  input \u0_uk_K_r8_reg[53]/NET0131  ;
  input \u0_uk_K_r8_reg[54]/NET0131  ;
  input \u0_uk_K_r8_reg[55]/NET0131  ;
  input \u0_uk_K_r8_reg[5]/NET0131  ;
  input \u0_uk_K_r8_reg[6]/NET0131  ;
  input \u0_uk_K_r8_reg[7]/NET0131  ;
  input \u0_uk_K_r8_reg[8]/NET0131  ;
  input \u0_uk_K_r8_reg[9]/P0001  ;
  input \u0_uk_K_r9_reg[0]/P0001  ;
  input \u0_uk_K_r9_reg[10]/NET0131  ;
  input \u0_uk_K_r9_reg[11]/NET0131  ;
  input \u0_uk_K_r9_reg[12]/NET0131  ;
  input \u0_uk_K_r9_reg[13]/NET0131  ;
  input \u0_uk_K_r9_reg[14]/NET0131  ;
  input \u0_uk_K_r9_reg[15]/NET0131  ;
  input \u0_uk_K_r9_reg[16]/NET0131  ;
  input \u0_uk_K_r9_reg[17]/NET0131  ;
  input \u0_uk_K_r9_reg[18]/NET0131  ;
  input \u0_uk_K_r9_reg[19]/NET0131  ;
  input \u0_uk_K_r9_reg[1]/NET0131  ;
  input \u0_uk_K_r9_reg[20]/NET0131  ;
  input \u0_uk_K_r9_reg[21]/NET0131  ;
  input \u0_uk_K_r9_reg[22]/NET0131  ;
  input \u0_uk_K_r9_reg[23]/P0001  ;
  input \u0_uk_K_r9_reg[25]/NET0131  ;
  input \u0_uk_K_r9_reg[26]/NET0131  ;
  input \u0_uk_K_r9_reg[27]/P0001  ;
  input \u0_uk_K_r9_reg[28]/NET0131  ;
  input \u0_uk_K_r9_reg[29]/NET0131  ;
  input \u0_uk_K_r9_reg[30]/NET0131  ;
  input \u0_uk_K_r9_reg[31]/P0001  ;
  input \u0_uk_K_r9_reg[32]/NET0131  ;
  input \u0_uk_K_r9_reg[33]/NET0131  ;
  input \u0_uk_K_r9_reg[34]/NET0131  ;
  input \u0_uk_K_r9_reg[35]/NET0131  ;
  input \u0_uk_K_r9_reg[36]/NET0131  ;
  input \u0_uk_K_r9_reg[37]/NET0131  ;
  input \u0_uk_K_r9_reg[38]/NET0131  ;
  input \u0_uk_K_r9_reg[39]/NET0131  ;
  input \u0_uk_K_r9_reg[3]/NET0131  ;
  input \u0_uk_K_r9_reg[40]/NET0131  ;
  input \u0_uk_K_r9_reg[41]/NET0131  ;
  input \u0_uk_K_r9_reg[42]/NET0131  ;
  input \u0_uk_K_r9_reg[43]/NET0131  ;
  input \u0_uk_K_r9_reg[44]/NET0131  ;
  input \u0_uk_K_r9_reg[45]/NET0131  ;
  input \u0_uk_K_r9_reg[46]/NET0131  ;
  input \u0_uk_K_r9_reg[47]/NET0131  ;
  input \u0_uk_K_r9_reg[48]/NET0131  ;
  input \u0_uk_K_r9_reg[49]/NET0131  ;
  input \u0_uk_K_r9_reg[4]/NET0131  ;
  input \u0_uk_K_r9_reg[50]/NET0131  ;
  input \u0_uk_K_r9_reg[51]/NET0131  ;
  input \u0_uk_K_r9_reg[52]/NET0131  ;
  input \u0_uk_K_r9_reg[53]/NET0131  ;
  input \u0_uk_K_r9_reg[54]/NET0131  ;
  input \u0_uk_K_r9_reg[55]/NET0131  ;
  input \u0_uk_K_r9_reg[5]/NET0131  ;
  input \u0_uk_K_r9_reg[6]/NET0131  ;
  input \u0_uk_K_r9_reg[7]/NET0131  ;
  input \u0_uk_K_r9_reg[8]/NET0131  ;
  input \u0_uk_K_r9_reg[9]/NET0131  ;
  input \u1_L0_reg[10]/NET0131  ;
  input \u1_L0_reg[11]/NET0131  ;
  input \u1_L0_reg[12]/NET0131  ;
  input \u1_L0_reg[13]/NET0131  ;
  input \u1_L0_reg[14]/NET0131  ;
  input \u1_L0_reg[15]/P0001  ;
  input \u1_L0_reg[16]/NET0131  ;
  input \u1_L0_reg[17]/NET0131  ;
  input \u1_L0_reg[18]/NET0131  ;
  input \u1_L0_reg[19]/NET0131  ;
  input \u1_L0_reg[1]/NET0131  ;
  input \u1_L0_reg[20]/NET0131  ;
  input \u1_L0_reg[21]/NET0131  ;
  input \u1_L0_reg[22]/NET0131  ;
  input \u1_L0_reg[23]/NET0131  ;
  input \u1_L0_reg[24]/NET0131  ;
  input \u1_L0_reg[25]/NET0131  ;
  input \u1_L0_reg[26]/NET0131  ;
  input \u1_L0_reg[27]/NET0131  ;
  input \u1_L0_reg[28]/NET0131  ;
  input \u1_L0_reg[29]/NET0131  ;
  input \u1_L0_reg[2]/NET0131  ;
  input \u1_L0_reg[30]/NET0131  ;
  input \u1_L0_reg[31]/NET0131  ;
  input \u1_L0_reg[32]/NET0131  ;
  input \u1_L0_reg[3]/NET0131  ;
  input \u1_L0_reg[4]/NET0131  ;
  input \u1_L0_reg[5]/NET0131  ;
  input \u1_L0_reg[6]/NET0131  ;
  input \u1_L0_reg[7]/NET0131  ;
  input \u1_L0_reg[8]/NET0131  ;
  input \u1_L0_reg[9]/NET0131  ;
  input \u1_L10_reg[10]/NET0131  ;
  input \u1_L10_reg[11]/NET0131  ;
  input \u1_L10_reg[12]/NET0131  ;
  input \u1_L10_reg[13]/NET0131  ;
  input \u1_L10_reg[14]/NET0131  ;
  input \u1_L10_reg[15]/P0001  ;
  input \u1_L10_reg[16]/NET0131  ;
  input \u1_L10_reg[17]/NET0131  ;
  input \u1_L10_reg[18]/P0001  ;
  input \u1_L10_reg[19]/P0001  ;
  input \u1_L10_reg[1]/NET0131  ;
  input \u1_L10_reg[20]/NET0131  ;
  input \u1_L10_reg[21]/NET0131  ;
  input \u1_L10_reg[22]/NET0131  ;
  input \u1_L10_reg[23]/NET0131  ;
  input \u1_L10_reg[24]/NET0131  ;
  input \u1_L10_reg[25]/NET0131  ;
  input \u1_L10_reg[26]/NET0131  ;
  input \u1_L10_reg[27]/NET0131  ;
  input \u1_L10_reg[28]/NET0131  ;
  input \u1_L10_reg[29]/NET0131  ;
  input \u1_L10_reg[2]/NET0131  ;
  input \u1_L10_reg[30]/NET0131  ;
  input \u1_L10_reg[31]/NET0131  ;
  input \u1_L10_reg[32]/NET0131  ;
  input \u1_L10_reg[3]/NET0131  ;
  input \u1_L10_reg[4]/NET0131  ;
  input \u1_L10_reg[5]/NET0131  ;
  input \u1_L10_reg[6]/NET0131  ;
  input \u1_L10_reg[7]/NET0131  ;
  input \u1_L10_reg[8]/NET0131  ;
  input \u1_L10_reg[9]/NET0131  ;
  input \u1_L11_reg[10]/NET0131  ;
  input \u1_L11_reg[11]/NET0131  ;
  input \u1_L11_reg[12]/NET0131  ;
  input \u1_L11_reg[13]/NET0131  ;
  input \u1_L11_reg[14]/NET0131  ;
  input \u1_L11_reg[15]/P0001  ;
  input \u1_L11_reg[16]/NET0131  ;
  input \u1_L11_reg[17]/NET0131  ;
  input \u1_L11_reg[18]/P0001  ;
  input \u1_L11_reg[19]/P0001  ;
  input \u1_L11_reg[1]/NET0131  ;
  input \u1_L11_reg[20]/NET0131  ;
  input \u1_L11_reg[21]/NET0131  ;
  input \u1_L11_reg[22]/NET0131  ;
  input \u1_L11_reg[23]/NET0131  ;
  input \u1_L11_reg[24]/NET0131  ;
  input \u1_L11_reg[25]/NET0131  ;
  input \u1_L11_reg[26]/NET0131  ;
  input \u1_L11_reg[27]/NET0131  ;
  input \u1_L11_reg[28]/NET0131  ;
  input \u1_L11_reg[29]/NET0131  ;
  input \u1_L11_reg[2]/NET0131  ;
  input \u1_L11_reg[30]/NET0131  ;
  input \u1_L11_reg[31]/NET0131  ;
  input \u1_L11_reg[32]/NET0131  ;
  input \u1_L11_reg[3]/NET0131  ;
  input \u1_L11_reg[4]/NET0131  ;
  input \u1_L11_reg[5]/NET0131  ;
  input \u1_L11_reg[6]/NET0131  ;
  input \u1_L11_reg[7]/NET0131  ;
  input \u1_L11_reg[8]/NET0131  ;
  input \u1_L11_reg[9]/NET0131  ;
  input \u1_L12_reg[10]/NET0131  ;
  input \u1_L12_reg[11]/NET0131  ;
  input \u1_L12_reg[12]/NET0131  ;
  input \u1_L12_reg[13]/NET0131  ;
  input \u1_L12_reg[14]/NET0131  ;
  input \u1_L12_reg[15]/P0001  ;
  input \u1_L12_reg[16]/NET0131  ;
  input \u1_L12_reg[17]/NET0131  ;
  input \u1_L12_reg[18]/P0001  ;
  input \u1_L12_reg[19]/NET0131  ;
  input \u1_L12_reg[1]/NET0131  ;
  input \u1_L12_reg[20]/NET0131  ;
  input \u1_L12_reg[21]/NET0131  ;
  input \u1_L12_reg[22]/NET0131  ;
  input \u1_L12_reg[23]/P0001  ;
  input \u1_L12_reg[24]/NET0131  ;
  input \u1_L12_reg[25]/NET0131  ;
  input \u1_L12_reg[26]/NET0131  ;
  input \u1_L12_reg[27]/NET0131  ;
  input \u1_L12_reg[28]/NET0131  ;
  input \u1_L12_reg[29]/NET0131  ;
  input \u1_L12_reg[2]/NET0131  ;
  input \u1_L12_reg[30]/NET0131  ;
  input \u1_L12_reg[31]/NET0131  ;
  input \u1_L12_reg[32]/NET0131  ;
  input \u1_L12_reg[3]/NET0131  ;
  input \u1_L12_reg[4]/NET0131  ;
  input \u1_L12_reg[5]/NET0131  ;
  input \u1_L12_reg[6]/NET0131  ;
  input \u1_L12_reg[7]/NET0131  ;
  input \u1_L12_reg[8]/NET0131  ;
  input \u1_L12_reg[9]/NET0131  ;
  input \u1_L13_reg[10]/NET0131  ;
  input \u1_L13_reg[11]/NET0131  ;
  input \u1_L13_reg[12]/NET0131  ;
  input \u1_L13_reg[13]/NET0131  ;
  input \u1_L13_reg[14]/NET0131  ;
  input \u1_L13_reg[15]/P0001  ;
  input \u1_L13_reg[16]/NET0131  ;
  input \u1_L13_reg[17]/NET0131  ;
  input \u1_L13_reg[18]/P0001  ;
  input \u1_L13_reg[19]/P0001  ;
  input \u1_L13_reg[1]/NET0131  ;
  input \u1_L13_reg[20]/NET0131  ;
  input \u1_L13_reg[21]/NET0131  ;
  input \u1_L13_reg[22]/NET0131  ;
  input \u1_L13_reg[23]/P0001  ;
  input \u1_L13_reg[24]/NET0131  ;
  input \u1_L13_reg[25]/NET0131  ;
  input \u1_L13_reg[26]/NET0131  ;
  input \u1_L13_reg[27]/NET0131  ;
  input \u1_L13_reg[28]/NET0131  ;
  input \u1_L13_reg[29]/NET0131  ;
  input \u1_L13_reg[2]/NET0131  ;
  input \u1_L13_reg[30]/NET0131  ;
  input \u1_L13_reg[31]/NET0131  ;
  input \u1_L13_reg[32]/NET0131  ;
  input \u1_L13_reg[3]/NET0131  ;
  input \u1_L13_reg[4]/NET0131  ;
  input \u1_L13_reg[5]/NET0131  ;
  input \u1_L13_reg[6]/NET0131  ;
  input \u1_L13_reg[7]/NET0131  ;
  input \u1_L13_reg[8]/NET0131  ;
  input \u1_L13_reg[9]/NET0131  ;
  input \u1_L14_reg[10]/P0001  ;
  input \u1_L14_reg[11]/P0001  ;
  input \u1_L14_reg[12]/P0001  ;
  input \u1_L14_reg[13]/P0001  ;
  input \u1_L14_reg[14]/P0001  ;
  input \u1_L14_reg[15]/P0001  ;
  input \u1_L14_reg[16]/P0001  ;
  input \u1_L14_reg[17]/P0001  ;
  input \u1_L14_reg[18]/P0001  ;
  input \u1_L14_reg[19]/P0001  ;
  input \u1_L14_reg[1]/P0001  ;
  input \u1_L14_reg[20]/P0001  ;
  input \u1_L14_reg[21]/P0001  ;
  input \u1_L14_reg[22]/P0001  ;
  input \u1_L14_reg[23]/P0001  ;
  input \u1_L14_reg[24]/P0001  ;
  input \u1_L14_reg[25]/P0001  ;
  input \u1_L14_reg[26]/P0001  ;
  input \u1_L14_reg[27]/P0001  ;
  input \u1_L14_reg[28]/P0001  ;
  input \u1_L14_reg[29]/P0001  ;
  input \u1_L14_reg[2]/P0001  ;
  input \u1_L14_reg[30]/P0001  ;
  input \u1_L14_reg[31]/P0001  ;
  input \u1_L14_reg[32]/P0001  ;
  input \u1_L14_reg[3]/P0001  ;
  input \u1_L14_reg[4]/P0001  ;
  input \u1_L14_reg[5]/P0001  ;
  input \u1_L14_reg[6]/P0001  ;
  input \u1_L14_reg[7]/P0001  ;
  input \u1_L14_reg[8]/P0001  ;
  input \u1_L14_reg[9]/P0001  ;
  input \u1_L1_reg[10]/NET0131  ;
  input \u1_L1_reg[11]/NET0131  ;
  input \u1_L1_reg[12]/NET0131  ;
  input \u1_L1_reg[13]/NET0131  ;
  input \u1_L1_reg[14]/NET0131  ;
  input \u1_L1_reg[15]/P0001  ;
  input \u1_L1_reg[16]/NET0131  ;
  input \u1_L1_reg[17]/NET0131  ;
  input \u1_L1_reg[18]/NET0131  ;
  input \u1_L1_reg[19]/P0001  ;
  input \u1_L1_reg[1]/NET0131  ;
  input \u1_L1_reg[20]/NET0131  ;
  input \u1_L1_reg[21]/NET0131  ;
  input \u1_L1_reg[22]/NET0131  ;
  input \u1_L1_reg[23]/NET0131  ;
  input \u1_L1_reg[24]/NET0131  ;
  input \u1_L1_reg[25]/NET0131  ;
  input \u1_L1_reg[26]/NET0131  ;
  input \u1_L1_reg[27]/NET0131  ;
  input \u1_L1_reg[28]/NET0131  ;
  input \u1_L1_reg[29]/NET0131  ;
  input \u1_L1_reg[2]/NET0131  ;
  input \u1_L1_reg[30]/NET0131  ;
  input \u1_L1_reg[31]/NET0131  ;
  input \u1_L1_reg[32]/NET0131  ;
  input \u1_L1_reg[3]/NET0131  ;
  input \u1_L1_reg[4]/NET0131  ;
  input \u1_L1_reg[5]/NET0131  ;
  input \u1_L1_reg[6]/NET0131  ;
  input \u1_L1_reg[7]/NET0131  ;
  input \u1_L1_reg[8]/NET0131  ;
  input \u1_L1_reg[9]/NET0131  ;
  input \u1_L2_reg[10]/NET0131  ;
  input \u1_L2_reg[11]/NET0131  ;
  input \u1_L2_reg[12]/NET0131  ;
  input \u1_L2_reg[13]/NET0131  ;
  input \u1_L2_reg[14]/NET0131  ;
  input \u1_L2_reg[15]/P0001  ;
  input \u1_L2_reg[16]/NET0131  ;
  input \u1_L2_reg[17]/NET0131  ;
  input \u1_L2_reg[18]/NET0131  ;
  input \u1_L2_reg[19]/NET0131  ;
  input \u1_L2_reg[1]/NET0131  ;
  input \u1_L2_reg[20]/NET0131  ;
  input \u1_L2_reg[21]/NET0131  ;
  input \u1_L2_reg[22]/NET0131  ;
  input \u1_L2_reg[23]/NET0131  ;
  input \u1_L2_reg[24]/NET0131  ;
  input \u1_L2_reg[25]/NET0131  ;
  input \u1_L2_reg[26]/NET0131  ;
  input \u1_L2_reg[27]/NET0131  ;
  input \u1_L2_reg[28]/NET0131  ;
  input \u1_L2_reg[29]/NET0131  ;
  input \u1_L2_reg[2]/NET0131  ;
  input \u1_L2_reg[30]/NET0131  ;
  input \u1_L2_reg[31]/NET0131  ;
  input \u1_L2_reg[32]/NET0131  ;
  input \u1_L2_reg[3]/NET0131  ;
  input \u1_L2_reg[4]/NET0131  ;
  input \u1_L2_reg[5]/NET0131  ;
  input \u1_L2_reg[6]/NET0131  ;
  input \u1_L2_reg[7]/NET0131  ;
  input \u1_L2_reg[8]/NET0131  ;
  input \u1_L2_reg[9]/NET0131  ;
  input \u1_L3_reg[10]/NET0131  ;
  input \u1_L3_reg[11]/NET0131  ;
  input \u1_L3_reg[12]/NET0131  ;
  input \u1_L3_reg[13]/NET0131  ;
  input \u1_L3_reg[14]/NET0131  ;
  input \u1_L3_reg[15]/P0001  ;
  input \u1_L3_reg[16]/NET0131  ;
  input \u1_L3_reg[17]/NET0131  ;
  input \u1_L3_reg[18]/NET0131  ;
  input \u1_L3_reg[19]/NET0131  ;
  input \u1_L3_reg[1]/NET0131  ;
  input \u1_L3_reg[20]/NET0131  ;
  input \u1_L3_reg[21]/NET0131  ;
  input \u1_L3_reg[22]/NET0131  ;
  input \u1_L3_reg[23]/NET0131  ;
  input \u1_L3_reg[24]/NET0131  ;
  input \u1_L3_reg[25]/NET0131  ;
  input \u1_L3_reg[26]/NET0131  ;
  input \u1_L3_reg[27]/NET0131  ;
  input \u1_L3_reg[28]/NET0131  ;
  input \u1_L3_reg[29]/NET0131  ;
  input \u1_L3_reg[2]/NET0131  ;
  input \u1_L3_reg[30]/NET0131  ;
  input \u1_L3_reg[31]/NET0131  ;
  input \u1_L3_reg[32]/NET0131  ;
  input \u1_L3_reg[3]/NET0131  ;
  input \u1_L3_reg[4]/NET0131  ;
  input \u1_L3_reg[5]/NET0131  ;
  input \u1_L3_reg[6]/NET0131  ;
  input \u1_L3_reg[7]/NET0131  ;
  input \u1_L3_reg[8]/NET0131  ;
  input \u1_L3_reg[9]/NET0131  ;
  input \u1_L4_reg[10]/NET0131  ;
  input \u1_L4_reg[11]/P0001  ;
  input \u1_L4_reg[12]/NET0131  ;
  input \u1_L4_reg[13]/NET0131  ;
  input \u1_L4_reg[14]/NET0131  ;
  input \u1_L4_reg[15]/P0001  ;
  input \u1_L4_reg[16]/NET0131  ;
  input \u1_L4_reg[17]/NET0131  ;
  input \u1_L4_reg[18]/NET0131  ;
  input \u1_L4_reg[19]/P0001  ;
  input \u1_L4_reg[1]/NET0131  ;
  input \u1_L4_reg[20]/NET0131  ;
  input \u1_L4_reg[21]/NET0131  ;
  input \u1_L4_reg[22]/NET0131  ;
  input \u1_L4_reg[23]/NET0131  ;
  input \u1_L4_reg[24]/NET0131  ;
  input \u1_L4_reg[25]/NET0131  ;
  input \u1_L4_reg[26]/NET0131  ;
  input \u1_L4_reg[27]/NET0131  ;
  input \u1_L4_reg[28]/NET0131  ;
  input \u1_L4_reg[29]/NET0131  ;
  input \u1_L4_reg[2]/NET0131  ;
  input \u1_L4_reg[30]/NET0131  ;
  input \u1_L4_reg[31]/NET0131  ;
  input \u1_L4_reg[32]/NET0131  ;
  input \u1_L4_reg[3]/NET0131  ;
  input \u1_L4_reg[4]/NET0131  ;
  input \u1_L4_reg[5]/NET0131  ;
  input \u1_L4_reg[6]/NET0131  ;
  input \u1_L4_reg[7]/NET0131  ;
  input \u1_L4_reg[8]/NET0131  ;
  input \u1_L4_reg[9]/NET0131  ;
  input \u1_L5_reg[10]/NET0131  ;
  input \u1_L5_reg[11]/NET0131  ;
  input \u1_L5_reg[12]/NET0131  ;
  input \u1_L5_reg[13]/NET0131  ;
  input \u1_L5_reg[14]/NET0131  ;
  input \u1_L5_reg[15]/P0001  ;
  input \u1_L5_reg[16]/NET0131  ;
  input \u1_L5_reg[17]/NET0131  ;
  input \u1_L5_reg[18]/NET0131  ;
  input \u1_L5_reg[19]/NET0131  ;
  input \u1_L5_reg[1]/NET0131  ;
  input \u1_L5_reg[20]/NET0131  ;
  input \u1_L5_reg[21]/NET0131  ;
  input \u1_L5_reg[22]/NET0131  ;
  input \u1_L5_reg[23]/NET0131  ;
  input \u1_L5_reg[24]/NET0131  ;
  input \u1_L5_reg[25]/NET0131  ;
  input \u1_L5_reg[26]/NET0131  ;
  input \u1_L5_reg[27]/NET0131  ;
  input \u1_L5_reg[28]/NET0131  ;
  input \u1_L5_reg[29]/NET0131  ;
  input \u1_L5_reg[2]/NET0131  ;
  input \u1_L5_reg[30]/NET0131  ;
  input \u1_L5_reg[31]/NET0131  ;
  input \u1_L5_reg[32]/NET0131  ;
  input \u1_L5_reg[3]/NET0131  ;
  input \u1_L5_reg[4]/NET0131  ;
  input \u1_L5_reg[5]/NET0131  ;
  input \u1_L5_reg[6]/NET0131  ;
  input \u1_L5_reg[7]/NET0131  ;
  input \u1_L5_reg[8]/NET0131  ;
  input \u1_L5_reg[9]/NET0131  ;
  input \u1_L6_reg[10]/NET0131  ;
  input \u1_L6_reg[11]/NET0131  ;
  input \u1_L6_reg[12]/NET0131  ;
  input \u1_L6_reg[13]/NET0131  ;
  input \u1_L6_reg[14]/NET0131  ;
  input \u1_L6_reg[15]/P0001  ;
  input \u1_L6_reg[16]/NET0131  ;
  input \u1_L6_reg[17]/NET0131  ;
  input \u1_L6_reg[18]/NET0131  ;
  input \u1_L6_reg[19]/NET0131  ;
  input \u1_L6_reg[1]/NET0131  ;
  input \u1_L6_reg[20]/NET0131  ;
  input \u1_L6_reg[21]/NET0131  ;
  input \u1_L6_reg[22]/NET0131  ;
  input \u1_L6_reg[23]/NET0131  ;
  input \u1_L6_reg[24]/NET0131  ;
  input \u1_L6_reg[25]/NET0131  ;
  input \u1_L6_reg[26]/NET0131  ;
  input \u1_L6_reg[27]/NET0131  ;
  input \u1_L6_reg[28]/NET0131  ;
  input \u1_L6_reg[29]/NET0131  ;
  input \u1_L6_reg[2]/NET0131  ;
  input \u1_L6_reg[30]/NET0131  ;
  input \u1_L6_reg[31]/NET0131  ;
  input \u1_L6_reg[32]/NET0131  ;
  input \u1_L6_reg[3]/NET0131  ;
  input \u1_L6_reg[4]/NET0131  ;
  input \u1_L6_reg[5]/NET0131  ;
  input \u1_L6_reg[6]/NET0131  ;
  input \u1_L6_reg[7]/NET0131  ;
  input \u1_L6_reg[8]/NET0131  ;
  input \u1_L6_reg[9]/NET0131  ;
  input \u1_L7_reg[10]/NET0131  ;
  input \u1_L7_reg[11]/NET0131  ;
  input \u1_L7_reg[12]/NET0131  ;
  input \u1_L7_reg[13]/NET0131  ;
  input \u1_L7_reg[14]/NET0131  ;
  input \u1_L7_reg[15]/P0001  ;
  input \u1_L7_reg[16]/NET0131  ;
  input \u1_L7_reg[17]/NET0131  ;
  input \u1_L7_reg[18]/NET0131  ;
  input \u1_L7_reg[19]/P0001  ;
  input \u1_L7_reg[1]/NET0131  ;
  input \u1_L7_reg[20]/NET0131  ;
  input \u1_L7_reg[21]/NET0131  ;
  input \u1_L7_reg[22]/NET0131  ;
  input \u1_L7_reg[23]/NET0131  ;
  input \u1_L7_reg[24]/NET0131  ;
  input \u1_L7_reg[25]/NET0131  ;
  input \u1_L7_reg[26]/NET0131  ;
  input \u1_L7_reg[27]/NET0131  ;
  input \u1_L7_reg[28]/NET0131  ;
  input \u1_L7_reg[29]/NET0131  ;
  input \u1_L7_reg[2]/NET0131  ;
  input \u1_L7_reg[30]/NET0131  ;
  input \u1_L7_reg[31]/NET0131  ;
  input \u1_L7_reg[32]/NET0131  ;
  input \u1_L7_reg[3]/NET0131  ;
  input \u1_L7_reg[4]/NET0131  ;
  input \u1_L7_reg[5]/NET0131  ;
  input \u1_L7_reg[6]/NET0131  ;
  input \u1_L7_reg[7]/NET0131  ;
  input \u1_L7_reg[8]/NET0131  ;
  input \u1_L7_reg[9]/NET0131  ;
  input \u1_L8_reg[10]/NET0131  ;
  input \u1_L8_reg[11]/NET0131  ;
  input \u1_L8_reg[12]/NET0131  ;
  input \u1_L8_reg[13]/NET0131  ;
  input \u1_L8_reg[14]/NET0131  ;
  input \u1_L8_reg[15]/P0001  ;
  input \u1_L8_reg[16]/NET0131  ;
  input \u1_L8_reg[17]/NET0131  ;
  input \u1_L8_reg[18]/NET0131  ;
  input \u1_L8_reg[19]/P0001  ;
  input \u1_L8_reg[1]/NET0131  ;
  input \u1_L8_reg[20]/NET0131  ;
  input \u1_L8_reg[21]/NET0131  ;
  input \u1_L8_reg[22]/NET0131  ;
  input \u1_L8_reg[23]/NET0131  ;
  input \u1_L8_reg[24]/NET0131  ;
  input \u1_L8_reg[25]/NET0131  ;
  input \u1_L8_reg[26]/NET0131  ;
  input \u1_L8_reg[27]/NET0131  ;
  input \u1_L8_reg[28]/NET0131  ;
  input \u1_L8_reg[29]/NET0131  ;
  input \u1_L8_reg[2]/NET0131  ;
  input \u1_L8_reg[30]/NET0131  ;
  input \u1_L8_reg[31]/NET0131  ;
  input \u1_L8_reg[32]/NET0131  ;
  input \u1_L8_reg[3]/NET0131  ;
  input \u1_L8_reg[4]/NET0131  ;
  input \u1_L8_reg[5]/NET0131  ;
  input \u1_L8_reg[6]/NET0131  ;
  input \u1_L8_reg[7]/NET0131  ;
  input \u1_L8_reg[8]/NET0131  ;
  input \u1_L8_reg[9]/NET0131  ;
  input \u1_L9_reg[10]/NET0131  ;
  input \u1_L9_reg[11]/NET0131  ;
  input \u1_L9_reg[12]/NET0131  ;
  input \u1_L9_reg[13]/NET0131  ;
  input \u1_L9_reg[14]/NET0131  ;
  input \u1_L9_reg[15]/P0001  ;
  input \u1_L9_reg[16]/NET0131  ;
  input \u1_L9_reg[17]/NET0131  ;
  input \u1_L9_reg[18]/P0001  ;
  input \u1_L9_reg[19]/NET0131  ;
  input \u1_L9_reg[1]/NET0131  ;
  input \u1_L9_reg[20]/NET0131  ;
  input \u1_L9_reg[21]/NET0131  ;
  input \u1_L9_reg[22]/NET0131  ;
  input \u1_L9_reg[23]/NET0131  ;
  input \u1_L9_reg[24]/NET0131  ;
  input \u1_L9_reg[25]/NET0131  ;
  input \u1_L9_reg[26]/NET0131  ;
  input \u1_L9_reg[27]/NET0131  ;
  input \u1_L9_reg[28]/NET0131  ;
  input \u1_L9_reg[29]/NET0131  ;
  input \u1_L9_reg[2]/NET0131  ;
  input \u1_L9_reg[30]/NET0131  ;
  input \u1_L9_reg[31]/NET0131  ;
  input \u1_L9_reg[32]/NET0131  ;
  input \u1_L9_reg[3]/NET0131  ;
  input \u1_L9_reg[4]/NET0131  ;
  input \u1_L9_reg[5]/NET0131  ;
  input \u1_L9_reg[6]/NET0131  ;
  input \u1_L9_reg[7]/NET0131  ;
  input \u1_L9_reg[8]/NET0131  ;
  input \u1_L9_reg[9]/NET0131  ;
  input \u1_R0_reg[10]/NET0131  ;
  input \u1_R0_reg[11]/NET0131  ;
  input \u1_R0_reg[12]/NET0131  ;
  input \u1_R0_reg[13]/NET0131  ;
  input \u1_R0_reg[14]/NET0131  ;
  input \u1_R0_reg[15]/NET0131  ;
  input \u1_R0_reg[16]/NET0131  ;
  input \u1_R0_reg[17]/NET0131  ;
  input \u1_R0_reg[18]/NET0131  ;
  input \u1_R0_reg[19]/NET0131  ;
  input \u1_R0_reg[1]/NET0131  ;
  input \u1_R0_reg[20]/NET0131  ;
  input \u1_R0_reg[21]/NET0131  ;
  input \u1_R0_reg[22]/NET0131  ;
  input \u1_R0_reg[23]/NET0131  ;
  input \u1_R0_reg[24]/NET0131  ;
  input \u1_R0_reg[25]/NET0131  ;
  input \u1_R0_reg[26]/NET0131  ;
  input \u1_R0_reg[27]/NET0131  ;
  input \u1_R0_reg[28]/NET0131  ;
  input \u1_R0_reg[29]/NET0131  ;
  input \u1_R0_reg[2]/NET0131  ;
  input \u1_R0_reg[30]/NET0131  ;
  input \u1_R0_reg[31]/P0001  ;
  input \u1_R0_reg[32]/NET0131  ;
  input \u1_R0_reg[3]/NET0131  ;
  input \u1_R0_reg[4]/NET0131  ;
  input \u1_R0_reg[5]/NET0131  ;
  input \u1_R0_reg[6]/NET0131  ;
  input \u1_R0_reg[7]/NET0131  ;
  input \u1_R0_reg[8]/NET0131  ;
  input \u1_R0_reg[9]/NET0131  ;
  input \u1_R10_reg[10]/NET0131  ;
  input \u1_R10_reg[11]/NET0131  ;
  input \u1_R10_reg[12]/NET0131  ;
  input \u1_R10_reg[13]/NET0131  ;
  input \u1_R10_reg[14]/NET0131  ;
  input \u1_R10_reg[15]/NET0131  ;
  input \u1_R10_reg[16]/NET0131  ;
  input \u1_R10_reg[17]/NET0131  ;
  input \u1_R10_reg[18]/NET0131  ;
  input \u1_R10_reg[19]/NET0131  ;
  input \u1_R10_reg[1]/NET0131  ;
  input \u1_R10_reg[20]/NET0131  ;
  input \u1_R10_reg[21]/NET0131  ;
  input \u1_R10_reg[22]/NET0131  ;
  input \u1_R10_reg[23]/NET0131  ;
  input \u1_R10_reg[24]/NET0131  ;
  input \u1_R10_reg[25]/NET0131  ;
  input \u1_R10_reg[26]/NET0131  ;
  input \u1_R10_reg[27]/NET0131  ;
  input \u1_R10_reg[28]/NET0131  ;
  input \u1_R10_reg[29]/NET0131  ;
  input \u1_R10_reg[2]/NET0131  ;
  input \u1_R10_reg[30]/NET0131  ;
  input \u1_R10_reg[31]/P0001  ;
  input \u1_R10_reg[32]/NET0131  ;
  input \u1_R10_reg[3]/NET0131  ;
  input \u1_R10_reg[4]/NET0131  ;
  input \u1_R10_reg[5]/NET0131  ;
  input \u1_R10_reg[6]/NET0131  ;
  input \u1_R10_reg[7]/NET0131  ;
  input \u1_R10_reg[8]/NET0131  ;
  input \u1_R10_reg[9]/NET0131  ;
  input \u1_R11_reg[10]/NET0131  ;
  input \u1_R11_reg[11]/NET0131  ;
  input \u1_R11_reg[12]/NET0131  ;
  input \u1_R11_reg[13]/NET0131  ;
  input \u1_R11_reg[14]/NET0131  ;
  input \u1_R11_reg[15]/NET0131  ;
  input \u1_R11_reg[16]/NET0131  ;
  input \u1_R11_reg[17]/NET0131  ;
  input \u1_R11_reg[18]/NET0131  ;
  input \u1_R11_reg[19]/NET0131  ;
  input \u1_R11_reg[1]/NET0131  ;
  input \u1_R11_reg[20]/NET0131  ;
  input \u1_R11_reg[21]/NET0131  ;
  input \u1_R11_reg[22]/NET0131  ;
  input \u1_R11_reg[23]/NET0131  ;
  input \u1_R11_reg[24]/NET0131  ;
  input \u1_R11_reg[25]/NET0131  ;
  input \u1_R11_reg[26]/NET0131  ;
  input \u1_R11_reg[27]/NET0131  ;
  input \u1_R11_reg[28]/NET0131  ;
  input \u1_R11_reg[29]/NET0131  ;
  input \u1_R11_reg[2]/NET0131  ;
  input \u1_R11_reg[30]/NET0131  ;
  input \u1_R11_reg[31]/NET0131  ;
  input \u1_R11_reg[32]/NET0131  ;
  input \u1_R11_reg[3]/NET0131  ;
  input \u1_R11_reg[4]/NET0131  ;
  input \u1_R11_reg[5]/NET0131  ;
  input \u1_R11_reg[6]/NET0131  ;
  input \u1_R11_reg[7]/NET0131  ;
  input \u1_R11_reg[8]/NET0131  ;
  input \u1_R11_reg[9]/NET0131  ;
  input \u1_R12_reg[10]/NET0131  ;
  input \u1_R12_reg[11]/NET0131  ;
  input \u1_R12_reg[12]/NET0131  ;
  input \u1_R12_reg[13]/NET0131  ;
  input \u1_R12_reg[14]/NET0131  ;
  input \u1_R12_reg[15]/NET0131  ;
  input \u1_R12_reg[16]/NET0131  ;
  input \u1_R12_reg[17]/NET0131  ;
  input \u1_R12_reg[18]/NET0131  ;
  input \u1_R12_reg[19]/NET0131  ;
  input \u1_R12_reg[1]/NET0131  ;
  input \u1_R12_reg[20]/NET0131  ;
  input \u1_R12_reg[21]/NET0131  ;
  input \u1_R12_reg[22]/NET0131  ;
  input \u1_R12_reg[23]/NET0131  ;
  input \u1_R12_reg[24]/NET0131  ;
  input \u1_R12_reg[25]/NET0131  ;
  input \u1_R12_reg[26]/NET0131  ;
  input \u1_R12_reg[27]/NET0131  ;
  input \u1_R12_reg[28]/NET0131  ;
  input \u1_R12_reg[29]/NET0131  ;
  input \u1_R12_reg[2]/NET0131  ;
  input \u1_R12_reg[30]/NET0131  ;
  input \u1_R12_reg[31]/NET0131  ;
  input \u1_R12_reg[32]/NET0131  ;
  input \u1_R12_reg[3]/NET0131  ;
  input \u1_R12_reg[4]/NET0131  ;
  input \u1_R12_reg[5]/NET0131  ;
  input \u1_R12_reg[6]/NET0131  ;
  input \u1_R12_reg[7]/NET0131  ;
  input \u1_R12_reg[8]/NET0131  ;
  input \u1_R12_reg[9]/NET0131  ;
  input \u1_R13_reg[10]/NET0131  ;
  input \u1_R13_reg[11]/P0001  ;
  input \u1_R13_reg[12]/NET0131  ;
  input \u1_R13_reg[13]/NET0131  ;
  input \u1_R13_reg[14]/NET0131  ;
  input \u1_R13_reg[15]/NET0131  ;
  input \u1_R13_reg[16]/NET0131  ;
  input \u1_R13_reg[17]/NET0131  ;
  input \u1_R13_reg[18]/NET0131  ;
  input \u1_R13_reg[19]/NET0131  ;
  input \u1_R13_reg[1]/NET0131  ;
  input \u1_R13_reg[20]/NET0131  ;
  input \u1_R13_reg[21]/NET0131  ;
  input \u1_R13_reg[22]/NET0131  ;
  input \u1_R13_reg[23]/P0001  ;
  input \u1_R13_reg[24]/NET0131  ;
  input \u1_R13_reg[25]/NET0131  ;
  input \u1_R13_reg[26]/NET0131  ;
  input \u1_R13_reg[27]/P0001  ;
  input \u1_R13_reg[28]/NET0131  ;
  input \u1_R13_reg[29]/NET0131  ;
  input \u1_R13_reg[2]/NET0131  ;
  input \u1_R13_reg[30]/NET0131  ;
  input \u1_R13_reg[31]/P0001  ;
  input \u1_R13_reg[32]/NET0131  ;
  input \u1_R13_reg[3]/NET0131  ;
  input \u1_R13_reg[4]/NET0131  ;
  input \u1_R13_reg[5]/NET0131  ;
  input \u1_R13_reg[6]/NET0131  ;
  input \u1_R13_reg[7]/NET0131  ;
  input \u1_R13_reg[8]/NET0131  ;
  input \u1_R13_reg[9]/NET0131  ;
  input \u1_R14_reg[10]/P0001  ;
  input \u1_R14_reg[11]/P0001  ;
  input \u1_R14_reg[12]/NET0131  ;
  input \u1_R14_reg[13]/NET0131  ;
  input \u1_R14_reg[14]/NET0131  ;
  input \u1_R14_reg[15]/NET0131  ;
  input \u1_R14_reg[16]/NET0131  ;
  input \u1_R14_reg[17]/NET0131  ;
  input \u1_R14_reg[18]/NET0131  ;
  input \u1_R14_reg[19]/P0001  ;
  input \u1_R14_reg[1]/NET0131  ;
  input \u1_R14_reg[20]/NET0131  ;
  input \u1_R14_reg[21]/NET0131  ;
  input \u1_R14_reg[22]/P0001  ;
  input \u1_R14_reg[23]/P0001  ;
  input \u1_R14_reg[24]/NET0131  ;
  input \u1_R14_reg[25]/NET0131  ;
  input \u1_R14_reg[26]/NET0131  ;
  input \u1_R14_reg[27]/P0001  ;
  input \u1_R14_reg[28]/NET0131  ;
  input \u1_R14_reg[29]/NET0131  ;
  input \u1_R14_reg[2]/NET0131  ;
  input \u1_R14_reg[30]/NET0131  ;
  input \u1_R14_reg[31]/P0001  ;
  input \u1_R14_reg[32]/NET0131  ;
  input \u1_R14_reg[3]/NET0131  ;
  input \u1_R14_reg[4]/NET0131  ;
  input \u1_R14_reg[5]/NET0131  ;
  input \u1_R14_reg[6]/NET0131  ;
  input \u1_R14_reg[7]/P0001  ;
  input \u1_R14_reg[8]/NET0131  ;
  input \u1_R14_reg[9]/NET0131  ;
  input \u1_R1_reg[10]/NET0131  ;
  input \u1_R1_reg[11]/NET0131  ;
  input \u1_R1_reg[12]/NET0131  ;
  input \u1_R1_reg[13]/NET0131  ;
  input \u1_R1_reg[14]/NET0131  ;
  input \u1_R1_reg[15]/NET0131  ;
  input \u1_R1_reg[16]/NET0131  ;
  input \u1_R1_reg[17]/NET0131  ;
  input \u1_R1_reg[18]/NET0131  ;
  input \u1_R1_reg[19]/NET0131  ;
  input \u1_R1_reg[1]/NET0131  ;
  input \u1_R1_reg[20]/NET0131  ;
  input \u1_R1_reg[21]/NET0131  ;
  input \u1_R1_reg[22]/NET0131  ;
  input \u1_R1_reg[23]/NET0131  ;
  input \u1_R1_reg[24]/NET0131  ;
  input \u1_R1_reg[25]/NET0131  ;
  input \u1_R1_reg[26]/NET0131  ;
  input \u1_R1_reg[27]/NET0131  ;
  input \u1_R1_reg[28]/NET0131  ;
  input \u1_R1_reg[29]/NET0131  ;
  input \u1_R1_reg[2]/NET0131  ;
  input \u1_R1_reg[30]/NET0131  ;
  input \u1_R1_reg[31]/P0001  ;
  input \u1_R1_reg[32]/NET0131  ;
  input \u1_R1_reg[3]/NET0131  ;
  input \u1_R1_reg[4]/NET0131  ;
  input \u1_R1_reg[5]/NET0131  ;
  input \u1_R1_reg[6]/NET0131  ;
  input \u1_R1_reg[7]/NET0131  ;
  input \u1_R1_reg[8]/NET0131  ;
  input \u1_R1_reg[9]/NET0131  ;
  input \u1_R2_reg[10]/NET0131  ;
  input \u1_R2_reg[11]/NET0131  ;
  input \u1_R2_reg[12]/NET0131  ;
  input \u1_R2_reg[13]/NET0131  ;
  input \u1_R2_reg[14]/NET0131  ;
  input \u1_R2_reg[15]/NET0131  ;
  input \u1_R2_reg[16]/NET0131  ;
  input \u1_R2_reg[17]/NET0131  ;
  input \u1_R2_reg[18]/NET0131  ;
  input \u1_R2_reg[19]/NET0131  ;
  input \u1_R2_reg[1]/NET0131  ;
  input \u1_R2_reg[20]/NET0131  ;
  input \u1_R2_reg[21]/NET0131  ;
  input \u1_R2_reg[22]/NET0131  ;
  input \u1_R2_reg[23]/NET0131  ;
  input \u1_R2_reg[24]/NET0131  ;
  input \u1_R2_reg[25]/NET0131  ;
  input \u1_R2_reg[26]/NET0131  ;
  input \u1_R2_reg[27]/NET0131  ;
  input \u1_R2_reg[28]/NET0131  ;
  input \u1_R2_reg[29]/NET0131  ;
  input \u1_R2_reg[2]/NET0131  ;
  input \u1_R2_reg[30]/NET0131  ;
  input \u1_R2_reg[31]/P0001  ;
  input \u1_R2_reg[32]/NET0131  ;
  input \u1_R2_reg[3]/NET0131  ;
  input \u1_R2_reg[4]/NET0131  ;
  input \u1_R2_reg[5]/NET0131  ;
  input \u1_R2_reg[6]/NET0131  ;
  input \u1_R2_reg[7]/NET0131  ;
  input \u1_R2_reg[8]/NET0131  ;
  input \u1_R2_reg[9]/NET0131  ;
  input \u1_R3_reg[10]/NET0131  ;
  input \u1_R3_reg[11]/NET0131  ;
  input \u1_R3_reg[12]/NET0131  ;
  input \u1_R3_reg[13]/NET0131  ;
  input \u1_R3_reg[14]/NET0131  ;
  input \u1_R3_reg[15]/NET0131  ;
  input \u1_R3_reg[16]/NET0131  ;
  input \u1_R3_reg[17]/NET0131  ;
  input \u1_R3_reg[18]/NET0131  ;
  input \u1_R3_reg[19]/NET0131  ;
  input \u1_R3_reg[1]/NET0131  ;
  input \u1_R3_reg[20]/NET0131  ;
  input \u1_R3_reg[21]/NET0131  ;
  input \u1_R3_reg[22]/NET0131  ;
  input \u1_R3_reg[23]/NET0131  ;
  input \u1_R3_reg[24]/NET0131  ;
  input \u1_R3_reg[25]/NET0131  ;
  input \u1_R3_reg[26]/NET0131  ;
  input \u1_R3_reg[27]/NET0131  ;
  input \u1_R3_reg[28]/NET0131  ;
  input \u1_R3_reg[29]/NET0131  ;
  input \u1_R3_reg[2]/NET0131  ;
  input \u1_R3_reg[30]/NET0131  ;
  input \u1_R3_reg[31]/P0001  ;
  input \u1_R3_reg[32]/NET0131  ;
  input \u1_R3_reg[3]/NET0131  ;
  input \u1_R3_reg[4]/NET0131  ;
  input \u1_R3_reg[5]/NET0131  ;
  input \u1_R3_reg[6]/NET0131  ;
  input \u1_R3_reg[7]/NET0131  ;
  input \u1_R3_reg[8]/NET0131  ;
  input \u1_R3_reg[9]/NET0131  ;
  input \u1_R4_reg[10]/NET0131  ;
  input \u1_R4_reg[11]/P0001  ;
  input \u1_R4_reg[12]/NET0131  ;
  input \u1_R4_reg[13]/NET0131  ;
  input \u1_R4_reg[14]/NET0131  ;
  input \u1_R4_reg[15]/NET0131  ;
  input \u1_R4_reg[16]/NET0131  ;
  input \u1_R4_reg[17]/NET0131  ;
  input \u1_R4_reg[18]/NET0131  ;
  input \u1_R4_reg[19]/NET0131  ;
  input \u1_R4_reg[1]/NET0131  ;
  input \u1_R4_reg[20]/NET0131  ;
  input \u1_R4_reg[21]/NET0131  ;
  input \u1_R4_reg[22]/NET0131  ;
  input \u1_R4_reg[23]/NET0131  ;
  input \u1_R4_reg[24]/NET0131  ;
  input \u1_R4_reg[25]/NET0131  ;
  input \u1_R4_reg[26]/NET0131  ;
  input \u1_R4_reg[27]/NET0131  ;
  input \u1_R4_reg[28]/NET0131  ;
  input \u1_R4_reg[29]/NET0131  ;
  input \u1_R4_reg[2]/NET0131  ;
  input \u1_R4_reg[30]/NET0131  ;
  input \u1_R4_reg[31]/P0001  ;
  input \u1_R4_reg[32]/NET0131  ;
  input \u1_R4_reg[3]/NET0131  ;
  input \u1_R4_reg[4]/NET0131  ;
  input \u1_R4_reg[5]/NET0131  ;
  input \u1_R4_reg[6]/NET0131  ;
  input \u1_R4_reg[7]/NET0131  ;
  input \u1_R4_reg[8]/NET0131  ;
  input \u1_R4_reg[9]/NET0131  ;
  input \u1_R5_reg[10]/NET0131  ;
  input \u1_R5_reg[11]/NET0131  ;
  input \u1_R5_reg[12]/NET0131  ;
  input \u1_R5_reg[13]/NET0131  ;
  input \u1_R5_reg[14]/NET0131  ;
  input \u1_R5_reg[15]/NET0131  ;
  input \u1_R5_reg[16]/NET0131  ;
  input \u1_R5_reg[17]/NET0131  ;
  input \u1_R5_reg[18]/NET0131  ;
  input \u1_R5_reg[19]/NET0131  ;
  input \u1_R5_reg[1]/NET0131  ;
  input \u1_R5_reg[20]/NET0131  ;
  input \u1_R5_reg[21]/NET0131  ;
  input \u1_R5_reg[22]/NET0131  ;
  input \u1_R5_reg[23]/NET0131  ;
  input \u1_R5_reg[24]/NET0131  ;
  input \u1_R5_reg[25]/NET0131  ;
  input \u1_R5_reg[26]/NET0131  ;
  input \u1_R5_reg[27]/NET0131  ;
  input \u1_R5_reg[28]/NET0131  ;
  input \u1_R5_reg[29]/NET0131  ;
  input \u1_R5_reg[2]/NET0131  ;
  input \u1_R5_reg[30]/NET0131  ;
  input \u1_R5_reg[31]/P0001  ;
  input \u1_R5_reg[32]/NET0131  ;
  input \u1_R5_reg[3]/NET0131  ;
  input \u1_R5_reg[4]/NET0131  ;
  input \u1_R5_reg[5]/NET0131  ;
  input \u1_R5_reg[6]/NET0131  ;
  input \u1_R5_reg[7]/NET0131  ;
  input \u1_R5_reg[8]/NET0131  ;
  input \u1_R5_reg[9]/NET0131  ;
  input \u1_R6_reg[10]/NET0131  ;
  input \u1_R6_reg[11]/NET0131  ;
  input \u1_R6_reg[12]/NET0131  ;
  input \u1_R6_reg[13]/NET0131  ;
  input \u1_R6_reg[14]/NET0131  ;
  input \u1_R6_reg[15]/NET0131  ;
  input \u1_R6_reg[16]/NET0131  ;
  input \u1_R6_reg[17]/NET0131  ;
  input \u1_R6_reg[18]/NET0131  ;
  input \u1_R6_reg[19]/NET0131  ;
  input \u1_R6_reg[1]/NET0131  ;
  input \u1_R6_reg[20]/NET0131  ;
  input \u1_R6_reg[21]/NET0131  ;
  input \u1_R6_reg[22]/NET0131  ;
  input \u1_R6_reg[23]/NET0131  ;
  input \u1_R6_reg[24]/NET0131  ;
  input \u1_R6_reg[25]/NET0131  ;
  input \u1_R6_reg[26]/NET0131  ;
  input \u1_R6_reg[27]/NET0131  ;
  input \u1_R6_reg[28]/NET0131  ;
  input \u1_R6_reg[29]/NET0131  ;
  input \u1_R6_reg[2]/NET0131  ;
  input \u1_R6_reg[30]/NET0131  ;
  input \u1_R6_reg[31]/P0001  ;
  input \u1_R6_reg[32]/NET0131  ;
  input \u1_R6_reg[3]/NET0131  ;
  input \u1_R6_reg[4]/NET0131  ;
  input \u1_R6_reg[5]/NET0131  ;
  input \u1_R6_reg[6]/NET0131  ;
  input \u1_R6_reg[7]/NET0131  ;
  input \u1_R6_reg[8]/NET0131  ;
  input \u1_R6_reg[9]/NET0131  ;
  input \u1_R7_reg[10]/NET0131  ;
  input \u1_R7_reg[11]/NET0131  ;
  input \u1_R7_reg[12]/NET0131  ;
  input \u1_R7_reg[13]/NET0131  ;
  input \u1_R7_reg[14]/NET0131  ;
  input \u1_R7_reg[15]/NET0131  ;
  input \u1_R7_reg[16]/NET0131  ;
  input \u1_R7_reg[17]/NET0131  ;
  input \u1_R7_reg[18]/NET0131  ;
  input \u1_R7_reg[19]/NET0131  ;
  input \u1_R7_reg[1]/NET0131  ;
  input \u1_R7_reg[20]/NET0131  ;
  input \u1_R7_reg[21]/NET0131  ;
  input \u1_R7_reg[22]/NET0131  ;
  input \u1_R7_reg[23]/NET0131  ;
  input \u1_R7_reg[24]/NET0131  ;
  input \u1_R7_reg[25]/NET0131  ;
  input \u1_R7_reg[26]/NET0131  ;
  input \u1_R7_reg[27]/NET0131  ;
  input \u1_R7_reg[28]/NET0131  ;
  input \u1_R7_reg[29]/NET0131  ;
  input \u1_R7_reg[2]/NET0131  ;
  input \u1_R7_reg[30]/NET0131  ;
  input \u1_R7_reg[31]/P0001  ;
  input \u1_R7_reg[32]/NET0131  ;
  input \u1_R7_reg[3]/NET0131  ;
  input \u1_R7_reg[4]/NET0131  ;
  input \u1_R7_reg[5]/NET0131  ;
  input \u1_R7_reg[6]/NET0131  ;
  input \u1_R7_reg[7]/NET0131  ;
  input \u1_R7_reg[8]/NET0131  ;
  input \u1_R7_reg[9]/NET0131  ;
  input \u1_R8_reg[10]/NET0131  ;
  input \u1_R8_reg[11]/NET0131  ;
  input \u1_R8_reg[12]/NET0131  ;
  input \u1_R8_reg[13]/NET0131  ;
  input \u1_R8_reg[14]/NET0131  ;
  input \u1_R8_reg[15]/NET0131  ;
  input \u1_R8_reg[16]/NET0131  ;
  input \u1_R8_reg[17]/NET0131  ;
  input \u1_R8_reg[18]/NET0131  ;
  input \u1_R8_reg[19]/NET0131  ;
  input \u1_R8_reg[1]/NET0131  ;
  input \u1_R8_reg[20]/NET0131  ;
  input \u1_R8_reg[21]/NET0131  ;
  input \u1_R8_reg[22]/NET0131  ;
  input \u1_R8_reg[23]/NET0131  ;
  input \u1_R8_reg[24]/NET0131  ;
  input \u1_R8_reg[25]/NET0131  ;
  input \u1_R8_reg[26]/NET0131  ;
  input \u1_R8_reg[27]/NET0131  ;
  input \u1_R8_reg[28]/NET0131  ;
  input \u1_R8_reg[29]/NET0131  ;
  input \u1_R8_reg[2]/NET0131  ;
  input \u1_R8_reg[30]/NET0131  ;
  input \u1_R8_reg[31]/P0001  ;
  input \u1_R8_reg[32]/NET0131  ;
  input \u1_R8_reg[3]/NET0131  ;
  input \u1_R8_reg[4]/NET0131  ;
  input \u1_R8_reg[5]/NET0131  ;
  input \u1_R8_reg[6]/NET0131  ;
  input \u1_R8_reg[7]/NET0131  ;
  input \u1_R8_reg[8]/NET0131  ;
  input \u1_R8_reg[9]/NET0131  ;
  input \u1_R9_reg[10]/NET0131  ;
  input \u1_R9_reg[11]/NET0131  ;
  input \u1_R9_reg[12]/NET0131  ;
  input \u1_R9_reg[13]/NET0131  ;
  input \u1_R9_reg[14]/NET0131  ;
  input \u1_R9_reg[15]/NET0131  ;
  input \u1_R9_reg[16]/NET0131  ;
  input \u1_R9_reg[17]/NET0131  ;
  input \u1_R9_reg[18]/NET0131  ;
  input \u1_R9_reg[19]/NET0131  ;
  input \u1_R9_reg[1]/NET0131  ;
  input \u1_R9_reg[20]/NET0131  ;
  input \u1_R9_reg[21]/NET0131  ;
  input \u1_R9_reg[22]/NET0131  ;
  input \u1_R9_reg[23]/NET0131  ;
  input \u1_R9_reg[24]/NET0131  ;
  input \u1_R9_reg[25]/NET0131  ;
  input \u1_R9_reg[26]/NET0131  ;
  input \u1_R9_reg[27]/NET0131  ;
  input \u1_R9_reg[28]/NET0131  ;
  input \u1_R9_reg[29]/NET0131  ;
  input \u1_R9_reg[2]/NET0131  ;
  input \u1_R9_reg[30]/NET0131  ;
  input \u1_R9_reg[31]/NET0131  ;
  input \u1_R9_reg[32]/NET0131  ;
  input \u1_R9_reg[3]/NET0131  ;
  input \u1_R9_reg[4]/NET0131  ;
  input \u1_R9_reg[5]/NET0131  ;
  input \u1_R9_reg[6]/NET0131  ;
  input \u1_R9_reg[7]/NET0131  ;
  input \u1_R9_reg[8]/NET0131  ;
  input \u1_R9_reg[9]/NET0131  ;
  input \u1_desIn_r_reg[0]/NET0131  ;
  input \u1_desIn_r_reg[10]/NET0131  ;
  input \u1_desIn_r_reg[11]/NET0131  ;
  input \u1_desIn_r_reg[12]/NET0131  ;
  input \u1_desIn_r_reg[13]/NET0131  ;
  input \u1_desIn_r_reg[14]/NET0131  ;
  input \u1_desIn_r_reg[15]/NET0131  ;
  input \u1_desIn_r_reg[16]/NET0131  ;
  input \u1_desIn_r_reg[17]/NET0131  ;
  input \u1_desIn_r_reg[18]/P0001  ;
  input \u1_desIn_r_reg[19]/NET0131  ;
  input \u1_desIn_r_reg[1]/NET0131  ;
  input \u1_desIn_r_reg[20]/NET0131  ;
  input \u1_desIn_r_reg[21]/NET0131  ;
  input \u1_desIn_r_reg[22]/NET0131  ;
  input \u1_desIn_r_reg[23]/NET0131  ;
  input \u1_desIn_r_reg[24]/NET0131  ;
  input \u1_desIn_r_reg[25]/NET0131  ;
  input \u1_desIn_r_reg[26]/NET0131  ;
  input \u1_desIn_r_reg[27]/NET0131  ;
  input \u1_desIn_r_reg[28]/NET0131  ;
  input \u1_desIn_r_reg[29]/NET0131  ;
  input \u1_desIn_r_reg[2]/NET0131  ;
  input \u1_desIn_r_reg[30]/NET0131  ;
  input \u1_desIn_r_reg[31]/NET0131  ;
  input \u1_desIn_r_reg[32]/NET0131  ;
  input \u1_desIn_r_reg[33]/NET0131  ;
  input \u1_desIn_r_reg[34]/NET0131  ;
  input \u1_desIn_r_reg[35]/NET0131  ;
  input \u1_desIn_r_reg[36]/NET0131  ;
  input \u1_desIn_r_reg[37]/NET0131  ;
  input \u1_desIn_r_reg[38]/NET0131  ;
  input \u1_desIn_r_reg[39]/NET0131  ;
  input \u1_desIn_r_reg[3]/NET0131  ;
  input \u1_desIn_r_reg[40]/NET0131  ;
  input \u1_desIn_r_reg[41]/NET0131  ;
  input \u1_desIn_r_reg[42]/NET0131  ;
  input \u1_desIn_r_reg[43]/NET0131  ;
  input \u1_desIn_r_reg[44]/NET0131  ;
  input \u1_desIn_r_reg[45]/NET0131  ;
  input \u1_desIn_r_reg[46]/NET0131  ;
  input \u1_desIn_r_reg[47]/NET0131  ;
  input \u1_desIn_r_reg[48]/NET0131  ;
  input \u1_desIn_r_reg[49]/NET0131  ;
  input \u1_desIn_r_reg[4]/NET0131  ;
  input \u1_desIn_r_reg[50]/NET0131  ;
  input \u1_desIn_r_reg[51]/NET0131  ;
  input \u1_desIn_r_reg[52]/P0001  ;
  input \u1_desIn_r_reg[53]/NET0131  ;
  input \u1_desIn_r_reg[54]/NET0131  ;
  input \u1_desIn_r_reg[55]/NET0131  ;
  input \u1_desIn_r_reg[56]/NET0131  ;
  input \u1_desIn_r_reg[57]/NET0131  ;
  input \u1_desIn_r_reg[58]/NET0131  ;
  input \u1_desIn_r_reg[59]/NET0131  ;
  input \u1_desIn_r_reg[5]/NET0131  ;
  input \u1_desIn_r_reg[60]/NET0131  ;
  input \u1_desIn_r_reg[61]/NET0131  ;
  input \u1_desIn_r_reg[62]/NET0131  ;
  input \u1_desIn_r_reg[63]/NET0131  ;
  input \u1_desIn_r_reg[6]/NET0131  ;
  input \u1_desIn_r_reg[7]/NET0131  ;
  input \u1_desIn_r_reg[8]/NET0131  ;
  input \u1_desIn_r_reg[9]/NET0131  ;
  input \u1_key_r_reg[0]/NET0131  ;
  input \u1_key_r_reg[10]/NET0131  ;
  input \u1_key_r_reg[11]/NET0131  ;
  input \u1_key_r_reg[12]/NET0131  ;
  input \u1_key_r_reg[13]/NET0131  ;
  input \u1_key_r_reg[14]/NET0131  ;
  input \u1_key_r_reg[15]/NET0131  ;
  input \u1_key_r_reg[16]/NET0131  ;
  input \u1_key_r_reg[17]/NET0131  ;
  input \u1_key_r_reg[18]/NET0131  ;
  input \u1_key_r_reg[19]/NET0131  ;
  input \u1_key_r_reg[1]/NET0131  ;
  input \u1_key_r_reg[20]/NET0131  ;
  input \u1_key_r_reg[21]/NET0131  ;
  input \u1_key_r_reg[22]/NET0131  ;
  input \u1_key_r_reg[23]/NET0131  ;
  input \u1_key_r_reg[24]/NET0131  ;
  input \u1_key_r_reg[25]/NET0131  ;
  input \u1_key_r_reg[26]/NET0131  ;
  input \u1_key_r_reg[27]/NET0131  ;
  input \u1_key_r_reg[28]/NET0131  ;
  input \u1_key_r_reg[29]/NET0131  ;
  input \u1_key_r_reg[2]/NET0131  ;
  input \u1_key_r_reg[30]/NET0131  ;
  input \u1_key_r_reg[31]/NET0131  ;
  input \u1_key_r_reg[32]/NET0131  ;
  input \u1_key_r_reg[33]/NET0131  ;
  input \u1_key_r_reg[34]/NET0131  ;
  input \u1_key_r_reg[35]/P0001  ;
  input \u1_key_r_reg[36]/NET0131  ;
  input \u1_key_r_reg[37]/NET0131  ;
  input \u1_key_r_reg[38]/NET0131  ;
  input \u1_key_r_reg[39]/P0001  ;
  input \u1_key_r_reg[3]/NET0131  ;
  input \u1_key_r_reg[40]/NET0131  ;
  input \u1_key_r_reg[41]/NET0131  ;
  input \u1_key_r_reg[42]/P0001  ;
  input \u1_key_r_reg[43]/NET0131  ;
  input \u1_key_r_reg[44]/NET0131  ;
  input \u1_key_r_reg[45]/NET0131  ;
  input \u1_key_r_reg[46]/NET0131  ;
  input \u1_key_r_reg[47]/NET0131  ;
  input \u1_key_r_reg[48]/NET0131  ;
  input \u1_key_r_reg[49]/NET0131  ;
  input \u1_key_r_reg[4]/NET0131  ;
  input \u1_key_r_reg[50]/NET0131  ;
  input \u1_key_r_reg[51]/NET0131  ;
  input \u1_key_r_reg[52]/NET0131  ;
  input \u1_key_r_reg[53]/NET0131  ;
  input \u1_key_r_reg[54]/NET0131  ;
  input \u1_key_r_reg[55]/NET0131  ;
  input \u1_key_r_reg[5]/NET0131  ;
  input \u1_key_r_reg[6]/NET0131  ;
  input \u1_key_r_reg[7]/NET0131  ;
  input \u1_key_r_reg[8]/NET0131  ;
  input \u1_key_r_reg[9]/NET0131  ;
  input \u1_uk_K_r0_reg[0]/NET0131  ;
  input \u1_uk_K_r0_reg[10]/NET0131  ;
  input \u1_uk_K_r0_reg[11]/NET0131  ;
  input \u1_uk_K_r0_reg[12]/NET0131  ;
  input \u1_uk_K_r0_reg[13]/NET0131  ;
  input \u1_uk_K_r0_reg[14]/NET0131  ;
  input \u1_uk_K_r0_reg[15]/NET0131  ;
  input \u1_uk_K_r0_reg[16]/NET0131  ;
  input \u1_uk_K_r0_reg[17]/NET0131  ;
  input \u1_uk_K_r0_reg[18]/NET0131  ;
  input \u1_uk_K_r0_reg[19]/NET0131  ;
  input \u1_uk_K_r0_reg[20]/NET0131  ;
  input \u1_uk_K_r0_reg[21]/NET0131  ;
  input \u1_uk_K_r0_reg[22]/NET0131  ;
  input \u1_uk_K_r0_reg[23]/NET0131  ;
  input \u1_uk_K_r0_reg[24]/NET0131  ;
  input \u1_uk_K_r0_reg[25]/P0001  ;
  input \u1_uk_K_r0_reg[26]/NET0131  ;
  input \u1_uk_K_r0_reg[27]/NET0131  ;
  input \u1_uk_K_r0_reg[28]/NET0131  ;
  input \u1_uk_K_r0_reg[29]/NET0131  ;
  input \u1_uk_K_r0_reg[2]/NET0131  ;
  input \u1_uk_K_r0_reg[30]/NET0131  ;
  input \u1_uk_K_r0_reg[31]/NET0131  ;
  input \u1_uk_K_r0_reg[32]/NET0131  ;
  input \u1_uk_K_r0_reg[33]/NET0131  ;
  input \u1_uk_K_r0_reg[34]/NET0131  ;
  input \u1_uk_K_r0_reg[35]/NET0131  ;
  input \u1_uk_K_r0_reg[36]/NET0131  ;
  input \u1_uk_K_r0_reg[37]/NET0131  ;
  input \u1_uk_K_r0_reg[38]/NET0131  ;
  input \u1_uk_K_r0_reg[39]/NET0131  ;
  input \u1_uk_K_r0_reg[3]/NET0131  ;
  input \u1_uk_K_r0_reg[40]/NET0131  ;
  input \u1_uk_K_r0_reg[41]/NET0131  ;
  input \u1_uk_K_r0_reg[42]/NET0131  ;
  input \u1_uk_K_r0_reg[43]/NET0131  ;
  input \u1_uk_K_r0_reg[44]/NET0131  ;
  input \u1_uk_K_r0_reg[45]/NET0131  ;
  input \u1_uk_K_r0_reg[46]/NET0131  ;
  input \u1_uk_K_r0_reg[47]/NET0131  ;
  input \u1_uk_K_r0_reg[48]/NET0131  ;
  input \u1_uk_K_r0_reg[49]/NET0131  ;
  input \u1_uk_K_r0_reg[4]/NET0131  ;
  input \u1_uk_K_r0_reg[50]/NET0131  ;
  input \u1_uk_K_r0_reg[51]/NET0131  ;
  input \u1_uk_K_r0_reg[52]/P0001  ;
  input \u1_uk_K_r0_reg[54]/NET0131  ;
  input \u1_uk_K_r0_reg[55]/NET0131  ;
  input \u1_uk_K_r0_reg[5]/NET0131  ;
  input \u1_uk_K_r0_reg[6]/NET0131  ;
  input \u1_uk_K_r0_reg[7]/NET0131  ;
  input \u1_uk_K_r0_reg[8]/NET0131  ;
  input \u1_uk_K_r0_reg[9]/NET0131  ;
  input \u1_uk_K_r10_reg[0]/NET0131  ;
  input \u1_uk_K_r10_reg[10]/NET0131  ;
  input \u1_uk_K_r10_reg[11]/NET0131  ;
  input \u1_uk_K_r10_reg[12]/NET0131  ;
  input \u1_uk_K_r10_reg[14]/NET0131  ;
  input \u1_uk_K_r10_reg[15]/NET0131  ;
  input \u1_uk_K_r10_reg[16]/NET0131  ;
  input \u1_uk_K_r10_reg[17]/NET0131  ;
  input \u1_uk_K_r10_reg[18]/NET0131  ;
  input \u1_uk_K_r10_reg[19]/NET0131  ;
  input \u1_uk_K_r10_reg[1]/NET0131  ;
  input \u1_uk_K_r10_reg[20]/NET0131  ;
  input \u1_uk_K_r10_reg[21]/NET0131  ;
  input \u1_uk_K_r10_reg[22]/NET0131  ;
  input \u1_uk_K_r10_reg[23]/NET0131  ;
  input \u1_uk_K_r10_reg[24]/NET0131  ;
  input \u1_uk_K_r10_reg[25]/NET0131  ;
  input \u1_uk_K_r10_reg[26]/NET0131  ;
  input \u1_uk_K_r10_reg[27]/NET0131  ;
  input \u1_uk_K_r10_reg[28]/NET0131  ;
  input \u1_uk_K_r10_reg[29]/NET0131  ;
  input \u1_uk_K_r10_reg[2]/NET0131  ;
  input \u1_uk_K_r10_reg[30]/NET0131  ;
  input \u1_uk_K_r10_reg[31]/NET0131  ;
  input \u1_uk_K_r10_reg[32]/NET0131  ;
  input \u1_uk_K_r10_reg[33]/NET0131  ;
  input \u1_uk_K_r10_reg[34]/NET0131  ;
  input \u1_uk_K_r10_reg[35]/NET0131  ;
  input \u1_uk_K_r10_reg[36]/NET0131  ;
  input \u1_uk_K_r10_reg[37]/NET0131  ;
  input \u1_uk_K_r10_reg[38]/NET0131  ;
  input \u1_uk_K_r10_reg[39]/NET0131  ;
  input \u1_uk_K_r10_reg[3]/NET0131  ;
  input \u1_uk_K_r10_reg[40]/NET0131  ;
  input \u1_uk_K_r10_reg[41]/P0001  ;
  input \u1_uk_K_r10_reg[42]/NET0131  ;
  input \u1_uk_K_r10_reg[43]/NET0131  ;
  input \u1_uk_K_r10_reg[44]/NET0131  ;
  input \u1_uk_K_r10_reg[45]/P0001  ;
  input \u1_uk_K_r10_reg[46]/NET0131  ;
  input \u1_uk_K_r10_reg[47]/NET0131  ;
  input \u1_uk_K_r10_reg[48]/NET0131  ;
  input \u1_uk_K_r10_reg[49]/NET0131  ;
  input \u1_uk_K_r10_reg[4]/NET0131  ;
  input \u1_uk_K_r10_reg[50]/NET0131  ;
  input \u1_uk_K_r10_reg[51]/NET0131  ;
  input \u1_uk_K_r10_reg[52]/NET0131  ;
  input \u1_uk_K_r10_reg[53]/NET0131  ;
  input \u1_uk_K_r10_reg[54]/NET0131  ;
  input \u1_uk_K_r10_reg[55]/NET0131  ;
  input \u1_uk_K_r10_reg[5]/NET0131  ;
  input \u1_uk_K_r10_reg[6]/NET0131  ;
  input \u1_uk_K_r10_reg[7]/NET0131  ;
  input \u1_uk_K_r10_reg[8]/NET0131  ;
  input \u1_uk_K_r10_reg[9]/NET0131  ;
  input \u1_uk_K_r11_reg[0]/NET0131  ;
  input \u1_uk_K_r11_reg[10]/NET0131  ;
  input \u1_uk_K_r11_reg[11]/NET0131  ;
  input \u1_uk_K_r11_reg[12]/NET0131  ;
  input \u1_uk_K_r11_reg[13]/NET0131  ;
  input \u1_uk_K_r11_reg[14]/NET0131  ;
  input \u1_uk_K_r11_reg[15]/NET0131  ;
  input \u1_uk_K_r11_reg[16]/NET0131  ;
  input \u1_uk_K_r11_reg[17]/NET0131  ;
  input \u1_uk_K_r11_reg[18]/NET0131  ;
  input \u1_uk_K_r11_reg[19]/NET0131  ;
  input \u1_uk_K_r11_reg[1]/NET0131  ;
  input \u1_uk_K_r11_reg[20]/NET0131  ;
  input \u1_uk_K_r11_reg[21]/NET0131  ;
  input \u1_uk_K_r11_reg[22]/NET0131  ;
  input \u1_uk_K_r11_reg[23]/NET0131  ;
  input \u1_uk_K_r11_reg[24]/NET0131  ;
  input \u1_uk_K_r11_reg[25]/NET0131  ;
  input \u1_uk_K_r11_reg[26]/NET0131  ;
  input \u1_uk_K_r11_reg[27]/P0001  ;
  input \u1_uk_K_r11_reg[28]/NET0131  ;
  input \u1_uk_K_r11_reg[29]/NET0131  ;
  input \u1_uk_K_r11_reg[2]/NET0131  ;
  input \u1_uk_K_r11_reg[31]/NET0131  ;
  input \u1_uk_K_r11_reg[32]/NET0131  ;
  input \u1_uk_K_r11_reg[33]/NET0131  ;
  input \u1_uk_K_r11_reg[34]/NET0131  ;
  input \u1_uk_K_r11_reg[35]/NET0131  ;
  input \u1_uk_K_r11_reg[36]/NET0131  ;
  input \u1_uk_K_r11_reg[37]/NET0131  ;
  input \u1_uk_K_r11_reg[38]/NET0131  ;
  input \u1_uk_K_r11_reg[39]/NET0131  ;
  input \u1_uk_K_r11_reg[3]/NET0131  ;
  input \u1_uk_K_r11_reg[40]/NET0131  ;
  input \u1_uk_K_r11_reg[41]/NET0131  ;
  input \u1_uk_K_r11_reg[42]/NET0131  ;
  input \u1_uk_K_r11_reg[43]/NET0131  ;
  input \u1_uk_K_r11_reg[44]/NET0131  ;
  input \u1_uk_K_r11_reg[45]/NET0131  ;
  input \u1_uk_K_r11_reg[46]/NET0131  ;
  input \u1_uk_K_r11_reg[47]/NET0131  ;
  input \u1_uk_K_r11_reg[48]/NET0131  ;
  input \u1_uk_K_r11_reg[49]/NET0131  ;
  input \u1_uk_K_r11_reg[4]/NET0131  ;
  input \u1_uk_K_r11_reg[50]/NET0131  ;
  input \u1_uk_K_r11_reg[51]/NET0131  ;
  input \u1_uk_K_r11_reg[52]/NET0131  ;
  input \u1_uk_K_r11_reg[53]/P0001  ;
  input \u1_uk_K_r11_reg[54]/NET0131  ;
  input \u1_uk_K_r11_reg[55]/NET0131  ;
  input \u1_uk_K_r11_reg[5]/NET0131  ;
  input \u1_uk_K_r11_reg[6]/NET0131  ;
  input \u1_uk_K_r11_reg[7]/NET0131  ;
  input \u1_uk_K_r11_reg[8]/NET0131  ;
  input \u1_uk_K_r11_reg[9]/NET0131  ;
  input \u1_uk_K_r12_reg[0]/NET0131  ;
  input \u1_uk_K_r12_reg[10]/P0001  ;
  input \u1_uk_K_r12_reg[11]/NET0131  ;
  input \u1_uk_K_r12_reg[12]/NET0131  ;
  input \u1_uk_K_r12_reg[13]/NET0131  ;
  input \u1_uk_K_r12_reg[14]/NET0131  ;
  input \u1_uk_K_r12_reg[15]/NET0131  ;
  input \u1_uk_K_r12_reg[16]/NET0131  ;
  input \u1_uk_K_r12_reg[17]/NET0131  ;
  input \u1_uk_K_r12_reg[18]/NET0131  ;
  input \u1_uk_K_r12_reg[19]/NET0131  ;
  input \u1_uk_K_r12_reg[1]/NET0131  ;
  input \u1_uk_K_r12_reg[20]/NET0131  ;
  input \u1_uk_K_r12_reg[21]/NET0131  ;
  input \u1_uk_K_r12_reg[22]/NET0131  ;
  input \u1_uk_K_r12_reg[23]/NET0131  ;
  input \u1_uk_K_r12_reg[24]/NET0131  ;
  input \u1_uk_K_r12_reg[25]/NET0131  ;
  input \u1_uk_K_r12_reg[26]/NET0131  ;
  input \u1_uk_K_r12_reg[27]/NET0131  ;
  input \u1_uk_K_r12_reg[28]/NET0131  ;
  input \u1_uk_K_r12_reg[29]/NET0131  ;
  input \u1_uk_K_r12_reg[2]/NET0131  ;
  input \u1_uk_K_r12_reg[30]/NET0131  ;
  input \u1_uk_K_r12_reg[31]/NET0131  ;
  input \u1_uk_K_r12_reg[32]/NET0131  ;
  input \u1_uk_K_r12_reg[33]/NET0131  ;
  input \u1_uk_K_r12_reg[34]/NET0131  ;
  input \u1_uk_K_r12_reg[35]/NET0131  ;
  input \u1_uk_K_r12_reg[36]/NET0131  ;
  input \u1_uk_K_r12_reg[37]/NET0131  ;
  input \u1_uk_K_r12_reg[38]/NET0131  ;
  input \u1_uk_K_r12_reg[3]/NET0131  ;
  input \u1_uk_K_r12_reg[40]/NET0131  ;
  input \u1_uk_K_r12_reg[41]/NET0131  ;
  input \u1_uk_K_r12_reg[42]/NET0131  ;
  input \u1_uk_K_r12_reg[43]/NET0131  ;
  input \u1_uk_K_r12_reg[44]/P0001  ;
  input \u1_uk_K_r12_reg[45]/NET0131  ;
  input \u1_uk_K_r12_reg[46]/NET0131  ;
  input \u1_uk_K_r12_reg[47]/NET0131  ;
  input \u1_uk_K_r12_reg[48]/NET0131  ;
  input \u1_uk_K_r12_reg[49]/NET0131  ;
  input \u1_uk_K_r12_reg[4]/NET0131  ;
  input \u1_uk_K_r12_reg[50]/NET0131  ;
  input \u1_uk_K_r12_reg[51]/NET0131  ;
  input \u1_uk_K_r12_reg[52]/NET0131  ;
  input \u1_uk_K_r12_reg[53]/NET0131  ;
  input \u1_uk_K_r12_reg[54]/NET0131  ;
  input \u1_uk_K_r12_reg[55]/NET0131  ;
  input \u1_uk_K_r12_reg[5]/NET0131  ;
  input \u1_uk_K_r12_reg[6]/NET0131  ;
  input \u1_uk_K_r12_reg[7]/P0001  ;
  input \u1_uk_K_r12_reg[8]/NET0131  ;
  input \u1_uk_K_r12_reg[9]/NET0131  ;
  input \u1_uk_K_r13_reg[0]/NET0131  ;
  input \u1_uk_K_r13_reg[10]/NET0131  ;
  input \u1_uk_K_r13_reg[11]/NET0131  ;
  input \u1_uk_K_r13_reg[12]/NET0131  ;
  input \u1_uk_K_r13_reg[13]/NET0131  ;
  input \u1_uk_K_r13_reg[14]/NET0131  ;
  input \u1_uk_K_r13_reg[15]/NET0131  ;
  input \u1_uk_K_r13_reg[16]/NET0131  ;
  input \u1_uk_K_r13_reg[17]/NET0131  ;
  input \u1_uk_K_r13_reg[18]/NET0131  ;
  input \u1_uk_K_r13_reg[19]/NET0131  ;
  input \u1_uk_K_r13_reg[20]/NET0131  ;
  input \u1_uk_K_r13_reg[21]/NET0131  ;
  input \u1_uk_K_r13_reg[22]/NET0131  ;
  input \u1_uk_K_r13_reg[23]/NET0131  ;
  input \u1_uk_K_r13_reg[24]/NET0131  ;
  input \u1_uk_K_r13_reg[25]/P0001  ;
  input \u1_uk_K_r13_reg[26]/NET0131  ;
  input \u1_uk_K_r13_reg[27]/NET0131  ;
  input \u1_uk_K_r13_reg[28]/NET0131  ;
  input \u1_uk_K_r13_reg[29]/NET0131  ;
  input \u1_uk_K_r13_reg[2]/NET0131  ;
  input \u1_uk_K_r13_reg[30]/NET0131  ;
  input \u1_uk_K_r13_reg[31]/NET0131  ;
  input \u1_uk_K_r13_reg[32]/NET0131  ;
  input \u1_uk_K_r13_reg[33]/NET0131  ;
  input \u1_uk_K_r13_reg[34]/NET0131  ;
  input \u1_uk_K_r13_reg[35]/NET0131  ;
  input \u1_uk_K_r13_reg[36]/NET0131  ;
  input \u1_uk_K_r13_reg[37]/NET0131  ;
  input \u1_uk_K_r13_reg[38]/NET0131  ;
  input \u1_uk_K_r13_reg[39]/NET0131  ;
  input \u1_uk_K_r13_reg[3]/NET0131  ;
  input \u1_uk_K_r13_reg[40]/NET0131  ;
  input \u1_uk_K_r13_reg[41]/NET0131  ;
  input \u1_uk_K_r13_reg[42]/NET0131  ;
  input \u1_uk_K_r13_reg[43]/NET0131  ;
  input \u1_uk_K_r13_reg[44]/NET0131  ;
  input \u1_uk_K_r13_reg[45]/NET0131  ;
  input \u1_uk_K_r13_reg[46]/NET0131  ;
  input \u1_uk_K_r13_reg[47]/NET0131  ;
  input \u1_uk_K_r13_reg[48]/NET0131  ;
  input \u1_uk_K_r13_reg[49]/NET0131  ;
  input \u1_uk_K_r13_reg[4]/NET0131  ;
  input \u1_uk_K_r13_reg[50]/NET0131  ;
  input \u1_uk_K_r13_reg[51]/NET0131  ;
  input \u1_uk_K_r13_reg[52]/P0001  ;
  input \u1_uk_K_r13_reg[54]/NET0131  ;
  input \u1_uk_K_r13_reg[55]/NET0131  ;
  input \u1_uk_K_r13_reg[5]/NET0131  ;
  input \u1_uk_K_r13_reg[6]/NET0131  ;
  input \u1_uk_K_r13_reg[7]/NET0131  ;
  input \u1_uk_K_r13_reg[8]/NET0131  ;
  input \u1_uk_K_r13_reg[9]/NET0131  ;
  input \u1_uk_K_r14_reg[0]/P0001  ;
  input \u1_uk_K_r14_reg[10]/P0001  ;
  input \u1_uk_K_r14_reg[11]/NET0131  ;
  input \u1_uk_K_r14_reg[12]/NET0131  ;
  input \u1_uk_K_r14_reg[13]/NET0131  ;
  input \u1_uk_K_r14_reg[14]/NET0131  ;
  input \u1_uk_K_r14_reg[15]/NET0131  ;
  input \u1_uk_K_r14_reg[16]/NET0131  ;
  input \u1_uk_K_r14_reg[17]/NET0131  ;
  input \u1_uk_K_r14_reg[18]/NET0131  ;
  input \u1_uk_K_r14_reg[19]/NET0131  ;
  input \u1_uk_K_r14_reg[1]/NET0131  ;
  input \u1_uk_K_r14_reg[20]/NET0131  ;
  input \u1_uk_K_r14_reg[21]/NET0131  ;
  input \u1_uk_K_r14_reg[22]/NET0131  ;
  input \u1_uk_K_r14_reg[23]/NET0131  ;
  input \u1_uk_K_r14_reg[24]/NET0131  ;
  input \u1_uk_K_r14_reg[25]/NET0131  ;
  input \u1_uk_K_r14_reg[26]/NET0131  ;
  input \u1_uk_K_r14_reg[27]/NET0131  ;
  input \u1_uk_K_r14_reg[28]/NET0131  ;
  input \u1_uk_K_r14_reg[29]/NET0131  ;
  input \u1_uk_K_r14_reg[2]/NET0131  ;
  input \u1_uk_K_r14_reg[30]/NET0131  ;
  input \u1_uk_K_r14_reg[31]/NET0131  ;
  input \u1_uk_K_r14_reg[32]/NET0131  ;
  input \u1_uk_K_r14_reg[33]/NET0131  ;
  input \u1_uk_K_r14_reg[34]/NET0131  ;
  input \u1_uk_K_r14_reg[35]/P0001  ;
  input \u1_uk_K_r14_reg[36]/NET0131  ;
  input \u1_uk_K_r14_reg[37]/NET0131  ;
  input \u1_uk_K_r14_reg[38]/NET0131  ;
  input \u1_uk_K_r14_reg[39]/P0001  ;
  input \u1_uk_K_r14_reg[3]/NET0131  ;
  input \u1_uk_K_r14_reg[40]/NET0131  ;
  input \u1_uk_K_r14_reg[41]/NET0131  ;
  input \u1_uk_K_r14_reg[42]/P0001  ;
  input \u1_uk_K_r14_reg[43]/NET0131  ;
  input \u1_uk_K_r14_reg[44]/NET0131  ;
  input \u1_uk_K_r14_reg[45]/NET0131  ;
  input \u1_uk_K_r14_reg[46]/NET0131  ;
  input \u1_uk_K_r14_reg[47]/NET0131  ;
  input \u1_uk_K_r14_reg[48]/NET0131  ;
  input \u1_uk_K_r14_reg[49]/NET0131  ;
  input \u1_uk_K_r14_reg[4]/NET0131  ;
  input \u1_uk_K_r14_reg[50]/NET0131  ;
  input \u1_uk_K_r14_reg[51]/NET0131  ;
  input \u1_uk_K_r14_reg[52]/NET0131  ;
  input \u1_uk_K_r14_reg[53]/NET0131  ;
  input \u1_uk_K_r14_reg[54]/NET0131  ;
  input \u1_uk_K_r14_reg[55]/NET0131  ;
  input \u1_uk_K_r14_reg[5]/NET0131  ;
  input \u1_uk_K_r14_reg[6]/NET0131  ;
  input \u1_uk_K_r14_reg[7]/NET0131  ;
  input \u1_uk_K_r14_reg[8]/P0001  ;
  input \u1_uk_K_r14_reg[9]/NET0131  ;
  input \u1_uk_K_r1_reg[0]/NET0131  ;
  input \u1_uk_K_r1_reg[10]/P0001  ;
  input \u1_uk_K_r1_reg[11]/NET0131  ;
  input \u1_uk_K_r1_reg[12]/NET0131  ;
  input \u1_uk_K_r1_reg[13]/NET0131  ;
  input \u1_uk_K_r1_reg[14]/NET0131  ;
  input \u1_uk_K_r1_reg[15]/NET0131  ;
  input \u1_uk_K_r1_reg[16]/NET0131  ;
  input \u1_uk_K_r1_reg[17]/NET0131  ;
  input \u1_uk_K_r1_reg[18]/NET0131  ;
  input \u1_uk_K_r1_reg[19]/NET0131  ;
  input \u1_uk_K_r1_reg[1]/NET0131  ;
  input \u1_uk_K_r1_reg[20]/NET0131  ;
  input \u1_uk_K_r1_reg[21]/NET0131  ;
  input \u1_uk_K_r1_reg[22]/NET0131  ;
  input \u1_uk_K_r1_reg[23]/NET0131  ;
  input \u1_uk_K_r1_reg[24]/NET0131  ;
  input \u1_uk_K_r1_reg[25]/NET0131  ;
  input \u1_uk_K_r1_reg[26]/NET0131  ;
  input \u1_uk_K_r1_reg[27]/NET0131  ;
  input \u1_uk_K_r1_reg[28]/NET0131  ;
  input \u1_uk_K_r1_reg[29]/NET0131  ;
  input \u1_uk_K_r1_reg[2]/NET0131  ;
  input \u1_uk_K_r1_reg[30]/NET0131  ;
  input \u1_uk_K_r1_reg[31]/NET0131  ;
  input \u1_uk_K_r1_reg[32]/NET0131  ;
  input \u1_uk_K_r1_reg[33]/NET0131  ;
  input \u1_uk_K_r1_reg[34]/NET0131  ;
  input \u1_uk_K_r1_reg[35]/NET0131  ;
  input \u1_uk_K_r1_reg[36]/NET0131  ;
  input \u1_uk_K_r1_reg[37]/NET0131  ;
  input \u1_uk_K_r1_reg[38]/NET0131  ;
  input \u1_uk_K_r1_reg[3]/NET0131  ;
  input \u1_uk_K_r1_reg[40]/NET0131  ;
  input \u1_uk_K_r1_reg[41]/NET0131  ;
  input \u1_uk_K_r1_reg[42]/NET0131  ;
  input \u1_uk_K_r1_reg[43]/NET0131  ;
  input \u1_uk_K_r1_reg[44]/P0001  ;
  input \u1_uk_K_r1_reg[45]/NET0131  ;
  input \u1_uk_K_r1_reg[46]/NET0131  ;
  input \u1_uk_K_r1_reg[47]/NET0131  ;
  input \u1_uk_K_r1_reg[48]/NET0131  ;
  input \u1_uk_K_r1_reg[49]/NET0131  ;
  input \u1_uk_K_r1_reg[4]/NET0131  ;
  input \u1_uk_K_r1_reg[50]/NET0131  ;
  input \u1_uk_K_r1_reg[51]/NET0131  ;
  input \u1_uk_K_r1_reg[52]/NET0131  ;
  input \u1_uk_K_r1_reg[53]/NET0131  ;
  input \u1_uk_K_r1_reg[54]/NET0131  ;
  input \u1_uk_K_r1_reg[55]/NET0131  ;
  input \u1_uk_K_r1_reg[5]/NET0131  ;
  input \u1_uk_K_r1_reg[6]/NET0131  ;
  input \u1_uk_K_r1_reg[7]/P0001  ;
  input \u1_uk_K_r1_reg[8]/NET0131  ;
  input \u1_uk_K_r1_reg[9]/NET0131  ;
  input \u1_uk_K_r2_reg[0]/NET0131  ;
  input \u1_uk_K_r2_reg[10]/NET0131  ;
  input \u1_uk_K_r2_reg[11]/NET0131  ;
  input \u1_uk_K_r2_reg[12]/NET0131  ;
  input \u1_uk_K_r2_reg[13]/NET0131  ;
  input \u1_uk_K_r2_reg[14]/NET0131  ;
  input \u1_uk_K_r2_reg[15]/NET0131  ;
  input \u1_uk_K_r2_reg[16]/NET0131  ;
  input \u1_uk_K_r2_reg[17]/NET0131  ;
  input \u1_uk_K_r2_reg[18]/NET0131  ;
  input \u1_uk_K_r2_reg[19]/NET0131  ;
  input \u1_uk_K_r2_reg[1]/NET0131  ;
  input \u1_uk_K_r2_reg[20]/NET0131  ;
  input \u1_uk_K_r2_reg[21]/NET0131  ;
  input \u1_uk_K_r2_reg[22]/NET0131  ;
  input \u1_uk_K_r2_reg[23]/NET0131  ;
  input \u1_uk_K_r2_reg[24]/NET0131  ;
  input \u1_uk_K_r2_reg[25]/NET0131  ;
  input \u1_uk_K_r2_reg[26]/NET0131  ;
  input \u1_uk_K_r2_reg[27]/NET0131  ;
  input \u1_uk_K_r2_reg[28]/NET0131  ;
  input \u1_uk_K_r2_reg[29]/NET0131  ;
  input \u1_uk_K_r2_reg[2]/NET0131  ;
  input \u1_uk_K_r2_reg[31]/NET0131  ;
  input \u1_uk_K_r2_reg[32]/NET0131  ;
  input \u1_uk_K_r2_reg[33]/NET0131  ;
  input \u1_uk_K_r2_reg[34]/NET0131  ;
  input \u1_uk_K_r2_reg[35]/NET0131  ;
  input \u1_uk_K_r2_reg[36]/NET0131  ;
  input \u1_uk_K_r2_reg[37]/NET0131  ;
  input \u1_uk_K_r2_reg[38]/NET0131  ;
  input \u1_uk_K_r2_reg[39]/NET0131  ;
  input \u1_uk_K_r2_reg[3]/NET0131  ;
  input \u1_uk_K_r2_reg[40]/NET0131  ;
  input \u1_uk_K_r2_reg[41]/NET0131  ;
  input \u1_uk_K_r2_reg[42]/NET0131  ;
  input \u1_uk_K_r2_reg[43]/NET0131  ;
  input \u1_uk_K_r2_reg[44]/NET0131  ;
  input \u1_uk_K_r2_reg[45]/NET0131  ;
  input \u1_uk_K_r2_reg[46]/NET0131  ;
  input \u1_uk_K_r2_reg[47]/NET0131  ;
  input \u1_uk_K_r2_reg[48]/NET0131  ;
  input \u1_uk_K_r2_reg[49]/NET0131  ;
  input \u1_uk_K_r2_reg[4]/NET0131  ;
  input \u1_uk_K_r2_reg[50]/NET0131  ;
  input \u1_uk_K_r2_reg[51]/NET0131  ;
  input \u1_uk_K_r2_reg[52]/NET0131  ;
  input \u1_uk_K_r2_reg[53]/P0001  ;
  input \u1_uk_K_r2_reg[54]/NET0131  ;
  input \u1_uk_K_r2_reg[55]/NET0131  ;
  input \u1_uk_K_r2_reg[5]/NET0131  ;
  input \u1_uk_K_r2_reg[6]/NET0131  ;
  input \u1_uk_K_r2_reg[7]/NET0131  ;
  input \u1_uk_K_r2_reg[8]/NET0131  ;
  input \u1_uk_K_r2_reg[9]/NET0131  ;
  input \u1_uk_K_r3_reg[0]/NET0131  ;
  input \u1_uk_K_r3_reg[10]/NET0131  ;
  input \u1_uk_K_r3_reg[11]/NET0131  ;
  input \u1_uk_K_r3_reg[12]/NET0131  ;
  input \u1_uk_K_r3_reg[14]/NET0131  ;
  input \u1_uk_K_r3_reg[15]/NET0131  ;
  input \u1_uk_K_r3_reg[16]/NET0131  ;
  input \u1_uk_K_r3_reg[17]/NET0131  ;
  input \u1_uk_K_r3_reg[18]/NET0131  ;
  input \u1_uk_K_r3_reg[19]/NET0131  ;
  input \u1_uk_K_r3_reg[1]/NET0131  ;
  input \u1_uk_K_r3_reg[20]/NET0131  ;
  input \u1_uk_K_r3_reg[21]/NET0131  ;
  input \u1_uk_K_r3_reg[22]/NET0131  ;
  input \u1_uk_K_r3_reg[23]/NET0131  ;
  input \u1_uk_K_r3_reg[24]/NET0131  ;
  input \u1_uk_K_r3_reg[25]/NET0131  ;
  input \u1_uk_K_r3_reg[26]/NET0131  ;
  input \u1_uk_K_r3_reg[27]/NET0131  ;
  input \u1_uk_K_r3_reg[28]/NET0131  ;
  input \u1_uk_K_r3_reg[29]/NET0131  ;
  input \u1_uk_K_r3_reg[2]/NET0131  ;
  input \u1_uk_K_r3_reg[30]/NET0131  ;
  input \u1_uk_K_r3_reg[31]/NET0131  ;
  input \u1_uk_K_r3_reg[32]/NET0131  ;
  input \u1_uk_K_r3_reg[33]/NET0131  ;
  input \u1_uk_K_r3_reg[34]/NET0131  ;
  input \u1_uk_K_r3_reg[35]/NET0131  ;
  input \u1_uk_K_r3_reg[36]/NET0131  ;
  input \u1_uk_K_r3_reg[37]/NET0131  ;
  input \u1_uk_K_r3_reg[38]/NET0131  ;
  input \u1_uk_K_r3_reg[39]/NET0131  ;
  input \u1_uk_K_r3_reg[3]/NET0131  ;
  input \u1_uk_K_r3_reg[40]/NET0131  ;
  input \u1_uk_K_r3_reg[41]/NET0131  ;
  input \u1_uk_K_r3_reg[42]/NET0131  ;
  input \u1_uk_K_r3_reg[43]/NET0131  ;
  input \u1_uk_K_r3_reg[44]/NET0131  ;
  input \u1_uk_K_r3_reg[45]/NET0131  ;
  input \u1_uk_K_r3_reg[46]/NET0131  ;
  input \u1_uk_K_r3_reg[47]/NET0131  ;
  input \u1_uk_K_r3_reg[48]/NET0131  ;
  input \u1_uk_K_r3_reg[49]/NET0131  ;
  input \u1_uk_K_r3_reg[4]/NET0131  ;
  input \u1_uk_K_r3_reg[50]/NET0131  ;
  input \u1_uk_K_r3_reg[51]/NET0131  ;
  input \u1_uk_K_r3_reg[52]/NET0131  ;
  input \u1_uk_K_r3_reg[53]/NET0131  ;
  input \u1_uk_K_r3_reg[54]/NET0131  ;
  input \u1_uk_K_r3_reg[55]/NET0131  ;
  input \u1_uk_K_r3_reg[5]/NET0131  ;
  input \u1_uk_K_r3_reg[6]/NET0131  ;
  input \u1_uk_K_r3_reg[7]/NET0131  ;
  input \u1_uk_K_r3_reg[8]/NET0131  ;
  input \u1_uk_K_r3_reg[9]/NET0131  ;
  input \u1_uk_K_r4_reg[0]/P0001  ;
  input \u1_uk_K_r4_reg[10]/NET0131  ;
  input \u1_uk_K_r4_reg[11]/NET0131  ;
  input \u1_uk_K_r4_reg[12]/NET0131  ;
  input \u1_uk_K_r4_reg[13]/NET0131  ;
  input \u1_uk_K_r4_reg[14]/NET0131  ;
  input \u1_uk_K_r4_reg[15]/NET0131  ;
  input \u1_uk_K_r4_reg[16]/NET0131  ;
  input \u1_uk_K_r4_reg[17]/NET0131  ;
  input \u1_uk_K_r4_reg[18]/NET0131  ;
  input \u1_uk_K_r4_reg[19]/NET0131  ;
  input \u1_uk_K_r4_reg[1]/NET0131  ;
  input \u1_uk_K_r4_reg[20]/NET0131  ;
  input \u1_uk_K_r4_reg[21]/NET0131  ;
  input \u1_uk_K_r4_reg[22]/NET0131  ;
  input \u1_uk_K_r4_reg[23]/P0001  ;
  input \u1_uk_K_r4_reg[25]/NET0131  ;
  input \u1_uk_K_r4_reg[26]/NET0131  ;
  input \u1_uk_K_r4_reg[27]/P0001  ;
  input \u1_uk_K_r4_reg[28]/NET0131  ;
  input \u1_uk_K_r4_reg[29]/NET0131  ;
  input \u1_uk_K_r4_reg[30]/NET0131  ;
  input \u1_uk_K_r4_reg[31]/P0001  ;
  input \u1_uk_K_r4_reg[32]/NET0131  ;
  input \u1_uk_K_r4_reg[33]/NET0131  ;
  input \u1_uk_K_r4_reg[34]/NET0131  ;
  input \u1_uk_K_r4_reg[35]/NET0131  ;
  input \u1_uk_K_r4_reg[36]/NET0131  ;
  input \u1_uk_K_r4_reg[37]/NET0131  ;
  input \u1_uk_K_r4_reg[38]/NET0131  ;
  input \u1_uk_K_r4_reg[39]/NET0131  ;
  input \u1_uk_K_r4_reg[3]/NET0131  ;
  input \u1_uk_K_r4_reg[40]/NET0131  ;
  input \u1_uk_K_r4_reg[41]/NET0131  ;
  input \u1_uk_K_r4_reg[42]/NET0131  ;
  input \u1_uk_K_r4_reg[43]/NET0131  ;
  input \u1_uk_K_r4_reg[44]/NET0131  ;
  input \u1_uk_K_r4_reg[45]/NET0131  ;
  input \u1_uk_K_r4_reg[46]/NET0131  ;
  input \u1_uk_K_r4_reg[47]/NET0131  ;
  input \u1_uk_K_r4_reg[48]/NET0131  ;
  input \u1_uk_K_r4_reg[49]/NET0131  ;
  input \u1_uk_K_r4_reg[4]/NET0131  ;
  input \u1_uk_K_r4_reg[50]/NET0131  ;
  input \u1_uk_K_r4_reg[51]/NET0131  ;
  input \u1_uk_K_r4_reg[52]/NET0131  ;
  input \u1_uk_K_r4_reg[53]/NET0131  ;
  input \u1_uk_K_r4_reg[54]/NET0131  ;
  input \u1_uk_K_r4_reg[55]/NET0131  ;
  input \u1_uk_K_r4_reg[5]/NET0131  ;
  input \u1_uk_K_r4_reg[6]/NET0131  ;
  input \u1_uk_K_r4_reg[7]/NET0131  ;
  input \u1_uk_K_r4_reg[8]/NET0131  ;
  input \u1_uk_K_r4_reg[9]/NET0131  ;
  input \u1_uk_K_r5_reg[0]/NET0131  ;
  input \u1_uk_K_r5_reg[10]/NET0131  ;
  input \u1_uk_K_r5_reg[11]/NET0131  ;
  input \u1_uk_K_r5_reg[12]/P0001  ;
  input \u1_uk_K_r5_reg[13]/P0001  ;
  input \u1_uk_K_r5_reg[14]/NET0131  ;
  input \u1_uk_K_r5_reg[15]/NET0131  ;
  input \u1_uk_K_r5_reg[16]/NET0131  ;
  input \u1_uk_K_r5_reg[17]/NET0131  ;
  input \u1_uk_K_r5_reg[18]/NET0131  ;
  input \u1_uk_K_r5_reg[19]/NET0131  ;
  input \u1_uk_K_r5_reg[1]/NET0131  ;
  input \u1_uk_K_r5_reg[20]/NET0131  ;
  input \u1_uk_K_r5_reg[21]/NET0131  ;
  input \u1_uk_K_r5_reg[22]/NET0131  ;
  input \u1_uk_K_r5_reg[23]/NET0131  ;
  input \u1_uk_K_r5_reg[24]/NET0131  ;
  input \u1_uk_K_r5_reg[25]/NET0131  ;
  input \u1_uk_K_r5_reg[26]/NET0131  ;
  input \u1_uk_K_r5_reg[27]/NET0131  ;
  input \u1_uk_K_r5_reg[28]/NET0131  ;
  input \u1_uk_K_r5_reg[29]/NET0131  ;
  input \u1_uk_K_r5_reg[2]/NET0131  ;
  input \u1_uk_K_r5_reg[30]/NET0131  ;
  input \u1_uk_K_r5_reg[31]/NET0131  ;
  input \u1_uk_K_r5_reg[32]/NET0131  ;
  input \u1_uk_K_r5_reg[33]/NET0131  ;
  input \u1_uk_K_r5_reg[34]/NET0131  ;
  input \u1_uk_K_r5_reg[35]/NET0131  ;
  input \u1_uk_K_r5_reg[36]/NET0131  ;
  input \u1_uk_K_r5_reg[37]/P0001  ;
  input \u1_uk_K_r5_reg[38]/NET0131  ;
  input \u1_uk_K_r5_reg[39]/NET0131  ;
  input \u1_uk_K_r5_reg[3]/NET0131  ;
  input \u1_uk_K_r5_reg[40]/NET0131  ;
  input \u1_uk_K_r5_reg[41]/NET0131  ;
  input \u1_uk_K_r5_reg[42]/NET0131  ;
  input \u1_uk_K_r5_reg[43]/NET0131  ;
  input \u1_uk_K_r5_reg[44]/NET0131  ;
  input \u1_uk_K_r5_reg[46]/NET0131  ;
  input \u1_uk_K_r5_reg[47]/NET0131  ;
  input \u1_uk_K_r5_reg[48]/NET0131  ;
  input \u1_uk_K_r5_reg[49]/NET0131  ;
  input \u1_uk_K_r5_reg[4]/NET0131  ;
  input \u1_uk_K_r5_reg[50]/NET0131  ;
  input \u1_uk_K_r5_reg[51]/NET0131  ;
  input \u1_uk_K_r5_reg[52]/NET0131  ;
  input \u1_uk_K_r5_reg[53]/NET0131  ;
  input \u1_uk_K_r5_reg[54]/NET0131  ;
  input \u1_uk_K_r5_reg[55]/NET0131  ;
  input \u1_uk_K_r5_reg[5]/NET0131  ;
  input \u1_uk_K_r5_reg[6]/NET0131  ;
  input \u1_uk_K_r5_reg[7]/NET0131  ;
  input \u1_uk_K_r5_reg[8]/NET0131  ;
  input \u1_uk_K_r5_reg[9]/NET0131  ;
  input \u1_uk_K_r6_reg[0]/NET0131  ;
  input \u1_uk_K_r6_reg[10]/NET0131  ;
  input \u1_uk_K_r6_reg[11]/NET0131  ;
  input \u1_uk_K_r6_reg[12]/NET0131  ;
  input \u1_uk_K_r6_reg[13]/NET0131  ;
  input \u1_uk_K_r6_reg[14]/NET0131  ;
  input \u1_uk_K_r6_reg[15]/NET0131  ;
  input \u1_uk_K_r6_reg[16]/NET0131  ;
  input \u1_uk_K_r6_reg[17]/NET0131  ;
  input \u1_uk_K_r6_reg[18]/NET0131  ;
  input \u1_uk_K_r6_reg[19]/NET0131  ;
  input \u1_uk_K_r6_reg[1]/NET0131  ;
  input \u1_uk_K_r6_reg[20]/NET0131  ;
  input \u1_uk_K_r6_reg[21]/NET0131  ;
  input \u1_uk_K_r6_reg[22]/NET0131  ;
  input \u1_uk_K_r6_reg[23]/P0001  ;
  input \u1_uk_K_r6_reg[24]/NET0131  ;
  input \u1_uk_K_r6_reg[25]/NET0131  ;
  input \u1_uk_K_r6_reg[26]/NET0131  ;
  input \u1_uk_K_r6_reg[27]/NET0131  ;
  input \u1_uk_K_r6_reg[28]/NET0131  ;
  input \u1_uk_K_r6_reg[29]/NET0131  ;
  input \u1_uk_K_r6_reg[2]/NET0131  ;
  input \u1_uk_K_r6_reg[30]/P0001  ;
  input \u1_uk_K_r6_reg[31]/NET0131  ;
  input \u1_uk_K_r6_reg[32]/NET0131  ;
  input \u1_uk_K_r6_reg[33]/NET0131  ;
  input \u1_uk_K_r6_reg[34]/NET0131  ;
  input \u1_uk_K_r6_reg[35]/NET0131  ;
  input \u1_uk_K_r6_reg[36]/NET0131  ;
  input \u1_uk_K_r6_reg[37]/NET0131  ;
  input \u1_uk_K_r6_reg[38]/NET0131  ;
  input \u1_uk_K_r6_reg[39]/NET0131  ;
  input \u1_uk_K_r6_reg[3]/NET0131  ;
  input \u1_uk_K_r6_reg[40]/NET0131  ;
  input \u1_uk_K_r6_reg[41]/NET0131  ;
  input \u1_uk_K_r6_reg[42]/NET0131  ;
  input \u1_uk_K_r6_reg[43]/NET0131  ;
  input \u1_uk_K_r6_reg[44]/NET0131  ;
  input \u1_uk_K_r6_reg[45]/NET0131  ;
  input \u1_uk_K_r6_reg[46]/NET0131  ;
  input \u1_uk_K_r6_reg[47]/NET0131  ;
  input \u1_uk_K_r6_reg[48]/NET0131  ;
  input \u1_uk_K_r6_reg[49]/NET0131  ;
  input \u1_uk_K_r6_reg[4]/NET0131  ;
  input \u1_uk_K_r6_reg[50]/NET0131  ;
  input \u1_uk_K_r6_reg[51]/NET0131  ;
  input \u1_uk_K_r6_reg[52]/NET0131  ;
  input \u1_uk_K_r6_reg[53]/NET0131  ;
  input \u1_uk_K_r6_reg[54]/NET0131  ;
  input \u1_uk_K_r6_reg[55]/P0001  ;
  input \u1_uk_K_r6_reg[5]/NET0131  ;
  input \u1_uk_K_r6_reg[6]/NET0131  ;
  input \u1_uk_K_r6_reg[7]/NET0131  ;
  input \u1_uk_K_r6_reg[8]/NET0131  ;
  input \u1_uk_K_r6_reg[9]/NET0131  ;
  input \u1_uk_K_r7_reg[0]/NET0131  ;
  input \u1_uk_K_r7_reg[10]/NET0131  ;
  input \u1_uk_K_r7_reg[11]/NET0131  ;
  input \u1_uk_K_r7_reg[12]/NET0131  ;
  input \u1_uk_K_r7_reg[13]/NET0131  ;
  input \u1_uk_K_r7_reg[14]/NET0131  ;
  input \u1_uk_K_r7_reg[15]/NET0131  ;
  input \u1_uk_K_r7_reg[16]/NET0131  ;
  input \u1_uk_K_r7_reg[17]/NET0131  ;
  input \u1_uk_K_r7_reg[18]/NET0131  ;
  input \u1_uk_K_r7_reg[19]/NET0131  ;
  input \u1_uk_K_r7_reg[1]/NET0131  ;
  input \u1_uk_K_r7_reg[20]/NET0131  ;
  input \u1_uk_K_r7_reg[21]/NET0131  ;
  input \u1_uk_K_r7_reg[22]/NET0131  ;
  input \u1_uk_K_r7_reg[23]/P0001  ;
  input \u1_uk_K_r7_reg[24]/NET0131  ;
  input \u1_uk_K_r7_reg[25]/NET0131  ;
  input \u1_uk_K_r7_reg[26]/P0001  ;
  input \u1_uk_K_r7_reg[27]/NET0131  ;
  input \u1_uk_K_r7_reg[28]/NET0131  ;
  input \u1_uk_K_r7_reg[29]/NET0131  ;
  input \u1_uk_K_r7_reg[2]/NET0131  ;
  input \u1_uk_K_r7_reg[30]/P0001  ;
  input \u1_uk_K_r7_reg[31]/NET0131  ;
  input \u1_uk_K_r7_reg[32]/NET0131  ;
  input \u1_uk_K_r7_reg[33]/NET0131  ;
  input \u1_uk_K_r7_reg[34]/NET0131  ;
  input \u1_uk_K_r7_reg[35]/NET0131  ;
  input \u1_uk_K_r7_reg[36]/NET0131  ;
  input \u1_uk_K_r7_reg[37]/NET0131  ;
  input \u1_uk_K_r7_reg[38]/NET0131  ;
  input \u1_uk_K_r7_reg[39]/NET0131  ;
  input \u1_uk_K_r7_reg[3]/NET0131  ;
  input \u1_uk_K_r7_reg[40]/NET0131  ;
  input \u1_uk_K_r7_reg[41]/NET0131  ;
  input \u1_uk_K_r7_reg[42]/NET0131  ;
  input \u1_uk_K_r7_reg[43]/NET0131  ;
  input \u1_uk_K_r7_reg[44]/NET0131  ;
  input \u1_uk_K_r7_reg[45]/NET0131  ;
  input \u1_uk_K_r7_reg[46]/NET0131  ;
  input \u1_uk_K_r7_reg[47]/NET0131  ;
  input \u1_uk_K_r7_reg[48]/NET0131  ;
  input \u1_uk_K_r7_reg[49]/NET0131  ;
  input \u1_uk_K_r7_reg[4]/NET0131  ;
  input \u1_uk_K_r7_reg[50]/NET0131  ;
  input \u1_uk_K_r7_reg[51]/NET0131  ;
  input \u1_uk_K_r7_reg[52]/NET0131  ;
  input \u1_uk_K_r7_reg[53]/NET0131  ;
  input \u1_uk_K_r7_reg[54]/NET0131  ;
  input \u1_uk_K_r7_reg[55]/P0001  ;
  input \u1_uk_K_r7_reg[5]/NET0131  ;
  input \u1_uk_K_r7_reg[6]/NET0131  ;
  input \u1_uk_K_r7_reg[7]/NET0131  ;
  input \u1_uk_K_r7_reg[8]/NET0131  ;
  input \u1_uk_K_r7_reg[9]/NET0131  ;
  input \u1_uk_K_r8_reg[0]/NET0131  ;
  input \u1_uk_K_r8_reg[10]/NET0131  ;
  input \u1_uk_K_r8_reg[11]/NET0131  ;
  input \u1_uk_K_r8_reg[12]/NET0131  ;
  input \u1_uk_K_r8_reg[13]/P0001  ;
  input \u1_uk_K_r8_reg[14]/NET0131  ;
  input \u1_uk_K_r8_reg[15]/NET0131  ;
  input \u1_uk_K_r8_reg[16]/NET0131  ;
  input \u1_uk_K_r8_reg[17]/NET0131  ;
  input \u1_uk_K_r8_reg[18]/NET0131  ;
  input \u1_uk_K_r8_reg[19]/NET0131  ;
  input \u1_uk_K_r8_reg[1]/NET0131  ;
  input \u1_uk_K_r8_reg[20]/NET0131  ;
  input \u1_uk_K_r8_reg[21]/NET0131  ;
  input \u1_uk_K_r8_reg[22]/NET0131  ;
  input \u1_uk_K_r8_reg[23]/NET0131  ;
  input \u1_uk_K_r8_reg[24]/NET0131  ;
  input \u1_uk_K_r8_reg[25]/NET0131  ;
  input \u1_uk_K_r8_reg[26]/NET0131  ;
  input \u1_uk_K_r8_reg[27]/NET0131  ;
  input \u1_uk_K_r8_reg[28]/NET0131  ;
  input \u1_uk_K_r8_reg[29]/NET0131  ;
  input \u1_uk_K_r8_reg[2]/NET0131  ;
  input \u1_uk_K_r8_reg[30]/NET0131  ;
  input \u1_uk_K_r8_reg[31]/NET0131  ;
  input \u1_uk_K_r8_reg[32]/NET0131  ;
  input \u1_uk_K_r8_reg[33]/NET0131  ;
  input \u1_uk_K_r8_reg[34]/NET0131  ;
  input \u1_uk_K_r8_reg[35]/NET0131  ;
  input \u1_uk_K_r8_reg[36]/NET0131  ;
  input \u1_uk_K_r8_reg[37]/P0001  ;
  input \u1_uk_K_r8_reg[38]/NET0131  ;
  input \u1_uk_K_r8_reg[39]/NET0131  ;
  input \u1_uk_K_r8_reg[3]/NET0131  ;
  input \u1_uk_K_r8_reg[40]/NET0131  ;
  input \u1_uk_K_r8_reg[41]/NET0131  ;
  input \u1_uk_K_r8_reg[42]/NET0131  ;
  input \u1_uk_K_r8_reg[43]/NET0131  ;
  input \u1_uk_K_r8_reg[44]/NET0131  ;
  input \u1_uk_K_r8_reg[46]/NET0131  ;
  input \u1_uk_K_r8_reg[47]/NET0131  ;
  input \u1_uk_K_r8_reg[48]/NET0131  ;
  input \u1_uk_K_r8_reg[49]/NET0131  ;
  input \u1_uk_K_r8_reg[4]/NET0131  ;
  input \u1_uk_K_r8_reg[50]/NET0131  ;
  input \u1_uk_K_r8_reg[51]/NET0131  ;
  input \u1_uk_K_r8_reg[52]/NET0131  ;
  input \u1_uk_K_r8_reg[53]/NET0131  ;
  input \u1_uk_K_r8_reg[54]/NET0131  ;
  input \u1_uk_K_r8_reg[55]/NET0131  ;
  input \u1_uk_K_r8_reg[5]/NET0131  ;
  input \u1_uk_K_r8_reg[6]/NET0131  ;
  input \u1_uk_K_r8_reg[7]/NET0131  ;
  input \u1_uk_K_r8_reg[8]/NET0131  ;
  input \u1_uk_K_r8_reg[9]/NET0131  ;
  input \u1_uk_K_r9_reg[0]/P0001  ;
  input \u1_uk_K_r9_reg[10]/NET0131  ;
  input \u1_uk_K_r9_reg[11]/NET0131  ;
  input \u1_uk_K_r9_reg[12]/NET0131  ;
  input \u1_uk_K_r9_reg[13]/NET0131  ;
  input \u1_uk_K_r9_reg[14]/NET0131  ;
  input \u1_uk_K_r9_reg[15]/NET0131  ;
  input \u1_uk_K_r9_reg[16]/NET0131  ;
  input \u1_uk_K_r9_reg[17]/NET0131  ;
  input \u1_uk_K_r9_reg[18]/NET0131  ;
  input \u1_uk_K_r9_reg[19]/NET0131  ;
  input \u1_uk_K_r9_reg[1]/NET0131  ;
  input \u1_uk_K_r9_reg[20]/NET0131  ;
  input \u1_uk_K_r9_reg[21]/NET0131  ;
  input \u1_uk_K_r9_reg[22]/NET0131  ;
  input \u1_uk_K_r9_reg[23]/NET0131  ;
  input \u1_uk_K_r9_reg[25]/NET0131  ;
  input \u1_uk_K_r9_reg[26]/NET0131  ;
  input \u1_uk_K_r9_reg[27]/P0001  ;
  input \u1_uk_K_r9_reg[28]/NET0131  ;
  input \u1_uk_K_r9_reg[29]/NET0131  ;
  input \u1_uk_K_r9_reg[30]/NET0131  ;
  input \u1_uk_K_r9_reg[31]/P0001  ;
  input \u1_uk_K_r9_reg[32]/NET0131  ;
  input \u1_uk_K_r9_reg[33]/NET0131  ;
  input \u1_uk_K_r9_reg[34]/NET0131  ;
  input \u1_uk_K_r9_reg[35]/NET0131  ;
  input \u1_uk_K_r9_reg[36]/NET0131  ;
  input \u1_uk_K_r9_reg[37]/NET0131  ;
  input \u1_uk_K_r9_reg[38]/NET0131  ;
  input \u1_uk_K_r9_reg[39]/NET0131  ;
  input \u1_uk_K_r9_reg[3]/NET0131  ;
  input \u1_uk_K_r9_reg[40]/NET0131  ;
  input \u1_uk_K_r9_reg[41]/NET0131  ;
  input \u1_uk_K_r9_reg[42]/NET0131  ;
  input \u1_uk_K_r9_reg[43]/NET0131  ;
  input \u1_uk_K_r9_reg[44]/NET0131  ;
  input \u1_uk_K_r9_reg[45]/NET0131  ;
  input \u1_uk_K_r9_reg[46]/NET0131  ;
  input \u1_uk_K_r9_reg[47]/NET0131  ;
  input \u1_uk_K_r9_reg[48]/NET0131  ;
  input \u1_uk_K_r9_reg[49]/NET0131  ;
  input \u1_uk_K_r9_reg[4]/NET0131  ;
  input \u1_uk_K_r9_reg[50]/NET0131  ;
  input \u1_uk_K_r9_reg[51]/NET0131  ;
  input \u1_uk_K_r9_reg[52]/NET0131  ;
  input \u1_uk_K_r9_reg[53]/NET0131  ;
  input \u1_uk_K_r9_reg[54]/NET0131  ;
  input \u1_uk_K_r9_reg[55]/NET0131  ;
  input \u1_uk_K_r9_reg[5]/NET0131  ;
  input \u1_uk_K_r9_reg[6]/NET0131  ;
  input \u1_uk_K_r9_reg[7]/NET0131  ;
  input \u1_uk_K_r9_reg[8]/NET0131  ;
  input \u1_uk_K_r9_reg[9]/NET0131  ;
  input \u2_L0_reg[10]/NET0131  ;
  input \u2_L0_reg[11]/NET0131  ;
  input \u2_L0_reg[12]/NET0131  ;
  input \u2_L0_reg[13]/NET0131  ;
  input \u2_L0_reg[14]/NET0131  ;
  input \u2_L0_reg[15]/NET0131  ;
  input \u2_L0_reg[16]/NET0131  ;
  input \u2_L0_reg[17]/NET0131  ;
  input \u2_L0_reg[18]/P0001  ;
  input \u2_L0_reg[19]/NET0131  ;
  input \u2_L0_reg[1]/NET0131  ;
  input \u2_L0_reg[20]/NET0131  ;
  input \u2_L0_reg[21]/NET0131  ;
  input \u2_L0_reg[22]/NET0131  ;
  input \u2_L0_reg[23]/NET0131  ;
  input \u2_L0_reg[24]/NET0131  ;
  input \u2_L0_reg[25]/NET0131  ;
  input \u2_L0_reg[26]/NET0131  ;
  input \u2_L0_reg[27]/NET0131  ;
  input \u2_L0_reg[28]/NET0131  ;
  input \u2_L0_reg[29]/NET0131  ;
  input \u2_L0_reg[2]/NET0131  ;
  input \u2_L0_reg[30]/NET0131  ;
  input \u2_L0_reg[31]/NET0131  ;
  input \u2_L0_reg[32]/NET0131  ;
  input \u2_L0_reg[3]/NET0131  ;
  input \u2_L0_reg[4]/NET0131  ;
  input \u2_L0_reg[5]/NET0131  ;
  input \u2_L0_reg[6]/NET0131  ;
  input \u2_L0_reg[7]/NET0131  ;
  input \u2_L0_reg[8]/NET0131  ;
  input \u2_L0_reg[9]/NET0131  ;
  input \u2_L10_reg[10]/NET0131  ;
  input \u2_L10_reg[11]/NET0131  ;
  input \u2_L10_reg[12]/NET0131  ;
  input \u2_L10_reg[13]/NET0131  ;
  input \u2_L10_reg[14]/NET0131  ;
  input \u2_L10_reg[15]/NET0131  ;
  input \u2_L10_reg[16]/NET0131  ;
  input \u2_L10_reg[17]/NET0131  ;
  input \u2_L10_reg[18]/P0001  ;
  input \u2_L10_reg[19]/NET0131  ;
  input \u2_L10_reg[1]/NET0131  ;
  input \u2_L10_reg[20]/NET0131  ;
  input \u2_L10_reg[21]/NET0131  ;
  input \u2_L10_reg[22]/NET0131  ;
  input \u2_L10_reg[23]/NET0131  ;
  input \u2_L10_reg[24]/NET0131  ;
  input \u2_L10_reg[25]/NET0131  ;
  input \u2_L10_reg[26]/NET0131  ;
  input \u2_L10_reg[27]/NET0131  ;
  input \u2_L10_reg[28]/NET0131  ;
  input \u2_L10_reg[29]/NET0131  ;
  input \u2_L10_reg[2]/NET0131  ;
  input \u2_L10_reg[30]/NET0131  ;
  input \u2_L10_reg[31]/NET0131  ;
  input \u2_L10_reg[32]/NET0131  ;
  input \u2_L10_reg[3]/NET0131  ;
  input \u2_L10_reg[4]/NET0131  ;
  input \u2_L10_reg[5]/NET0131  ;
  input \u2_L10_reg[6]/NET0131  ;
  input \u2_L10_reg[7]/NET0131  ;
  input \u2_L10_reg[8]/NET0131  ;
  input \u2_L10_reg[9]/NET0131  ;
  input \u2_L11_reg[10]/NET0131  ;
  input \u2_L11_reg[11]/NET0131  ;
  input \u2_L11_reg[12]/NET0131  ;
  input \u2_L11_reg[13]/NET0131  ;
  input \u2_L11_reg[14]/NET0131  ;
  input \u2_L11_reg[15]/NET0131  ;
  input \u2_L11_reg[16]/NET0131  ;
  input \u2_L11_reg[17]/NET0131  ;
  input \u2_L11_reg[18]/P0001  ;
  input \u2_L11_reg[19]/NET0131  ;
  input \u2_L11_reg[1]/NET0131  ;
  input \u2_L11_reg[20]/NET0131  ;
  input \u2_L11_reg[21]/NET0131  ;
  input \u2_L11_reg[22]/NET0131  ;
  input \u2_L11_reg[23]/NET0131  ;
  input \u2_L11_reg[24]/NET0131  ;
  input \u2_L11_reg[25]/NET0131  ;
  input \u2_L11_reg[26]/NET0131  ;
  input \u2_L11_reg[27]/NET0131  ;
  input \u2_L11_reg[28]/NET0131  ;
  input \u2_L11_reg[29]/NET0131  ;
  input \u2_L11_reg[2]/NET0131  ;
  input \u2_L11_reg[30]/NET0131  ;
  input \u2_L11_reg[31]/NET0131  ;
  input \u2_L11_reg[32]/NET0131  ;
  input \u2_L11_reg[3]/NET0131  ;
  input \u2_L11_reg[4]/NET0131  ;
  input \u2_L11_reg[5]/NET0131  ;
  input \u2_L11_reg[6]/NET0131  ;
  input \u2_L11_reg[7]/NET0131  ;
  input \u2_L11_reg[8]/NET0131  ;
  input \u2_L11_reg[9]/NET0131  ;
  input \u2_L12_reg[10]/NET0131  ;
  input \u2_L12_reg[11]/NET0131  ;
  input \u2_L12_reg[12]/NET0131  ;
  input \u2_L12_reg[13]/NET0131  ;
  input \u2_L12_reg[14]/NET0131  ;
  input \u2_L12_reg[15]/NET0131  ;
  input \u2_L12_reg[16]/NET0131  ;
  input \u2_L12_reg[17]/NET0131  ;
  input \u2_L12_reg[18]/P0001  ;
  input \u2_L12_reg[19]/NET0131  ;
  input \u2_L12_reg[1]/NET0131  ;
  input \u2_L12_reg[20]/NET0131  ;
  input \u2_L12_reg[21]/NET0131  ;
  input \u2_L12_reg[22]/NET0131  ;
  input \u2_L12_reg[23]/NET0131  ;
  input \u2_L12_reg[24]/NET0131  ;
  input \u2_L12_reg[25]/NET0131  ;
  input \u2_L12_reg[26]/NET0131  ;
  input \u2_L12_reg[27]/NET0131  ;
  input \u2_L12_reg[28]/NET0131  ;
  input \u2_L12_reg[29]/NET0131  ;
  input \u2_L12_reg[2]/NET0131  ;
  input \u2_L12_reg[30]/NET0131  ;
  input \u2_L12_reg[31]/NET0131  ;
  input \u2_L12_reg[32]/NET0131  ;
  input \u2_L12_reg[3]/NET0131  ;
  input \u2_L12_reg[4]/NET0131  ;
  input \u2_L12_reg[5]/NET0131  ;
  input \u2_L12_reg[6]/NET0131  ;
  input \u2_L12_reg[7]/NET0131  ;
  input \u2_L12_reg[8]/NET0131  ;
  input \u2_L12_reg[9]/NET0131  ;
  input \u2_L13_reg[10]/NET0131  ;
  input \u2_L13_reg[11]/NET0131  ;
  input \u2_L13_reg[12]/NET0131  ;
  input \u2_L13_reg[13]/NET0131  ;
  input \u2_L13_reg[14]/NET0131  ;
  input \u2_L13_reg[15]/NET0131  ;
  input \u2_L13_reg[16]/NET0131  ;
  input \u2_L13_reg[17]/NET0131  ;
  input \u2_L13_reg[18]/P0001  ;
  input \u2_L13_reg[19]/P0001  ;
  input \u2_L13_reg[1]/NET0131  ;
  input \u2_L13_reg[20]/NET0131  ;
  input \u2_L13_reg[21]/NET0131  ;
  input \u2_L13_reg[22]/NET0131  ;
  input \u2_L13_reg[23]/P0001  ;
  input \u2_L13_reg[24]/NET0131  ;
  input \u2_L13_reg[25]/NET0131  ;
  input \u2_L13_reg[26]/NET0131  ;
  input \u2_L13_reg[27]/NET0131  ;
  input \u2_L13_reg[28]/NET0131  ;
  input \u2_L13_reg[29]/NET0131  ;
  input \u2_L13_reg[2]/NET0131  ;
  input \u2_L13_reg[30]/NET0131  ;
  input \u2_L13_reg[31]/NET0131  ;
  input \u2_L13_reg[32]/NET0131  ;
  input \u2_L13_reg[3]/NET0131  ;
  input \u2_L13_reg[4]/NET0131  ;
  input \u2_L13_reg[5]/NET0131  ;
  input \u2_L13_reg[6]/NET0131  ;
  input \u2_L13_reg[7]/NET0131  ;
  input \u2_L13_reg[8]/NET0131  ;
  input \u2_L13_reg[9]/NET0131  ;
  input \u2_L14_reg[10]/P0001  ;
  input \u2_L14_reg[11]/P0001  ;
  input \u2_L14_reg[12]/P0001  ;
  input \u2_L14_reg[13]/P0001  ;
  input \u2_L14_reg[14]/P0001  ;
  input \u2_L14_reg[15]/P0001  ;
  input \u2_L14_reg[16]/P0001  ;
  input \u2_L14_reg[17]/P0001  ;
  input \u2_L14_reg[18]/P0001  ;
  input \u2_L14_reg[19]/P0001  ;
  input \u2_L14_reg[1]/P0001  ;
  input \u2_L14_reg[20]/P0001  ;
  input \u2_L14_reg[21]/P0001  ;
  input \u2_L14_reg[22]/P0001  ;
  input \u2_L14_reg[23]/P0001  ;
  input \u2_L14_reg[24]/P0001  ;
  input \u2_L14_reg[25]/P0001  ;
  input \u2_L14_reg[26]/P0001  ;
  input \u2_L14_reg[27]/P0001  ;
  input \u2_L14_reg[28]/P0001  ;
  input \u2_L14_reg[29]/P0001  ;
  input \u2_L14_reg[2]/P0001  ;
  input \u2_L14_reg[30]/P0001  ;
  input \u2_L14_reg[31]/P0001  ;
  input \u2_L14_reg[32]/P0001  ;
  input \u2_L14_reg[3]/P0001  ;
  input \u2_L14_reg[4]/P0001  ;
  input \u2_L14_reg[5]/P0001  ;
  input \u2_L14_reg[6]/P0001  ;
  input \u2_L14_reg[7]/P0001  ;
  input \u2_L14_reg[8]/P0001  ;
  input \u2_L14_reg[9]/P0001  ;
  input \u2_L1_reg[10]/NET0131  ;
  input \u2_L1_reg[11]/NET0131  ;
  input \u2_L1_reg[12]/NET0131  ;
  input \u2_L1_reg[13]/NET0131  ;
  input \u2_L1_reg[14]/NET0131  ;
  input \u2_L1_reg[15]/NET0131  ;
  input \u2_L1_reg[16]/NET0131  ;
  input \u2_L1_reg[17]/NET0131  ;
  input \u2_L1_reg[18]/P0001  ;
  input \u2_L1_reg[19]/NET0131  ;
  input \u2_L1_reg[1]/NET0131  ;
  input \u2_L1_reg[20]/NET0131  ;
  input \u2_L1_reg[21]/NET0131  ;
  input \u2_L1_reg[22]/NET0131  ;
  input \u2_L1_reg[23]/NET0131  ;
  input \u2_L1_reg[24]/NET0131  ;
  input \u2_L1_reg[25]/NET0131  ;
  input \u2_L1_reg[26]/NET0131  ;
  input \u2_L1_reg[27]/NET0131  ;
  input \u2_L1_reg[28]/NET0131  ;
  input \u2_L1_reg[29]/NET0131  ;
  input \u2_L1_reg[2]/NET0131  ;
  input \u2_L1_reg[30]/NET0131  ;
  input \u2_L1_reg[31]/NET0131  ;
  input \u2_L1_reg[32]/NET0131  ;
  input \u2_L1_reg[3]/NET0131  ;
  input \u2_L1_reg[4]/NET0131  ;
  input \u2_L1_reg[5]/NET0131  ;
  input \u2_L1_reg[6]/NET0131  ;
  input \u2_L1_reg[7]/NET0131  ;
  input \u2_L1_reg[8]/NET0131  ;
  input \u2_L1_reg[9]/NET0131  ;
  input \u2_L2_reg[10]/NET0131  ;
  input \u2_L2_reg[11]/NET0131  ;
  input \u2_L2_reg[12]/NET0131  ;
  input \u2_L2_reg[13]/NET0131  ;
  input \u2_L2_reg[14]/NET0131  ;
  input \u2_L2_reg[15]/NET0131  ;
  input \u2_L2_reg[16]/NET0131  ;
  input \u2_L2_reg[17]/NET0131  ;
  input \u2_L2_reg[18]/P0001  ;
  input \u2_L2_reg[19]/NET0131  ;
  input \u2_L2_reg[1]/NET0131  ;
  input \u2_L2_reg[20]/NET0131  ;
  input \u2_L2_reg[21]/NET0131  ;
  input \u2_L2_reg[22]/NET0131  ;
  input \u2_L2_reg[23]/NET0131  ;
  input \u2_L2_reg[24]/NET0131  ;
  input \u2_L2_reg[25]/NET0131  ;
  input \u2_L2_reg[26]/NET0131  ;
  input \u2_L2_reg[27]/NET0131  ;
  input \u2_L2_reg[28]/NET0131  ;
  input \u2_L2_reg[29]/NET0131  ;
  input \u2_L2_reg[2]/NET0131  ;
  input \u2_L2_reg[30]/NET0131  ;
  input \u2_L2_reg[31]/NET0131  ;
  input \u2_L2_reg[32]/NET0131  ;
  input \u2_L2_reg[3]/NET0131  ;
  input \u2_L2_reg[4]/NET0131  ;
  input \u2_L2_reg[5]/NET0131  ;
  input \u2_L2_reg[6]/NET0131  ;
  input \u2_L2_reg[7]/NET0131  ;
  input \u2_L2_reg[8]/NET0131  ;
  input \u2_L2_reg[9]/NET0131  ;
  input \u2_L3_reg[10]/NET0131  ;
  input \u2_L3_reg[11]/NET0131  ;
  input \u2_L3_reg[12]/NET0131  ;
  input \u2_L3_reg[13]/NET0131  ;
  input \u2_L3_reg[14]/NET0131  ;
  input \u2_L3_reg[15]/NET0131  ;
  input \u2_L3_reg[16]/NET0131  ;
  input \u2_L3_reg[17]/NET0131  ;
  input \u2_L3_reg[18]/P0001  ;
  input \u2_L3_reg[19]/NET0131  ;
  input \u2_L3_reg[1]/NET0131  ;
  input \u2_L3_reg[20]/NET0131  ;
  input \u2_L3_reg[21]/NET0131  ;
  input \u2_L3_reg[22]/NET0131  ;
  input \u2_L3_reg[23]/NET0131  ;
  input \u2_L3_reg[24]/NET0131  ;
  input \u2_L3_reg[25]/NET0131  ;
  input \u2_L3_reg[26]/NET0131  ;
  input \u2_L3_reg[27]/NET0131  ;
  input \u2_L3_reg[28]/NET0131  ;
  input \u2_L3_reg[29]/NET0131  ;
  input \u2_L3_reg[2]/NET0131  ;
  input \u2_L3_reg[30]/NET0131  ;
  input \u2_L3_reg[31]/NET0131  ;
  input \u2_L3_reg[32]/NET0131  ;
  input \u2_L3_reg[3]/NET0131  ;
  input \u2_L3_reg[4]/NET0131  ;
  input \u2_L3_reg[5]/NET0131  ;
  input \u2_L3_reg[6]/NET0131  ;
  input \u2_L3_reg[7]/NET0131  ;
  input \u2_L3_reg[8]/NET0131  ;
  input \u2_L3_reg[9]/NET0131  ;
  input \u2_L4_reg[10]/NET0131  ;
  input \u2_L4_reg[11]/NET0131  ;
  input \u2_L4_reg[12]/NET0131  ;
  input \u2_L4_reg[13]/NET0131  ;
  input \u2_L4_reg[14]/NET0131  ;
  input \u2_L4_reg[15]/NET0131  ;
  input \u2_L4_reg[16]/NET0131  ;
  input \u2_L4_reg[17]/NET0131  ;
  input \u2_L4_reg[18]/P0001  ;
  input \u2_L4_reg[19]/NET0131  ;
  input \u2_L4_reg[1]/NET0131  ;
  input \u2_L4_reg[20]/NET0131  ;
  input \u2_L4_reg[21]/NET0131  ;
  input \u2_L4_reg[22]/NET0131  ;
  input \u2_L4_reg[23]/NET0131  ;
  input \u2_L4_reg[24]/NET0131  ;
  input \u2_L4_reg[25]/NET0131  ;
  input \u2_L4_reg[26]/NET0131  ;
  input \u2_L4_reg[27]/NET0131  ;
  input \u2_L4_reg[28]/NET0131  ;
  input \u2_L4_reg[29]/NET0131  ;
  input \u2_L4_reg[2]/NET0131  ;
  input \u2_L4_reg[30]/NET0131  ;
  input \u2_L4_reg[31]/NET0131  ;
  input \u2_L4_reg[32]/NET0131  ;
  input \u2_L4_reg[3]/NET0131  ;
  input \u2_L4_reg[4]/NET0131  ;
  input \u2_L4_reg[5]/NET0131  ;
  input \u2_L4_reg[6]/NET0131  ;
  input \u2_L4_reg[7]/NET0131  ;
  input \u2_L4_reg[8]/NET0131  ;
  input \u2_L4_reg[9]/NET0131  ;
  input \u2_L5_reg[10]/NET0131  ;
  input \u2_L5_reg[11]/NET0131  ;
  input \u2_L5_reg[12]/NET0131  ;
  input \u2_L5_reg[13]/NET0131  ;
  input \u2_L5_reg[14]/NET0131  ;
  input \u2_L5_reg[15]/NET0131  ;
  input \u2_L5_reg[16]/NET0131  ;
  input \u2_L5_reg[17]/NET0131  ;
  input \u2_L5_reg[18]/NET0131  ;
  input \u2_L5_reg[19]/NET0131  ;
  input \u2_L5_reg[1]/NET0131  ;
  input \u2_L5_reg[20]/NET0131  ;
  input \u2_L5_reg[21]/NET0131  ;
  input \u2_L5_reg[22]/NET0131  ;
  input \u2_L5_reg[23]/NET0131  ;
  input \u2_L5_reg[24]/NET0131  ;
  input \u2_L5_reg[25]/NET0131  ;
  input \u2_L5_reg[26]/NET0131  ;
  input \u2_L5_reg[27]/NET0131  ;
  input \u2_L5_reg[28]/NET0131  ;
  input \u2_L5_reg[29]/NET0131  ;
  input \u2_L5_reg[2]/NET0131  ;
  input \u2_L5_reg[30]/NET0131  ;
  input \u2_L5_reg[31]/NET0131  ;
  input \u2_L5_reg[32]/NET0131  ;
  input \u2_L5_reg[3]/NET0131  ;
  input \u2_L5_reg[4]/NET0131  ;
  input \u2_L5_reg[5]/NET0131  ;
  input \u2_L5_reg[6]/NET0131  ;
  input \u2_L5_reg[7]/NET0131  ;
  input \u2_L5_reg[8]/NET0131  ;
  input \u2_L5_reg[9]/NET0131  ;
  input \u2_L6_reg[10]/NET0131  ;
  input \u2_L6_reg[11]/NET0131  ;
  input \u2_L6_reg[12]/NET0131  ;
  input \u2_L6_reg[13]/NET0131  ;
  input \u2_L6_reg[14]/NET0131  ;
  input \u2_L6_reg[15]/NET0131  ;
  input \u2_L6_reg[16]/NET0131  ;
  input \u2_L6_reg[17]/NET0131  ;
  input \u2_L6_reg[18]/P0001  ;
  input \u2_L6_reg[19]/NET0131  ;
  input \u2_L6_reg[1]/NET0131  ;
  input \u2_L6_reg[20]/NET0131  ;
  input \u2_L6_reg[21]/NET0131  ;
  input \u2_L6_reg[22]/NET0131  ;
  input \u2_L6_reg[23]/NET0131  ;
  input \u2_L6_reg[24]/NET0131  ;
  input \u2_L6_reg[25]/NET0131  ;
  input \u2_L6_reg[26]/NET0131  ;
  input \u2_L6_reg[27]/NET0131  ;
  input \u2_L6_reg[28]/NET0131  ;
  input \u2_L6_reg[29]/NET0131  ;
  input \u2_L6_reg[2]/NET0131  ;
  input \u2_L6_reg[30]/NET0131  ;
  input \u2_L6_reg[31]/NET0131  ;
  input \u2_L6_reg[32]/NET0131  ;
  input \u2_L6_reg[3]/NET0131  ;
  input \u2_L6_reg[4]/NET0131  ;
  input \u2_L6_reg[5]/NET0131  ;
  input \u2_L6_reg[6]/NET0131  ;
  input \u2_L6_reg[7]/NET0131  ;
  input \u2_L6_reg[8]/NET0131  ;
  input \u2_L6_reg[9]/NET0131  ;
  input \u2_L7_reg[10]/NET0131  ;
  input \u2_L7_reg[11]/NET0131  ;
  input \u2_L7_reg[12]/NET0131  ;
  input \u2_L7_reg[13]/NET0131  ;
  input \u2_L7_reg[14]/NET0131  ;
  input \u2_L7_reg[15]/NET0131  ;
  input \u2_L7_reg[16]/NET0131  ;
  input \u2_L7_reg[17]/NET0131  ;
  input \u2_L7_reg[18]/P0001  ;
  input \u2_L7_reg[19]/NET0131  ;
  input \u2_L7_reg[1]/NET0131  ;
  input \u2_L7_reg[20]/NET0131  ;
  input \u2_L7_reg[21]/NET0131  ;
  input \u2_L7_reg[22]/NET0131  ;
  input \u2_L7_reg[23]/NET0131  ;
  input \u2_L7_reg[24]/NET0131  ;
  input \u2_L7_reg[25]/NET0131  ;
  input \u2_L7_reg[26]/NET0131  ;
  input \u2_L7_reg[27]/NET0131  ;
  input \u2_L7_reg[28]/NET0131  ;
  input \u2_L7_reg[29]/NET0131  ;
  input \u2_L7_reg[2]/NET0131  ;
  input \u2_L7_reg[30]/NET0131  ;
  input \u2_L7_reg[31]/NET0131  ;
  input \u2_L7_reg[32]/NET0131  ;
  input \u2_L7_reg[3]/NET0131  ;
  input \u2_L7_reg[4]/NET0131  ;
  input \u2_L7_reg[5]/NET0131  ;
  input \u2_L7_reg[6]/NET0131  ;
  input \u2_L7_reg[7]/NET0131  ;
  input \u2_L7_reg[8]/NET0131  ;
  input \u2_L7_reg[9]/NET0131  ;
  input \u2_L8_reg[10]/NET0131  ;
  input \u2_L8_reg[11]/NET0131  ;
  input \u2_L8_reg[12]/NET0131  ;
  input \u2_L8_reg[13]/NET0131  ;
  input \u2_L8_reg[14]/NET0131  ;
  input \u2_L8_reg[15]/NET0131  ;
  input \u2_L8_reg[16]/NET0131  ;
  input \u2_L8_reg[17]/NET0131  ;
  input \u2_L8_reg[18]/P0001  ;
  input \u2_L8_reg[19]/NET0131  ;
  input \u2_L8_reg[1]/NET0131  ;
  input \u2_L8_reg[20]/NET0131  ;
  input \u2_L8_reg[21]/NET0131  ;
  input \u2_L8_reg[22]/NET0131  ;
  input \u2_L8_reg[23]/NET0131  ;
  input \u2_L8_reg[24]/NET0131  ;
  input \u2_L8_reg[25]/NET0131  ;
  input \u2_L8_reg[26]/NET0131  ;
  input \u2_L8_reg[27]/NET0131  ;
  input \u2_L8_reg[28]/NET0131  ;
  input \u2_L8_reg[29]/NET0131  ;
  input \u2_L8_reg[2]/NET0131  ;
  input \u2_L8_reg[30]/NET0131  ;
  input \u2_L8_reg[31]/NET0131  ;
  input \u2_L8_reg[32]/NET0131  ;
  input \u2_L8_reg[3]/NET0131  ;
  input \u2_L8_reg[4]/NET0131  ;
  input \u2_L8_reg[5]/NET0131  ;
  input \u2_L8_reg[6]/NET0131  ;
  input \u2_L8_reg[7]/NET0131  ;
  input \u2_L8_reg[8]/NET0131  ;
  input \u2_L8_reg[9]/NET0131  ;
  input \u2_L9_reg[10]/NET0131  ;
  input \u2_L9_reg[11]/NET0131  ;
  input \u2_L9_reg[12]/NET0131  ;
  input \u2_L9_reg[13]/NET0131  ;
  input \u2_L9_reg[14]/NET0131  ;
  input \u2_L9_reg[15]/NET0131  ;
  input \u2_L9_reg[16]/NET0131  ;
  input \u2_L9_reg[17]/NET0131  ;
  input \u2_L9_reg[18]/P0001  ;
  input \u2_L9_reg[19]/NET0131  ;
  input \u2_L9_reg[1]/NET0131  ;
  input \u2_L9_reg[20]/NET0131  ;
  input \u2_L9_reg[21]/NET0131  ;
  input \u2_L9_reg[22]/NET0131  ;
  input \u2_L9_reg[23]/NET0131  ;
  input \u2_L9_reg[24]/NET0131  ;
  input \u2_L9_reg[25]/NET0131  ;
  input \u2_L9_reg[26]/NET0131  ;
  input \u2_L9_reg[27]/NET0131  ;
  input \u2_L9_reg[28]/NET0131  ;
  input \u2_L9_reg[29]/NET0131  ;
  input \u2_L9_reg[2]/NET0131  ;
  input \u2_L9_reg[30]/NET0131  ;
  input \u2_L9_reg[31]/NET0131  ;
  input \u2_L9_reg[32]/NET0131  ;
  input \u2_L9_reg[3]/NET0131  ;
  input \u2_L9_reg[4]/NET0131  ;
  input \u2_L9_reg[5]/NET0131  ;
  input \u2_L9_reg[6]/NET0131  ;
  input \u2_L9_reg[7]/NET0131  ;
  input \u2_L9_reg[8]/NET0131  ;
  input \u2_L9_reg[9]/NET0131  ;
  input \u2_R0_reg[10]/NET0131  ;
  input \u2_R0_reg[11]/P0001  ;
  input \u2_R0_reg[12]/NET0131  ;
  input \u2_R0_reg[13]/NET0131  ;
  input \u2_R0_reg[14]/NET0131  ;
  input \u2_R0_reg[15]/NET0131  ;
  input \u2_R0_reg[16]/NET0131  ;
  input \u2_R0_reg[17]/NET0131  ;
  input \u2_R0_reg[18]/NET0131  ;
  input \u2_R0_reg[19]/NET0131  ;
  input \u2_R0_reg[1]/NET0131  ;
  input \u2_R0_reg[20]/NET0131  ;
  input \u2_R0_reg[21]/NET0131  ;
  input \u2_R0_reg[22]/NET0131  ;
  input \u2_R0_reg[23]/NET0131  ;
  input \u2_R0_reg[24]/NET0131  ;
  input \u2_R0_reg[25]/NET0131  ;
  input \u2_R0_reg[26]/NET0131  ;
  input \u2_R0_reg[27]/NET0131  ;
  input \u2_R0_reg[28]/NET0131  ;
  input \u2_R0_reg[29]/NET0131  ;
  input \u2_R0_reg[2]/NET0131  ;
  input \u2_R0_reg[30]/NET0131  ;
  input \u2_R0_reg[31]/P0001  ;
  input \u2_R0_reg[32]/NET0131  ;
  input \u2_R0_reg[3]/NET0131  ;
  input \u2_R0_reg[4]/NET0131  ;
  input \u2_R0_reg[5]/NET0131  ;
  input \u2_R0_reg[6]/NET0131  ;
  input \u2_R0_reg[7]/NET0131  ;
  input \u2_R0_reg[8]/NET0131  ;
  input \u2_R0_reg[9]/NET0131  ;
  input \u2_R10_reg[10]/NET0131  ;
  input \u2_R10_reg[11]/NET0131  ;
  input \u2_R10_reg[12]/NET0131  ;
  input \u2_R10_reg[13]/NET0131  ;
  input \u2_R10_reg[14]/NET0131  ;
  input \u2_R10_reg[15]/NET0131  ;
  input \u2_R10_reg[16]/NET0131  ;
  input \u2_R10_reg[17]/NET0131  ;
  input \u2_R10_reg[18]/NET0131  ;
  input \u2_R10_reg[19]/NET0131  ;
  input \u2_R10_reg[1]/NET0131  ;
  input \u2_R10_reg[20]/NET0131  ;
  input \u2_R10_reg[21]/NET0131  ;
  input \u2_R10_reg[22]/NET0131  ;
  input \u2_R10_reg[23]/NET0131  ;
  input \u2_R10_reg[24]/NET0131  ;
  input \u2_R10_reg[25]/NET0131  ;
  input \u2_R10_reg[26]/NET0131  ;
  input \u2_R10_reg[27]/NET0131  ;
  input \u2_R10_reg[28]/NET0131  ;
  input \u2_R10_reg[29]/NET0131  ;
  input \u2_R10_reg[2]/NET0131  ;
  input \u2_R10_reg[30]/NET0131  ;
  input \u2_R10_reg[31]/P0001  ;
  input \u2_R10_reg[32]/NET0131  ;
  input \u2_R10_reg[3]/NET0131  ;
  input \u2_R10_reg[4]/NET0131  ;
  input \u2_R10_reg[5]/NET0131  ;
  input \u2_R10_reg[6]/NET0131  ;
  input \u2_R10_reg[7]/NET0131  ;
  input \u2_R10_reg[8]/NET0131  ;
  input \u2_R10_reg[9]/NET0131  ;
  input \u2_R11_reg[10]/NET0131  ;
  input \u2_R11_reg[11]/NET0131  ;
  input \u2_R11_reg[12]/NET0131  ;
  input \u2_R11_reg[13]/NET0131  ;
  input \u2_R11_reg[14]/NET0131  ;
  input \u2_R11_reg[15]/NET0131  ;
  input \u2_R11_reg[16]/NET0131  ;
  input \u2_R11_reg[17]/NET0131  ;
  input \u2_R11_reg[18]/NET0131  ;
  input \u2_R11_reg[19]/NET0131  ;
  input \u2_R11_reg[1]/NET0131  ;
  input \u2_R11_reg[20]/NET0131  ;
  input \u2_R11_reg[21]/NET0131  ;
  input \u2_R11_reg[22]/NET0131  ;
  input \u2_R11_reg[23]/NET0131  ;
  input \u2_R11_reg[24]/NET0131  ;
  input \u2_R11_reg[25]/NET0131  ;
  input \u2_R11_reg[26]/NET0131  ;
  input \u2_R11_reg[27]/NET0131  ;
  input \u2_R11_reg[28]/NET0131  ;
  input \u2_R11_reg[29]/NET0131  ;
  input \u2_R11_reg[2]/NET0131  ;
  input \u2_R11_reg[30]/NET0131  ;
  input \u2_R11_reg[31]/P0001  ;
  input \u2_R11_reg[32]/NET0131  ;
  input \u2_R11_reg[3]/NET0131  ;
  input \u2_R11_reg[4]/NET0131  ;
  input \u2_R11_reg[5]/NET0131  ;
  input \u2_R11_reg[6]/NET0131  ;
  input \u2_R11_reg[7]/NET0131  ;
  input \u2_R11_reg[8]/NET0131  ;
  input \u2_R11_reg[9]/NET0131  ;
  input \u2_R12_reg[10]/NET0131  ;
  input \u2_R12_reg[11]/NET0131  ;
  input \u2_R12_reg[12]/NET0131  ;
  input \u2_R12_reg[13]/NET0131  ;
  input \u2_R12_reg[14]/NET0131  ;
  input \u2_R12_reg[15]/NET0131  ;
  input \u2_R12_reg[16]/NET0131  ;
  input \u2_R12_reg[17]/NET0131  ;
  input \u2_R12_reg[18]/NET0131  ;
  input \u2_R12_reg[19]/NET0131  ;
  input \u2_R12_reg[1]/NET0131  ;
  input \u2_R12_reg[20]/NET0131  ;
  input \u2_R12_reg[21]/NET0131  ;
  input \u2_R12_reg[22]/NET0131  ;
  input \u2_R12_reg[23]/NET0131  ;
  input \u2_R12_reg[24]/NET0131  ;
  input \u2_R12_reg[25]/NET0131  ;
  input \u2_R12_reg[26]/NET0131  ;
  input \u2_R12_reg[27]/NET0131  ;
  input \u2_R12_reg[28]/NET0131  ;
  input \u2_R12_reg[29]/NET0131  ;
  input \u2_R12_reg[2]/NET0131  ;
  input \u2_R12_reg[30]/NET0131  ;
  input \u2_R12_reg[31]/P0001  ;
  input \u2_R12_reg[32]/NET0131  ;
  input \u2_R12_reg[3]/NET0131  ;
  input \u2_R12_reg[4]/NET0131  ;
  input \u2_R12_reg[5]/NET0131  ;
  input \u2_R12_reg[6]/NET0131  ;
  input \u2_R12_reg[7]/NET0131  ;
  input \u2_R12_reg[8]/NET0131  ;
  input \u2_R12_reg[9]/NET0131  ;
  input \u2_R13_reg[10]/NET0131  ;
  input \u2_R13_reg[11]/NET0131  ;
  input \u2_R13_reg[12]/NET0131  ;
  input \u2_R13_reg[13]/NET0131  ;
  input \u2_R13_reg[14]/NET0131  ;
  input \u2_R13_reg[15]/NET0131  ;
  input \u2_R13_reg[16]/NET0131  ;
  input \u2_R13_reg[17]/NET0131  ;
  input \u2_R13_reg[18]/NET0131  ;
  input \u2_R13_reg[19]/NET0131  ;
  input \u2_R13_reg[1]/NET0131  ;
  input \u2_R13_reg[20]/NET0131  ;
  input \u2_R13_reg[21]/NET0131  ;
  input \u2_R13_reg[22]/NET0131  ;
  input \u2_R13_reg[23]/NET0131  ;
  input \u2_R13_reg[24]/NET0131  ;
  input \u2_R13_reg[25]/NET0131  ;
  input \u2_R13_reg[26]/NET0131  ;
  input \u2_R13_reg[27]/P0001  ;
  input \u2_R13_reg[28]/NET0131  ;
  input \u2_R13_reg[29]/NET0131  ;
  input \u2_R13_reg[2]/NET0131  ;
  input \u2_R13_reg[30]/NET0131  ;
  input \u2_R13_reg[31]/P0001  ;
  input \u2_R13_reg[32]/NET0131  ;
  input \u2_R13_reg[3]/NET0131  ;
  input \u2_R13_reg[4]/NET0131  ;
  input \u2_R13_reg[5]/NET0131  ;
  input \u2_R13_reg[6]/NET0131  ;
  input \u2_R13_reg[7]/NET0131  ;
  input \u2_R13_reg[8]/NET0131  ;
  input \u2_R13_reg[9]/NET0131  ;
  input \u2_R14_reg[10]/P0001  ;
  input \u2_R14_reg[11]/P0001  ;
  input \u2_R14_reg[12]/NET0131  ;
  input \u2_R14_reg[13]/NET0131  ;
  input \u2_R14_reg[14]/NET0131  ;
  input \u2_R14_reg[15]/NET0131  ;
  input \u2_R14_reg[16]/NET0131  ;
  input \u2_R14_reg[17]/NET0131  ;
  input \u2_R14_reg[18]/NET0131  ;
  input \u2_R14_reg[19]/P0001  ;
  input \u2_R14_reg[1]/NET0131  ;
  input \u2_R14_reg[20]/NET0131  ;
  input \u2_R14_reg[21]/NET0131  ;
  input \u2_R14_reg[22]/P0001  ;
  input \u2_R14_reg[23]/P0001  ;
  input \u2_R14_reg[24]/NET0131  ;
  input \u2_R14_reg[25]/NET0131  ;
  input \u2_R14_reg[26]/P0001  ;
  input \u2_R14_reg[27]/P0001  ;
  input \u2_R14_reg[28]/NET0131  ;
  input \u2_R14_reg[29]/NET0131  ;
  input \u2_R14_reg[2]/NET0131  ;
  input \u2_R14_reg[30]/NET0131  ;
  input \u2_R14_reg[31]/P0001  ;
  input \u2_R14_reg[32]/NET0131  ;
  input \u2_R14_reg[3]/NET0131  ;
  input \u2_R14_reg[4]/NET0131  ;
  input \u2_R14_reg[5]/NET0131  ;
  input \u2_R14_reg[6]/NET0131  ;
  input \u2_R14_reg[7]/P0001  ;
  input \u2_R14_reg[8]/NET0131  ;
  input \u2_R14_reg[9]/NET0131  ;
  input \u2_R1_reg[10]/NET0131  ;
  input \u2_R1_reg[11]/P0001  ;
  input \u2_R1_reg[12]/NET0131  ;
  input \u2_R1_reg[13]/NET0131  ;
  input \u2_R1_reg[14]/NET0131  ;
  input \u2_R1_reg[15]/NET0131  ;
  input \u2_R1_reg[16]/NET0131  ;
  input \u2_R1_reg[17]/NET0131  ;
  input \u2_R1_reg[18]/NET0131  ;
  input \u2_R1_reg[19]/NET0131  ;
  input \u2_R1_reg[1]/NET0131  ;
  input \u2_R1_reg[20]/NET0131  ;
  input \u2_R1_reg[21]/NET0131  ;
  input \u2_R1_reg[22]/NET0131  ;
  input \u2_R1_reg[23]/NET0131  ;
  input \u2_R1_reg[24]/NET0131  ;
  input \u2_R1_reg[25]/NET0131  ;
  input \u2_R1_reg[26]/NET0131  ;
  input \u2_R1_reg[27]/NET0131  ;
  input \u2_R1_reg[28]/NET0131  ;
  input \u2_R1_reg[29]/NET0131  ;
  input \u2_R1_reg[2]/NET0131  ;
  input \u2_R1_reg[30]/NET0131  ;
  input \u2_R1_reg[31]/P0001  ;
  input \u2_R1_reg[32]/NET0131  ;
  input \u2_R1_reg[3]/NET0131  ;
  input \u2_R1_reg[4]/NET0131  ;
  input \u2_R1_reg[5]/NET0131  ;
  input \u2_R1_reg[6]/NET0131  ;
  input \u2_R1_reg[7]/NET0131  ;
  input \u2_R1_reg[8]/NET0131  ;
  input \u2_R1_reg[9]/NET0131  ;
  input \u2_R2_reg[10]/NET0131  ;
  input \u2_R2_reg[11]/NET0131  ;
  input \u2_R2_reg[12]/NET0131  ;
  input \u2_R2_reg[13]/NET0131  ;
  input \u2_R2_reg[14]/NET0131  ;
  input \u2_R2_reg[15]/NET0131  ;
  input \u2_R2_reg[16]/NET0131  ;
  input \u2_R2_reg[17]/NET0131  ;
  input \u2_R2_reg[18]/NET0131  ;
  input \u2_R2_reg[19]/NET0131  ;
  input \u2_R2_reg[1]/NET0131  ;
  input \u2_R2_reg[20]/NET0131  ;
  input \u2_R2_reg[21]/NET0131  ;
  input \u2_R2_reg[22]/NET0131  ;
  input \u2_R2_reg[23]/NET0131  ;
  input \u2_R2_reg[24]/NET0131  ;
  input \u2_R2_reg[25]/NET0131  ;
  input \u2_R2_reg[26]/NET0131  ;
  input \u2_R2_reg[27]/NET0131  ;
  input \u2_R2_reg[28]/NET0131  ;
  input \u2_R2_reg[29]/NET0131  ;
  input \u2_R2_reg[2]/NET0131  ;
  input \u2_R2_reg[30]/NET0131  ;
  input \u2_R2_reg[31]/P0001  ;
  input \u2_R2_reg[32]/NET0131  ;
  input \u2_R2_reg[3]/NET0131  ;
  input \u2_R2_reg[4]/NET0131  ;
  input \u2_R2_reg[5]/NET0131  ;
  input \u2_R2_reg[6]/NET0131  ;
  input \u2_R2_reg[7]/NET0131  ;
  input \u2_R2_reg[8]/NET0131  ;
  input \u2_R2_reg[9]/NET0131  ;
  input \u2_R3_reg[10]/NET0131  ;
  input \u2_R3_reg[11]/P0001  ;
  input \u2_R3_reg[12]/NET0131  ;
  input \u2_R3_reg[13]/NET0131  ;
  input \u2_R3_reg[14]/NET0131  ;
  input \u2_R3_reg[15]/NET0131  ;
  input \u2_R3_reg[16]/NET0131  ;
  input \u2_R3_reg[17]/NET0131  ;
  input \u2_R3_reg[18]/NET0131  ;
  input \u2_R3_reg[19]/NET0131  ;
  input \u2_R3_reg[1]/NET0131  ;
  input \u2_R3_reg[20]/NET0131  ;
  input \u2_R3_reg[21]/NET0131  ;
  input \u2_R3_reg[22]/NET0131  ;
  input \u2_R3_reg[23]/NET0131  ;
  input \u2_R3_reg[24]/NET0131  ;
  input \u2_R3_reg[25]/NET0131  ;
  input \u2_R3_reg[26]/NET0131  ;
  input \u2_R3_reg[27]/NET0131  ;
  input \u2_R3_reg[28]/NET0131  ;
  input \u2_R3_reg[29]/NET0131  ;
  input \u2_R3_reg[2]/NET0131  ;
  input \u2_R3_reg[30]/NET0131  ;
  input \u2_R3_reg[31]/P0001  ;
  input \u2_R3_reg[32]/NET0131  ;
  input \u2_R3_reg[3]/NET0131  ;
  input \u2_R3_reg[4]/NET0131  ;
  input \u2_R3_reg[5]/NET0131  ;
  input \u2_R3_reg[6]/NET0131  ;
  input \u2_R3_reg[7]/NET0131  ;
  input \u2_R3_reg[8]/NET0131  ;
  input \u2_R3_reg[9]/NET0131  ;
  input \u2_R4_reg[10]/NET0131  ;
  input \u2_R4_reg[11]/NET0131  ;
  input \u2_R4_reg[12]/NET0131  ;
  input \u2_R4_reg[13]/NET0131  ;
  input \u2_R4_reg[14]/NET0131  ;
  input \u2_R4_reg[15]/NET0131  ;
  input \u2_R4_reg[16]/NET0131  ;
  input \u2_R4_reg[17]/NET0131  ;
  input \u2_R4_reg[18]/NET0131  ;
  input \u2_R4_reg[19]/NET0131  ;
  input \u2_R4_reg[1]/NET0131  ;
  input \u2_R4_reg[20]/NET0131  ;
  input \u2_R4_reg[21]/NET0131  ;
  input \u2_R4_reg[22]/NET0131  ;
  input \u2_R4_reg[23]/NET0131  ;
  input \u2_R4_reg[24]/NET0131  ;
  input \u2_R4_reg[25]/NET0131  ;
  input \u2_R4_reg[26]/NET0131  ;
  input \u2_R4_reg[27]/NET0131  ;
  input \u2_R4_reg[28]/NET0131  ;
  input \u2_R4_reg[29]/NET0131  ;
  input \u2_R4_reg[2]/NET0131  ;
  input \u2_R4_reg[30]/NET0131  ;
  input \u2_R4_reg[31]/P0001  ;
  input \u2_R4_reg[32]/NET0131  ;
  input \u2_R4_reg[3]/NET0131  ;
  input \u2_R4_reg[4]/NET0131  ;
  input \u2_R4_reg[5]/NET0131  ;
  input \u2_R4_reg[6]/NET0131  ;
  input \u2_R4_reg[7]/NET0131  ;
  input \u2_R4_reg[8]/NET0131  ;
  input \u2_R4_reg[9]/NET0131  ;
  input \u2_R5_reg[10]/NET0131  ;
  input \u2_R5_reg[11]/NET0131  ;
  input \u2_R5_reg[12]/NET0131  ;
  input \u2_R5_reg[13]/NET0131  ;
  input \u2_R5_reg[14]/NET0131  ;
  input \u2_R5_reg[15]/NET0131  ;
  input \u2_R5_reg[16]/NET0131  ;
  input \u2_R5_reg[17]/NET0131  ;
  input \u2_R5_reg[18]/NET0131  ;
  input \u2_R5_reg[19]/NET0131  ;
  input \u2_R5_reg[1]/NET0131  ;
  input \u2_R5_reg[20]/NET0131  ;
  input \u2_R5_reg[21]/NET0131  ;
  input \u2_R5_reg[22]/NET0131  ;
  input \u2_R5_reg[23]/NET0131  ;
  input \u2_R5_reg[24]/NET0131  ;
  input \u2_R5_reg[25]/NET0131  ;
  input \u2_R5_reg[26]/NET0131  ;
  input \u2_R5_reg[27]/NET0131  ;
  input \u2_R5_reg[28]/NET0131  ;
  input \u2_R5_reg[29]/NET0131  ;
  input \u2_R5_reg[2]/NET0131  ;
  input \u2_R5_reg[30]/NET0131  ;
  input \u2_R5_reg[31]/P0001  ;
  input \u2_R5_reg[32]/NET0131  ;
  input \u2_R5_reg[3]/NET0131  ;
  input \u2_R5_reg[4]/NET0131  ;
  input \u2_R5_reg[5]/NET0131  ;
  input \u2_R5_reg[6]/NET0131  ;
  input \u2_R5_reg[7]/NET0131  ;
  input \u2_R5_reg[8]/NET0131  ;
  input \u2_R5_reg[9]/NET0131  ;
  input \u2_R6_reg[10]/NET0131  ;
  input \u2_R6_reg[11]/NET0131  ;
  input \u2_R6_reg[12]/NET0131  ;
  input \u2_R6_reg[13]/NET0131  ;
  input \u2_R6_reg[14]/NET0131  ;
  input \u2_R6_reg[15]/NET0131  ;
  input \u2_R6_reg[16]/NET0131  ;
  input \u2_R6_reg[17]/NET0131  ;
  input \u2_R6_reg[18]/NET0131  ;
  input \u2_R6_reg[19]/NET0131  ;
  input \u2_R6_reg[1]/NET0131  ;
  input \u2_R6_reg[20]/NET0131  ;
  input \u2_R6_reg[21]/NET0131  ;
  input \u2_R6_reg[22]/NET0131  ;
  input \u2_R6_reg[23]/NET0131  ;
  input \u2_R6_reg[24]/NET0131  ;
  input \u2_R6_reg[25]/NET0131  ;
  input \u2_R6_reg[26]/NET0131  ;
  input \u2_R6_reg[27]/NET0131  ;
  input \u2_R6_reg[28]/NET0131  ;
  input \u2_R6_reg[29]/NET0131  ;
  input \u2_R6_reg[2]/NET0131  ;
  input \u2_R6_reg[30]/NET0131  ;
  input \u2_R6_reg[31]/P0001  ;
  input \u2_R6_reg[32]/NET0131  ;
  input \u2_R6_reg[3]/NET0131  ;
  input \u2_R6_reg[4]/NET0131  ;
  input \u2_R6_reg[5]/NET0131  ;
  input \u2_R6_reg[6]/NET0131  ;
  input \u2_R6_reg[7]/NET0131  ;
  input \u2_R6_reg[8]/NET0131  ;
  input \u2_R6_reg[9]/NET0131  ;
  input \u2_R7_reg[10]/NET0131  ;
  input \u2_R7_reg[11]/NET0131  ;
  input \u2_R7_reg[12]/NET0131  ;
  input \u2_R7_reg[13]/NET0131  ;
  input \u2_R7_reg[14]/NET0131  ;
  input \u2_R7_reg[15]/NET0131  ;
  input \u2_R7_reg[16]/NET0131  ;
  input \u2_R7_reg[17]/NET0131  ;
  input \u2_R7_reg[18]/NET0131  ;
  input \u2_R7_reg[19]/NET0131  ;
  input \u2_R7_reg[1]/NET0131  ;
  input \u2_R7_reg[20]/NET0131  ;
  input \u2_R7_reg[21]/NET0131  ;
  input \u2_R7_reg[22]/NET0131  ;
  input \u2_R7_reg[23]/NET0131  ;
  input \u2_R7_reg[24]/NET0131  ;
  input \u2_R7_reg[25]/NET0131  ;
  input \u2_R7_reg[26]/NET0131  ;
  input \u2_R7_reg[27]/NET0131  ;
  input \u2_R7_reg[28]/NET0131  ;
  input \u2_R7_reg[29]/NET0131  ;
  input \u2_R7_reg[2]/NET0131  ;
  input \u2_R7_reg[30]/NET0131  ;
  input \u2_R7_reg[31]/P0001  ;
  input \u2_R7_reg[32]/NET0131  ;
  input \u2_R7_reg[3]/NET0131  ;
  input \u2_R7_reg[4]/NET0131  ;
  input \u2_R7_reg[5]/NET0131  ;
  input \u2_R7_reg[6]/NET0131  ;
  input \u2_R7_reg[7]/NET0131  ;
  input \u2_R7_reg[8]/NET0131  ;
  input \u2_R7_reg[9]/NET0131  ;
  input \u2_R8_reg[10]/NET0131  ;
  input \u2_R8_reg[11]/NET0131  ;
  input \u2_R8_reg[12]/NET0131  ;
  input \u2_R8_reg[13]/NET0131  ;
  input \u2_R8_reg[14]/NET0131  ;
  input \u2_R8_reg[15]/NET0131  ;
  input \u2_R8_reg[16]/NET0131  ;
  input \u2_R8_reg[17]/NET0131  ;
  input \u2_R8_reg[18]/NET0131  ;
  input \u2_R8_reg[19]/NET0131  ;
  input \u2_R8_reg[1]/NET0131  ;
  input \u2_R8_reg[20]/NET0131  ;
  input \u2_R8_reg[21]/NET0131  ;
  input \u2_R8_reg[22]/NET0131  ;
  input \u2_R8_reg[23]/NET0131  ;
  input \u2_R8_reg[24]/NET0131  ;
  input \u2_R8_reg[25]/NET0131  ;
  input \u2_R8_reg[26]/NET0131  ;
  input \u2_R8_reg[27]/NET0131  ;
  input \u2_R8_reg[28]/NET0131  ;
  input \u2_R8_reg[29]/NET0131  ;
  input \u2_R8_reg[2]/NET0131  ;
  input \u2_R8_reg[30]/NET0131  ;
  input \u2_R8_reg[31]/P0001  ;
  input \u2_R8_reg[32]/NET0131  ;
  input \u2_R8_reg[3]/NET0131  ;
  input \u2_R8_reg[4]/NET0131  ;
  input \u2_R8_reg[5]/NET0131  ;
  input \u2_R8_reg[6]/NET0131  ;
  input \u2_R8_reg[7]/NET0131  ;
  input \u2_R8_reg[8]/NET0131  ;
  input \u2_R8_reg[9]/NET0131  ;
  input \u2_R9_reg[10]/NET0131  ;
  input \u2_R9_reg[11]/NET0131  ;
  input \u2_R9_reg[12]/NET0131  ;
  input \u2_R9_reg[13]/NET0131  ;
  input \u2_R9_reg[14]/NET0131  ;
  input \u2_R9_reg[15]/NET0131  ;
  input \u2_R9_reg[16]/NET0131  ;
  input \u2_R9_reg[17]/NET0131  ;
  input \u2_R9_reg[18]/NET0131  ;
  input \u2_R9_reg[19]/NET0131  ;
  input \u2_R9_reg[1]/NET0131  ;
  input \u2_R9_reg[20]/NET0131  ;
  input \u2_R9_reg[21]/NET0131  ;
  input \u2_R9_reg[22]/NET0131  ;
  input \u2_R9_reg[23]/NET0131  ;
  input \u2_R9_reg[24]/NET0131  ;
  input \u2_R9_reg[25]/NET0131  ;
  input \u2_R9_reg[26]/NET0131  ;
  input \u2_R9_reg[27]/NET0131  ;
  input \u2_R9_reg[28]/NET0131  ;
  input \u2_R9_reg[29]/NET0131  ;
  input \u2_R9_reg[2]/NET0131  ;
  input \u2_R9_reg[30]/NET0131  ;
  input \u2_R9_reg[31]/P0001  ;
  input \u2_R9_reg[32]/NET0131  ;
  input \u2_R9_reg[3]/NET0131  ;
  input \u2_R9_reg[4]/NET0131  ;
  input \u2_R9_reg[5]/NET0131  ;
  input \u2_R9_reg[6]/NET0131  ;
  input \u2_R9_reg[7]/NET0131  ;
  input \u2_R9_reg[8]/NET0131  ;
  input \u2_R9_reg[9]/NET0131  ;
  input \u2_desIn_r_reg[0]/NET0131  ;
  input \u2_desIn_r_reg[10]/P0001  ;
  input \u2_desIn_r_reg[11]/NET0131  ;
  input \u2_desIn_r_reg[12]/NET0131  ;
  input \u2_desIn_r_reg[13]/NET0131  ;
  input \u2_desIn_r_reg[14]/NET0131  ;
  input \u2_desIn_r_reg[15]/NET0131  ;
  input \u2_desIn_r_reg[16]/NET0131  ;
  input \u2_desIn_r_reg[17]/NET0131  ;
  input \u2_desIn_r_reg[18]/NET0131  ;
  input \u2_desIn_r_reg[19]/NET0131  ;
  input \u2_desIn_r_reg[1]/NET0131  ;
  input \u2_desIn_r_reg[20]/NET0131  ;
  input \u2_desIn_r_reg[21]/NET0131  ;
  input \u2_desIn_r_reg[22]/NET0131  ;
  input \u2_desIn_r_reg[23]/NET0131  ;
  input \u2_desIn_r_reg[24]/NET0131  ;
  input \u2_desIn_r_reg[25]/NET0131  ;
  input \u2_desIn_r_reg[26]/NET0131  ;
  input \u2_desIn_r_reg[27]/NET0131  ;
  input \u2_desIn_r_reg[28]/NET0131  ;
  input \u2_desIn_r_reg[29]/NET0131  ;
  input \u2_desIn_r_reg[2]/NET0131  ;
  input \u2_desIn_r_reg[30]/NET0131  ;
  input \u2_desIn_r_reg[31]/NET0131  ;
  input \u2_desIn_r_reg[32]/NET0131  ;
  input \u2_desIn_r_reg[33]/NET0131  ;
  input \u2_desIn_r_reg[34]/NET0131  ;
  input \u2_desIn_r_reg[35]/NET0131  ;
  input \u2_desIn_r_reg[36]/NET0131  ;
  input \u2_desIn_r_reg[37]/NET0131  ;
  input \u2_desIn_r_reg[38]/NET0131  ;
  input \u2_desIn_r_reg[39]/NET0131  ;
  input \u2_desIn_r_reg[3]/NET0131  ;
  input \u2_desIn_r_reg[40]/NET0131  ;
  input \u2_desIn_r_reg[41]/NET0131  ;
  input \u2_desIn_r_reg[42]/NET0131  ;
  input \u2_desIn_r_reg[43]/NET0131  ;
  input \u2_desIn_r_reg[44]/NET0131  ;
  input \u2_desIn_r_reg[45]/NET0131  ;
  input \u2_desIn_r_reg[46]/NET0131  ;
  input \u2_desIn_r_reg[47]/NET0131  ;
  input \u2_desIn_r_reg[48]/NET0131  ;
  input \u2_desIn_r_reg[49]/NET0131  ;
  input \u2_desIn_r_reg[4]/NET0131  ;
  input \u2_desIn_r_reg[50]/NET0131  ;
  input \u2_desIn_r_reg[51]/NET0131  ;
  input \u2_desIn_r_reg[52]/NET0131  ;
  input \u2_desIn_r_reg[53]/NET0131  ;
  input \u2_desIn_r_reg[54]/NET0131  ;
  input \u2_desIn_r_reg[55]/NET0131  ;
  input \u2_desIn_r_reg[56]/NET0131  ;
  input \u2_desIn_r_reg[57]/NET0131  ;
  input \u2_desIn_r_reg[58]/NET0131  ;
  input \u2_desIn_r_reg[59]/NET0131  ;
  input \u2_desIn_r_reg[5]/NET0131  ;
  input \u2_desIn_r_reg[60]/NET0131  ;
  input \u2_desIn_r_reg[61]/NET0131  ;
  input \u2_desIn_r_reg[62]/NET0131  ;
  input \u2_desIn_r_reg[63]/NET0131  ;
  input \u2_desIn_r_reg[6]/NET0131  ;
  input \u2_desIn_r_reg[7]/NET0131  ;
  input \u2_desIn_r_reg[8]/NET0131  ;
  input \u2_desIn_r_reg[9]/NET0131  ;
  input \u2_key_r_reg[0]/NET0131  ;
  input \u2_key_r_reg[10]/NET0131  ;
  input \u2_key_r_reg[11]/NET0131  ;
  input \u2_key_r_reg[12]/NET0131  ;
  input \u2_key_r_reg[13]/NET0131  ;
  input \u2_key_r_reg[14]/NET0131  ;
  input \u2_key_r_reg[15]/NET0131  ;
  input \u2_key_r_reg[16]/NET0131  ;
  input \u2_key_r_reg[17]/NET0131  ;
  input \u2_key_r_reg[18]/NET0131  ;
  input \u2_key_r_reg[19]/NET0131  ;
  input \u2_key_r_reg[1]/NET0131  ;
  input \u2_key_r_reg[20]/NET0131  ;
  input \u2_key_r_reg[21]/NET0131  ;
  input \u2_key_r_reg[22]/NET0131  ;
  input \u2_key_r_reg[23]/NET0131  ;
  input \u2_key_r_reg[24]/NET0131  ;
  input \u2_key_r_reg[25]/NET0131  ;
  input \u2_key_r_reg[26]/NET0131  ;
  input \u2_key_r_reg[27]/NET0131  ;
  input \u2_key_r_reg[28]/NET0131  ;
  input \u2_key_r_reg[29]/NET0131  ;
  input \u2_key_r_reg[2]/NET0131  ;
  input \u2_key_r_reg[30]/NET0131  ;
  input \u2_key_r_reg[31]/NET0131  ;
  input \u2_key_r_reg[32]/NET0131  ;
  input \u2_key_r_reg[33]/NET0131  ;
  input \u2_key_r_reg[34]/NET0131  ;
  input \u2_key_r_reg[35]/P0001  ;
  input \u2_key_r_reg[36]/NET0131  ;
  input \u2_key_r_reg[37]/NET0131  ;
  input \u2_key_r_reg[38]/NET0131  ;
  input \u2_key_r_reg[39]/P0001  ;
  input \u2_key_r_reg[3]/NET0131  ;
  input \u2_key_r_reg[40]/NET0131  ;
  input \u2_key_r_reg[41]/NET0131  ;
  input \u2_key_r_reg[42]/P0001  ;
  input \u2_key_r_reg[43]/NET0131  ;
  input \u2_key_r_reg[44]/NET0131  ;
  input \u2_key_r_reg[45]/NET0131  ;
  input \u2_key_r_reg[46]/NET0131  ;
  input \u2_key_r_reg[47]/NET0131  ;
  input \u2_key_r_reg[48]/NET0131  ;
  input \u2_key_r_reg[49]/NET0131  ;
  input \u2_key_r_reg[4]/NET0131  ;
  input \u2_key_r_reg[50]/NET0131  ;
  input \u2_key_r_reg[51]/NET0131  ;
  input \u2_key_r_reg[52]/NET0131  ;
  input \u2_key_r_reg[53]/NET0131  ;
  input \u2_key_r_reg[54]/NET0131  ;
  input \u2_key_r_reg[55]/NET0131  ;
  input \u2_key_r_reg[5]/NET0131  ;
  input \u2_key_r_reg[6]/NET0131  ;
  input \u2_key_r_reg[7]/NET0131  ;
  input \u2_key_r_reg[8]/NET0131  ;
  input \u2_key_r_reg[9]/NET0131  ;
  input \u2_uk_K_r0_reg[0]/NET0131  ;
  input \u2_uk_K_r0_reg[10]/NET0131  ;
  input \u2_uk_K_r0_reg[11]/NET0131  ;
  input \u2_uk_K_r0_reg[12]/NET0131  ;
  input \u2_uk_K_r0_reg[13]/NET0131  ;
  input \u2_uk_K_r0_reg[14]/NET0131  ;
  input \u2_uk_K_r0_reg[15]/NET0131  ;
  input \u2_uk_K_r0_reg[16]/NET0131  ;
  input \u2_uk_K_r0_reg[17]/NET0131  ;
  input \u2_uk_K_r0_reg[18]/NET0131  ;
  input \u2_uk_K_r0_reg[19]/NET0131  ;
  input \u2_uk_K_r0_reg[20]/NET0131  ;
  input \u2_uk_K_r0_reg[21]/NET0131  ;
  input \u2_uk_K_r0_reg[22]/NET0131  ;
  input \u2_uk_K_r0_reg[23]/NET0131  ;
  input \u2_uk_K_r0_reg[24]/P0001  ;
  input \u2_uk_K_r0_reg[25]/P0001  ;
  input \u2_uk_K_r0_reg[26]/NET0131  ;
  input \u2_uk_K_r0_reg[27]/NET0131  ;
  input \u2_uk_K_r0_reg[28]/NET0131  ;
  input \u2_uk_K_r0_reg[29]/NET0131  ;
  input \u2_uk_K_r0_reg[2]/NET0131  ;
  input \u2_uk_K_r0_reg[30]/NET0131  ;
  input \u2_uk_K_r0_reg[31]/NET0131  ;
  input \u2_uk_K_r0_reg[32]/NET0131  ;
  input \u2_uk_K_r0_reg[33]/NET0131  ;
  input \u2_uk_K_r0_reg[34]/NET0131  ;
  input \u2_uk_K_r0_reg[35]/NET0131  ;
  input \u2_uk_K_r0_reg[36]/NET0131  ;
  input \u2_uk_K_r0_reg[37]/NET0131  ;
  input \u2_uk_K_r0_reg[38]/NET0131  ;
  input \u2_uk_K_r0_reg[39]/NET0131  ;
  input \u2_uk_K_r0_reg[3]/NET0131  ;
  input \u2_uk_K_r0_reg[40]/NET0131  ;
  input \u2_uk_K_r0_reg[41]/NET0131  ;
  input \u2_uk_K_r0_reg[42]/NET0131  ;
  input \u2_uk_K_r0_reg[43]/NET0131  ;
  input \u2_uk_K_r0_reg[44]/NET0131  ;
  input \u2_uk_K_r0_reg[45]/NET0131  ;
  input \u2_uk_K_r0_reg[46]/NET0131  ;
  input \u2_uk_K_r0_reg[47]/NET0131  ;
  input \u2_uk_K_r0_reg[48]/NET0131  ;
  input \u2_uk_K_r0_reg[49]/NET0131  ;
  input \u2_uk_K_r0_reg[4]/NET0131  ;
  input \u2_uk_K_r0_reg[50]/NET0131  ;
  input \u2_uk_K_r0_reg[51]/NET0131  ;
  input \u2_uk_K_r0_reg[52]/P0001  ;
  input \u2_uk_K_r0_reg[54]/NET0131  ;
  input \u2_uk_K_r0_reg[55]/NET0131  ;
  input \u2_uk_K_r0_reg[5]/NET0131  ;
  input \u2_uk_K_r0_reg[6]/NET0131  ;
  input \u2_uk_K_r0_reg[7]/NET0131  ;
  input \u2_uk_K_r0_reg[8]/NET0131  ;
  input \u2_uk_K_r0_reg[9]/NET0131  ;
  input \u2_uk_K_r10_reg[0]/NET0131  ;
  input \u2_uk_K_r10_reg[10]/NET0131  ;
  input \u2_uk_K_r10_reg[11]/NET0131  ;
  input \u2_uk_K_r10_reg[12]/NET0131  ;
  input \u2_uk_K_r10_reg[14]/NET0131  ;
  input \u2_uk_K_r10_reg[15]/NET0131  ;
  input \u2_uk_K_r10_reg[16]/NET0131  ;
  input \u2_uk_K_r10_reg[17]/NET0131  ;
  input \u2_uk_K_r10_reg[18]/NET0131  ;
  input \u2_uk_K_r10_reg[19]/NET0131  ;
  input \u2_uk_K_r10_reg[1]/NET0131  ;
  input \u2_uk_K_r10_reg[20]/NET0131  ;
  input \u2_uk_K_r10_reg[21]/NET0131  ;
  input \u2_uk_K_r10_reg[22]/NET0131  ;
  input \u2_uk_K_r10_reg[23]/NET0131  ;
  input \u2_uk_K_r10_reg[24]/NET0131  ;
  input \u2_uk_K_r10_reg[25]/NET0131  ;
  input \u2_uk_K_r10_reg[26]/NET0131  ;
  input \u2_uk_K_r10_reg[27]/NET0131  ;
  input \u2_uk_K_r10_reg[28]/NET0131  ;
  input \u2_uk_K_r10_reg[29]/NET0131  ;
  input \u2_uk_K_r10_reg[2]/NET0131  ;
  input \u2_uk_K_r10_reg[30]/NET0131  ;
  input \u2_uk_K_r10_reg[31]/NET0131  ;
  input \u2_uk_K_r10_reg[32]/NET0131  ;
  input \u2_uk_K_r10_reg[33]/NET0131  ;
  input \u2_uk_K_r10_reg[34]/NET0131  ;
  input \u2_uk_K_r10_reg[35]/NET0131  ;
  input \u2_uk_K_r10_reg[36]/NET0131  ;
  input \u2_uk_K_r10_reg[37]/NET0131  ;
  input \u2_uk_K_r10_reg[38]/NET0131  ;
  input \u2_uk_K_r10_reg[39]/NET0131  ;
  input \u2_uk_K_r10_reg[3]/NET0131  ;
  input \u2_uk_K_r10_reg[40]/NET0131  ;
  input \u2_uk_K_r10_reg[41]/NET0131  ;
  input \u2_uk_K_r10_reg[42]/NET0131  ;
  input \u2_uk_K_r10_reg[43]/NET0131  ;
  input \u2_uk_K_r10_reg[44]/NET0131  ;
  input \u2_uk_K_r10_reg[45]/P0001  ;
  input \u2_uk_K_r10_reg[46]/NET0131  ;
  input \u2_uk_K_r10_reg[47]/NET0131  ;
  input \u2_uk_K_r10_reg[48]/NET0131  ;
  input \u2_uk_K_r10_reg[49]/NET0131  ;
  input \u2_uk_K_r10_reg[4]/NET0131  ;
  input \u2_uk_K_r10_reg[50]/NET0131  ;
  input \u2_uk_K_r10_reg[51]/NET0131  ;
  input \u2_uk_K_r10_reg[52]/NET0131  ;
  input \u2_uk_K_r10_reg[53]/NET0131  ;
  input \u2_uk_K_r10_reg[54]/NET0131  ;
  input \u2_uk_K_r10_reg[55]/NET0131  ;
  input \u2_uk_K_r10_reg[5]/NET0131  ;
  input \u2_uk_K_r10_reg[6]/NET0131  ;
  input \u2_uk_K_r10_reg[7]/NET0131  ;
  input \u2_uk_K_r10_reg[8]/NET0131  ;
  input \u2_uk_K_r10_reg[9]/NET0131  ;
  input \u2_uk_K_r11_reg[0]/NET0131  ;
  input \u2_uk_K_r11_reg[10]/NET0131  ;
  input \u2_uk_K_r11_reg[11]/NET0131  ;
  input \u2_uk_K_r11_reg[12]/NET0131  ;
  input \u2_uk_K_r11_reg[13]/NET0131  ;
  input \u2_uk_K_r11_reg[14]/NET0131  ;
  input \u2_uk_K_r11_reg[15]/NET0131  ;
  input \u2_uk_K_r11_reg[16]/NET0131  ;
  input \u2_uk_K_r11_reg[17]/NET0131  ;
  input \u2_uk_K_r11_reg[18]/NET0131  ;
  input \u2_uk_K_r11_reg[19]/NET0131  ;
  input \u2_uk_K_r11_reg[1]/NET0131  ;
  input \u2_uk_K_r11_reg[20]/NET0131  ;
  input \u2_uk_K_r11_reg[21]/NET0131  ;
  input \u2_uk_K_r11_reg[22]/NET0131  ;
  input \u2_uk_K_r11_reg[23]/NET0131  ;
  input \u2_uk_K_r11_reg[24]/NET0131  ;
  input \u2_uk_K_r11_reg[25]/NET0131  ;
  input \u2_uk_K_r11_reg[26]/NET0131  ;
  input \u2_uk_K_r11_reg[27]/NET0131  ;
  input \u2_uk_K_r11_reg[28]/NET0131  ;
  input \u2_uk_K_r11_reg[29]/NET0131  ;
  input \u2_uk_K_r11_reg[2]/NET0131  ;
  input \u2_uk_K_r11_reg[31]/NET0131  ;
  input \u2_uk_K_r11_reg[32]/NET0131  ;
  input \u2_uk_K_r11_reg[33]/NET0131  ;
  input \u2_uk_K_r11_reg[34]/NET0131  ;
  input \u2_uk_K_r11_reg[35]/NET0131  ;
  input \u2_uk_K_r11_reg[36]/NET0131  ;
  input \u2_uk_K_r11_reg[37]/NET0131  ;
  input \u2_uk_K_r11_reg[38]/NET0131  ;
  input \u2_uk_K_r11_reg[39]/NET0131  ;
  input \u2_uk_K_r11_reg[3]/NET0131  ;
  input \u2_uk_K_r11_reg[40]/NET0131  ;
  input \u2_uk_K_r11_reg[41]/NET0131  ;
  input \u2_uk_K_r11_reg[42]/NET0131  ;
  input \u2_uk_K_r11_reg[43]/NET0131  ;
  input \u2_uk_K_r11_reg[44]/NET0131  ;
  input \u2_uk_K_r11_reg[45]/NET0131  ;
  input \u2_uk_K_r11_reg[46]/NET0131  ;
  input \u2_uk_K_r11_reg[47]/NET0131  ;
  input \u2_uk_K_r11_reg[48]/NET0131  ;
  input \u2_uk_K_r11_reg[49]/NET0131  ;
  input \u2_uk_K_r11_reg[4]/NET0131  ;
  input \u2_uk_K_r11_reg[50]/NET0131  ;
  input \u2_uk_K_r11_reg[51]/NET0131  ;
  input \u2_uk_K_r11_reg[52]/NET0131  ;
  input \u2_uk_K_r11_reg[53]/P0001  ;
  input \u2_uk_K_r11_reg[54]/NET0131  ;
  input \u2_uk_K_r11_reg[55]/NET0131  ;
  input \u2_uk_K_r11_reg[5]/NET0131  ;
  input \u2_uk_K_r11_reg[6]/NET0131  ;
  input \u2_uk_K_r11_reg[7]/NET0131  ;
  input \u2_uk_K_r11_reg[8]/NET0131  ;
  input \u2_uk_K_r11_reg[9]/NET0131  ;
  input \u2_uk_K_r12_reg[0]/NET0131  ;
  input \u2_uk_K_r12_reg[10]/P0001  ;
  input \u2_uk_K_r12_reg[11]/NET0131  ;
  input \u2_uk_K_r12_reg[12]/NET0131  ;
  input \u2_uk_K_r12_reg[13]/NET0131  ;
  input \u2_uk_K_r12_reg[14]/NET0131  ;
  input \u2_uk_K_r12_reg[15]/NET0131  ;
  input \u2_uk_K_r12_reg[16]/NET0131  ;
  input \u2_uk_K_r12_reg[17]/NET0131  ;
  input \u2_uk_K_r12_reg[18]/NET0131  ;
  input \u2_uk_K_r12_reg[19]/NET0131  ;
  input \u2_uk_K_r12_reg[1]/NET0131  ;
  input \u2_uk_K_r12_reg[20]/NET0131  ;
  input \u2_uk_K_r12_reg[21]/NET0131  ;
  input \u2_uk_K_r12_reg[22]/NET0131  ;
  input \u2_uk_K_r12_reg[23]/NET0131  ;
  input \u2_uk_K_r12_reg[24]/NET0131  ;
  input \u2_uk_K_r12_reg[25]/NET0131  ;
  input \u2_uk_K_r12_reg[26]/NET0131  ;
  input \u2_uk_K_r12_reg[27]/NET0131  ;
  input \u2_uk_K_r12_reg[28]/NET0131  ;
  input \u2_uk_K_r12_reg[29]/NET0131  ;
  input \u2_uk_K_r12_reg[2]/NET0131  ;
  input \u2_uk_K_r12_reg[30]/NET0131  ;
  input \u2_uk_K_r12_reg[31]/NET0131  ;
  input \u2_uk_K_r12_reg[32]/NET0131  ;
  input \u2_uk_K_r12_reg[33]/NET0131  ;
  input \u2_uk_K_r12_reg[34]/NET0131  ;
  input \u2_uk_K_r12_reg[35]/NET0131  ;
  input \u2_uk_K_r12_reg[36]/NET0131  ;
  input \u2_uk_K_r12_reg[37]/NET0131  ;
  input \u2_uk_K_r12_reg[38]/NET0131  ;
  input \u2_uk_K_r12_reg[3]/NET0131  ;
  input \u2_uk_K_r12_reg[40]/NET0131  ;
  input \u2_uk_K_r12_reg[41]/NET0131  ;
  input \u2_uk_K_r12_reg[42]/NET0131  ;
  input \u2_uk_K_r12_reg[43]/NET0131  ;
  input \u2_uk_K_r12_reg[44]/P0001  ;
  input \u2_uk_K_r12_reg[45]/NET0131  ;
  input \u2_uk_K_r12_reg[46]/NET0131  ;
  input \u2_uk_K_r12_reg[47]/NET0131  ;
  input \u2_uk_K_r12_reg[48]/NET0131  ;
  input \u2_uk_K_r12_reg[49]/NET0131  ;
  input \u2_uk_K_r12_reg[4]/NET0131  ;
  input \u2_uk_K_r12_reg[50]/NET0131  ;
  input \u2_uk_K_r12_reg[51]/NET0131  ;
  input \u2_uk_K_r12_reg[52]/NET0131  ;
  input \u2_uk_K_r12_reg[53]/NET0131  ;
  input \u2_uk_K_r12_reg[54]/NET0131  ;
  input \u2_uk_K_r12_reg[55]/NET0131  ;
  input \u2_uk_K_r12_reg[5]/NET0131  ;
  input \u2_uk_K_r12_reg[6]/NET0131  ;
  input \u2_uk_K_r12_reg[7]/P0001  ;
  input \u2_uk_K_r12_reg[8]/NET0131  ;
  input \u2_uk_K_r12_reg[9]/NET0131  ;
  input \u2_uk_K_r13_reg[0]/NET0131  ;
  input \u2_uk_K_r13_reg[10]/NET0131  ;
  input \u2_uk_K_r13_reg[11]/NET0131  ;
  input \u2_uk_K_r13_reg[12]/NET0131  ;
  input \u2_uk_K_r13_reg[13]/NET0131  ;
  input \u2_uk_K_r13_reg[14]/NET0131  ;
  input \u2_uk_K_r13_reg[15]/NET0131  ;
  input \u2_uk_K_r13_reg[16]/NET0131  ;
  input \u2_uk_K_r13_reg[17]/NET0131  ;
  input \u2_uk_K_r13_reg[18]/NET0131  ;
  input \u2_uk_K_r13_reg[19]/NET0131  ;
  input \u2_uk_K_r13_reg[20]/NET0131  ;
  input \u2_uk_K_r13_reg[21]/NET0131  ;
  input \u2_uk_K_r13_reg[22]/NET0131  ;
  input \u2_uk_K_r13_reg[23]/NET0131  ;
  input \u2_uk_K_r13_reg[24]/NET0131  ;
  input \u2_uk_K_r13_reg[25]/P0001  ;
  input \u2_uk_K_r13_reg[26]/NET0131  ;
  input \u2_uk_K_r13_reg[27]/NET0131  ;
  input \u2_uk_K_r13_reg[28]/NET0131  ;
  input \u2_uk_K_r13_reg[29]/NET0131  ;
  input \u2_uk_K_r13_reg[2]/NET0131  ;
  input \u2_uk_K_r13_reg[30]/NET0131  ;
  input \u2_uk_K_r13_reg[31]/NET0131  ;
  input \u2_uk_K_r13_reg[32]/NET0131  ;
  input \u2_uk_K_r13_reg[33]/NET0131  ;
  input \u2_uk_K_r13_reg[34]/NET0131  ;
  input \u2_uk_K_r13_reg[35]/NET0131  ;
  input \u2_uk_K_r13_reg[36]/NET0131  ;
  input \u2_uk_K_r13_reg[37]/NET0131  ;
  input \u2_uk_K_r13_reg[38]/NET0131  ;
  input \u2_uk_K_r13_reg[39]/NET0131  ;
  input \u2_uk_K_r13_reg[3]/NET0131  ;
  input \u2_uk_K_r13_reg[40]/NET0131  ;
  input \u2_uk_K_r13_reg[41]/NET0131  ;
  input \u2_uk_K_r13_reg[42]/NET0131  ;
  input \u2_uk_K_r13_reg[43]/NET0131  ;
  input \u2_uk_K_r13_reg[44]/NET0131  ;
  input \u2_uk_K_r13_reg[45]/NET0131  ;
  input \u2_uk_K_r13_reg[46]/NET0131  ;
  input \u2_uk_K_r13_reg[47]/NET0131  ;
  input \u2_uk_K_r13_reg[48]/NET0131  ;
  input \u2_uk_K_r13_reg[49]/NET0131  ;
  input \u2_uk_K_r13_reg[4]/NET0131  ;
  input \u2_uk_K_r13_reg[50]/NET0131  ;
  input \u2_uk_K_r13_reg[51]/NET0131  ;
  input \u2_uk_K_r13_reg[52]/NET0131  ;
  input \u2_uk_K_r13_reg[54]/NET0131  ;
  input \u2_uk_K_r13_reg[55]/NET0131  ;
  input \u2_uk_K_r13_reg[5]/NET0131  ;
  input \u2_uk_K_r13_reg[6]/NET0131  ;
  input \u2_uk_K_r13_reg[7]/NET0131  ;
  input \u2_uk_K_r13_reg[8]/NET0131  ;
  input \u2_uk_K_r13_reg[9]/NET0131  ;
  input \u2_uk_K_r14_reg[0]/NET0131  ;
  input \u2_uk_K_r14_reg[10]/P0001  ;
  input \u2_uk_K_r14_reg[11]/NET0131  ;
  input \u2_uk_K_r14_reg[12]/NET0131  ;
  input \u2_uk_K_r14_reg[13]/NET0131  ;
  input \u2_uk_K_r14_reg[14]/NET0131  ;
  input \u2_uk_K_r14_reg[15]/NET0131  ;
  input \u2_uk_K_r14_reg[16]/NET0131  ;
  input \u2_uk_K_r14_reg[17]/NET0131  ;
  input \u2_uk_K_r14_reg[18]/NET0131  ;
  input \u2_uk_K_r14_reg[19]/NET0131  ;
  input \u2_uk_K_r14_reg[1]/NET0131  ;
  input \u2_uk_K_r14_reg[20]/NET0131  ;
  input \u2_uk_K_r14_reg[21]/NET0131  ;
  input \u2_uk_K_r14_reg[22]/NET0131  ;
  input \u2_uk_K_r14_reg[23]/NET0131  ;
  input \u2_uk_K_r14_reg[24]/NET0131  ;
  input \u2_uk_K_r14_reg[25]/NET0131  ;
  input \u2_uk_K_r14_reg[26]/NET0131  ;
  input \u2_uk_K_r14_reg[27]/NET0131  ;
  input \u2_uk_K_r14_reg[28]/NET0131  ;
  input \u2_uk_K_r14_reg[29]/NET0131  ;
  input \u2_uk_K_r14_reg[2]/NET0131  ;
  input \u2_uk_K_r14_reg[30]/NET0131  ;
  input \u2_uk_K_r14_reg[31]/NET0131  ;
  input \u2_uk_K_r14_reg[32]/NET0131  ;
  input \u2_uk_K_r14_reg[33]/NET0131  ;
  input \u2_uk_K_r14_reg[34]/NET0131  ;
  input \u2_uk_K_r14_reg[35]/P0001  ;
  input \u2_uk_K_r14_reg[36]/NET0131  ;
  input \u2_uk_K_r14_reg[37]/NET0131  ;
  input \u2_uk_K_r14_reg[38]/NET0131  ;
  input \u2_uk_K_r14_reg[39]/P0001  ;
  input \u2_uk_K_r14_reg[3]/NET0131  ;
  input \u2_uk_K_r14_reg[40]/NET0131  ;
  input \u2_uk_K_r14_reg[41]/NET0131  ;
  input \u2_uk_K_r14_reg[42]/P0001  ;
  input \u2_uk_K_r14_reg[43]/NET0131  ;
  input \u2_uk_K_r14_reg[44]/NET0131  ;
  input \u2_uk_K_r14_reg[45]/NET0131  ;
  input \u2_uk_K_r14_reg[46]/NET0131  ;
  input \u2_uk_K_r14_reg[47]/NET0131  ;
  input \u2_uk_K_r14_reg[48]/NET0131  ;
  input \u2_uk_K_r14_reg[49]/P0001  ;
  input \u2_uk_K_r14_reg[4]/NET0131  ;
  input \u2_uk_K_r14_reg[50]/NET0131  ;
  input \u2_uk_K_r14_reg[51]/NET0131  ;
  input \u2_uk_K_r14_reg[52]/NET0131  ;
  input \u2_uk_K_r14_reg[53]/NET0131  ;
  input \u2_uk_K_r14_reg[54]/NET0131  ;
  input \u2_uk_K_r14_reg[55]/NET0131  ;
  input \u2_uk_K_r14_reg[5]/NET0131  ;
  input \u2_uk_K_r14_reg[6]/NET0131  ;
  input \u2_uk_K_r14_reg[7]/NET0131  ;
  input \u2_uk_K_r14_reg[8]/NET0131  ;
  input \u2_uk_K_r14_reg[9]/NET0131  ;
  input \u2_uk_K_r1_reg[0]/NET0131  ;
  input \u2_uk_K_r1_reg[10]/P0001  ;
  input \u2_uk_K_r1_reg[11]/NET0131  ;
  input \u2_uk_K_r1_reg[12]/NET0131  ;
  input \u2_uk_K_r1_reg[13]/NET0131  ;
  input \u2_uk_K_r1_reg[14]/NET0131  ;
  input \u2_uk_K_r1_reg[15]/NET0131  ;
  input \u2_uk_K_r1_reg[16]/NET0131  ;
  input \u2_uk_K_r1_reg[17]/NET0131  ;
  input \u2_uk_K_r1_reg[18]/NET0131  ;
  input \u2_uk_K_r1_reg[19]/NET0131  ;
  input \u2_uk_K_r1_reg[1]/NET0131  ;
  input \u2_uk_K_r1_reg[20]/NET0131  ;
  input \u2_uk_K_r1_reg[21]/NET0131  ;
  input \u2_uk_K_r1_reg[22]/NET0131  ;
  input \u2_uk_K_r1_reg[23]/NET0131  ;
  input \u2_uk_K_r1_reg[24]/NET0131  ;
  input \u2_uk_K_r1_reg[25]/NET0131  ;
  input \u2_uk_K_r1_reg[26]/NET0131  ;
  input \u2_uk_K_r1_reg[27]/NET0131  ;
  input \u2_uk_K_r1_reg[28]/NET0131  ;
  input \u2_uk_K_r1_reg[29]/NET0131  ;
  input \u2_uk_K_r1_reg[2]/NET0131  ;
  input \u2_uk_K_r1_reg[30]/NET0131  ;
  input \u2_uk_K_r1_reg[31]/NET0131  ;
  input \u2_uk_K_r1_reg[32]/NET0131  ;
  input \u2_uk_K_r1_reg[33]/NET0131  ;
  input \u2_uk_K_r1_reg[34]/NET0131  ;
  input \u2_uk_K_r1_reg[35]/NET0131  ;
  input \u2_uk_K_r1_reg[36]/NET0131  ;
  input \u2_uk_K_r1_reg[37]/NET0131  ;
  input \u2_uk_K_r1_reg[38]/NET0131  ;
  input \u2_uk_K_r1_reg[3]/NET0131  ;
  input \u2_uk_K_r1_reg[40]/NET0131  ;
  input \u2_uk_K_r1_reg[41]/NET0131  ;
  input \u2_uk_K_r1_reg[42]/NET0131  ;
  input \u2_uk_K_r1_reg[43]/NET0131  ;
  input \u2_uk_K_r1_reg[44]/P0001  ;
  input \u2_uk_K_r1_reg[45]/NET0131  ;
  input \u2_uk_K_r1_reg[46]/NET0131  ;
  input \u2_uk_K_r1_reg[47]/NET0131  ;
  input \u2_uk_K_r1_reg[48]/NET0131  ;
  input \u2_uk_K_r1_reg[49]/NET0131  ;
  input \u2_uk_K_r1_reg[4]/NET0131  ;
  input \u2_uk_K_r1_reg[50]/NET0131  ;
  input \u2_uk_K_r1_reg[51]/NET0131  ;
  input \u2_uk_K_r1_reg[52]/NET0131  ;
  input \u2_uk_K_r1_reg[53]/NET0131  ;
  input \u2_uk_K_r1_reg[54]/NET0131  ;
  input \u2_uk_K_r1_reg[55]/NET0131  ;
  input \u2_uk_K_r1_reg[5]/NET0131  ;
  input \u2_uk_K_r1_reg[6]/NET0131  ;
  input \u2_uk_K_r1_reg[7]/P0001  ;
  input \u2_uk_K_r1_reg[8]/NET0131  ;
  input \u2_uk_K_r1_reg[9]/NET0131  ;
  input \u2_uk_K_r2_reg[0]/NET0131  ;
  input \u2_uk_K_r2_reg[10]/NET0131  ;
  input \u2_uk_K_r2_reg[11]/NET0131  ;
  input \u2_uk_K_r2_reg[12]/NET0131  ;
  input \u2_uk_K_r2_reg[13]/NET0131  ;
  input \u2_uk_K_r2_reg[14]/NET0131  ;
  input \u2_uk_K_r2_reg[15]/NET0131  ;
  input \u2_uk_K_r2_reg[16]/NET0131  ;
  input \u2_uk_K_r2_reg[17]/NET0131  ;
  input \u2_uk_K_r2_reg[18]/NET0131  ;
  input \u2_uk_K_r2_reg[19]/NET0131  ;
  input \u2_uk_K_r2_reg[1]/NET0131  ;
  input \u2_uk_K_r2_reg[20]/NET0131  ;
  input \u2_uk_K_r2_reg[21]/NET0131  ;
  input \u2_uk_K_r2_reg[22]/NET0131  ;
  input \u2_uk_K_r2_reg[23]/NET0131  ;
  input \u2_uk_K_r2_reg[24]/NET0131  ;
  input \u2_uk_K_r2_reg[25]/NET0131  ;
  input \u2_uk_K_r2_reg[26]/NET0131  ;
  input \u2_uk_K_r2_reg[27]/NET0131  ;
  input \u2_uk_K_r2_reg[28]/NET0131  ;
  input \u2_uk_K_r2_reg[29]/NET0131  ;
  input \u2_uk_K_r2_reg[2]/NET0131  ;
  input \u2_uk_K_r2_reg[31]/NET0131  ;
  input \u2_uk_K_r2_reg[32]/NET0131  ;
  input \u2_uk_K_r2_reg[33]/NET0131  ;
  input \u2_uk_K_r2_reg[34]/NET0131  ;
  input \u2_uk_K_r2_reg[35]/NET0131  ;
  input \u2_uk_K_r2_reg[36]/NET0131  ;
  input \u2_uk_K_r2_reg[37]/NET0131  ;
  input \u2_uk_K_r2_reg[38]/NET0131  ;
  input \u2_uk_K_r2_reg[39]/NET0131  ;
  input \u2_uk_K_r2_reg[3]/NET0131  ;
  input \u2_uk_K_r2_reg[40]/NET0131  ;
  input \u2_uk_K_r2_reg[41]/NET0131  ;
  input \u2_uk_K_r2_reg[42]/NET0131  ;
  input \u2_uk_K_r2_reg[43]/NET0131  ;
  input \u2_uk_K_r2_reg[44]/NET0131  ;
  input \u2_uk_K_r2_reg[45]/NET0131  ;
  input \u2_uk_K_r2_reg[46]/NET0131  ;
  input \u2_uk_K_r2_reg[47]/NET0131  ;
  input \u2_uk_K_r2_reg[48]/NET0131  ;
  input \u2_uk_K_r2_reg[49]/NET0131  ;
  input \u2_uk_K_r2_reg[4]/NET0131  ;
  input \u2_uk_K_r2_reg[50]/NET0131  ;
  input \u2_uk_K_r2_reg[51]/NET0131  ;
  input \u2_uk_K_r2_reg[52]/NET0131  ;
  input \u2_uk_K_r2_reg[53]/P0001  ;
  input \u2_uk_K_r2_reg[54]/NET0131  ;
  input \u2_uk_K_r2_reg[55]/NET0131  ;
  input \u2_uk_K_r2_reg[5]/NET0131  ;
  input \u2_uk_K_r2_reg[6]/NET0131  ;
  input \u2_uk_K_r2_reg[7]/NET0131  ;
  input \u2_uk_K_r2_reg[8]/NET0131  ;
  input \u2_uk_K_r2_reg[9]/NET0131  ;
  input \u2_uk_K_r3_reg[0]/NET0131  ;
  input \u2_uk_K_r3_reg[10]/NET0131  ;
  input \u2_uk_K_r3_reg[11]/NET0131  ;
  input \u2_uk_K_r3_reg[12]/NET0131  ;
  input \u2_uk_K_r3_reg[14]/NET0131  ;
  input \u2_uk_K_r3_reg[15]/NET0131  ;
  input \u2_uk_K_r3_reg[16]/NET0131  ;
  input \u2_uk_K_r3_reg[17]/NET0131  ;
  input \u2_uk_K_r3_reg[18]/NET0131  ;
  input \u2_uk_K_r3_reg[19]/NET0131  ;
  input \u2_uk_K_r3_reg[1]/NET0131  ;
  input \u2_uk_K_r3_reg[20]/NET0131  ;
  input \u2_uk_K_r3_reg[21]/NET0131  ;
  input \u2_uk_K_r3_reg[22]/NET0131  ;
  input \u2_uk_K_r3_reg[23]/NET0131  ;
  input \u2_uk_K_r3_reg[24]/NET0131  ;
  input \u2_uk_K_r3_reg[25]/NET0131  ;
  input \u2_uk_K_r3_reg[26]/NET0131  ;
  input \u2_uk_K_r3_reg[27]/NET0131  ;
  input \u2_uk_K_r3_reg[28]/NET0131  ;
  input \u2_uk_K_r3_reg[29]/NET0131  ;
  input \u2_uk_K_r3_reg[2]/NET0131  ;
  input \u2_uk_K_r3_reg[30]/NET0131  ;
  input \u2_uk_K_r3_reg[31]/NET0131  ;
  input \u2_uk_K_r3_reg[32]/NET0131  ;
  input \u2_uk_K_r3_reg[33]/NET0131  ;
  input \u2_uk_K_r3_reg[34]/NET0131  ;
  input \u2_uk_K_r3_reg[35]/NET0131  ;
  input \u2_uk_K_r3_reg[36]/NET0131  ;
  input \u2_uk_K_r3_reg[37]/NET0131  ;
  input \u2_uk_K_r3_reg[38]/NET0131  ;
  input \u2_uk_K_r3_reg[39]/NET0131  ;
  input \u2_uk_K_r3_reg[3]/NET0131  ;
  input \u2_uk_K_r3_reg[40]/NET0131  ;
  input \u2_uk_K_r3_reg[41]/NET0131  ;
  input \u2_uk_K_r3_reg[42]/NET0131  ;
  input \u2_uk_K_r3_reg[43]/NET0131  ;
  input \u2_uk_K_r3_reg[44]/NET0131  ;
  input \u2_uk_K_r3_reg[45]/P0001  ;
  input \u2_uk_K_r3_reg[46]/NET0131  ;
  input \u2_uk_K_r3_reg[47]/NET0131  ;
  input \u2_uk_K_r3_reg[48]/NET0131  ;
  input \u2_uk_K_r3_reg[49]/NET0131  ;
  input \u2_uk_K_r3_reg[4]/NET0131  ;
  input \u2_uk_K_r3_reg[50]/NET0131  ;
  input \u2_uk_K_r3_reg[51]/NET0131  ;
  input \u2_uk_K_r3_reg[52]/NET0131  ;
  input \u2_uk_K_r3_reg[53]/NET0131  ;
  input \u2_uk_K_r3_reg[54]/NET0131  ;
  input \u2_uk_K_r3_reg[55]/NET0131  ;
  input \u2_uk_K_r3_reg[5]/NET0131  ;
  input \u2_uk_K_r3_reg[6]/NET0131  ;
  input \u2_uk_K_r3_reg[7]/NET0131  ;
  input \u2_uk_K_r3_reg[8]/NET0131  ;
  input \u2_uk_K_r3_reg[9]/NET0131  ;
  input \u2_uk_K_r4_reg[0]/P0001  ;
  input \u2_uk_K_r4_reg[10]/NET0131  ;
  input \u2_uk_K_r4_reg[11]/NET0131  ;
  input \u2_uk_K_r4_reg[12]/NET0131  ;
  input \u2_uk_K_r4_reg[13]/NET0131  ;
  input \u2_uk_K_r4_reg[14]/NET0131  ;
  input \u2_uk_K_r4_reg[15]/NET0131  ;
  input \u2_uk_K_r4_reg[16]/NET0131  ;
  input \u2_uk_K_r4_reg[17]/NET0131  ;
  input \u2_uk_K_r4_reg[18]/NET0131  ;
  input \u2_uk_K_r4_reg[19]/NET0131  ;
  input \u2_uk_K_r4_reg[1]/NET0131  ;
  input \u2_uk_K_r4_reg[20]/NET0131  ;
  input \u2_uk_K_r4_reg[21]/NET0131  ;
  input \u2_uk_K_r4_reg[22]/NET0131  ;
  input \u2_uk_K_r4_reg[23]/NET0131  ;
  input \u2_uk_K_r4_reg[25]/NET0131  ;
  input \u2_uk_K_r4_reg[26]/NET0131  ;
  input \u2_uk_K_r4_reg[27]/P0001  ;
  input \u2_uk_K_r4_reg[28]/NET0131  ;
  input \u2_uk_K_r4_reg[29]/NET0131  ;
  input \u2_uk_K_r4_reg[30]/NET0131  ;
  input \u2_uk_K_r4_reg[31]/P0001  ;
  input \u2_uk_K_r4_reg[32]/NET0131  ;
  input \u2_uk_K_r4_reg[33]/NET0131  ;
  input \u2_uk_K_r4_reg[34]/NET0131  ;
  input \u2_uk_K_r4_reg[35]/NET0131  ;
  input \u2_uk_K_r4_reg[36]/NET0131  ;
  input \u2_uk_K_r4_reg[37]/NET0131  ;
  input \u2_uk_K_r4_reg[38]/NET0131  ;
  input \u2_uk_K_r4_reg[39]/NET0131  ;
  input \u2_uk_K_r4_reg[3]/NET0131  ;
  input \u2_uk_K_r4_reg[40]/NET0131  ;
  input \u2_uk_K_r4_reg[41]/NET0131  ;
  input \u2_uk_K_r4_reg[42]/NET0131  ;
  input \u2_uk_K_r4_reg[43]/NET0131  ;
  input \u2_uk_K_r4_reg[44]/NET0131  ;
  input \u2_uk_K_r4_reg[45]/NET0131  ;
  input \u2_uk_K_r4_reg[46]/NET0131  ;
  input \u2_uk_K_r4_reg[47]/NET0131  ;
  input \u2_uk_K_r4_reg[48]/NET0131  ;
  input \u2_uk_K_r4_reg[49]/NET0131  ;
  input \u2_uk_K_r4_reg[4]/NET0131  ;
  input \u2_uk_K_r4_reg[50]/NET0131  ;
  input \u2_uk_K_r4_reg[51]/NET0131  ;
  input \u2_uk_K_r4_reg[52]/NET0131  ;
  input \u2_uk_K_r4_reg[53]/NET0131  ;
  input \u2_uk_K_r4_reg[54]/NET0131  ;
  input \u2_uk_K_r4_reg[55]/NET0131  ;
  input \u2_uk_K_r4_reg[5]/NET0131  ;
  input \u2_uk_K_r4_reg[6]/NET0131  ;
  input \u2_uk_K_r4_reg[7]/NET0131  ;
  input \u2_uk_K_r4_reg[8]/NET0131  ;
  input \u2_uk_K_r4_reg[9]/NET0131  ;
  input \u2_uk_K_r5_reg[0]/NET0131  ;
  input \u2_uk_K_r5_reg[10]/NET0131  ;
  input \u2_uk_K_r5_reg[11]/NET0131  ;
  input \u2_uk_K_r5_reg[12]/NET0131  ;
  input \u2_uk_K_r5_reg[13]/P0001  ;
  input \u2_uk_K_r5_reg[14]/NET0131  ;
  input \u2_uk_K_r5_reg[15]/NET0131  ;
  input \u2_uk_K_r5_reg[16]/NET0131  ;
  input \u2_uk_K_r5_reg[17]/NET0131  ;
  input \u2_uk_K_r5_reg[18]/NET0131  ;
  input \u2_uk_K_r5_reg[19]/NET0131  ;
  input \u2_uk_K_r5_reg[1]/NET0131  ;
  input \u2_uk_K_r5_reg[20]/NET0131  ;
  input \u2_uk_K_r5_reg[21]/NET0131  ;
  input \u2_uk_K_r5_reg[22]/NET0131  ;
  input \u2_uk_K_r5_reg[23]/NET0131  ;
  input \u2_uk_K_r5_reg[24]/NET0131  ;
  input \u2_uk_K_r5_reg[25]/NET0131  ;
  input \u2_uk_K_r5_reg[26]/NET0131  ;
  input \u2_uk_K_r5_reg[27]/NET0131  ;
  input \u2_uk_K_r5_reg[28]/NET0131  ;
  input \u2_uk_K_r5_reg[29]/NET0131  ;
  input \u2_uk_K_r5_reg[2]/NET0131  ;
  input \u2_uk_K_r5_reg[30]/NET0131  ;
  input \u2_uk_K_r5_reg[31]/NET0131  ;
  input \u2_uk_K_r5_reg[32]/NET0131  ;
  input \u2_uk_K_r5_reg[33]/NET0131  ;
  input \u2_uk_K_r5_reg[34]/NET0131  ;
  input \u2_uk_K_r5_reg[35]/NET0131  ;
  input \u2_uk_K_r5_reg[36]/NET0131  ;
  input \u2_uk_K_r5_reg[37]/P0001  ;
  input \u2_uk_K_r5_reg[38]/NET0131  ;
  input \u2_uk_K_r5_reg[39]/NET0131  ;
  input \u2_uk_K_r5_reg[3]/NET0131  ;
  input \u2_uk_K_r5_reg[40]/NET0131  ;
  input \u2_uk_K_r5_reg[41]/NET0131  ;
  input \u2_uk_K_r5_reg[42]/NET0131  ;
  input \u2_uk_K_r5_reg[43]/NET0131  ;
  input \u2_uk_K_r5_reg[44]/NET0131  ;
  input \u2_uk_K_r5_reg[46]/NET0131  ;
  input \u2_uk_K_r5_reg[47]/NET0131  ;
  input \u2_uk_K_r5_reg[48]/NET0131  ;
  input \u2_uk_K_r5_reg[49]/NET0131  ;
  input \u2_uk_K_r5_reg[4]/NET0131  ;
  input \u2_uk_K_r5_reg[50]/NET0131  ;
  input \u2_uk_K_r5_reg[51]/NET0131  ;
  input \u2_uk_K_r5_reg[52]/NET0131  ;
  input \u2_uk_K_r5_reg[53]/NET0131  ;
  input \u2_uk_K_r5_reg[54]/NET0131  ;
  input \u2_uk_K_r5_reg[55]/NET0131  ;
  input \u2_uk_K_r5_reg[5]/NET0131  ;
  input \u2_uk_K_r5_reg[6]/NET0131  ;
  input \u2_uk_K_r5_reg[7]/NET0131  ;
  input \u2_uk_K_r5_reg[8]/NET0131  ;
  input \u2_uk_K_r5_reg[9]/P0001  ;
  input \u2_uk_K_r6_reg[0]/NET0131  ;
  input \u2_uk_K_r6_reg[10]/NET0131  ;
  input \u2_uk_K_r6_reg[11]/NET0131  ;
  input \u2_uk_K_r6_reg[12]/NET0131  ;
  input \u2_uk_K_r6_reg[13]/NET0131  ;
  input \u2_uk_K_r6_reg[14]/NET0131  ;
  input \u2_uk_K_r6_reg[15]/NET0131  ;
  input \u2_uk_K_r6_reg[16]/NET0131  ;
  input \u2_uk_K_r6_reg[17]/NET0131  ;
  input \u2_uk_K_r6_reg[18]/NET0131  ;
  input \u2_uk_K_r6_reg[19]/NET0131  ;
  input \u2_uk_K_r6_reg[1]/NET0131  ;
  input \u2_uk_K_r6_reg[20]/NET0131  ;
  input \u2_uk_K_r6_reg[21]/NET0131  ;
  input \u2_uk_K_r6_reg[22]/NET0131  ;
  input \u2_uk_K_r6_reg[23]/P0001  ;
  input \u2_uk_K_r6_reg[24]/NET0131  ;
  input \u2_uk_K_r6_reg[25]/NET0131  ;
  input \u2_uk_K_r6_reg[26]/NET0131  ;
  input \u2_uk_K_r6_reg[27]/NET0131  ;
  input \u2_uk_K_r6_reg[28]/NET0131  ;
  input \u2_uk_K_r6_reg[29]/NET0131  ;
  input \u2_uk_K_r6_reg[2]/NET0131  ;
  input \u2_uk_K_r6_reg[30]/P0001  ;
  input \u2_uk_K_r6_reg[31]/NET0131  ;
  input \u2_uk_K_r6_reg[32]/NET0131  ;
  input \u2_uk_K_r6_reg[33]/NET0131  ;
  input \u2_uk_K_r6_reg[34]/NET0131  ;
  input \u2_uk_K_r6_reg[35]/NET0131  ;
  input \u2_uk_K_r6_reg[36]/NET0131  ;
  input \u2_uk_K_r6_reg[37]/NET0131  ;
  input \u2_uk_K_r6_reg[38]/NET0131  ;
  input \u2_uk_K_r6_reg[39]/NET0131  ;
  input \u2_uk_K_r6_reg[3]/NET0131  ;
  input \u2_uk_K_r6_reg[40]/NET0131  ;
  input \u2_uk_K_r6_reg[41]/NET0131  ;
  input \u2_uk_K_r6_reg[42]/NET0131  ;
  input \u2_uk_K_r6_reg[43]/NET0131  ;
  input \u2_uk_K_r6_reg[44]/NET0131  ;
  input \u2_uk_K_r6_reg[45]/NET0131  ;
  input \u2_uk_K_r6_reg[46]/NET0131  ;
  input \u2_uk_K_r6_reg[47]/NET0131  ;
  input \u2_uk_K_r6_reg[48]/NET0131  ;
  input \u2_uk_K_r6_reg[49]/NET0131  ;
  input \u2_uk_K_r6_reg[4]/NET0131  ;
  input \u2_uk_K_r6_reg[50]/NET0131  ;
  input \u2_uk_K_r6_reg[51]/NET0131  ;
  input \u2_uk_K_r6_reg[52]/NET0131  ;
  input \u2_uk_K_r6_reg[53]/NET0131  ;
  input \u2_uk_K_r6_reg[54]/NET0131  ;
  input \u2_uk_K_r6_reg[55]/P0001  ;
  input \u2_uk_K_r6_reg[5]/NET0131  ;
  input \u2_uk_K_r6_reg[6]/NET0131  ;
  input \u2_uk_K_r6_reg[7]/NET0131  ;
  input \u2_uk_K_r6_reg[8]/NET0131  ;
  input \u2_uk_K_r6_reg[9]/NET0131  ;
  input \u2_uk_K_r7_reg[0]/NET0131  ;
  input \u2_uk_K_r7_reg[10]/NET0131  ;
  input \u2_uk_K_r7_reg[11]/NET0131  ;
  input \u2_uk_K_r7_reg[12]/NET0131  ;
  input \u2_uk_K_r7_reg[13]/NET0131  ;
  input \u2_uk_K_r7_reg[14]/NET0131  ;
  input \u2_uk_K_r7_reg[15]/NET0131  ;
  input \u2_uk_K_r7_reg[16]/NET0131  ;
  input \u2_uk_K_r7_reg[17]/NET0131  ;
  input \u2_uk_K_r7_reg[18]/NET0131  ;
  input \u2_uk_K_r7_reg[19]/NET0131  ;
  input \u2_uk_K_r7_reg[1]/NET0131  ;
  input \u2_uk_K_r7_reg[20]/NET0131  ;
  input \u2_uk_K_r7_reg[21]/NET0131  ;
  input \u2_uk_K_r7_reg[22]/NET0131  ;
  input \u2_uk_K_r7_reg[23]/P0001  ;
  input \u2_uk_K_r7_reg[24]/NET0131  ;
  input \u2_uk_K_r7_reg[25]/NET0131  ;
  input \u2_uk_K_r7_reg[26]/NET0131  ;
  input \u2_uk_K_r7_reg[27]/NET0131  ;
  input \u2_uk_K_r7_reg[28]/NET0131  ;
  input \u2_uk_K_r7_reg[29]/NET0131  ;
  input \u2_uk_K_r7_reg[2]/NET0131  ;
  input \u2_uk_K_r7_reg[30]/P0001  ;
  input \u2_uk_K_r7_reg[31]/NET0131  ;
  input \u2_uk_K_r7_reg[32]/NET0131  ;
  input \u2_uk_K_r7_reg[33]/NET0131  ;
  input \u2_uk_K_r7_reg[34]/NET0131  ;
  input \u2_uk_K_r7_reg[35]/NET0131  ;
  input \u2_uk_K_r7_reg[36]/NET0131  ;
  input \u2_uk_K_r7_reg[37]/NET0131  ;
  input \u2_uk_K_r7_reg[38]/NET0131  ;
  input \u2_uk_K_r7_reg[39]/NET0131  ;
  input \u2_uk_K_r7_reg[3]/NET0131  ;
  input \u2_uk_K_r7_reg[40]/NET0131  ;
  input \u2_uk_K_r7_reg[41]/NET0131  ;
  input \u2_uk_K_r7_reg[42]/NET0131  ;
  input \u2_uk_K_r7_reg[43]/NET0131  ;
  input \u2_uk_K_r7_reg[44]/NET0131  ;
  input \u2_uk_K_r7_reg[45]/NET0131  ;
  input \u2_uk_K_r7_reg[46]/NET0131  ;
  input \u2_uk_K_r7_reg[47]/NET0131  ;
  input \u2_uk_K_r7_reg[48]/NET0131  ;
  input \u2_uk_K_r7_reg[49]/NET0131  ;
  input \u2_uk_K_r7_reg[4]/NET0131  ;
  input \u2_uk_K_r7_reg[50]/NET0131  ;
  input \u2_uk_K_r7_reg[51]/NET0131  ;
  input \u2_uk_K_r7_reg[52]/NET0131  ;
  input \u2_uk_K_r7_reg[53]/NET0131  ;
  input \u2_uk_K_r7_reg[54]/NET0131  ;
  input \u2_uk_K_r7_reg[55]/P0001  ;
  input \u2_uk_K_r7_reg[5]/NET0131  ;
  input \u2_uk_K_r7_reg[6]/NET0131  ;
  input \u2_uk_K_r7_reg[7]/NET0131  ;
  input \u2_uk_K_r7_reg[8]/NET0131  ;
  input \u2_uk_K_r7_reg[9]/NET0131  ;
  input \u2_uk_K_r8_reg[0]/NET0131  ;
  input \u2_uk_K_r8_reg[10]/NET0131  ;
  input \u2_uk_K_r8_reg[11]/NET0131  ;
  input \u2_uk_K_r8_reg[12]/NET0131  ;
  input \u2_uk_K_r8_reg[13]/P0001  ;
  input \u2_uk_K_r8_reg[14]/NET0131  ;
  input \u2_uk_K_r8_reg[15]/NET0131  ;
  input \u2_uk_K_r8_reg[16]/NET0131  ;
  input \u2_uk_K_r8_reg[17]/NET0131  ;
  input \u2_uk_K_r8_reg[18]/NET0131  ;
  input \u2_uk_K_r8_reg[19]/NET0131  ;
  input \u2_uk_K_r8_reg[1]/NET0131  ;
  input \u2_uk_K_r8_reg[20]/NET0131  ;
  input \u2_uk_K_r8_reg[21]/NET0131  ;
  input \u2_uk_K_r8_reg[22]/NET0131  ;
  input \u2_uk_K_r8_reg[23]/NET0131  ;
  input \u2_uk_K_r8_reg[24]/NET0131  ;
  input \u2_uk_K_r8_reg[25]/NET0131  ;
  input \u2_uk_K_r8_reg[26]/NET0131  ;
  input \u2_uk_K_r8_reg[27]/NET0131  ;
  input \u2_uk_K_r8_reg[28]/NET0131  ;
  input \u2_uk_K_r8_reg[29]/NET0131  ;
  input \u2_uk_K_r8_reg[2]/NET0131  ;
  input \u2_uk_K_r8_reg[30]/NET0131  ;
  input \u2_uk_K_r8_reg[31]/NET0131  ;
  input \u2_uk_K_r8_reg[32]/NET0131  ;
  input \u2_uk_K_r8_reg[33]/NET0131  ;
  input \u2_uk_K_r8_reg[34]/NET0131  ;
  input \u2_uk_K_r8_reg[35]/NET0131  ;
  input \u2_uk_K_r8_reg[36]/NET0131  ;
  input \u2_uk_K_r8_reg[37]/P0001  ;
  input \u2_uk_K_r8_reg[38]/NET0131  ;
  input \u2_uk_K_r8_reg[39]/NET0131  ;
  input \u2_uk_K_r8_reg[3]/NET0131  ;
  input \u2_uk_K_r8_reg[40]/NET0131  ;
  input \u2_uk_K_r8_reg[41]/NET0131  ;
  input \u2_uk_K_r8_reg[42]/NET0131  ;
  input \u2_uk_K_r8_reg[43]/NET0131  ;
  input \u2_uk_K_r8_reg[44]/NET0131  ;
  input \u2_uk_K_r8_reg[46]/NET0131  ;
  input \u2_uk_K_r8_reg[47]/NET0131  ;
  input \u2_uk_K_r8_reg[48]/NET0131  ;
  input \u2_uk_K_r8_reg[49]/NET0131  ;
  input \u2_uk_K_r8_reg[4]/NET0131  ;
  input \u2_uk_K_r8_reg[50]/NET0131  ;
  input \u2_uk_K_r8_reg[51]/NET0131  ;
  input \u2_uk_K_r8_reg[52]/NET0131  ;
  input \u2_uk_K_r8_reg[53]/NET0131  ;
  input \u2_uk_K_r8_reg[54]/NET0131  ;
  input \u2_uk_K_r8_reg[55]/NET0131  ;
  input \u2_uk_K_r8_reg[5]/NET0131  ;
  input \u2_uk_K_r8_reg[6]/NET0131  ;
  input \u2_uk_K_r8_reg[7]/NET0131  ;
  input \u2_uk_K_r8_reg[8]/NET0131  ;
  input \u2_uk_K_r8_reg[9]/NET0131  ;
  input \u2_uk_K_r9_reg[0]/P0001  ;
  input \u2_uk_K_r9_reg[10]/NET0131  ;
  input \u2_uk_K_r9_reg[11]/NET0131  ;
  input \u2_uk_K_r9_reg[12]/NET0131  ;
  input \u2_uk_K_r9_reg[13]/NET0131  ;
  input \u2_uk_K_r9_reg[14]/NET0131  ;
  input \u2_uk_K_r9_reg[15]/NET0131  ;
  input \u2_uk_K_r9_reg[16]/NET0131  ;
  input \u2_uk_K_r9_reg[17]/NET0131  ;
  input \u2_uk_K_r9_reg[18]/NET0131  ;
  input \u2_uk_K_r9_reg[19]/NET0131  ;
  input \u2_uk_K_r9_reg[1]/NET0131  ;
  input \u2_uk_K_r9_reg[20]/NET0131  ;
  input \u2_uk_K_r9_reg[21]/NET0131  ;
  input \u2_uk_K_r9_reg[22]/NET0131  ;
  input \u2_uk_K_r9_reg[23]/NET0131  ;
  input \u2_uk_K_r9_reg[25]/NET0131  ;
  input \u2_uk_K_r9_reg[26]/NET0131  ;
  input \u2_uk_K_r9_reg[27]/NET0131  ;
  input \u2_uk_K_r9_reg[28]/NET0131  ;
  input \u2_uk_K_r9_reg[29]/NET0131  ;
  input \u2_uk_K_r9_reg[30]/NET0131  ;
  input \u2_uk_K_r9_reg[31]/P0001  ;
  input \u2_uk_K_r9_reg[32]/NET0131  ;
  input \u2_uk_K_r9_reg[33]/NET0131  ;
  input \u2_uk_K_r9_reg[34]/NET0131  ;
  input \u2_uk_K_r9_reg[35]/NET0131  ;
  input \u2_uk_K_r9_reg[36]/NET0131  ;
  input \u2_uk_K_r9_reg[37]/NET0131  ;
  input \u2_uk_K_r9_reg[38]/NET0131  ;
  input \u2_uk_K_r9_reg[39]/NET0131  ;
  input \u2_uk_K_r9_reg[3]/NET0131  ;
  input \u2_uk_K_r9_reg[40]/NET0131  ;
  input \u2_uk_K_r9_reg[41]/NET0131  ;
  input \u2_uk_K_r9_reg[42]/NET0131  ;
  input \u2_uk_K_r9_reg[43]/NET0131  ;
  input \u2_uk_K_r9_reg[44]/NET0131  ;
  input \u2_uk_K_r9_reg[45]/NET0131  ;
  input \u2_uk_K_r9_reg[46]/NET0131  ;
  input \u2_uk_K_r9_reg[47]/NET0131  ;
  input \u2_uk_K_r9_reg[48]/NET0131  ;
  input \u2_uk_K_r9_reg[49]/NET0131  ;
  input \u2_uk_K_r9_reg[4]/NET0131  ;
  input \u2_uk_K_r9_reg[50]/NET0131  ;
  input \u2_uk_K_r9_reg[51]/NET0131  ;
  input \u2_uk_K_r9_reg[52]/NET0131  ;
  input \u2_uk_K_r9_reg[53]/NET0131  ;
  input \u2_uk_K_r9_reg[54]/NET0131  ;
  input \u2_uk_K_r9_reg[55]/NET0131  ;
  input \u2_uk_K_r9_reg[5]/NET0131  ;
  input \u2_uk_K_r9_reg[6]/NET0131  ;
  input \u2_uk_K_r9_reg[7]/NET0131  ;
  input \u2_uk_K_r9_reg[8]/NET0131  ;
  input \u2_uk_K_r9_reg[9]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g16/_0_  ;
  output \g191647/_3_  ;
  output \g191648/_3_  ;
  output \g191819/_3_  ;
  output \g191821/_0_  ;
  output \g191940/_3_  ;
  output \g191941/_0_  ;
  output \g191942/_0_  ;
  output \g191944/_0_  ;
  output \g191945/_0_  ;
  output \g191946/_0_  ;
  output \g191947/_3_  ;
  output \g191948/_0_  ;
  output \g191949/_0_  ;
  output \g191950/_0_  ;
  output \g191951/_3_  ;
  output \g191952/_0_  ;
  output \g192015/_3_  ;
  output \g192016/_3_  ;
  output \g192017/_3_  ;
  output \g192018/_3_  ;
  output \g192019/_3_  ;
  output \g192020/_0_  ;
  output \g192021/_3_  ;
  output \g192022/_0_  ;
  output \g192047/_0_  ;
  output \g192048/_0_  ;
  output \g192049/_0_  ;
  output \g192050/_0_  ;
  output \g192051/_0_  ;
  output \g192081/_0_  ;
  output \g193428/_3_  ;
  output \g193720/_0_  ;
  output \g193721/_0_  ;
  output \g193877/_0_  ;
  output \g193878/_0_  ;
  output \g193879/_0_  ;
  output \g193880/_3_  ;
  output \g193881/_0_  ;
  output \g193882/_0_  ;
  output \g193998/_0_  ;
  output \g193999/_0_  ;
  output \g194000/_3_  ;
  output \g194001/_0_  ;
  output \g194002/_0_  ;
  output \g194003/_0_  ;
  output \g194004/_0_  ;
  output \g194005/_0_  ;
  output \g194006/_0_  ;
  output \g194007/_0_  ;
  output \g194008/_0_  ;
  output \g194009/_0_  ;
  output \g194010/_0_  ;
  output \g194055/_3_  ;
  output \g194056/_3_  ;
  output \g194057/_0_  ;
  output \g194058/_0_  ;
  output \g194059/_0_  ;
  output \g194060/_0_  ;
  output \g194090/_0_  ;
  output \g194091/_0_  ;
  output \g194092/_0_  ;
  output \g194093/_0_  ;
  output \g195671/_0_  ;
  output \g195672/_3_  ;
  output \g195868/_0_  ;
  output \g195869/_0_  ;
  output \g195870/_0_  ;
  output \g196010/_0_  ;
  output \g196011/_0_  ;
  output \g196012/_0_  ;
  output \g196013/_0_  ;
  output \g196014/_0_  ;
  output \g196015/_0_  ;
  output \g196016/_0_  ;
  output \g196017/_0_  ;
  output \g196018/_0_  ;
  output \g196019/_3_  ;
  output \g196020/_0_  ;
  output \g196021/_0_  ;
  output \g196022/_0_  ;
  output \g196096/_3_  ;
  output \g196097/_0_  ;
  output \g196098/_0_  ;
  output \g196099/_0_  ;
  output \g196100/_3_  ;
  output \g196101/_0_  ;
  output \g196102/_0_  ;
  output \g196103/_0_  ;
  output \g196136/_0_  ;
  output \g196137/_0_  ;
  output \g196138/_0_  ;
  output \g196139/_0_  ;
  output \g196140/_0_  ;
  output \g196170/_0_  ;
  output \g197520/_3_  ;
  output \g197821/_0_  ;
  output \g197923/_0_  ;
  output \g197996/_0_  ;
  output \g197997/_3_  ;
  output \g197998/_0_  ;
  output \g197999/_0_  ;
  output \g198000/_0_  ;
  output \g198071/_0_  ;
  output \g198123/_0_  ;
  output \g198124/_0_  ;
  output \g198125/_0_  ;
  output \g198126/_0_  ;
  output \g198127/_0_  ;
  output \g198128/_0_  ;
  output \g198129/_0_  ;
  output \g198130/_0_  ;
  output \g198131/_0_  ;
  output \g198132/_0_  ;
  output \g198133/_0_  ;
  output \g198134/_3_  ;
  output \g198135/_0_  ;
  output \g198182/_0_  ;
  output \g198183/_3_  ;
  output \g198184/_0_  ;
  output \g198185/_0_  ;
  output \g198186/_0_  ;
  output \g198187/_0_  ;
  output \g198219/_0_  ;
  output \g198220/_0_  ;
  output \g198221/_0_  ;
  output \g198222/_0_  ;
  output \g199794/_0_  ;
  output \g199795/_3_  ;
  output \g200006/_0_  ;
  output \g200007/_0_  ;
  output \g200008/_0_  ;
  output \g200139/_0_  ;
  output \g200140/_0_  ;
  output \g200141/_0_  ;
  output \g200142/_0_  ;
  output \g200143/_0_  ;
  output \g200144/_0_  ;
  output \g200145/_0_  ;
  output \g200146/_0_  ;
  output \g200147/_0_  ;
  output \g200148/_0_  ;
  output \g200149/_0_  ;
  output \g200150/_3_  ;
  output \g200151/_0_  ;
  output \g200228/_3_  ;
  output \g200229/_0_  ;
  output \g200230/_0_  ;
  output \g200231/_0_  ;
  output \g200232/_3_  ;
  output \g200233/_0_  ;
  output \g200234/_0_  ;
  output \g200235/_0_  ;
  output \g200268/_0_  ;
  output \g200269/_0_  ;
  output \g200270/_0_  ;
  output \g200271/_0_  ;
  output \g200272/_0_  ;
  output \g200299/_0_  ;
  output \g201655/_3_  ;
  output \g201960/_0_  ;
  output \g201961/_0_  ;
  output \g202131/_0_  ;
  output \g202132/_0_  ;
  output \g202133/_3_  ;
  output \g202134/_0_  ;
  output \g202135/_0_  ;
  output \g202136/_0_  ;
  output \g202257/_0_  ;
  output \g202258/_0_  ;
  output \g202259/_3_  ;
  output \g202260/_0_  ;
  output \g202261/_0_  ;
  output \g202262/_0_  ;
  output \g202263/_0_  ;
  output \g202264/_0_  ;
  output \g202265/_0_  ;
  output \g202266/_0_  ;
  output \g202267/_0_  ;
  output \g202268/_0_  ;
  output \g202269/_0_  ;
  output \g202317/_0_  ;
  output \g202318/_3_  ;
  output \g202319/_0_  ;
  output \g202320/_0_  ;
  output \g202321/_0_  ;
  output \g202322/_0_  ;
  output \g202354/_0_  ;
  output \g202355/_0_  ;
  output \g202356/_0_  ;
  output \g202357/_0_  ;
  output \g203927/_0_  ;
  output \g203928/_3_  ;
  output \g204142/_0_  ;
  output \g204143/_0_  ;
  output \g204144/_0_  ;
  output \g204275/_0_  ;
  output \g204276/_0_  ;
  output \g204277/_0_  ;
  output \g204278/_0_  ;
  output \g204279/_0_  ;
  output \g204280/_0_  ;
  output \g204281/_0_  ;
  output \g204282/_0_  ;
  output \g204283/_0_  ;
  output \g204284/_0_  ;
  output \g204285/_0_  ;
  output \g204286/_3_  ;
  output \g204287/_0_  ;
  output \g204363/_3_  ;
  output \g204364/_0_  ;
  output \g204365/_0_  ;
  output \g204366/_0_  ;
  output \g204367/_3_  ;
  output \g204368/_0_  ;
  output \g204369/_0_  ;
  output \g204370/_0_  ;
  output \g204403/_0_  ;
  output \g204404/_0_  ;
  output \g204405/_0_  ;
  output \g204406/_0_  ;
  output \g204407/_0_  ;
  output \g204434/_0_  ;
  output \g205833/_3_  ;
  output \g206103/_0_  ;
  output \g206104/_0_  ;
  output \g206266/_0_  ;
  output \g206267/_0_  ;
  output \g206268/_0_  ;
  output \g206269/_3_  ;
  output \g206270/_0_  ;
  output \g206271/_0_  ;
  output \g206387/_0_  ;
  output \g206388/_0_  ;
  output \g206389/_3_  ;
  output \g206390/_0_  ;
  output \g206391/_0_  ;
  output \g206392/_0_  ;
  output \g206393/_0_  ;
  output \g206394/_0_  ;
  output \g206395/_0_  ;
  output \g206396/_0_  ;
  output \g206397/_0_  ;
  output \g206398/_0_  ;
  output \g206399/_0_  ;
  output \g206446/_0_  ;
  output \g206447/_3_  ;
  output \g206448/_0_  ;
  output \g206449/_0_  ;
  output \g206450/_0_  ;
  output \g206451/_0_  ;
  output \g206483/_0_  ;
  output \g206484/_0_  ;
  output \g206485/_0_  ;
  output \g206486/_0_  ;
  output \g208069/_0_  ;
  output \g208070/_3_  ;
  output \g208253/_0_  ;
  output \g208254/_0_  ;
  output \g208255/_0_  ;
  output \g208406/_0_  ;
  output \g208407/_0_  ;
  output \g208408/_0_  ;
  output \g208409/_0_  ;
  output \g208410/_0_  ;
  output \g208411/_0_  ;
  output \g208412/_0_  ;
  output \g208413/_0_  ;
  output \g208414/_0_  ;
  output \g208415/_3_  ;
  output \g208416/_0_  ;
  output \g208417/_0_  ;
  output \g208418/_0_  ;
  output \g208493/_3_  ;
  output \g208494/_0_  ;
  output \g208495/_0_  ;
  output \g208496/_0_  ;
  output \g208497/_3_  ;
  output \g208498/_0_  ;
  output \g208499/_0_  ;
  output \g208500/_0_  ;
  output \g208533/_0_  ;
  output \g208534/_0_  ;
  output \g208535/_0_  ;
  output \g208536/_0_  ;
  output \g208537/_0_  ;
  output \g208564/_0_  ;
  output \g209938/_3_  ;
  output \g210205/_0_  ;
  output \g210206/_0_  ;
  output \g210380/_0_  ;
  output \g210381/_0_  ;
  output \g210382/_0_  ;
  output \g210383/_3_  ;
  output \g210384/_0_  ;
  output \g210385/_0_  ;
  output \g210499/_0_  ;
  output \g210500/_0_  ;
  output \g210501/_3_  ;
  output \g210502/_0_  ;
  output \g210503/_0_  ;
  output \g210504/_0_  ;
  output \g210505/_0_  ;
  output \g210506/_0_  ;
  output \g210507/_0_  ;
  output \g210508/_0_  ;
  output \g210509/_0_  ;
  output \g210510/_0_  ;
  output \g210511/_0_  ;
  output \g210558/_0_  ;
  output \g210559/_3_  ;
  output \g210560/_0_  ;
  output \g210561/_0_  ;
  output \g210562/_0_  ;
  output \g210563/_0_  ;
  output \g210595/_0_  ;
  output \g210596/_0_  ;
  output \g210597/_0_  ;
  output \g210598/_0_  ;
  output \g212159/_0_  ;
  output \g212160/_3_  ;
  output \g212384/_0_  ;
  output \g212385/_0_  ;
  output \g212386/_0_  ;
  output \g212536/_0_  ;
  output \g212537/_0_  ;
  output \g212538/_0_  ;
  output \g212539/_0_  ;
  output \g212540/_0_  ;
  output \g212541/_0_  ;
  output \g212542/_0_  ;
  output \g212543/_0_  ;
  output \g212544/_0_  ;
  output \g212545/_0_  ;
  output \g212546/_3_  ;
  output \g212547/_0_  ;
  output \g212623/_3_  ;
  output \g212624/_0_  ;
  output \g212625/_0_  ;
  output \g212626/_0_  ;
  output \g212627/_0_  ;
  output \g212628/_3_  ;
  output \g212629/_0_  ;
  output \g212630/_0_  ;
  output \g212631/_0_  ;
  output \g212667/_0_  ;
  output \g212668/_0_  ;
  output \g212669/_0_  ;
  output \g212670/_0_  ;
  output \g212671/_0_  ;
  output \g212699/_0_  ;
  output \g214033/_3_  ;
  output \g214309/_3_  ;
  output \g214310/_0_  ;
  output \g214494/_0_  ;
  output \g214495/_0_  ;
  output \g214496/_0_  ;
  output \g214497/_3_  ;
  output \g214632/_0_  ;
  output \g214633/_0_  ;
  output \g214634/_3_  ;
  output \g214635/_0_  ;
  output \g214636/_0_  ;
  output \g214637/_0_  ;
  output \g214638/_0_  ;
  output \g214639/_0_  ;
  output \g214640/_0_  ;
  output \g214641/_0_  ;
  output \g214642/_0_  ;
  output \g214643/_0_  ;
  output \g214691/_0_  ;
  output \g214692/_0_  ;
  output \g214693/_3_  ;
  output \g214694/_0_  ;
  output \g214695/_0_  ;
  output \g214696/_0_  ;
  output \g214697/_0_  ;
  output \g214729/_0_  ;
  output \g214730/_0_  ;
  output \g214731/_0_  ;
  output \g214732/_0_  ;
  output \g214733/_0_  ;
  output \g216157/_0_  ;
  output \g216158/_3_  ;
  output \g216492/_0_  ;
  output \g216493/_0_  ;
  output \g216671/_0_  ;
  output \g216672/_0_  ;
  output \g216673/_0_  ;
  output \g216674/_0_  ;
  output \g216675/_0_  ;
  output \g216676/_3_  ;
  output \g216677/_0_  ;
  output \g216735/_0_  ;
  output \g216736/_3_  ;
  output \g216737/_0_  ;
  output \g216738/_0_  ;
  output \g216739/_0_  ;
  output \g216740/_0_  ;
  output \g216741/_0_  ;
  output \g216742/_0_  ;
  output \g216743/_0_  ;
  output \g216744/_0_  ;
  output \g216745/_0_  ;
  output \g216746/_3_  ;
  output \g216747/_0_  ;
  output \g216748/_0_  ;
  output \g216749/_0_  ;
  output \g216788/_0_  ;
  output \g216789/_0_  ;
  output \g216790/_0_  ;
  output \g216791/_0_  ;
  output \g216792/_0_  ;
  output \g216829/_0_  ;
  output \g218407/_3_  ;
  output \g218408/_0_  ;
  output \g218423/_3_  ;
  output \g218601/_0_  ;
  output \g218602/_0_  ;
  output \g218603/_0_  ;
  output \g218604/_0_  ;
  output \g218724/_0_  ;
  output \g218725/_0_  ;
  output \g218726/_0_  ;
  output \g218727/_0_  ;
  output \g218728/_0_  ;
  output \g218729/_0_  ;
  output \g218730/_0_  ;
  output \g218731/_0_  ;
  output \g218732/_0_  ;
  output \g218733/_0_  ;
  output \g218734/_0_  ;
  output \g218735/_3_  ;
  output \g218736/_0_  ;
  output \g218808/_3_  ;
  output \g218809/_0_  ;
  output \g218810/_0_  ;
  output \g218811/_3_  ;
  output \g218812/_0_  ;
  output \g218813/_0_  ;
  output \g218814/_0_  ;
  output \g218846/_0_  ;
  output \g218847/_0_  ;
  output \g218848/_0_  ;
  output \g218849/_0_  ;
  output \g218877/_0_  ;
  output \g22/_0_  ;
  output \g220545/_0_  ;
  output \g220546/_3_  ;
  output \g220725/_3_  ;
  output \g220726/_0_  ;
  output \g220793/_0_  ;
  output \g220794/_0_  ;
  output \g220795/_0_  ;
  output \g220796/_0_  ;
  output \g220797/_0_  ;
  output \g220798/_0_  ;
  output \g220799/_0_  ;
  output \g220800/_0_  ;
  output \g220801/_0_  ;
  output \g220802/_0_  ;
  output \g220803/_0_  ;
  output \g220804/_3_  ;
  output \g220805/_0_  ;
  output \g220806/_0_  ;
  output \g220807/_0_  ;
  output \g220872/_3_  ;
  output \g220873/_0_  ;
  output \g220874/_3_  ;
  output \g220875/_0_  ;
  output \g220876/_0_  ;
  output \g220877/_0_  ;
  output \g220921/_0_  ;
  output \g220922/_0_  ;
  output \g220923/_0_  ;
  output \g220924/_0_  ;
  output \g220925/_0_  ;
  output \g220926/_0_  ;
  output \g220969/_0_  ;
  output \g221011/_3_  ;
  output \g221039/_3_  ;
  output \g221086/_3_  ;
  output \g221131/_0_  ;
  output \g224010/_3_  ;
  output \g224368/_3_  ;
  output \g224369/_3_  ;
  output \g224532/_0_  ;
  output \g224533/_0_  ;
  output \g224534/_0_  ;
  output \g224535/_3_  ;
  output \g224536/_0_  ;
  output \g224537/_0_  ;
  output \g224640/_3_  ;
  output \g224641/_0_  ;
  output \g224642/_0_  ;
  output \g224643/_3_  ;
  output \g224644/_0_  ;
  output \g224645/_0_  ;
  output \g224646/_3_  ;
  output \g224647/_0_  ;
  output \g224648/_3_  ;
  output \g224649/_0_  ;
  output \g224650/_0_  ;
  output \g224651/_0_  ;
  output \g224652/_0_  ;
  output \g224690/_0_  ;
  output \g224691/_3_  ;
  output \g224692/_3_  ;
  output \g224693/_0_  ;
  output \g224694/_0_  ;
  output \g224695/_3_  ;
  output \g224723/_0_  ;
  output \g224724/_0_  ;
  output \g224725/_0_  ;
  output \g224726/_0_  ;
  output \g226372/_0_  ;
  output \g226373/_3_  ;
  output \g226549/_3_  ;
  output \g226550/_0_  ;
  output \g226616/_0_  ;
  output \g226635/_0_  ;
  output \g226636/_0_  ;
  output \g226637/_0_  ;
  output \g226638/_0_  ;
  output \g226639/_0_  ;
  output \g226640/_0_  ;
  output \g226641/_3_  ;
  output \g226642/_0_  ;
  output \g226643/_0_  ;
  output \g226644/_0_  ;
  output \g226645/_0_  ;
  output \g226646/_0_  ;
  output \g226692/_3_  ;
  output \g226693/_0_  ;
  output \g226694/_3_  ;
  output \g226695/_3_  ;
  output \g226696/_3_  ;
  output \g226697/_0_  ;
  output \g226698/_0_  ;
  output \g226699/_0_  ;
  output \g226728/_0_  ;
  output \g226729/_0_  ;
  output \g226730/_0_  ;
  output \g226731/_0_  ;
  output \g226732/_0_  ;
  output \g226759/_0_  ;
  output \g228250/_0_  ;
  output \g228396/_0_  ;
  output \g228397/_0_  ;
  output \g228566/_0_  ;
  output \g228567/_0_  ;
  output \g228568/_0_  ;
  output \g228609/_0_  ;
  output \g228610/_3_  ;
  output \g228688/_0_  ;
  output \g228689/_0_  ;
  output \g228690/_3_  ;
  output \g228691/_0_  ;
  output \g228692/_0_  ;
  output \g228693/_0_  ;
  output \g228694/_0_  ;
  output \g228695/_0_  ;
  output \g228696/_0_  ;
  output \g228697/_0_  ;
  output \g228698/_0_  ;
  output \g228699/_0_  ;
  output \g228700/_0_  ;
  output \g228748/_0_  ;
  output \g228749/_3_  ;
  output \g228750/_0_  ;
  output \g228751/_0_  ;
  output \g228752/_0_  ;
  output \g228753/_0_  ;
  output \g228784/_0_  ;
  output \g228785/_0_  ;
  output \g228786/_0_  ;
  output \g228787/_3_  ;
  output \g230339/_0_  ;
  output \g230340/_0_  ;
  output \g230546/_0_  ;
  output \g230580/_0_  ;
  output \g230679/_0_  ;
  output \g230680/_0_  ;
  output \g230681/_0_  ;
  output \g230682/_0_  ;
  output \g230683/_0_  ;
  output \g230684/_0_  ;
  output \g230685/_0_  ;
  output \g230686/_0_  ;
  output \g230687/_0_  ;
  output \g230688/_0_  ;
  output \g230689/_3_  ;
  output \g230690/_0_  ;
  output \g230710/_0_  ;
  output \g230766/_0_  ;
  output \g230767/_0_  ;
  output \g230768/_0_  ;
  output \g230769/_3_  ;
  output \g230770/_0_  ;
  output \g230771/_0_  ;
  output \g230772/_0_  ;
  output \g230773/_3_  ;
  output \g230810/_0_  ;
  output \g230811/_0_  ;
  output \g230812/_0_  ;
  output \g230813/_0_  ;
  output \g230814/_0_  ;
  output \g230840/_3_  ;
  output \g232196/_3_  ;
  output \g232469/_0_  ;
  output \g232470/_0_  ;
  output \g232633/_0_  ;
  output \g232635/_3_  ;
  output \g232636/_0_  ;
  output \g232637/_0_  ;
  output \g232691/_0_  ;
  output \g232747/_0_  ;
  output \g232748/_0_  ;
  output \g232749/_3_  ;
  output \g232750/_0_  ;
  output \g232751/_0_  ;
  output \g232752/_0_  ;
  output \g232753/_0_  ;
  output \g232754/_0_  ;
  output \g232755/_0_  ;
  output \g232756/_0_  ;
  output \g232757/_0_  ;
  output \g232758/_0_  ;
  output \g232759/_0_  ;
  output \g232804/_0_  ;
  output \g232805/_0_  ;
  output \g232806/_0_  ;
  output \g232807/_0_  ;
  output \g232808/_3_  ;
  output \g232809/_0_  ;
  output \g232841/_0_  ;
  output \g232842/_3_  ;
  output \g232843/_0_  ;
  output \g232844/_0_  ;
  output \g234520/_0_  ;
  output \g234687/_0_  ;
  output \g234688/_0_  ;
  output \g234689/_0_  ;
  output \g234764/_0_  ;
  output \g234765/_0_  ;
  output \g234766/_0_  ;
  output \g234767/_3_  ;
  output \g234768/_0_  ;
  output \g234769/_0_  ;
  output \g234770/_0_  ;
  output \g234771/_0_  ;
  output \g234772/_0_  ;
  output \g234773/_0_  ;
  output \g234774/_3_  ;
  output \g234775/_0_  ;
  output \g234776/_0_  ;
  output \g234824/_3_  ;
  output \g234825/_0_  ;
  output \g234826/_0_  ;
  output \g234827/_0_  ;
  output \g234828/_3_  ;
  output \g234829/_0_  ;
  output \g234830/_0_  ;
  output \g234831/_0_  ;
  output \g234867/_0_  ;
  output \g234868/_0_  ;
  output \g234869/_0_  ;
  output \g234870/_0_  ;
  output \g234896/_0_  ;
  output \g236294/_3_  ;
  output \g236541/_0_  ;
  output \g236542/_0_  ;
  output \g236724/_0_  ;
  output \g236725/_0_  ;
  output \g236726/_0_  ;
  output \g236727/_3_  ;
  output \g236728/_0_  ;
  output \g236729/_0_  ;
  output \g236821/_0_  ;
  output \g236822/_3_  ;
  output \g236823/_0_  ;
  output \g236824/_3_  ;
  output \g236825/_0_  ;
  output \g236826/_0_  ;
  output \g236827/_0_  ;
  output \g236828/_0_  ;
  output \g236829/_0_  ;
  output \g236830/_0_  ;
  output \g236831/_0_  ;
  output \g236832/_0_  ;
  output \g236877/_0_  ;
  output \g236878/_3_  ;
  output \g236879/_0_  ;
  output \g236880/_0_  ;
  output \g236881/_0_  ;
  output \g236882/_0_  ;
  output \g236914/_0_  ;
  output \g236915/_0_  ;
  output \g236916/_0_  ;
  output \g236917/_0_  ;
  output \g238530/_0_  ;
  output \g238531/_3_  ;
  output \g238723/_0_  ;
  output \g238724/_0_  ;
  output \g238725/_0_  ;
  output \g238840/_0_  ;
  output \g238841/_0_  ;
  output \g238842/_0_  ;
  output \g238843/_3_  ;
  output \g238844/_0_  ;
  output \g238845/_0_  ;
  output \g238846/_0_  ;
  output \g238847/_0_  ;
  output \g238848/_0_  ;
  output \g238849/_0_  ;
  output \g238850/_0_  ;
  output \g238851/_3_  ;
  output \g238852/_0_  ;
  output \g238924/_0_  ;
  output \g238925/_0_  ;
  output \g238926/_0_  ;
  output \g238927/_3_  ;
  output \g238928/_0_  ;
  output \g238929/_0_  ;
  output \g238930/_0_  ;
  output \g238965/_0_  ;
  output \g238966/_0_  ;
  output \g238967/_0_  ;
  output \g238968/_0_  ;
  output \g238969/_0_  ;
  output \g238996/_0_  ;
  output \g240353/_3_  ;
  output \g240640/_0_  ;
  output \g240641/_0_  ;
  output \g240813/_0_  ;
  output \g240814/_0_  ;
  output \g240815/_3_  ;
  output \g240816/_0_  ;
  output \g240817/_0_  ;
  output \g240818/_0_  ;
  output \g240925/_0_  ;
  output \g240926/_0_  ;
  output \g240927/_3_  ;
  output \g240928/_0_  ;
  output \g240929/_3_  ;
  output \g240930/_0_  ;
  output \g240931/_0_  ;
  output \g240932/_0_  ;
  output \g240933/_0_  ;
  output \g240934/_0_  ;
  output \g240935/_0_  ;
  output \g240936/_0_  ;
  output \g240937/_0_  ;
  output \g240984/_0_  ;
  output \g240985/_3_  ;
  output \g240986/_0_  ;
  output \g240987/_0_  ;
  output \g240988/_0_  ;
  output \g240989/_0_  ;
  output \g241021/_0_  ;
  output \g241022/_0_  ;
  output \g241023/_0_  ;
  output \g241024/_0_  ;
  output \g242616/_0_  ;
  output \g242617/_3_  ;
  output \g242815/_0_  ;
  output \g242816/_0_  ;
  output \g242817/_0_  ;
  output \g242955/_0_  ;
  output \g242956/_0_  ;
  output \g242957/_0_  ;
  output \g242958/_3_  ;
  output \g242959/_0_  ;
  output \g242960/_0_  ;
  output \g242961/_0_  ;
  output \g242962/_0_  ;
  output \g242963/_3_  ;
  output \g242964/_0_  ;
  output \g242965/_0_  ;
  output \g242966/_0_  ;
  output \g242967/_0_  ;
  output \g243037/_3_  ;
  output \g243038/_0_  ;
  output \g243039/_0_  ;
  output \g243040/_0_  ;
  output \g243041/_3_  ;
  output \g243042/_0_  ;
  output \g243043/_0_  ;
  output \g243044/_0_  ;
  output \g243078/_0_  ;
  output \g243079/_0_  ;
  output \g243080/_0_  ;
  output \g243081/_0_  ;
  output \g243082/_0_  ;
  output \g243109/_0_  ;
  output \g244465/_3_  ;
  output \g244753/_3_  ;
  output \g244754/_0_  ;
  output \g244924/_0_  ;
  output \g244925/_0_  ;
  output \g244926/_3_  ;
  output \g244927/_0_  ;
  output \g244928/_0_  ;
  output \g245035/_0_  ;
  output \g245036/_0_  ;
  output \g245037/_0_  ;
  output \g245038/_3_  ;
  output \g245039/_3_  ;
  output \g245040/_0_  ;
  output \g245041/_0_  ;
  output \g245043/_0_  ;
  output \g245045/_0_  ;
  output \g245046/_0_  ;
  output \g245047/_0_  ;
  output \g245092/_0_  ;
  output \g245093/_3_  ;
  output \g245094/_0_  ;
  output \g245095/_0_  ;
  output \g245096/_0_  ;
  output \g245097/_0_  ;
  output \g245129/_0_  ;
  output \g245130/_0_  ;
  output \g245131/_0_  ;
  output \g245132/_0_  ;
  output \g246715/_0_  ;
  output \g246716/_3_  ;
  output \g246911/_0_  ;
  output \g246912/_0_  ;
  output \g246913/_0_  ;
  output \g247057/_0_  ;
  output \g247058/_0_  ;
  output \g247059/_0_  ;
  output \g247060/_0_  ;
  output \g247061/_0_  ;
  output \g247062/_3_  ;
  output \g247063/_0_  ;
  output \g247064/_0_  ;
  output \g247065/_0_  ;
  output \g247066/_0_  ;
  output \g247067/_3_  ;
  output \g247068/_0_  ;
  output \g247069/_0_  ;
  output \g247137/_3_  ;
  output \g247138/_0_  ;
  output \g247139/_0_  ;
  output \g247140/_0_  ;
  output \g247141/_3_  ;
  output \g247142/_0_  ;
  output \g247143/_0_  ;
  output \g247144/_0_  ;
  output \g247179/_0_  ;
  output \g247180/_0_  ;
  output \g247181/_0_  ;
  output \g247182/_0_  ;
  output \g247183/_0_  ;
  output \g247210/_0_  ;
  output \g248581/_3_  ;
  output \g248828/_0_  ;
  output \g248829/_0_  ;
  output \g249033/_0_  ;
  output \g249035/_0_  ;
  output \g249036/_3_  ;
  output \g249037/_0_  ;
  output \g249038/_0_  ;
  output \g249147/_0_  ;
  output \g249148/_0_  ;
  output \g249149/_3_  ;
  output \g249150/_0_  ;
  output \g249152/_0_  ;
  output \g249153/_0_  ;
  output \g249155/_0_  ;
  output \g249156/_0_  ;
  output \g249157/_0_  ;
  output \g249200/_3_  ;
  output \g249201/_0_  ;
  output \g249202/_0_  ;
  output \g249203/_3_  ;
  output \g249204/_0_  ;
  output \g249205/_0_  ;
  output \g249206/_0_  ;
  output \g249207/_0_  ;
  output \g249239/_0_  ;
  output \g249240/_0_  ;
  output \g249241/_0_  ;
  output \g249242/_0_  ;
  output \g250815/_0_  ;
  output \g251006/_0_  ;
  output \g251007/_0_  ;
  output \g251008/_0_  ;
  output \g251009/_3_  ;
  output \g251160/_0_  ;
  output \g251161/_0_  ;
  output \g251162/_0_  ;
  output \g251163/_3_  ;
  output \g251164/_0_  ;
  output \g251165/_0_  ;
  output \g251166/_0_  ;
  output \g251167/_0_  ;
  output \g251168/_0_  ;
  output \g251169/_0_  ;
  output \g251170/_3_  ;
  output \g251171/_0_  ;
  output \g251245/_3_  ;
  output \g251246/_0_  ;
  output \g251247/_0_  ;
  output \g251248/_0_  ;
  output \g251249/_3_  ;
  output \g251250/_0_  ;
  output \g251251/_0_  ;
  output \g251252/_0_  ;
  output \g251286/_0_  ;
  output \g251287/_0_  ;
  output \g251288/_0_  ;
  output \g251289/_0_  ;
  output \g251290/_0_  ;
  output \g251291/_0_  ;
  output \g251318/_0_  ;
  output \g252698/_3_  ;
  output \g252942/_0_  ;
  output \g252943/_0_  ;
  output \g253118/_0_  ;
  output \g253119/_0_  ;
  output \g253120/_0_  ;
  output \g253121/_0_  ;
  output \g253122/_3_  ;
  output \g253123/_0_  ;
  output \g253236/_0_  ;
  output \g253237/_3_  ;
  output \g253238/_3_  ;
  output \g253239/_0_  ;
  output \g253240/_0_  ;
  output \g253241/_0_  ;
  output \g253242/_0_  ;
  output \g253243/_0_  ;
  output \g253244/_0_  ;
  output \g253245/_0_  ;
  output \g253246/_0_  ;
  output \g253247/_0_  ;
  output \g253248/_0_  ;
  output \g253306/_0_  ;
  output \g253307/_3_  ;
  output \g253308/_0_  ;
  output \g253309/_0_  ;
  output \g253310/_0_  ;
  output \g253311/_0_  ;
  output \g253356/_0_  ;
  output \g253357/_0_  ;
  output \g253358/_0_  ;
  output \g253359/_0_  ;
  output \g253436/_3_  ;
  output \g253437/_0_  ;
  output \g253438/_0_  ;
  output \g253469/_3_  ;
  output \g253470/_3_  ;
  output \g253471/_3_  ;
  output \g253521/_0_  ;
  output \g253522/_0_  ;
  output \g253523/_0_  ;
  output \g253524/_3_  ;
  output \g256730/_3_  ;
  output \g256731/_3_  ;
  output \g256927/_0_  ;
  output \g256928/_0_  ;
  output \g256929/_3_  ;
  output \g257049/_0_  ;
  output \g257050/_0_  ;
  output \g257051/_3_  ;
  output \g257052/_0_  ;
  output \g257053/_0_  ;
  output \g257054/_0_  ;
  output \g257055/_3_  ;
  output \g257056/_0_  ;
  output \g257057/_0_  ;
  output \g257058/_3_  ;
  output \g257059/_0_  ;
  output \g257060/_0_  ;
  output \g257082/_0_  ;
  output \g257125/_3_  ;
  output \g257126/_0_  ;
  output \g257127/_0_  ;
  output \g257128/_3_  ;
  output \g257129/_3_  ;
  output \g257130/_0_  ;
  output \g257131/_0_  ;
  output \g257132/_0_  ;
  output \g257163/_0_  ;
  output \g257164/_0_  ;
  output \g257165/_0_  ;
  output \g257166/_0_  ;
  output \g257167/_0_  ;
  output \g257194/_0_  ;
  output \g258552/_0_  ;
  output \g258850/_0_  ;
  output \g258851/_3_  ;
  output \g258993/_0_  ;
  output \g258994/_0_  ;
  output \g258995/_0_  ;
  output \g258996/_0_  ;
  output \g259026/_3_  ;
  output \g259027/_0_  ;
  output \g259105/_0_  ;
  output \g259106/_0_  ;
  output \g259107/_3_  ;
  output \g259108/_0_  ;
  output \g259109/_3_  ;
  output \g259110/_0_  ;
  output \g259111/_0_  ;
  output \g259112/_0_  ;
  output \g259113/_0_  ;
  output \g259114/_0_  ;
  output \g259115/_0_  ;
  output \g259116/_0_  ;
  output \g259117/_0_  ;
  output \g259163/_3_  ;
  output \g259164/_3_  ;
  output \g259165/_0_  ;
  output \g259166/_0_  ;
  output \g259167/_0_  ;
  output \g259168/_0_  ;
  output \g259197/_0_  ;
  output \g259198/_0_  ;
  output \g259199/_0_  ;
  output \g259200/_0_  ;
  output \g260774/_0_  ;
  output \g260792/_3_  ;
  output \g260991/_0_  ;
  output \g261013/_0_  ;
  output \g261070/_0_  ;
  output \g261125/_0_  ;
  output \g261126/_0_  ;
  output \g261128/_0_  ;
  output \g261129/_0_  ;
  output \g261130/_0_  ;
  output \g261131/_0_  ;
  output \g261132/_0_  ;
  output \g261133/_0_  ;
  output \g261134/_3_  ;
  output \g261135/_0_  ;
  output \g261136/_0_  ;
  output \g261158/_3_  ;
  output \g261206/_0_  ;
  output \g261207/_0_  ;
  output \g261208/_0_  ;
  output \g261209/_0_  ;
  output \g261210/_3_  ;
  output \g261211/_0_  ;
  output \g261212/_3_  ;
  output \g261213/_0_  ;
  output \g261248/_0_  ;
  output \g261249/_0_  ;
  output \g261250/_0_  ;
  output \g261251/_0_  ;
  output \g261252/_0_  ;
  output \g261279/_0_  ;
  output \g262658/_3_  ;
  output \g262949/_0_  ;
  output \g263008/_3_  ;
  output \g263092/_0_  ;
  output \g263093/_0_  ;
  output \g263099/_0_  ;
  output \g263100/_0_  ;
  output \g263101/_0_  ;
  output \g263159/_3_  ;
  output \g263204/_3_  ;
  output \g263205/_0_  ;
  output \g263206/_0_  ;
  output \g263208/_0_  ;
  output \g263209/_0_  ;
  output \g263210/_0_  ;
  output \g263211/_0_  ;
  output \g263212/_0_  ;
  output \g263213/_0_  ;
  output \g263214/_0_  ;
  output \g263215/_3_  ;
  output \g263216/_0_  ;
  output \g263260/_0_  ;
  output \g263261/_0_  ;
  output \g263262/_3_  ;
  output \g263263/_0_  ;
  output \g263264/_0_  ;
  output \g263265/_0_  ;
  output \g263297/_0_  ;
  output \g263298/_0_  ;
  output \g263299/_0_  ;
  output \g263300/_0_  ;
  output \g264930/_0_  ;
  output \g264946/_3_  ;
  output \g265143/_0_  ;
  output \g265144/_0_  ;
  output \g265152/_0_  ;
  output \g265222/_0_  ;
  output \g265223/_0_  ;
  output \g265224/_0_  ;
  output \g265225/_0_  ;
  output \g265226/_0_  ;
  output \g265227/_3_  ;
  output \g265228/_0_  ;
  output \g265229/_0_  ;
  output \g265230/_0_  ;
  output \g265231/_0_  ;
  output \g265232/_0_  ;
  output \g265233/_3_  ;
  output \g265234/_0_  ;
  output \g265306/_0_  ;
  output \g265307/_0_  ;
  output \g265308/_3_  ;
  output \g265309/_3_  ;
  output \g265310/_0_  ;
  output \g265311/_0_  ;
  output \g265312/_0_  ;
  output \g265313/_0_  ;
  output \g265348/_0_  ;
  output \g265349/_0_  ;
  output \g265350/_0_  ;
  output \g265351/_0_  ;
  output \g265379/_0_  ;
  output \g266965/_3_  ;
  output \g267049/_3_  ;
  output \g267050/_0_  ;
  output \g267215/_0_  ;
  output \g267216/_0_  ;
  output \g267263/_0_  ;
  output \g267264/_3_  ;
  output \g267265/_0_  ;
  output \g267266/_0_  ;
  output \g267314/_3_  ;
  output \g267315/_0_  ;
  output \g267316/_0_  ;
  output \g267317/_0_  ;
  output \g267318/_0_  ;
  output \g267319/_0_  ;
  output \g267320/_3_  ;
  output \g267321/_0_  ;
  output \g267322/_0_  ;
  output \g267324/_0_  ;
  output \g267325/_0_  ;
  output \g267326/_0_  ;
  output \g267372/_0_  ;
  output \g267373/_3_  ;
  output \g267374/_0_  ;
  output \g267375/_0_  ;
  output \g267376/_0_  ;
  output \g267377/_0_  ;
  output \g267409/_0_  ;
  output \g267410/_0_  ;
  output \g267411/_0_  ;
  output \g267412/_0_  ;
  output \g269004/_0_  ;
  output \g269099/_3_  ;
  output \g269202/_0_  ;
  output \g269226/_0_  ;
  output \g269333/_3_  ;
  output \g269334/_0_  ;
  output \g269335/_0_  ;
  output \g269355/_0_  ;
  output \g269356/_0_  ;
  output \g269357/_3_  ;
  output \g269358/_0_  ;
  output \g269359/_0_  ;
  output \g269360/_0_  ;
  output \g269361/_0_  ;
  output \g269362/_0_  ;
  output \g269363/_0_  ;
  output \g269364/_0_  ;
  output \g269414/_0_  ;
  output \g269415/_0_  ;
  output \g269416/_0_  ;
  output \g269417/_0_  ;
  output \g269418/_3_  ;
  output \g269419/_0_  ;
  output \g269420/_3_  ;
  output \g269421/_0_  ;
  output \g269456/_0_  ;
  output \g269457/_0_  ;
  output \g269458/_0_  ;
  output \g269459/_0_  ;
  output \g269460/_0_  ;
  output \g269487/_0_  ;
  output \g271006/_3_  ;
  output \g271186/_3_  ;
  output \g271187/_0_  ;
  output \g271299/_0_  ;
  output \g271300/_0_  ;
  output \g271301/_3_  ;
  output \g271302/_0_  ;
  output \g271303/_0_  ;
  output \g271352/_0_  ;
  output \g271410/_0_  ;
  output \g271411/_0_  ;
  output \g271412/_0_  ;
  output \g271413/_0_  ;
  output \g271414/_0_  ;
  output \g271415/_0_  ;
  output \g271416/_0_  ;
  output \g271417/_3_  ;
  output \g271418/_3_  ;
  output \g271419/_0_  ;
  output \g271420/_0_  ;
  output \g271421/_0_  ;
  output \g271422/_0_  ;
  output \g271468/_3_  ;
  output \g271469/_0_  ;
  output \g271470/_0_  ;
  output \g271471/_0_  ;
  output \g271472/_0_  ;
  output \g271473/_0_  ;
  output \g271505/_0_  ;
  output \g271506/_0_  ;
  output \g271507/_0_  ;
  output \g271508/_0_  ;
  output \g273135/_0_  ;
  output \g273136/_3_  ;
  output \g273362/_0_  ;
  output \g273373/_0_  ;
  output \g273374/_0_  ;
  output \g273431/_0_  ;
  output \g273432/_0_  ;
  output \g273433/_3_  ;
  output \g273434/_0_  ;
  output \g273435/_0_  ;
  output \g273436/_0_  ;
  output \g273437/_3_  ;
  output \g273438/_0_  ;
  output \g273439/_0_  ;
  output \g273441/_0_  ;
  output \g273442/_0_  ;
  output \g273443/_0_  ;
  output \g273515/_3_  ;
  output \g273516/_0_  ;
  output \g273517/_0_  ;
  output \g273518/_3_  ;
  output \g273519/_0_  ;
  output \g273520/_0_  ;
  output \g273521/_0_  ;
  output \g273522/_0_  ;
  output \g273557/_0_  ;
  output \g273558/_0_  ;
  output \g273559/_0_  ;
  output \g273560/_0_  ;
  output \g273561/_0_  ;
  output \g273588/_0_  ;
  output \g274960/_3_  ;
  output \g275266/_3_  ;
  output \g275327/_0_  ;
  output \g275396/_0_  ;
  output \g275397/_3_  ;
  output \g275398/_0_  ;
  output \g275455/_0_  ;
  output \g275456/_0_  ;
  output \g275463/_0_  ;
  output \g275510/_3_  ;
  output \g275511/_0_  ;
  output \g275512/_0_  ;
  output \g275513/_0_  ;
  output \g275514/_3_  ;
  output \g275515/_0_  ;
  output \g275516/_0_  ;
  output \g275517/_0_  ;
  output \g275518/_0_  ;
  output \g275519/_0_  ;
  output \g275520/_0_  ;
  output \g275521/_0_  ;
  output \g275522/_0_  ;
  output \g275568/_0_  ;
  output \g275569/_0_  ;
  output \g275570/_0_  ;
  output \g275571/_0_  ;
  output \g275572/_3_  ;
  output \g275573/_0_  ;
  output \g275605/_0_  ;
  output \g275606/_0_  ;
  output \g275607/_0_  ;
  output \g275608/_0_  ;
  output \g277189/_0_  ;
  output \g277294/_3_  ;
  output \g277367/_0_  ;
  output \g277456/_0_  ;
  output \g277457/_0_  ;
  output \g277512/_0_  ;
  output \g277513/_0_  ;
  output \g277514/_3_  ;
  output \g277515/_0_  ;
  output \g277516/_0_  ;
  output \g277517/_3_  ;
  output \g277518/_0_  ;
  output \g277519/_0_  ;
  output \g277520/_0_  ;
  output \g277521/_0_  ;
  output \g277594/_0_  ;
  output \g277595/_0_  ;
  output \g277596/_3_  ;
  output \g277597/_0_  ;
  output \g277598/_0_  ;
  output \g277599/_0_  ;
  output \g277600/_0_  ;
  output \g277601/_3_  ;
  output \g277635/_0_  ;
  output \g277636/_0_  ;
  output \g277637/_0_  ;
  output \g277638/_0_  ;
  output \g277639/_0_  ;
  output \g277666/_0_  ;
  output \g279090/_3_  ;
  output \g279330/_0_  ;
  output \g279331/_0_  ;
  output \g279493/_3_  ;
  output \g279494/_0_  ;
  output \g279495/_0_  ;
  output \g279502/_0_  ;
  output \g279503/_0_  ;
  output \g279504/_0_  ;
  output \g279590/_0_  ;
  output \g279591/_0_  ;
  output \g279592/_0_  ;
  output \g279593/_0_  ;
  output \g279594/_3_  ;
  output \g279595/_3_  ;
  output \g279596/_0_  ;
  output \g279597/_0_  ;
  output \g279598/_0_  ;
  output \g279599/_0_  ;
  output \g279600/_0_  ;
  output \g279601/_0_  ;
  output \g279602/_0_  ;
  output \g279649/_0_  ;
  output \g279650/_0_  ;
  output \g279651/_0_  ;
  output \g279652/_0_  ;
  output \g279653/_0_  ;
  output \g279654/_3_  ;
  output \g279686/_0_  ;
  output \g279687/_0_  ;
  output \g279688/_0_  ;
  output \g279689/_0_  ;
  output \g281329/_0_  ;
  output \g281394/_0_  ;
  output \g281483/_0_  ;
  output \g281498/_0_  ;
  output \g281532/_0_  ;
  output \g281616/_0_  ;
  output \g281617/_0_  ;
  output \g281618/_0_  ;
  output \g281619/_0_  ;
  output \g281620/_0_  ;
  output \g281621/_0_  ;
  output \g281622/_0_  ;
  output \g281623/_3_  ;
  output \g281624/_0_  ;
  output \g281642/_0_  ;
  output \g281643/_0_  ;
  output \g281644/_3_  ;
  output \g281645/_0_  ;
  output \g281696/_0_  ;
  output \g281697/_3_  ;
  output \g281698/_0_  ;
  output \g281699/_0_  ;
  output \g281700/_0_  ;
  output \g281701/_0_  ;
  output \g281702/_3_  ;
  output \g281703/_0_  ;
  output \g281799/_0_  ;
  output \g281800/_0_  ;
  output \g281801/_0_  ;
  output \g281802/_0_  ;
  output \g281803/_0_  ;
  output \g281965/_0_  ;
  output \g287377/_0_  ;
  output \g287867/_0_  ;
  output \g287899/_0_  ;
  output \g288304/_0_  ;
  output \g288334/_0_  ;
  output \g288350/_0_  ;
  output \g288351/_0_  ;
  output \g288352/_3_  ;
  output \g288353/_0_  ;
  output \g288668/_0_  ;
  output \g288669/_0_  ;
  output \g288670/_0_  ;
  output \g288671/_0_  ;
  output \g288673/_0_  ;
  output \g288674/_3_  ;
  output \g288675/_0_  ;
  output \g288676/_0_  ;
  output \g288677/_0_  ;
  output \g288678/_0_  ;
  output \g288679/_0_  ;
  output \g288680/_3_  ;
  output \g288889/_0_  ;
  output \g288890/_0_  ;
  output \g288891/_0_  ;
  output \g288892/_0_  ;
  output \g288893/_3_  ;
  output \g288894/_0_  ;
  output \g288895/_0_  ;
  output \g288984/_0_  ;
  output \g288985/_0_  ;
  output \g288986/_0_  ;
  output \g294974/_0_  ;
  output \g295054/_0_  ;
  output \g295601/_0_  ;
  output \g295607/_0_  ;
  output \g296036/_0_  ;
  output \g296037/_0_  ;
  output \g296038/_0_  ;
  output \g296039/_0_  ;
  output \g296040/_0_  ;
  output \g296041/_0_  ;
  output \g296042/_0_  ;
  output \g296043/_3_  ;
  output \g296044/_0_  ;
  output \g296045/_0_  ;
  output \g296046/_0_  ;
  output \g296047/_0_  ;
  output \g296048/_0_  ;
  output \g296049/_3_  ;
  output \g296522/_3_  ;
  output \g296523/_3_  ;
  output \g296524/_0_  ;
  output \g296525/_0_  ;
  output \g296526/_0_  ;
  output \g296527/_0_  ;
  output \g296528/_3_  ;
  output \g296529/_0_  ;
  output \g296530/_0_  ;
  output \g296531/_0_  ;
  output \g297026/_0_  ;
  output \g297027/_0_  ;
  output \g305620/_3_  ;
  output \g305621/_3_  ;
  output \g305622/_3_  ;
  output \g305623/_3_  ;
  output \g305624/_3_  ;
  output \g305625/_3_  ;
  output \g305626/_3_  ;
  output \g305627/_3_  ;
  output \g305628/_3_  ;
  output \g305629/_3_  ;
  output \g305630/_3_  ;
  output \g305631/_3_  ;
  output \g305632/_3_  ;
  output \g305633/_3_  ;
  output \g305634/_3_  ;
  output \g305635/_3_  ;
  output \g305636/_3_  ;
  output \g305637/_3_  ;
  output \g305638/_3_  ;
  output \g305639/_3_  ;
  output \g305640/_3_  ;
  output \g305641/_3_  ;
  output \g305642/_3_  ;
  output \g305643/_3_  ;
  output \g305644/_3_  ;
  output \g305645/_3_  ;
  output \g305646/_3_  ;
  output \g305647/_3_  ;
  output \g305648/_3_  ;
  output \g305649/_3_  ;
  output \g305650/_3_  ;
  output \g305651/_3_  ;
  output \g305652/_3_  ;
  output \g305653/_3_  ;
  output \g305654/_3_  ;
  output \g305655/_3_  ;
  output \g305656/_3_  ;
  output \g305657/_3_  ;
  output \g305658/_3_  ;
  output \g305659/_3_  ;
  output \g305660/_3_  ;
  output \g305661/_3_  ;
  output \g305662/_3_  ;
  output \g305663/_3_  ;
  output \g305664/_3_  ;
  output \g305665/_3_  ;
  output \g305666/_3_  ;
  output \g305667/_3_  ;
  output \g305668/_3_  ;
  output \g305669/_3_  ;
  output \g305670/_3_  ;
  output \g305671/_3_  ;
  output \g305672/_3_  ;
  output \g305673/_3_  ;
  output \g305674/_3_  ;
  output \g305675/_3_  ;
  output \g305676/_3_  ;
  output \g305677/_3_  ;
  output \g305678/_3_  ;
  output \g305679/_3_  ;
  output \g305680/_3_  ;
  output \g305681/_3_  ;
  output \g305682/_3_  ;
  output \g305683/_3_  ;
  output \g305684/_3_  ;
  output \g305685/_3_  ;
  output \g305686/_3_  ;
  output \g305687/_3_  ;
  output \g305688/_3_  ;
  output \g305689/_3_  ;
  output \g305690/_3_  ;
  output \g305691/_3_  ;
  output \g305692/_3_  ;
  output \g305693/_3_  ;
  output \g305694/_3_  ;
  output \g305695/_3_  ;
  output \g305696/_3_  ;
  output \g305697/_3_  ;
  output \g305698/_3_  ;
  output \g305699/_3_  ;
  output \g305700/_3_  ;
  output \g305701/_3_  ;
  output \g305702/_3_  ;
  output \g305703/_3_  ;
  output \g305704/_3_  ;
  output \g305705/_3_  ;
  output \g305706/_3_  ;
  output \g305707/_3_  ;
  output \g305708/_3_  ;
  output \g305709/_3_  ;
  output \g305710/_3_  ;
  output \g305711/_3_  ;
  output \g305712/_3_  ;
  output \g305713/_3_  ;
  output \g305714/_3_  ;
  output \g305715/_3_  ;
  output \g305716/_3_  ;
  output \g305717/_3_  ;
  output \g305718/_3_  ;
  output \g305719/_3_  ;
  output \g305720/_3_  ;
  output \g305721/_3_  ;
  output \g305722/_3_  ;
  output \g305723/_3_  ;
  output \g305724/_3_  ;
  output \g305725/_3_  ;
  output \g305726/_3_  ;
  output \g305727/_3_  ;
  output \g305728/_3_  ;
  output \g305729/_3_  ;
  output \g305730/_3_  ;
  output \g305731/_3_  ;
  output \g321371/_0_  ;
  output \g321424/_0_  ;
  output \g321474/_3_  ;
  output \g321637/_3_  ;
  output \g321688/_0_  ;
  output \g321712/_0_  ;
  output \g321772/_3_  ;
  output \g321832/_0_  ;
  output \g321999/_0_  ;
  output \g322013/_3_  ;
  output \g322109/_0_  ;
  output \g322184/_0_  ;
  output \g322250/_0_  ;
  output \g322274/_0_  ;
  output \g322293/_3_  ;
  output \g322437/_0_  ;
  output \g322537/_3_  ;
  output \g322584/_0_  ;
  output \g322830/_0_  ;
  output \g322871/_0_  ;
  output \g322882/_0_  ;
  output \g322933/_0_  ;
  output \g323004/_0_  ;
  output \g323104/_0_  ;
  output \g323125/_0_  ;
  output \g323138/_3_  ;
  output \g323273/_0_  ;
  output \u0_desOut_reg[0]/_05_  ;
  output \u0_desOut_reg[12]/_05_  ;
  output \u0_desOut_reg[14]/_05_  ;
  output \u0_desOut_reg[18]/_05_  ;
  output \u0_desOut_reg[20]/_05_  ;
  output \u0_desOut_reg[24]/_05_  ;
  output \u0_desOut_reg[26]/_05_  ;
  output \u0_desOut_reg[28]/_05_  ;
  output \u0_desOut_reg[2]/_05_  ;
  output \u0_desOut_reg[30]/_05_  ;
  output \u0_desOut_reg[32]/_05_  ;
  output \u0_desOut_reg[34]/_05_  ;
  output \u0_desOut_reg[36]/_05_  ;
  output \u0_desOut_reg[42]/_05_  ;
  output \u0_desOut_reg[44]/_05_  ;
  output \u0_desOut_reg[46]/_05_  ;
  output \u0_desOut_reg[48]/_05_  ;
  output \u0_desOut_reg[54]/_05_  ;
  output \u0_desOut_reg[56]/_05_  ;
  output \u0_desOut_reg[62]/_05_  ;
  output \u0_desOut_reg[6]/_05_  ;
  output \u0_desOut_reg[8]/_05_  ;
  output \u1_desOut_reg[0]/_05_  ;
  output \u1_desOut_reg[12]/_05_  ;
  output \u1_desOut_reg[14]/_05_  ;
  output \u1_desOut_reg[16]/_05_  ;
  output \u1_desOut_reg[18]/_05_  ;
  output \u1_desOut_reg[20]/_05_  ;
  output \u1_desOut_reg[22]/_05_  ;
  output \u1_desOut_reg[24]/_05_  ;
  output \u1_desOut_reg[26]/_05_  ;
  output \u1_desOut_reg[28]/_05_  ;
  output \u1_desOut_reg[2]/_05_  ;
  output \u1_desOut_reg[30]/_05_  ;
  output \u1_desOut_reg[32]/_05_  ;
  output \u1_desOut_reg[34]/_05_  ;
  output \u1_desOut_reg[36]/_05_  ;
  output \u1_desOut_reg[38]/_05_  ;
  output \u1_desOut_reg[42]/_05_  ;
  output \u1_desOut_reg[44]/_05_  ;
  output \u1_desOut_reg[46]/_05_  ;
  output \u1_desOut_reg[48]/_05_  ;
  output \u1_desOut_reg[4]/_05_  ;
  output \u1_desOut_reg[54]/_05_  ;
  output \u1_desOut_reg[56]/_05_  ;
  output \u1_desOut_reg[58]/_05_  ;
  output \u1_desOut_reg[60]/_05_  ;
  output \u1_desOut_reg[62]/_05_  ;
  output \u1_desOut_reg[6]/_05_  ;
  output \u1_desOut_reg[8]/_05_  ;
  output \u2_desOut_reg[0]/_05_  ;
  output \u2_desOut_reg[10]/_05_  ;
  output \u2_desOut_reg[12]/_05_  ;
  output \u2_desOut_reg[14]/_05_  ;
  output \u2_desOut_reg[16]/_05_  ;
  output \u2_desOut_reg[18]/_05_  ;
  output \u2_desOut_reg[20]/_05_  ;
  output \u2_desOut_reg[22]/_05_  ;
  output \u2_desOut_reg[24]/_05_  ;
  output \u2_desOut_reg[26]/_05_  ;
  output \u2_desOut_reg[28]/_05_  ;
  output \u2_desOut_reg[2]/_05_  ;
  output \u2_desOut_reg[30]/_05_  ;
  output \u2_desOut_reg[32]/_05_  ;
  output \u2_desOut_reg[34]/_05_  ;
  output \u2_desOut_reg[36]/_05_  ;
  output \u2_desOut_reg[38]/_05_  ;
  output \u2_desOut_reg[40]/_05_  ;
  output \u2_desOut_reg[42]/_05_  ;
  output \u2_desOut_reg[44]/_05_  ;
  output \u2_desOut_reg[46]/_05_  ;
  output \u2_desOut_reg[48]/_05_  ;
  output \u2_desOut_reg[4]/_05_  ;
  output \u2_desOut_reg[50]/_05_  ;
  output \u2_desOut_reg[52]/_05_  ;
  output \u2_desOut_reg[54]/_05_  ;
  output \u2_desOut_reg[56]/_05_  ;
  output \u2_desOut_reg[58]/_05_  ;
  output \u2_desOut_reg[60]/_05_  ;
  output \u2_desOut_reg[62]/_05_  ;
  output \u2_desOut_reg[6]/_05_  ;
  output \u2_desOut_reg[8]/_05_  ;
  wire n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , n57647 , n57648 , n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , n57657 , n57658 , n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , n57677 , n57678 , n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , n57687 , n57688 , n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , n57697 , n57698 , n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , n57707 , n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , n57717 , n57718 , n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , n57727 , n57728 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , n57737 , n57738 , n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , n57747 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , n57787 , n57788 , n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , n57797 , n57798 , n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , n57807 , n57808 , n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , n57817 , n57818 , n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , n57827 , n57828 , n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , n57837 , n57838 , n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , n57847 , n57848 , n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , n57857 , n57858 , n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , n57867 , n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , n57877 , n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , n57887 , n57888 , n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , n57897 , n57898 , n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , n57907 , n57908 , n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , n57917 , n57918 , n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , n57927 , n57928 , n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , n57937 , n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , n57947 , n57948 , n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , n57957 , n57958 , n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , n57967 , n57968 , n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , n57977 , n57978 , n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , n57987 , n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , n57997 , n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , n58007 , n58008 , n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , n58017 , n58018 , n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , n58027 , n58028 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , n58037 , n58038 , n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , n58047 , n58048 , n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , n58057 , n58058 , n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , n58067 , n58068 , n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , n58077 , n58078 , n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , n58087 , n58088 , n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , n58097 , n58098 , n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , n58107 , n58108 , n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , n58117 , n58118 , n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , n58127 , n58128 , n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , n58137 , n58138 , n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , n58147 , n58148 , n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , n58157 , n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , n58167 , n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , n58177 , n58178 , n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , n58187 , n58188 , n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , n58197 , n58198 , n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , n58207 , n58208 , n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , n58217 , n58218 , n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , n58227 , n58228 , n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , n58237 , n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , n58247 , n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , n58257 , n58258 , n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , n58267 , n58268 , n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , n58277 , n58278 , n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , n58287 , n58288 , n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , n58297 , n58298 , n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , n58307 , n58308 , n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , n58317 , n58318 , n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , n58327 , n58328 , n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , n58337 , n58338 , n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , n58347 , n58348 , n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , n58357 , n58358 , n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , n58367 , n58368 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , n58377 , n58378 , n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , n58387 , n58388 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , n58397 , n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , n58407 , n58408 , n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , n58417 , n58418 , n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , n58427 , n58428 , n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , n58437 , n58438 , n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , n58447 , n58448 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , n58487 , n58488 , n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , n58537 , n58538 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , n58557 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , n58587 , n58588 , n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , n58607 , n58608 , n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , n58617 , n58618 , n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , n58627 , n58628 , n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , n58637 , n58638 , n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , n58647 , n58648 , n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , n58657 , n58658 , n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , n58667 , n58668 , n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , n58677 , n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , n58687 , n58688 , n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , n58697 , n58698 , n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , n58707 , n58708 , n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , n58717 , n58718 , n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , n58727 , n58728 , n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , n58737 , n58738 , n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , n58747 , n58748 , n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , n58757 , n58758 , n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , n58767 , n58768 , n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , n58777 , n58778 , n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , n58787 , n58788 , n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , n58797 , n58798 , n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , n58807 , n58808 , n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , n58817 , n58818 , n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , n58827 , n58828 , n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , n58837 , n58838 , n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , n58847 , n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , n58857 , n58858 , n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , n58867 , n58868 , n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , n58877 , n58878 , n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , n58887 , n58888 , n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , n58897 , n58898 , n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , n58907 , n58908 , n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , n58917 , n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , n58937 , n58938 , n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , n58947 , n58948 , n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , n58957 , n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , n58967 , n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , n58977 , n58978 , n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , n58987 , n58988 , n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , n58997 , n58998 , n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , n59007 , n59008 , n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , n59017 , n59018 , n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , n59027 , n59028 , n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , n59037 , n59038 , n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , n59047 , n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , n59057 , n59058 , n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , n59067 , n59068 , n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , n59077 , n59078 , n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , n59087 , n59088 , n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , n59097 , n59098 , n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , n59107 , n59108 , n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , n59127 , n59128 , n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , n59137 , n59138 , n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , n59147 , n59148 , n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , n59157 , n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , n59167 , n59168 , n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , n59177 , n59178 , n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , n59187 , n59188 , n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , n59197 , n59198 , n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , n59207 , n59208 , n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , n59217 , n59218 , n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , n59227 , n59228 , n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , n59237 , n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , n59247 , n59248 , n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , n59257 , n59258 , n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , n59267 , n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , n59277 , n59278 , n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , n59287 , n59288 , n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , n59297 , n59298 , n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , n59307 , n59308 , n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , n59317 , n59318 , n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , n59327 , n59328 , n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , n59337 , n59338 , n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , n59347 , n59348 , n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , n59357 , n59358 , n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , n59367 , n59368 , n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , n59377 , n59378 , n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , n59387 , n59388 , n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , n59397 , n59398 , n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , n59407 , n59408 , n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , n59417 , n59418 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , n59437 , n59438 , n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , n59447 , n59448 , n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , n59457 , n59458 , n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , n59467 , n59468 , n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , n59477 , n59478 , n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , n59487 , n59488 , n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , n59497 , n59498 , n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , n59507 , n59508 , n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , n59517 , n59518 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , n59527 , n59528 , n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , n59537 , n59538 , n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , n59547 , n59548 , n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , n59557 , n59558 , n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , n59567 , n59568 , n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , n59577 , n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , n59587 , n59588 , n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , n59597 , n59598 , n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , n59607 , n59608 , n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , n59617 , n59618 , n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , n59627 , n59628 , n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , n59637 , n59638 , n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , n59647 , n59648 , n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , n59657 , n59658 , n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , n59667 , n59668 , n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , n59687 , n59688 , n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , n59697 , n59698 , n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , n59707 , n59708 , n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , n59717 , n59718 , n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , n59727 , n59728 , n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , n59737 , n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , n59747 , n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , n59757 , n59758 , n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , n59767 , n59768 , n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , n59777 , n59778 , n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , n59787 , n59788 , n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , n59797 , n59798 , n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , n59807 , n59808 , n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , n59817 , n59818 , n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , n59827 , n59828 , n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , n59837 , n59838 , n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , n59847 , n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , n59857 , n59858 , n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , n59887 , n59888 , n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , n59897 , n59898 , n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , n59907 , n59908 , n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , n59917 , n59918 , n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , n59927 , n59928 , n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , n59937 , n59938 , n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , n59947 , n59948 , n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , n59957 , n59958 , n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , n59967 , n59968 , n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , n59977 , n59978 , n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , n59987 , n59988 , n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , n59997 , n59998 , n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , n60007 , n60008 , n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , n60017 , n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , n60027 , n60028 , n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , n60037 , n60038 , n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , n60047 , n60048 , n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , n60077 , n60078 , n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , n60087 , n60088 , n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , n60097 , n60098 , n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , n60107 , n60108 , n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , n60117 , n60118 , n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , n60127 , n60128 , n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , n60137 , n60138 , n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , n60147 , n60148 , n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , n60157 , n60158 , n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , n60167 , n60168 , n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , n60177 , n60178 , n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , n60187 , n60188 , n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , n60197 , n60198 , n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , n60207 , n60208 , n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , n60217 , n60218 , n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , n60227 , n60228 , n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , n60237 , n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , n60247 , n60248 , n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , n60257 , n60258 , n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , n60267 , n60268 , n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , n60277 , n60278 , n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , n60287 , n60288 , n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , n60297 , n60298 , n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , n60307 , n60308 , n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , n60317 , n60318 , n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , n60327 , n60328 , n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , n60337 , n60338 , n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , n60347 , n60348 , n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , n60357 , n60358 , n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , n60367 , n60368 , n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , n60377 , n60378 , n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , n60397 , n60398 , n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , n60447 , n60448 , n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , n60467 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , n60487 , n60488 , n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , n60497 , n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , n60517 , n60518 , n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , n60527 , n60528 , n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , n60537 , n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , n60547 , n60548 , n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , n60557 , n60558 , n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , n60567 , n60568 , n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , n60577 , n60578 , n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , n60587 , n60588 , n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , n60597 , n60598 , n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , n60607 , n60608 , n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , n60637 , n60638 , n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , n60647 , n60648 , n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , n60657 , n60658 , n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , n60667 , n60668 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , n60677 , n60678 , n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , n60687 , n60688 , n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , n60697 , n60698 , n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , n60707 , n60708 , n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , n60717 , n60718 , n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , n60727 , n60728 , n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , n60737 , n60738 , n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , n60747 , n60748 , n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , n60757 , n60758 , n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , n60767 , n60768 , n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , n60777 , n60778 , n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , n60787 , n60788 , n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , n60797 , n60798 , n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , n60807 , n60808 , n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , n60817 , n60818 , n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , n60827 , n60828 , n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , n60837 , n60838 , n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , n60847 , n60848 , n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , n60857 , n60858 , n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , n60867 , n60868 , n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , n60887 , n60888 , n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , n60897 , n60898 , n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , n60907 , n60908 , n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , n60917 , n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , n60927 , n60928 , n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , n60937 , n60938 , n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , n60947 , n60948 , n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , n60957 , n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , n60967 , n60968 , n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , n60977 , n60978 , n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , n60987 , n60988 , n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , n60997 , n60998 , n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , n61007 , n61008 , n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , n61037 , n61038 , n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , n61047 , n61048 , n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , n61057 , n61058 , n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , n61067 , n61068 , n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , n61077 , n61078 , n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , n61087 , n61088 , n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , n61107 , n61108 , n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , n61117 , n61118 , n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , n61127 , n61128 , n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , n61137 , n61138 , n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , n61147 , n61148 , n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , n61157 , n61158 , n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , n61167 , n61168 , n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , n61177 , n61178 , n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , n61187 , n61188 , n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , n61207 , n61208 , n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , n61217 , n61218 , n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , n61227 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , n61247 , n61248 , n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , n61257 , n61258 , n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , n61267 , n61268 , n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , n61277 , n61278 , n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , n61287 , n61288 , n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , n61297 , n61298 , n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , n61307 , n61308 , n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , n61317 , n61318 , n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , n61327 , n61328 , n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , n61337 , n61338 , n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , n61347 , n61348 , n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , n61357 , n61358 , n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , n61367 , n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , n61377 , n61378 , n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , n61387 , n61388 , n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , n61397 , n61398 , n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , n61407 , n61408 , n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , n61417 , n61418 , n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , n61427 , n61428 , n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , n61437 , n61438 , n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , n61447 , n61448 , n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , n61457 , n61458 , n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , n61467 , n61468 , n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , n61477 , n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , n61497 , n61498 , n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , n61507 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , n61527 , n61528 , n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , n61537 , n61538 , n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , n61547 , n61548 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , n61557 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , n61577 , n61578 , n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , n61587 , n61588 , n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , n61597 , n61598 , n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , n61607 , n61608 , n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , n61617 , n61618 , n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , n61627 , n61628 , n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , n61637 , n61638 , n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , n61647 , n61648 , n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , n61657 , n61658 , n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , n61667 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , n61677 , n61678 , n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , n61687 , n61688 , n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , n61697 , n61698 , n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , n61707 , n61708 , n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , n61717 , n61718 , n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , n61727 , n61728 , n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , n61737 , n61738 , n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , n61747 , n61748 , n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , n61757 , n61758 , n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , n61767 , n61768 , n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , n61787 , n61788 , n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , n61797 , n61798 , n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , n61807 , n61808 , n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , n61817 , n61818 , n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , n61827 , n61828 , n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , n61837 , n61838 , n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , n61847 , n61848 , n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , n61857 , n61858 , n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , n61867 , n61868 , n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , n61877 , n61878 , n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , n61887 , n61888 , n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , n61897 , n61898 , n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , n61907 , n61908 , n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , n61917 , n61918 , n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , n61927 , n61928 , n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , n61937 , n61938 , n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , n61947 , n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , n61957 , n61958 , n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , n61967 , n61968 , n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , n61977 , n61978 , n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , n61987 , n61988 , n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , n61997 , n61998 , n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , n62007 , n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , n62017 , n62018 , n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , n62037 , n62038 , n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , n62047 , n62048 , n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , n62057 , n62058 , n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , n62067 , n62068 , n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , n62077 , n62078 , n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , n62087 , n62088 , n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , n62097 , n62098 , n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , n62107 , n62108 , n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , n62117 , n62118 , n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , n62127 , n62128 , n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , n62137 , n62138 , n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , n62147 , n62148 , n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , n62157 , n62158 , n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , n62167 , n62168 , n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , n62177 , n62178 , n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , n62187 , n62188 , n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , n62197 , n62198 , n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , n62207 , n62208 , n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , n62217 , n62218 , n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , n62227 , n62228 , n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , n62237 , n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , n62247 , n62248 , n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , n62257 , n62258 , n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , n62267 , n62268 , n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , n62277 , n62278 , n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , n62287 , n62288 , n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , n62297 , n62298 , n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , n62307 , n62308 , n62309 , n62310 , n62311 , n62312 , n62313 , n62314 , n62315 , n62316 , n62317 , n62318 , n62319 , n62320 , n62321 , n62322 , n62323 , n62324 , n62325 , n62326 , n62327 , n62328 , n62329 , n62330 , n62331 , n62332 , n62333 , n62334 , n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , n62341 , n62342 , n62343 , n62344 , n62345 , n62346 , n62347 , n62348 , n62349 , n62350 , n62351 , n62352 , n62353 , n62354 , n62355 , n62356 , n62357 , n62358 , n62359 , n62360 , n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , n62367 , n62368 , n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , n62375 , n62376 , n62377 , n62378 , n62379 , n62380 , n62381 , n62382 , n62383 , n62384 , n62385 , n62386 , n62387 , n62388 , n62389 , n62390 , n62391 , n62392 , n62393 , n62394 , n62395 , n62396 , n62397 , n62398 , n62399 , n62400 , n62401 , n62402 , n62403 , n62404 , n62405 , n62406 , n62407 , n62408 , n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , n62415 , n62416 , n62417 , n62418 , n62419 , n62420 , n62421 , n62422 , n62423 , n62424 , n62425 , n62426 , n62427 , n62428 , n62429 , n62430 , n62431 , n62432 , n62433 , n62434 , n62435 , n62436 , n62437 , n62438 , n62439 , n62440 , n62441 , n62442 , n62443 , n62444 , n62445 , n62446 , n62447 , n62448 , n62449 , n62450 , n62451 , n62452 , n62453 , n62454 , n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , n62468 , n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , n62477 , n62478 , n62479 , n62480 , n62481 , n62482 , n62483 , n62484 , n62485 , n62486 , n62487 , n62488 , n62489 , n62490 , n62491 , n62492 , n62493 , n62494 , n62495 , n62496 , n62497 , n62498 , n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , n62505 , n62506 , n62507 , n62508 , n62509 , n62510 , n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , n62517 , n62518 , n62519 , n62520 , n62521 , n62522 , n62523 , n62524 , n62525 , n62526 , n62527 , n62528 , n62529 , n62530 , n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , n62537 , n62538 , n62539 , n62540 , n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , n62547 , n62548 , n62549 , n62550 , n62551 , n62552 , n62553 , n62554 , n62555 , n62556 , n62557 , n62558 , n62559 , n62560 , n62561 , n62562 , n62563 , n62564 , n62565 , n62566 , n62567 , n62568 , n62569 , n62570 , n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , n62581 , n62582 , n62583 , n62584 , n62585 , n62586 , n62587 , n62588 , n62589 , n62590 , n62591 , n62592 , n62593 , n62594 , n62595 , n62596 , n62597 , n62598 , n62599 , n62600 , n62601 , n62602 , n62603 , n62604 , n62605 , n62606 , n62607 , n62608 , n62609 , n62610 , n62611 , n62612 , n62613 , n62614 , n62615 , n62616 , n62617 , n62618 , n62619 , n62620 , n62621 , n62622 , n62623 , n62624 , n62625 , n62626 , n62627 , n62628 , n62629 , n62630 , n62631 , n62632 , n62633 , n62634 , n62635 , n62636 , n62637 , n62638 , n62639 , n62640 , n62641 , n62642 , n62643 , n62644 , n62645 , n62646 , n62647 , n62648 , n62649 , n62650 , n62651 , n62652 , n62653 , n62654 , n62655 , n62656 , n62657 , n62658 , n62659 , n62660 , n62661 , n62662 , n62663 , n62664 , n62665 , n62666 , n62667 , n62668 , n62669 , n62670 , n62671 , n62672 , n62673 , n62674 , n62675 , n62676 , n62677 , n62678 , n62679 , n62680 , n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , n62687 , n62688 , n62689 , n62690 , n62691 , n62692 , n62693 , n62694 , n62695 , n62696 , n62697 , n62698 , n62699 , n62700 , n62701 , n62702 , n62703 , n62704 , n62705 , n62706 , n62707 , n62708 , n62709 , n62710 , n62711 , n62712 , n62713 , n62714 , n62715 , n62716 , n62717 , n62718 , n62719 , n62720 , n62721 , n62722 , n62723 , n62724 , n62725 , n62726 , n62727 , n62728 , n62729 , n62730 , n62731 , n62732 , n62733 , n62734 , n62735 , n62736 , n62737 , n62738 , n62739 , n62740 , n62741 , n62742 , n62743 , n62744 , n62745 , n62746 , n62747 , n62748 , n62749 , n62750 , n62751 , n62752 , n62753 , n62754 , n62755 , n62756 , n62757 , n62758 , n62759 , n62760 , n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , n62767 , n62768 , n62769 , n62770 , n62771 , n62772 , n62773 , n62774 , n62775 , n62776 , n62777 , n62778 , n62779 , n62780 , n62781 , n62782 , n62783 , n62784 , n62785 , n62786 , n62787 , n62788 , n62789 , n62790 , n62791 , n62792 , n62793 , n62794 , n62795 , n62796 , n62797 , n62798 , n62799 , n62800 , n62801 , n62802 , n62803 , n62804 , n62805 , n62806 , n62807 , n62808 , n62809 , n62810 , n62811 , n62812 , n62813 , n62814 , n62815 , n62816 , n62817 , n62818 , n62819 , n62820 , n62821 , n62822 , n62823 , n62824 , n62825 , n62826 , n62827 , n62828 , n62829 , n62830 , n62831 , n62832 , n62833 , n62834 , n62835 , n62836 , n62837 , n62838 , n62839 , n62840 , n62841 , n62842 , n62843 , n62844 , n62845 , n62846 , n62847 , n62848 , n62849 , n62850 , n62851 , n62852 , n62853 , n62854 , n62855 , n62856 , n62857 , n62858 , n62859 , n62860 , n62861 , n62862 , n62863 , n62864 , n62865 , n62866 , n62867 , n62868 , n62869 , n62870 , n62871 , n62872 , n62873 , n62874 , n62875 , n62876 , n62877 , n62878 , n62879 , n62880 , n62881 , n62882 , n62883 , n62884 , n62885 , n62886 , n62887 , n62888 , n62889 , n62890 , n62891 , n62892 , n62893 , n62894 , n62895 , n62896 , n62897 , n62898 , n62899 , n62900 , n62901 , n62902 , n62903 , n62904 , n62905 , n62906 , n62907 , n62908 , n62909 , n62910 , n62911 , n62912 , n62913 , n62914 , n62915 , n62916 , n62917 , n62918 , n62919 , n62920 , n62921 , n62922 , n62923 , n62924 , n62925 , n62926 , n62927 , n62928 , n62929 , n62930 , n62931 , n62932 , n62933 , n62934 , n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , n62941 , n62942 , n62943 , n62944 , n62945 , n62946 , n62947 , n62948 , n62949 , n62950 , n62951 , n62952 , n62953 , n62954 , n62955 , n62956 , n62957 , n62958 , n62959 , n62960 , n62961 , n62962 , n62963 , n62964 , n62965 , n62966 , n62967 , n62968 , n62969 , n62970 , n62971 , n62972 , n62973 , n62974 , n62975 , n62976 , n62977 , n62978 , n62979 , n62980 , n62981 , n62982 , n62983 , n62984 , n62985 , n62986 , n62987 , n62988 , n62989 , n62990 , n62991 , n62992 , n62993 , n62994 , n62995 , n62996 , n62997 , n62998 , n62999 , n63000 , n63001 , n63002 , n63003 , n63004 , n63005 , n63006 , n63007 , n63008 , n63009 , n63010 , n63011 , n63012 , n63013 , n63014 , n63015 , n63016 , n63017 , n63018 , n63019 , n63020 , n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , n63027 , n63028 , n63029 , n63030 , n63031 , n63032 , n63033 , n63034 , n63035 , n63036 , n63037 , n63038 , n63039 , n63040 , n63041 , n63042 , n63043 , n63044 , n63045 , n63046 , n63047 , n63048 , n63049 , n63050 , n63051 , n63052 , n63053 , n63054 , n63055 , n63056 , n63057 , n63058 , n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , n63067 , n63068 , n63069 , n63070 , n63071 , n63072 , n63073 , n63074 , n63075 , n63076 , n63077 , n63078 , n63079 , n63080 , n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , n63087 , n63088 , n63089 , n63090 , n63091 , n63092 , n63093 , n63094 , n63095 , n63096 , n63097 , n63098 , n63099 , n63100 , n63101 , n63102 , n63103 , n63104 , n63105 , n63106 , n63107 , n63108 , n63109 , n63110 , n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , n63117 , n63118 , n63119 , n63120 , n63121 , n63122 , n63123 , n63124 , n63125 , n63126 , n63127 , n63128 , n63129 , n63130 , n63131 , n63132 , n63133 , n63134 , n63135 , n63136 , n63137 , n63138 , n63139 , n63140 , n63141 , n63142 , n63143 , n63144 , n63145 , n63146 , n63147 , n63148 , n63149 , n63150 , n63151 , n63152 , n63153 , n63154 , n63155 , n63156 , n63157 , n63158 , n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , n63167 , n63168 , n63169 , n63170 , n63171 , n63172 , n63173 , n63174 , n63175 , n63176 , n63177 , n63178 , n63179 , n63180 , n63181 , n63182 , n63183 , n63184 , n63185 , n63186 , n63187 , n63188 , n63189 , n63190 , n63191 , n63192 , n63193 , n63194 , n63195 , n63196 , n63197 , n63198 , n63199 , n63200 , n63201 , n63202 , n63203 , n63204 , n63205 , n63206 , n63207 , n63208 , n63209 , n63210 , n63211 , n63212 , n63213 , n63214 , n63215 , n63216 , n63217 , n63218 , n63219 , n63220 , n63221 , n63222 , n63223 , n63224 , n63225 , n63226 , n63227 , n63228 , n63229 , n63230 , n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , n63237 , n63238 , n63239 , n63240 , n63241 , n63242 , n63243 , n63244 , n63245 , n63246 , n63247 , n63248 , n63249 , n63250 , n63251 , n63252 , n63253 , n63254 , n63255 , n63256 , n63257 , n63258 , n63259 , n63260 , n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , n63267 , n63268 , n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , n63275 , n63276 , n63277 , n63278 , n63279 , n63280 , n63281 , n63282 , n63283 , n63284 , n63285 , n63286 , n63287 , n63288 , n63289 , n63290 , n63291 , n63292 , n63293 , n63294 , n63295 , n63296 , n63297 , n63298 , n63299 , n63300 , n63301 , n63302 , n63303 , n63304 , n63305 , n63306 , n63307 , n63308 , n63309 , n63310 , n63311 , n63312 , n63313 , n63314 , n63315 , n63316 , n63317 , n63318 , n63319 , n63320 , n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , n63327 , n63328 , n63329 , n63330 , n63331 , n63332 , n63333 , n63334 , n63335 , n63336 , n63337 , n63338 , n63339 , n63340 , n63341 , n63342 , n63343 , n63344 , n63345 , n63346 , n63347 , n63348 , n63349 , n63350 , n63351 , n63352 , n63353 , n63354 , n63355 , n63356 , n63357 , n63358 , n63359 , n63360 , n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , n63367 , n63368 , n63369 , n63370 , n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , n63385 , n63386 , n63387 , n63388 , n63389 , n63390 , n63391 , n63392 , n63393 , n63394 , n63395 , n63396 , n63397 , n63398 , n63399 , n63400 , n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , n63407 , n63408 , n63409 , n63410 , n63411 , n63412 , n63413 , n63414 , n63415 , n63416 , n63417 , n63418 , n63419 , n63420 , n63421 , n63422 , n63423 , n63424 , n63425 , n63426 , n63427 , n63428 , n63429 , n63430 , n63431 , n63432 , n63433 , n63434 , n63435 , n63436 , n63437 , n63438 , n63439 , n63440 , n63441 , n63442 , n63443 , n63444 , n63445 , n63446 , n63447 , n63448 , n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , n63457 , n63458 , n63459 , n63460 , n63461 , n63462 , n63463 , n63464 , n63465 , n63466 , n63467 , n63468 , n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , n63477 , n63478 , n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , n63487 , n63488 , n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , n63497 , n63498 , n63499 , n63500 , n63501 , n63502 , n63503 , n63504 , n63505 , n63506 , n63507 , n63508 , n63509 , n63510 , n63511 , n63512 , n63513 , n63514 , n63515 , n63516 , n63517 , n63518 , n63519 , n63520 , n63521 , n63522 , n63523 , n63524 , n63525 , n63526 , n63527 , n63528 , n63529 , n63530 , n63531 , n63532 , n63533 , n63534 , n63535 , n63536 , n63537 , n63538 , n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , n63545 , n63546 , n63547 , n63548 , n63549 , n63550 , n63551 , n63552 , n63553 , n63554 , n63555 , n63556 , n63557 , n63558 , n63559 , n63560 , n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , n63567 , n63568 , n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , n63577 , n63578 , n63579 , n63580 , n63581 , n63582 , n63583 , n63584 , n63585 , n63586 , n63587 , n63588 , n63589 , n63590 , n63591 , n63592 , n63593 , n63594 , n63595 , n63596 , n63597 , n63598 , n63599 , n63600 , n63601 , n63602 , n63603 , n63604 , n63605 , n63606 , n63607 , n63608 , n63609 , n63610 , n63611 , n63612 , n63613 , n63614 , n63615 , n63616 , n63617 , n63618 , n63619 , n63620 , n63621 , n63622 , n63623 , n63624 , n63625 , n63626 , n63627 , n63628 , n63629 , n63630 , n63631 , n63632 , n63633 , n63634 , n63635 , n63636 , n63637 , n63638 , n63639 , n63640 , n63641 , n63642 , n63643 , n63644 , n63645 , n63646 , n63647 , n63648 , n63649 , n63650 , n63651 , n63652 , n63653 , n63654 , n63655 , n63656 , n63657 , n63658 , n63659 , n63660 , n63661 , n63662 , n63663 , n63664 , n63665 , n63666 , n63667 , n63668 , n63669 , n63670 , n63671 , n63672 , n63673 , n63674 , n63675 , n63676 , n63677 , n63678 , n63679 , n63680 , n63681 , n63682 , n63683 , n63684 , n63685 , n63686 , n63687 , n63688 , n63689 , n63690 , n63691 , n63692 , n63693 , n63694 , n63695 , n63696 , n63697 , n63698 , n63699 , n63700 , n63701 , n63702 , n63703 , n63704 , n63705 , n63706 , n63707 , n63708 , n63709 , n63710 , n63711 , n63712 , n63713 , n63714 , n63715 , n63716 , n63717 , n63718 , n63719 , n63720 , n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , n63727 , n63728 , n63729 , n63730 , n63731 , n63732 , n63733 , n63734 , n63735 , n63736 , n63737 , n63738 , n63739 , n63740 , n63741 , n63742 , n63743 , n63744 , n63745 , n63746 , n63747 , n63748 , n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , n63757 , n63758 , n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , n63767 , n63768 , n63769 , n63770 , n63771 , n63772 , n63773 , n63774 , n63775 , n63776 , n63777 , n63778 , n63779 , n63780 , n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , n63805 , n63806 , n63807 , n63808 , n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , n63817 , n63818 , n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , n63827 , n63828 , n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , n63837 , n63838 , n63839 , n63840 , n63841 , n63842 , n63843 , n63844 , n63845 , n63846 , n63847 , n63848 , n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , n63857 , n63858 , n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , n63867 , n63868 , n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , n63888 , n63889 , n63890 , n63891 , n63892 , n63893 , n63894 , n63895 , n63896 , n63897 , n63898 , n63899 , n63900 , n63901 , n63902 , n63903 , n63904 , n63905 , n63906 , n63907 , n63908 , n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , n63915 , n63916 , n63917 , n63918 , n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , n63927 , n63928 , n63929 , n63930 , n63931 , n63932 , n63933 , n63934 , n63935 , n63936 , n63937 , n63938 , n63939 , n63940 , n63941 , n63942 , n63943 , n63944 , n63945 , n63946 , n63947 , n63948 , n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , n63957 , n63958 , n63959 , n63960 , n63961 , n63962 , n63963 , n63964 , n63965 , n63966 , n63967 , n63968 , n63969 , n63970 , n63971 , n63972 , n63973 , n63974 , n63975 , n63976 , n63977 , n63978 , n63979 , n63980 , n63981 , n63982 , n63983 , n63984 , n63985 , n63986 , n63987 , n63988 , n63989 , n63990 , n63991 , n63992 , n63993 , n63994 , n63995 , n63996 , n63997 , n63998 , n63999 , n64000 , n64001 , n64002 , n64003 , n64004 , n64005 , n64006 , n64007 , n64008 , n64009 , n64010 , n64011 , n64012 , n64013 , n64014 , n64015 , n64016 , n64017 , n64018 , n64019 , n64020 , n64021 , n64022 , n64023 , n64024 , n64025 , n64026 , n64027 , n64028 , n64029 , n64030 , n64031 , n64032 , n64033 , n64034 , n64035 , n64036 , n64037 , n64038 , n64039 , n64040 , n64041 , n64042 , n64043 , n64044 , n64045 , n64046 , n64047 , n64048 , n64049 , n64050 , n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , n64061 , n64062 , n64063 , n64064 , n64065 , n64066 , n64067 , n64068 , n64069 , n64070 , n64071 , n64072 , n64073 , n64074 , n64075 , n64076 , n64077 , n64078 , n64079 , n64080 , n64081 , n64082 , n64083 , n64084 , n64085 , n64086 , n64087 , n64088 , n64089 , n64090 , n64091 , n64092 , n64093 , n64094 , n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , n64107 , n64108 , n64109 , n64110 , n64111 , n64112 , n64113 , n64114 , n64115 , n64116 , n64117 , n64118 , n64119 , n64120 , n64121 , n64122 , n64123 , n64124 , n64125 , n64126 , n64127 , n64128 , n64129 , n64130 , n64131 , n64132 , n64133 , n64134 , n64135 , n64136 , n64137 , n64138 , n64139 , n64140 , n64141 , n64142 , n64143 , n64144 , n64145 , n64146 , n64147 , n64148 , n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , n64155 , n64156 , n64157 , n64158 , n64159 , n64160 , n64161 , n64162 , n64163 , n64164 , n64165 , n64166 , n64167 , n64168 , n64169 , n64170 , n64171 , n64172 , n64173 , n64174 , n64175 , n64176 , n64177 , n64178 , n64179 , n64180 , n64181 , n64182 , n64183 , n64184 , n64185 , n64186 , n64187 , n64188 , n64189 , n64190 , n64191 , n64192 , n64193 , n64194 , n64195 , n64196 , n64197 , n64198 , n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , n64205 , n64206 , n64207 , n64208 , n64209 , n64210 , n64211 , n64212 , n64213 , n64214 , n64215 , n64216 , n64217 , n64218 , n64219 , n64220 , n64221 , n64222 , n64223 , n64224 , n64225 , n64226 , n64227 , n64228 , n64229 , n64230 , n64231 , n64232 , n64233 , n64234 , n64235 , n64236 , n64237 , n64238 , n64239 , n64240 , n64241 , n64242 , n64243 , n64244 , n64245 , n64246 , n64247 , n64248 , n64249 , n64250 , n64251 , n64252 , n64253 , n64254 , n64255 , n64256 , n64257 , n64258 , n64259 , n64260 , n64261 , n64262 , n64263 , n64264 , n64265 , n64266 , n64267 , n64268 , n64269 , n64270 , n64271 , n64272 , n64273 , n64274 , n64275 , n64276 , n64277 , n64278 , n64279 , n64280 , n64281 , n64282 , n64283 , n64284 , n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , n64295 , n64296 , n64297 , n64298 , n64299 , n64300 , n64301 , n64302 , n64303 , n64304 , n64305 , n64306 , n64307 , n64308 , n64309 , n64310 , n64311 , n64312 , n64313 , n64314 , n64315 , n64316 , n64317 , n64318 , n64319 , n64320 , n64321 , n64322 , n64323 , n64324 , n64325 , n64326 , n64327 , n64328 , n64329 , n64330 , n64331 , n64332 , n64333 , n64334 , n64335 , n64336 , n64337 , n64338 , n64339 , n64340 , n64341 , n64342 , n64343 , n64344 , n64345 , n64346 , n64347 , n64348 , n64349 , n64350 , n64351 , n64352 , n64353 , n64354 , n64355 , n64356 , n64357 , n64358 , n64359 , n64360 , n64361 , n64362 , n64363 , n64364 , n64365 , n64366 , n64367 , n64368 , n64369 , n64370 , n64371 , n64372 , n64373 , n64374 , n64375 , n64376 , n64377 , n64378 , n64379 , n64380 , n64381 , n64382 , n64383 , n64384 , n64385 , n64386 , n64387 , n64388 , n64389 , n64390 , n64391 , n64392 , n64393 , n64394 , n64395 , n64396 , n64397 , n64398 , n64399 , n64400 , n64401 , n64402 , n64403 , n64404 , n64405 , n64406 , n64407 , n64408 , n64409 , n64410 , n64411 , n64412 , n64413 , n64414 , n64415 , n64416 , n64417 , n64418 , n64419 , n64420 , n64421 , n64422 , n64423 , n64424 , n64425 , n64426 , n64427 , n64428 , n64429 , n64430 , n64431 , n64432 , n64433 , n64434 , n64435 , n64436 , n64437 , n64438 , n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , n64445 , n64446 , n64447 , n64448 , n64449 , n64450 , n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , n64457 , n64458 , n64459 , n64460 , n64461 , n64462 , n64463 , n64464 , n64465 , n64466 , n64467 , n64468 , n64469 , n64470 , n64471 , n64472 , n64473 , n64474 , n64475 , n64476 , n64477 , n64478 , n64479 , n64480 , n64481 , n64482 , n64483 , n64484 , n64485 , n64486 , n64487 , n64488 , n64489 , n64490 , n64491 , n64492 , n64493 , n64494 , n64495 , n64496 , n64497 , n64498 , n64499 , n64500 , n64501 , n64502 , n64503 , n64504 , n64505 , n64506 , n64507 , n64508 , n64509 , n64510 , n64511 , n64512 , n64513 , n64514 , n64515 , n64516 , n64517 , n64518 , n64519 , n64520 , n64521 , n64522 , n64523 , n64524 , n64525 , n64526 , n64527 , n64528 , n64529 , n64530 , n64531 , n64532 , n64533 , n64534 , n64535 , n64536 , n64537 , n64538 , n64539 , n64540 , n64541 , n64542 , n64543 , n64544 , n64545 , n64546 , n64547 , n64548 , n64549 , n64550 , n64551 , n64552 , n64553 , n64554 , n64555 , n64556 , n64557 , n64558 , n64559 , n64560 , n64561 , n64562 , n64563 , n64564 , n64565 , n64566 , n64567 , n64568 , n64569 , n64570 , n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , n64577 , n64578 , n64579 , n64580 , n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , n64587 , n64588 , n64589 , n64590 , n64591 , n64592 , n64593 , n64594 , n64595 , n64596 , n64597 , n64598 , n64599 , n64600 , n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , n64607 , n64608 , n64609 , n64610 , n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , n64617 , n64618 , n64619 , n64620 , n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , n64627 , n64628 , n64629 , n64630 , n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , n64637 , n64638 , n64639 , n64640 , n64641 , n64642 , n64643 , n64644 , n64645 , n64646 , n64647 , n64648 , n64649 , n64650 , n64651 , n64652 , n64653 , n64654 , n64655 , n64656 , n64657 , n64658 , n64659 , n64660 , n64661 , n64662 , n64663 , n64664 , n64665 , n64666 , n64667 , n64668 , n64669 , n64670 , n64671 , n64672 , n64673 , n64674 , n64675 , n64676 , n64677 , n64678 , n64679 , n64680 , n64681 , n64682 , n64683 , n64684 , n64685 , n64686 , n64687 , n64688 , n64689 , n64690 , n64691 , n64692 , n64693 , n64694 , n64695 , n64696 , n64697 , n64698 , n64699 , n64700 , n64701 , n64702 , n64703 , n64704 , n64705 , n64706 , n64707 , n64708 , n64709 , n64710 , n64711 , n64712 , n64713 , n64714 , n64715 , n64716 , n64717 , n64718 , n64719 , n64720 , n64721 , n64722 , n64723 , n64724 , n64725 , n64726 , n64727 , n64728 , n64729 , n64730 , n64731 , n64732 , n64733 , n64734 , n64735 , n64736 , n64737 , n64738 , n64739 , n64740 , n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , n64747 , n64748 , n64749 , n64750 , n64751 , n64752 , n64753 , n64754 , n64755 , n64756 , n64757 , n64758 , n64759 , n64760 , n64761 , n64762 , n64763 , n64764 , n64765 , n64766 , n64767 , n64768 , n64769 , n64770 , n64771 , n64772 , n64773 , n64774 , n64775 , n64776 , n64777 , n64778 , n64779 , n64780 , n64781 , n64782 , n64783 , n64784 , n64785 , n64786 , n64787 , n64788 , n64789 , n64790 , n64791 , n64792 , n64793 , n64794 , n64795 , n64796 , n64797 , n64798 , n64799 , n64800 , n64801 , n64802 , n64803 , n64804 , n64805 , n64806 , n64807 , n64808 , n64809 , n64810 , n64811 , n64812 , n64813 , n64814 , n64815 , n64816 , n64817 , n64818 , n64819 , n64820 , n64821 , n64822 , n64823 , n64824 , n64825 , n64826 , n64827 , n64828 , n64829 , n64830 , n64831 , n64832 , n64833 , n64834 , n64835 , n64836 , n64837 , n64838 , n64839 , n64840 , n64841 , n64842 , n64843 , n64844 , n64845 , n64846 , n64847 , n64848 , n64849 , n64850 , n64851 , n64852 , n64853 , n64854 , n64855 , n64856 , n64857 , n64858 , n64859 , n64860 , n64861 , n64862 , n64863 , n64864 , n64865 , n64866 , n64867 , n64868 , n64869 , n64870 , n64871 , n64872 , n64873 , n64874 , n64875 , n64876 , n64877 , n64878 , n64879 , n64880 , n64881 , n64882 , n64883 , n64884 , n64885 , n64886 , n64887 , n64888 , n64889 , n64890 , n64891 , n64892 , n64893 , n64894 , n64895 , n64896 , n64897 , n64898 , n64899 , n64900 , n64901 , n64902 , n64903 , n64904 , n64905 , n64906 , n64907 , n64908 , n64909 , n64910 , n64911 , n64912 , n64913 , n64914 , n64915 , n64916 , n64917 , n64918 , n64919 , n64920 , n64921 , n64922 , n64923 , n64924 , n64925 , n64926 , n64927 , n64928 , n64929 , n64930 , n64931 , n64932 , n64933 , n64934 , n64935 , n64936 , n64937 , n64938 , n64939 , n64940 , n64941 , n64942 , n64943 , n64944 , n64945 , n64946 , n64947 , n64948 , n64949 , n64950 , n64951 , n64952 , n64953 , n64954 , n64955 , n64956 , n64957 , n64958 , n64959 , n64960 , n64961 , n64962 , n64963 , n64964 , n64965 , n64966 , n64967 , n64968 , n64969 , n64970 , n64971 , n64972 , n64973 , n64974 , n64975 , n64976 , n64977 , n64978 , n64979 , n64980 , n64981 , n64982 , n64983 , n64984 , n64985 , n64986 , n64987 , n64988 , n64989 , n64990 , n64991 , n64992 , n64993 , n64994 , n64995 , n64996 , n64997 , n64998 , n64999 , n65000 , n65001 , n65002 , n65003 , n65004 , n65005 , n65006 , n65007 , n65008 , n65009 , n65010 , n65011 , n65012 , n65013 , n65014 , n65015 , n65016 , n65017 , n65018 , n65019 , n65020 , n65021 , n65022 , n65023 , n65024 , n65025 , n65026 , n65027 , n65028 , n65029 , n65030 , n65031 , n65032 , n65033 , n65034 , n65035 , n65036 , n65037 , n65038 , n65039 , n65040 , n65041 , n65042 , n65043 , n65044 , n65045 , n65046 , n65047 , n65048 , n65049 , n65050 , n65051 , n65052 , n65053 , n65054 , n65055 , n65056 , n65057 , n65058 , n65059 , n65060 , n65061 , n65062 , n65063 , n65064 , n65065 , n65066 , n65067 , n65068 , n65069 , n65070 , n65071 , n65072 , n65073 , n65074 , n65075 , n65076 , n65077 , n65078 , n65079 , n65080 , n65081 , n65082 , n65083 , n65084 , n65085 , n65086 , n65087 , n65088 , n65089 , n65090 , n65091 , n65092 , n65093 , n65094 , n65095 , n65096 , n65097 , n65098 , n65099 , n65100 , n65101 , n65102 , n65103 , n65104 , n65105 , n65106 , n65107 , n65108 , n65109 , n65110 , n65111 , n65112 , n65113 , n65114 , n65115 , n65116 , n65117 , n65118 , n65119 , n65120 , n65121 , n65122 , n65123 , n65124 , n65125 , n65126 , n65127 , n65128 , n65129 , n65130 , n65131 , n65132 , n65133 , n65134 , n65135 , n65136 , n65137 , n65138 , n65139 , n65140 , n65141 , n65142 , n65143 , n65144 , n65145 , n65146 , n65147 , n65148 , n65149 , n65150 , n65151 , n65152 , n65153 , n65154 , n65155 , n65156 , n65157 , n65158 , n65159 , n65160 , n65161 , n65162 , n65163 , n65164 , n65165 , n65166 , n65167 , n65168 , n65169 , n65170 , n65171 , n65172 , n65173 , n65174 , n65175 , n65176 , n65177 , n65178 , n65179 , n65180 , n65181 , n65182 , n65183 , n65184 , n65185 , n65186 , n65187 , n65188 , n65189 , n65190 , n65191 , n65192 , n65193 , n65194 , n65195 , n65196 , n65197 , n65198 , n65199 , n65200 , n65201 , n65202 , n65203 , n65204 , n65205 , n65206 , n65207 , n65208 , n65209 , n65210 , n65211 , n65212 , n65213 , n65214 , n65215 , n65216 , n65217 , n65218 , n65219 , n65220 , n65221 , n65222 , n65223 , n65224 , n65225 , n65226 , n65227 , n65228 , n65229 , n65230 , n65231 , n65232 , n65233 , n65234 , n65235 , n65236 , n65237 , n65238 , n65239 , n65240 , n65241 , n65242 , n65243 , n65244 , n65245 , n65246 , n65247 , n65248 , n65249 , n65250 , n65251 , n65252 , n65253 , n65254 , n65255 , n65256 , n65257 , n65258 , n65259 , n65260 , n65261 , n65262 , n65263 , n65264 , n65265 , n65266 , n65267 , n65268 , n65269 , n65270 , n65271 , n65272 , n65273 , n65274 , n65275 , n65276 , n65277 , n65278 , n65279 , n65280 , n65281 , n65282 , n65283 , n65284 , n65285 , n65286 , n65287 , n65288 , n65289 , n65290 , n65291 , n65292 , n65293 , n65294 , n65295 , n65296 , n65297 , n65298 , n65299 , n65300 , n65301 , n65302 , n65303 , n65304 , n65305 , n65306 , n65307 , n65308 , n65309 , n65310 , n65311 , n65312 , n65313 , n65314 , n65315 , n65316 , n65317 , n65318 , n65319 , n65320 , n65321 , n65322 , n65323 , n65324 , n65325 , n65326 , n65327 , n65328 , n65329 , n65330 , n65331 , n65332 , n65333 , n65334 , n65335 , n65336 , n65337 , n65338 , n65339 , n65340 , n65341 , n65342 , n65343 , n65344 , n65345 , n65346 , n65347 , n65348 , n65349 , n65350 , n65351 , n65352 , n65353 , n65354 , n65355 , n65356 , n65357 , n65358 , n65359 , n65360 , n65361 , n65362 , n65363 , n65364 , n65365 , n65366 , n65367 , n65368 , n65369 , n65370 , n65371 , n65372 , n65373 , n65374 , n65375 , n65376 , n65377 , n65378 , n65379 , n65380 , n65381 , n65382 , n65383 , n65384 , n65385 , n65386 , n65387 , n65388 , n65389 , n65390 , n65391 , n65392 , n65393 , n65394 , n65395 , n65396 , n65397 , n65398 , n65399 , n65400 , n65401 , n65402 , n65403 , n65404 , n65405 , n65406 , n65407 , n65408 , n65409 , n65410 , n65411 , n65412 , n65413 , n65414 , n65415 , n65416 , n65417 , n65418 , n65419 , n65420 , n65421 , n65422 , n65423 , n65424 , n65425 , n65426 , n65427 , n65428 , n65429 , n65430 , n65431 , n65432 , n65433 , n65434 , n65435 , n65436 , n65437 , n65438 , n65439 , n65440 , n65441 , n65442 , n65443 , n65444 , n65445 , n65446 , n65447 , n65448 , n65449 , n65450 , n65451 , n65452 , n65453 , n65454 , n65455 , n65456 , n65457 , n65458 , n65459 , n65460 , n65461 , n65462 , n65463 , n65464 , n65465 , n65466 , n65467 , n65468 , n65469 , n65470 , n65471 , n65472 , n65473 , n65474 , n65475 , n65476 , n65477 , n65478 , n65479 , n65480 , n65481 , n65482 , n65483 , n65484 , n65485 , n65486 , n65487 , n65488 , n65489 , n65490 , n65491 , n65492 , n65493 , n65494 , n65495 , n65496 , n65497 , n65498 , n65499 , n65500 , n65501 , n65502 , n65503 , n65504 , n65505 , n65506 , n65507 , n65508 , n65509 , n65510 , n65511 , n65512 , n65513 , n65514 , n65515 , n65516 , n65517 , n65518 , n65519 , n65520 , n65521 , n65522 , n65523 , n65524 , n65525 , n65526 , n65527 , n65528 , n65529 , n65530 , n65531 , n65532 , n65533 , n65534 , n65535 , n65536 , n65537 , n65538 , n65539 , n65540 , n65541 , n65542 , n65543 , n65544 , n65545 , n65546 , n65547 , n65548 , n65549 , n65550 , n65551 , n65552 , n65553 , n65554 , n65555 , n65556 , n65557 , n65558 , n65559 , n65560 , n65561 , n65562 , n65563 , n65564 , n65565 , n65566 , n65567 , n65568 , n65569 , n65570 , n65571 , n65572 , n65573 , n65574 , n65575 , n65576 , n65577 , n65578 , n65579 , n65580 , n65581 , n65582 , n65583 , n65584 , n65585 , n65586 , n65587 , n65588 , n65589 , n65590 , n65591 , n65592 , n65593 , n65594 , n65595 , n65596 , n65597 , n65598 , n65599 , n65600 , n65601 , n65602 , n65603 , n65604 , n65605 , n65606 , n65607 , n65608 , n65609 , n65610 , n65611 , n65612 , n65613 , n65614 , n65615 , n65616 , n65617 , n65618 , n65619 , n65620 , n65621 , n65622 , n65623 , n65624 , n65625 , n65626 , n65627 , n65628 , n65629 , n65630 , n65631 , n65632 , n65633 , n65634 , n65635 , n65636 , n65637 , n65638 , n65639 , n65640 , n65641 , n65642 , n65643 , n65644 , n65645 , n65646 , n65647 , n65648 , n65649 , n65650 , n65651 , n65652 , n65653 , n65654 , n65655 , n65656 , n65657 , n65658 , n65659 , n65660 , n65661 , n65662 , n65663 , n65664 , n65665 , n65666 , n65667 , n65668 , n65669 , n65670 , n65671 , n65672 , n65673 , n65674 , n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , n65681 , n65682 , n65683 , n65684 , n65685 , n65686 , n65687 , n65688 , n65689 , n65690 , n65691 , n65692 , n65693 , n65694 , n65695 , n65696 , n65697 , n65698 , n65699 , n65700 , n65701 , n65702 , n65703 , n65704 , n65705 , n65706 , n65707 , n65708 , n65709 , n65710 , n65711 , n65712 , n65713 , n65714 , n65715 , n65716 , n65717 , n65718 , n65719 , n65720 , n65721 , n65722 , n65723 , n65724 , n65725 , n65726 , n65727 , n65728 , n65729 , n65730 , n65731 , n65732 , n65733 , n65734 , n65735 , n65736 , n65737 , n65738 , n65739 , n65740 , n65741 , n65742 , n65743 , n65744 , n65745 , n65746 , n65747 , n65748 , n65749 , n65750 , n65751 , n65752 , n65753 , n65754 , n65755 , n65756 , n65757 , n65758 , n65759 , n65760 , n65761 , n65762 , n65763 , n65764 , n65765 , n65766 , n65767 , n65768 , n65769 , n65770 , n65771 , n65772 , n65773 , n65774 , n65775 , n65776 , n65777 , n65778 , n65779 , n65780 , n65781 , n65782 , n65783 , n65784 , n65785 , n65786 , n65787 , n65788 , n65789 , n65790 , n65791 , n65792 , n65793 , n65794 , n65795 , n65796 , n65797 , n65798 , n65799 , n65800 , n65801 , n65802 , n65803 , n65804 , n65805 , n65806 , n65807 , n65808 , n65809 , n65810 , n65811 , n65812 , n65813 , n65814 , n65815 , n65816 , n65817 , n65818 , n65819 , n65820 , n65821 , n65822 , n65823 , n65824 , n65825 , n65826 , n65827 , n65828 , n65829 , n65830 , n65831 , n65832 , n65833 , n65834 , n65835 , n65836 , n65837 , n65838 , n65839 , n65840 , n65841 , n65842 , n65843 , n65844 , n65845 , n65846 , n65847 , n65848 , n65849 , n65850 , n65851 , n65852 , n65853 , n65854 , n65855 , n65856 , n65857 , n65858 , n65859 , n65860 , n65861 , n65862 , n65863 , n65864 , n65865 , n65866 , n65867 , n65868 , n65869 , n65870 , n65871 , n65872 , n65873 , n65874 , n65875 , n65876 , n65877 , n65878 , n65879 , n65880 , n65881 , n65882 , n65883 , n65884 , n65885 , n65886 , n65887 , n65888 , n65889 , n65890 , n65891 , n65892 , n65893 , n65894 , n65895 , n65896 , n65897 , n65898 , n65899 , n65900 , n65901 , n65902 , n65903 , n65904 , n65905 , n65906 , n65907 , n65908 , n65909 , n65910 , n65911 , n65912 , n65913 , n65914 , n65915 , n65916 , n65917 , n65918 , n65919 , n65920 , n65921 , n65922 , n65923 , n65924 , n65925 , n65926 , n65927 , n65928 , n65929 , n65930 , n65931 , n65932 , n65933 , n65934 , n65935 , n65936 , n65937 , n65938 , n65939 , n65940 , n65941 , n65942 , n65943 , n65944 , n65945 , n65946 , n65947 , n65948 , n65949 , n65950 , n65951 , n65952 , n65953 , n65954 , n65955 , n65956 , n65957 , n65958 , n65959 , n65960 , n65961 , n65962 , n65963 , n65964 , n65965 , n65966 , n65967 , n65968 , n65969 , n65970 , n65971 , n65972 , n65973 , n65974 , n65975 , n65976 , n65977 , n65978 , n65979 , n65980 , n65981 , n65982 , n65983 , n65984 , n65985 , n65986 , n65987 , n65988 , n65989 , n65990 , n65991 , n65992 , n65993 , n65994 , n65995 , n65996 , n65997 , n65998 , n65999 , n66000 , n66001 , n66002 , n66003 , n66004 , n66005 , n66006 , n66007 , n66008 , n66009 , n66010 , n66011 , n66012 , n66013 , n66014 , n66015 , n66016 , n66017 , n66018 , n66019 , n66020 , n66021 , n66022 , n66023 , n66024 , n66025 , n66026 , n66027 , n66028 , n66029 , n66030 , n66031 , n66032 , n66033 , n66034 , n66035 , n66036 , n66037 , n66038 , n66039 , n66040 , n66041 , n66042 , n66043 , n66044 , n66045 , n66046 , n66047 , n66048 , n66049 , n66050 , n66051 , n66052 , n66053 , n66054 , n66055 , n66056 , n66057 , n66058 , n66059 , n66060 , n66061 , n66062 , n66063 , n66064 , n66065 , n66066 , n66067 , n66068 , n66069 , n66070 , n66071 , n66072 , n66073 , n66074 , n66075 , n66076 , n66077 , n66078 , n66079 , n66080 , n66081 , n66082 , n66083 , n66084 , n66085 , n66086 , n66087 , n66088 , n66089 , n66090 , n66091 , n66092 , n66093 , n66094 , n66095 , n66096 , n66097 , n66098 , n66099 , n66100 , n66101 , n66102 , n66103 , n66104 , n66105 , n66106 , n66107 , n66108 , n66109 , n66110 , n66111 , n66112 , n66113 , n66114 , n66115 , n66116 , n66117 , n66118 , n66119 , n66120 , n66121 , n66122 , n66123 , n66124 , n66125 , n66126 , n66127 , n66128 , n66129 , n66130 , n66131 , n66132 , n66133 , n66134 , n66135 , n66136 , n66137 , n66138 , n66139 , n66140 , n66141 , n66142 , n66143 , n66144 , n66145 , n66146 , n66147 , n66148 , n66149 , n66150 , n66151 , n66152 , n66153 , n66154 , n66155 , n66156 , n66157 , n66158 , n66159 , n66160 , n66161 , n66162 , n66163 , n66164 , n66165 , n66166 , n66167 , n66168 , n66169 , n66170 , n66171 , n66172 , n66173 , n66174 , n66175 , n66176 , n66177 , n66178 , n66179 , n66180 , n66181 , n66182 , n66183 , n66184 , n66185 , n66186 , n66187 , n66188 , n66189 , n66190 , n66191 , n66192 , n66193 , n66194 , n66195 , n66196 , n66197 , n66198 , n66199 , n66200 , n66201 , n66202 , n66203 , n66204 , n66205 , n66206 , n66207 , n66208 , n66209 , n66210 , n66211 , n66212 , n66213 , n66214 , n66215 , n66216 , n66217 , n66218 , n66219 , n66220 , n66221 , n66222 , n66223 , n66224 , n66225 , n66226 , n66227 , n66228 , n66229 , n66230 , n66231 , n66232 , n66233 , n66234 , n66235 , n66236 , n66237 , n66238 , n66239 , n66240 , n66241 , n66242 , n66243 , n66244 , n66245 , n66246 , n66247 , n66248 , n66249 , n66250 , n66251 , n66252 , n66253 , n66254 , n66255 , n66256 , n66257 , n66258 , n66259 , n66260 , n66261 , n66262 , n66263 , n66264 , n66265 , n66266 , n66267 , n66268 , n66269 , n66270 , n66271 , n66272 , n66273 , n66274 , n66275 , n66276 , n66277 , n66278 , n66279 , n66280 , n66281 , n66282 , n66283 , n66284 , n66285 , n66286 , n66287 , n66288 , n66289 , n66290 , n66291 , n66292 , n66293 , n66294 , n66295 , n66296 , n66297 , n66298 , n66299 , n66300 , n66301 , n66302 , n66303 , n66304 , n66305 , n66306 , n66307 , n66308 , n66309 , n66310 , n66311 , n66312 , n66313 , n66314 , n66315 , n66316 , n66317 , n66318 , n66319 , n66320 , n66321 , n66322 , n66323 , n66324 , n66325 , n66326 , n66327 , n66328 , n66329 , n66330 , n66331 , n66332 , n66333 , n66334 , n66335 , n66336 , n66337 , n66338 , n66339 , n66340 , n66341 , n66342 , n66343 , n66344 , n66345 , n66346 , n66347 , n66348 , n66349 , n66350 , n66351 , n66352 , n66353 , n66354 , n66355 , n66356 , n66357 , n66358 , n66359 , n66360 , n66361 , n66362 , n66363 , n66364 , n66365 , n66366 , n66367 , n66368 , n66369 , n66370 , n66371 , n66372 , n66373 , n66374 , n66375 , n66376 , n66377 , n66378 , n66379 , n66380 , n66381 , n66382 , n66383 , n66384 , n66385 , n66386 , n66387 , n66388 , n66389 , n66390 , n66391 , n66392 , n66393 , n66394 , n66395 , n66396 , n66397 , n66398 , n66399 , n66400 , n66401 , n66402 , n66403 , n66404 , n66405 , n66406 , n66407 , n66408 , n66409 , n66410 , n66411 , n66412 , n66413 , n66414 , n66415 , n66416 , n66417 , n66418 , n66419 , n66420 , n66421 , n66422 , n66423 , n66424 , n66425 , n66426 , n66427 , n66428 , n66429 , n66430 , n66431 , n66432 , n66433 , n66434 , n66435 , n66436 , n66437 , n66438 , n66439 , n66440 , n66441 , n66442 , n66443 , n66444 , n66445 , n66446 , n66447 , n66448 , n66449 , n66450 , n66451 , n66452 , n66453 , n66454 , n66455 , n66456 , n66457 , n66458 , n66459 , n66460 , n66461 , n66462 , n66463 , n66464 , n66465 , n66466 , n66467 , n66468 , n66469 , n66470 , n66471 , n66472 , n66473 , n66474 , n66475 , n66476 , n66477 , n66478 , n66479 , n66480 , n66481 , n66482 , n66483 , n66484 , n66485 , n66486 , n66487 , n66488 , n66489 , n66490 , n66491 , n66492 , n66493 , n66494 , n66495 , n66496 , n66497 , n66498 , n66499 , n66500 , n66501 , n66502 , n66503 , n66504 , n66505 , n66506 , n66507 , n66508 , n66509 , n66510 , n66511 , n66512 , n66513 , n66514 , n66515 , n66516 , n66517 , n66518 , n66519 , n66520 , n66521 , n66522 , n66523 , n66524 , n66525 , n66526 , n66527 , n66528 , n66529 , n66530 , n66531 , n66532 , n66533 , n66534 , n66535 , n66536 , n66537 , n66538 , n66539 , n66540 , n66541 , n66542 , n66543 , n66544 , n66545 , n66546 , n66547 , n66548 , n66549 , n66550 , n66551 , n66552 , n66553 , n66554 , n66555 , n66556 , n66557 , n66558 , n66559 , n66560 , n66561 , n66562 , n66563 , n66564 , n66565 , n66566 , n66567 , n66568 , n66569 , n66570 , n66571 , n66572 , n66573 , n66574 , n66575 , n66576 , n66577 , n66578 , n66579 , n66580 , n66581 , n66582 , n66583 , n66584 , n66585 , n66586 , n66587 , n66588 , n66589 , n66590 , n66591 , n66592 , n66593 , n66594 , n66595 , n66596 , n66597 , n66598 , n66599 , n66600 , n66601 , n66602 , n66603 , n66604 , n66605 , n66606 , n66607 , n66608 , n66609 , n66610 , n66611 , n66612 , n66613 , n66614 , n66615 , n66616 , n66617 , n66618 , n66619 , n66620 , n66621 , n66622 , n66623 , n66624 , n66625 , n66626 , n66627 , n66628 , n66629 , n66630 , n66631 , n66632 , n66633 , n66634 , n66635 , n66636 , n66637 , n66638 , n66639 , n66640 , n66641 , n66642 , n66643 , n66644 , n66645 , n66646 , n66647 , n66648 , n66649 , n66650 , n66651 , n66652 , n66653 , n66654 , n66655 , n66656 , n66657 , n66658 , n66659 , n66660 , n66661 , n66662 , n66663 , n66664 , n66665 , n66666 , n66667 , n66668 , n66669 , n66670 , n66671 , n66672 , n66673 , n66674 , n66675 , n66676 , n66677 , n66678 , n66679 , n66680 , n66681 , n66682 , n66683 , n66684 , n66685 , n66686 , n66687 , n66688 , n66689 , n66690 , n66691 , n66692 , n66693 , n66694 , n66695 , n66696 , n66697 , n66698 , n66699 , n66700 , n66701 , n66702 , n66703 , n66704 , n66705 , n66706 , n66707 , n66708 , n66709 , n66710 , n66711 , n66712 , n66713 , n66714 , n66715 , n66716 , n66717 , n66718 , n66719 , n66720 , n66721 , n66722 , n66723 , n66724 , n66725 , n66726 , n66727 , n66728 , n66729 , n66730 , n66731 , n66732 , n66733 , n66734 , n66735 , n66736 , n66737 , n66738 , n66739 , n66740 , n66741 , n66742 , n66743 , n66744 , n66745 , n66746 , n66747 , n66748 , n66749 , n66750 , n66751 , n66752 , n66753 , n66754 , n66755 , n66756 , n66757 , n66758 , n66759 , n66760 , n66761 , n66762 , n66763 , n66764 , n66765 , n66766 , n66767 , n66768 , n66769 , n66770 , n66771 , n66772 , n66773 , n66774 , n66775 , n66776 , n66777 , n66778 , n66779 , n66780 , n66781 , n66782 , n66783 , n66784 , n66785 , n66786 , n66787 , n66788 , n66789 , n66790 , n66791 , n66792 , n66793 , n66794 , n66795 , n66796 , n66797 , n66798 , n66799 , n66800 , n66801 , n66802 , n66803 , n66804 , n66805 , n66806 , n66807 , n66808 , n66809 , n66810 , n66811 , n66812 , n66813 , n66814 , n66815 , n66816 , n66817 , n66818 , n66819 , n66820 , n66821 , n66822 , n66823 , n66824 , n66825 , n66826 , n66827 , n66828 , n66829 , n66830 , n66831 , n66832 , n66833 , n66834 , n66835 , n66836 , n66837 , n66838 , n66839 , n66840 , n66841 , n66842 , n66843 , n66844 , n66845 , n66846 , n66847 , n66848 , n66849 , n66850 , n66851 , n66852 , n66853 , n66854 , n66855 , n66856 , n66857 , n66858 , n66859 , n66860 , n66861 , n66862 , n66863 , n66864 , n66865 , n66866 , n66867 , n66868 , n66869 , n66870 , n66871 , n66872 , n66873 , n66874 , n66875 , n66876 , n66877 , n66878 , n66879 , n66880 , n66881 , n66882 , n66883 , n66884 , n66885 , n66886 , n66887 , n66888 , n66889 , n66890 , n66891 , n66892 , n66893 , n66894 , n66895 , n66896 , n66897 , n66898 , n66899 , n66900 , n66901 , n66902 , n66903 , n66904 , n66905 , n66906 , n66907 , n66908 , n66909 , n66910 , n66911 , n66912 , n66913 , n66914 , n66915 , n66916 , n66917 , n66918 , n66919 , n66920 , n66921 , n66922 , n66923 , n66924 , n66925 , n66926 , n66927 , n66928 , n66929 , n66930 , n66931 , n66932 , n66933 , n66934 , n66935 , n66936 , n66937 , n66938 , n66939 , n66940 , n66941 , n66942 , n66943 , n66944 , n66945 , n66946 , n66947 , n66948 , n66949 , n66950 , n66951 , n66952 , n66953 , n66954 , n66955 , n66956 , n66957 , n66958 , n66959 , n66960 , n66961 , n66962 , n66963 , n66964 , n66965 , n66966 , n66967 , n66968 , n66969 , n66970 , n66971 , n66972 , n66973 , n66974 , n66975 , n66976 , n66977 , n66978 , n66979 , n66980 , n66981 , n66982 , n66983 , n66984 , n66985 , n66986 , n66987 , n66988 , n66989 , n66990 , n66991 , n66992 , n66993 , n66994 , n66995 , n66996 , n66997 , n66998 , n66999 , n67000 , n67001 , n67002 , n67003 , n67004 , n67005 , n67006 , n67007 , n67008 , n67009 , n67010 , n67011 , n67012 , n67013 , n67014 , n67015 , n67016 , n67017 , n67018 , n67019 , n67020 , n67021 , n67022 , n67023 , n67024 , n67025 , n67026 , n67027 , n67028 , n67029 , n67030 , n67031 , n67032 , n67033 , n67034 , n67035 , n67036 , n67037 , n67038 , n67039 , n67040 , n67041 , n67042 , n67043 , n67044 , n67045 , n67046 , n67047 , n67048 , n67049 , n67050 , n67051 , n67052 , n67053 , n67054 , n67055 , n67056 , n67057 , n67058 , n67059 , n67060 , n67061 , n67062 , n67063 , n67064 , n67065 , n67066 , n67067 , n67068 , n67069 , n67070 , n67071 , n67072 , n67073 , n67074 , n67075 , n67076 , n67077 , n67078 , n67079 , n67080 , n67081 , n67082 , n67083 , n67084 , n67085 , n67086 , n67087 , n67088 , n67089 , n67090 , n67091 , n67092 , n67093 , n67094 , n67095 , n67096 , n67097 , n67098 , n67099 , n67100 , n67101 , n67102 , n67103 , n67104 , n67105 , n67106 , n67107 , n67108 , n67109 , n67110 , n67111 , n67112 , n67113 , n67114 , n67115 , n67116 , n67117 , n67118 , n67119 , n67120 , n67121 , n67122 , n67123 , n67124 , n67125 , n67126 , n67127 , n67128 , n67129 , n67130 , n67131 , n67132 , n67133 , n67134 , n67135 , n67136 , n67137 , n67138 , n67139 , n67140 , n67141 , n67142 , n67143 , n67144 , n67145 , n67146 , n67147 , n67148 , n67149 , n67150 , n67151 , n67152 , n67153 , n67154 , n67155 , n67156 , n67157 , n67158 , n67159 , n67160 , n67161 , n67162 , n67163 , n67164 , n67165 , n67166 , n67167 , n67168 , n67169 , n67170 , n67171 , n67172 , n67173 , n67174 , n67175 , n67176 , n67177 , n67178 , n67179 , n67180 , n67181 , n67182 , n67183 , n67184 , n67185 , n67186 , n67187 , n67188 , n67189 , n67190 , n67191 , n67192 , n67193 , n67194 , n67195 , n67196 , n67197 , n67198 , n67199 , n67200 , n67201 , n67202 , n67203 , n67204 , n67205 , n67206 , n67207 , n67208 , n67209 , n67210 , n67211 , n67212 , n67213 , n67214 , n67215 , n67216 , n67217 , n67218 , n67219 , n67220 , n67221 , n67222 , n67223 , n67224 , n67225 , n67226 , n67227 , n67228 , n67229 , n67230 , n67231 , n67232 , n67233 , n67234 , n67235 , n67236 , n67237 , n67238 , n67239 , n67240 , n67241 , n67242 , n67243 , n67244 , n67245 , n67246 , n67247 , n67248 , n67249 , n67250 , n67251 , n67252 , n67253 , n67254 , n67255 , n67256 , n67257 , n67258 , n67259 , n67260 , n67261 , n67262 , n67263 , n67264 , n67265 , n67266 , n67267 , n67268 , n67269 , n67270 , n67271 , n67272 , n67273 , n67274 , n67275 , n67276 , n67277 , n67278 , n67279 , n67280 , n67281 , n67282 , n67283 , n67284 , n67285 , n67286 , n67287 , n67288 , n67289 , n67290 , n67291 , n67292 , n67293 , n67294 , n67295 , n67296 , n67297 , n67298 , n67299 , n67300 , n67301 , n67302 , n67303 , n67304 , n67305 , n67306 , n67307 , n67308 , n67309 , n67310 , n67311 , n67312 , n67313 , n67314 , n67315 , n67316 , n67317 , n67318 , n67319 , n67320 , n67321 , n67322 , n67323 , n67324 , n67325 , n67326 , n67327 , n67328 , n67329 , n67330 , n67331 , n67332 , n67333 , n67334 , n67335 , n67336 , n67337 , n67338 , n67339 , n67340 , n67341 , n67342 , n67343 , n67344 , n67345 , n67346 , n67347 , n67348 , n67349 , n67350 , n67351 , n67352 , n67353 , n67354 , n67355 , n67356 , n67357 , n67358 , n67359 , n67360 , n67361 , n67362 , n67363 , n67364 , n67365 , n67366 , n67367 , n67368 , n67369 , n67370 , n67371 , n67372 , n67373 , n67374 , n67375 , n67376 , n67377 , n67378 , n67379 , n67380 , n67381 , n67382 , n67383 , n67384 , n67385 , n67386 , n67387 , n67388 , n67389 , n67390 , n67391 , n67392 , n67393 , n67394 , n67395 , n67396 , n67397 , n67398 , n67399 , n67400 , n67401 , n67402 , n67403 , n67404 , n67405 , n67406 , n67407 , n67408 , n67409 , n67410 , n67411 , n67412 , n67413 , n67414 , n67415 , n67416 , n67417 , n67418 , n67419 , n67420 , n67421 , n67422 , n67423 , n67424 , n67425 , n67426 , n67427 , n67428 , n67429 , n67430 , n67431 , n67432 , n67433 , n67434 , n67435 , n67436 , n67437 , n67438 , n67439 , n67440 , n67441 , n67442 , n67443 , n67444 , n67445 , n67446 , n67447 , n67448 , n67449 , n67450 , n67451 , n67452 , n67453 , n67454 , n67455 , n67456 , n67457 , n67458 , n67459 , n67460 , n67461 , n67462 , n67463 , n67464 , n67465 , n67466 , n67467 , n67468 , n67469 , n67470 , n67471 , n67472 , n67473 , n67474 , n67475 , n67476 , n67477 , n67478 , n67479 , n67480 , n67481 , n67482 , n67483 , n67484 , n67485 , n67486 , n67487 , n67488 , n67489 , n67490 , n67491 , n67492 , n67493 , n67494 , n67495 , n67496 , n67497 , n67498 , n67499 , n67500 , n67501 , n67502 , n67503 , n67504 , n67505 , n67506 , n67507 , n67508 , n67509 , n67510 , n67511 , n67512 , n67513 , n67514 , n67515 , n67516 , n67517 , n67518 , n67519 , n67520 , n67521 , n67522 , n67523 , n67524 , n67525 , n67526 , n67527 , n67528 , n67529 , n67530 , n67531 , n67532 , n67533 , n67534 , n67535 , n67536 , n67537 , n67538 , n67539 , n67540 , n67541 , n67542 , n67543 , n67544 , n67545 , n67546 , n67547 , n67548 , n67549 , n67550 , n67551 , n67552 , n67553 , n67554 , n67555 , n67556 , n67557 , n67558 , n67559 , n67560 , n67561 , n67562 , n67563 , n67564 , n67565 , n67566 , n67567 , n67568 , n67569 , n67570 , n67571 , n67572 , n67573 , n67574 , n67575 , n67576 , n67577 , n67578 , n67579 , n67580 , n67581 , n67582 , n67583 , n67584 , n67585 , n67586 , n67587 , n67588 , n67589 , n67590 , n67591 , n67592 , n67593 , n67594 , n67595 , n67596 , n67597 , n67598 , n67599 , n67600 , n67601 , n67602 , n67603 , n67604 , n67605 , n67606 , n67607 , n67608 , n67609 , n67610 , n67611 , n67612 , n67613 , n67614 , n67615 , n67616 , n67617 , n67618 , n67619 , n67620 , n67621 , n67622 , n67623 , n67624 , n67625 , n67626 , n67627 , n67628 , n67629 , n67630 , n67631 , n67632 , n67633 , n67634 , n67635 , n67636 , n67637 , n67638 , n67639 , n67640 , n67641 , n67642 , n67643 , n67644 , n67645 , n67646 , n67647 , n67648 , n67649 , n67650 , n67651 , n67652 , n67653 , n67654 , n67655 , n67656 , n67657 , n67658 , n67659 , n67660 , n67661 , n67662 , n67663 , n67664 , n67665 , n67666 , n67667 , n67668 , n67669 , n67670 , n67671 , n67672 , n67673 , n67674 , n67675 , n67676 , n67677 , n67678 , n67679 , n67680 , n67681 , n67682 , n67683 , n67684 , n67685 , n67686 , n67687 , n67688 , n67689 , n67690 , n67691 , n67692 , n67693 , n67694 , n67695 , n67696 , n67697 , n67698 , n67699 , n67700 , n67701 , n67702 , n67703 , n67704 , n67705 , n67706 , n67707 , n67708 , n67709 , n67710 , n67711 , n67712 , n67713 , n67714 , n67715 , n67716 , n67717 , n67718 , n67719 , n67720 , n67721 , n67722 , n67723 , n67724 , n67725 , n67726 , n67727 , n67728 , n67729 , n67730 , n67731 , n67732 , n67733 , n67734 , n67735 , n67736 , n67737 , n67738 , n67739 , n67740 , n67741 , n67742 , n67743 , n67744 , n67745 , n67746 , n67747 , n67748 , n67749 , n67750 , n67751 , n67752 , n67753 , n67754 , n67755 , n67756 , n67757 , n67758 , n67759 , n67760 , n67761 , n67762 , n67763 , n67764 , n67765 , n67766 , n67767 , n67768 , n67769 , n67770 , n67771 , n67772 , n67773 , n67774 , n67775 , n67776 , n67777 , n67778 , n67779 , n67780 , n67781 , n67782 , n67783 , n67784 , n67785 , n67786 , n67787 , n67788 , n67789 , n67790 , n67791 , n67792 , n67793 , n67794 , n67795 , n67796 , n67797 , n67798 , n67799 , n67800 , n67801 , n67802 , n67803 , n67804 , n67805 , n67806 , n67807 , n67808 , n67809 , n67810 , n67811 , n67812 , n67813 , n67814 , n67815 , n67816 , n67817 , n67818 , n67819 , n67820 , n67821 , n67822 , n67823 , n67824 , n67825 , n67826 , n67827 , n67828 , n67829 , n67830 , n67831 , n67832 , n67833 , n67834 , n67835 , n67836 , n67837 , n67838 , n67839 , n67840 , n67841 , n67842 , n67843 , n67844 , n67845 , n67846 , n67847 , n67848 , n67849 , n67850 , n67851 , n67852 , n67853 , n67854 , n67855 , n67856 , n67857 , n67858 , n67859 , n67860 , n67861 , n67862 , n67863 , n67864 , n67865 , n67866 , n67867 , n67868 , n67869 , n67870 , n67871 , n67872 , n67873 , n67874 , n67875 , n67876 , n67877 , n67878 , n67879 , n67880 , n67881 , n67882 , n67883 , n67884 , n67885 , n67886 , n67887 , n67888 , n67889 , n67890 , n67891 , n67892 , n67893 , n67894 , n67895 , n67896 , n67897 , n67898 , n67899 , n67900 , n67901 , n67902 , n67903 , n67904 , n67905 , n67906 , n67907 , n67908 , n67909 , n67910 , n67911 , n67912 , n67913 , n67914 , n67915 , n67916 , n67917 , n67918 , n67919 , n67920 , n67921 , n67922 , n67923 , n67924 , n67925 , n67926 , n67927 , n67928 , n67929 , n67930 , n67931 , n67932 , n67933 , n67934 , n67935 , n67936 , n67937 , n67938 , n67939 , n67940 , n67941 , n67942 , n67943 , n67944 , n67945 , n67946 , n67947 , n67948 , n67949 , n67950 , n67951 , n67952 , n67953 , n67954 , n67955 , n67956 , n67957 , n67958 , n67959 , n67960 , n67961 , n67962 , n67963 , n67964 , n67965 , n67966 , n67967 , n67968 , n67969 , n67970 , n67971 , n67972 , n67973 , n67974 , n67975 , n67976 , n67977 , n67978 , n67979 , n67980 , n67981 , n67982 , n67983 , n67984 , n67985 , n67986 , n67987 , n67988 , n67989 , n67990 , n67991 , n67992 , n67993 , n67994 , n67995 , n67996 , n67997 , n67998 , n67999 , n68000 , n68001 , n68002 , n68003 , n68004 , n68005 , n68006 , n68007 , n68008 , n68009 , n68010 , n68011 , n68012 , n68013 , n68014 , n68015 , n68016 , n68017 , n68018 , n68019 , n68020 , n68021 , n68022 , n68023 , n68024 , n68025 , n68026 , n68027 , n68028 , n68029 , n68030 , n68031 , n68032 , n68033 , n68034 , n68035 , n68036 , n68037 , n68038 , n68039 , n68040 , n68041 , n68042 , n68043 , n68044 , n68045 , n68046 , n68047 , n68048 , n68049 , n68050 , n68051 , n68052 , n68053 , n68054 , n68055 , n68056 , n68057 , n68058 , n68059 , n68060 , n68061 , n68062 , n68063 , n68064 , n68065 , n68066 , n68067 , n68068 , n68069 , n68070 , n68071 , n68072 , n68073 , n68074 , n68075 , n68076 , n68077 , n68078 , n68079 , n68080 , n68081 , n68082 , n68083 , n68084 , n68085 , n68086 , n68087 , n68088 , n68089 , n68090 , n68091 , n68092 , n68093 , n68094 , n68095 , n68096 , n68097 , n68098 , n68099 , n68100 , n68101 , n68102 , n68103 , n68104 , n68105 , n68106 , n68107 , n68108 , n68109 , n68110 , n68111 , n68112 , n68113 , n68114 , n68115 , n68116 , n68117 , n68118 , n68119 , n68120 , n68121 , n68122 , n68123 , n68124 , n68125 , n68126 , n68127 , n68128 , n68129 , n68130 , n68131 , n68132 , n68133 , n68134 , n68135 , n68136 , n68137 , n68138 , n68139 , n68140 , n68141 , n68142 , n68143 , n68144 , n68145 , n68146 , n68147 , n68148 , n68149 , n68150 , n68151 , n68152 , n68153 , n68154 , n68155 , n68156 , n68157 , n68158 , n68159 , n68160 , n68161 , n68162 , n68163 , n68164 , n68165 , n68166 , n68167 , n68168 , n68169 , n68170 , n68171 , n68172 , n68173 , n68174 , n68175 , n68176 , n68177 , n68178 , n68179 , n68180 , n68181 , n68182 , n68183 , n68184 , n68185 , n68186 , n68187 , n68188 , n68189 , n68190 , n68191 , n68192 , n68193 , n68194 , n68195 , n68196 , n68197 , n68198 , n68199 , n68200 , n68201 , n68202 , n68203 , n68204 , n68205 , n68206 , n68207 , n68208 , n68209 , n68210 , n68211 , n68212 , n68213 , n68214 , n68215 , n68216 , n68217 , n68218 , n68219 , n68220 , n68221 , n68222 , n68223 , n68224 , n68225 , n68226 , n68227 , n68228 , n68229 , n68230 , n68231 , n68232 , n68233 , n68234 , n68235 , n68236 , n68237 , n68238 , n68239 , n68240 , n68241 , n68242 , n68243 , n68244 , n68245 , n68246 , n68247 , n68248 , n68249 , n68250 , n68251 , n68252 , n68253 , n68254 , n68255 , n68256 , n68257 , n68258 , n68259 , n68260 , n68261 , n68262 , n68263 , n68264 , n68265 , n68266 , n68267 , n68268 , n68269 , n68270 , n68271 , n68272 , n68273 , n68274 , n68275 , n68276 , n68277 , n68278 , n68279 , n68280 , n68281 , n68282 , n68283 , n68284 , n68285 , n68286 , n68287 , n68288 , n68289 , n68290 , n68291 , n68292 , n68293 , n68294 , n68295 , n68296 , n68297 , n68298 , n68299 , n68300 , n68301 , n68302 , n68303 , n68304 , n68305 , n68306 , n68307 , n68308 , n68309 , n68310 , n68311 , n68312 , n68313 , n68314 , n68315 , n68316 , n68317 , n68318 , n68319 , n68320 , n68321 , n68322 , n68323 , n68324 , n68325 , n68326 , n68327 , n68328 , n68329 , n68330 , n68331 , n68332 , n68333 , n68334 , n68335 , n68336 , n68337 , n68338 , n68339 , n68340 , n68341 , n68342 , n68343 , n68344 , n68345 , n68346 , n68347 , n68348 , n68349 , n68350 , n68351 , n68352 , n68353 , n68354 , n68355 , n68356 , n68357 , n68358 , n68359 , n68360 , n68361 , n68362 , n68363 , n68364 , n68365 , n68366 , n68367 , n68368 , n68369 , n68370 , n68371 , n68372 , n68373 , n68374 , n68375 , n68376 , n68377 , n68378 , n68379 , n68380 , n68381 , n68382 , n68383 , n68384 , n68385 , n68386 , n68387 , n68388 , n68389 , n68390 , n68391 , n68392 , n68393 , n68394 , n68395 , n68396 , n68397 , n68398 , n68399 , n68400 , n68401 , n68402 , n68403 , n68404 , n68405 , n68406 , n68407 , n68408 , n68409 , n68410 , n68411 , n68412 , n68413 , n68414 , n68415 , n68416 , n68417 , n68418 , n68419 , n68420 , n68421 , n68422 , n68423 , n68424 , n68425 , n68426 , n68427 , n68428 , n68429 , n68430 , n68431 , n68432 , n68433 , n68434 , n68435 , n68436 , n68437 , n68438 , n68439 , n68440 , n68441 , n68442 , n68443 , n68444 , n68445 , n68446 , n68447 , n68448 , n68449 , n68450 , n68451 , n68452 , n68453 , n68454 , n68455 , n68456 , n68457 , n68458 , n68459 , n68460 , n68461 , n68462 , n68463 , n68464 , n68465 , n68466 , n68467 , n68468 , n68469 , n68470 , n68471 , n68472 , n68473 , n68474 , n68475 , n68476 , n68477 , n68478 , n68479 , n68480 , n68481 , n68482 , n68483 , n68484 , n68485 , n68486 , n68487 , n68488 , n68489 , n68490 , n68491 , n68492 , n68493 , n68494 , n68495 , n68496 , n68497 , n68498 , n68499 , n68500 , n68501 , n68502 , n68503 , n68504 , n68505 , n68506 , n68507 , n68508 , n68509 , n68510 , n68511 , n68512 , n68513 , n68514 , n68515 , n68516 , n68517 , n68518 , n68519 , n68520 , n68521 , n68522 , n68523 , n68524 , n68525 , n68526 , n68527 , n68528 , n68529 , n68530 , n68531 , n68532 , n68533 , n68534 , n68535 , n68536 , n68537 , n68538 , n68539 , n68540 , n68541 , n68542 , n68543 , n68544 , n68545 , n68546 , n68547 , n68548 , n68549 , n68550 , n68551 , n68552 , n68553 , n68554 , n68555 , n68556 , n68557 , n68558 , n68559 , n68560 , n68561 , n68562 , n68563 , n68564 , n68565 , n68566 , n68567 , n68568 , n68569 , n68570 , n68571 , n68572 , n68573 , n68574 , n68575 , n68576 , n68577 , n68578 , n68579 , n68580 , n68581 , n68582 , n68583 , n68584 , n68585 , n68586 , n68587 , n68588 , n68589 , n68590 , n68591 , n68592 , n68593 , n68594 , n68595 , n68596 , n68597 , n68598 , n68599 , n68600 , n68601 , n68602 , n68603 , n68604 , n68605 , n68606 , n68607 , n68608 , n68609 , n68610 , n68611 , n68612 , n68613 , n68614 , n68615 , n68616 , n68617 , n68618 , n68619 , n68620 , n68621 , n68622 , n68623 , n68624 , n68625 , n68626 , n68627 , n68628 , n68629 , n68630 , n68631 , n68632 , n68633 , n68634 , n68635 , n68636 , n68637 , n68638 , n68639 , n68640 , n68641 , n68642 , n68643 , n68644 , n68645 , n68646 , n68647 , n68648 , n68649 , n68650 , n68651 , n68652 , n68653 , n68654 , n68655 , n68656 , n68657 , n68658 , n68659 , n68660 , n68661 , n68662 , n68663 , n68664 , n68665 , n68666 , n68667 , n68668 , n68669 , n68670 , n68671 , n68672 , n68673 , n68674 , n68675 , n68676 , n68677 , n68678 , n68679 , n68680 , n68681 , n68682 , n68683 , n68684 , n68685 , n68686 , n68687 , n68688 , n68689 , n68690 , n68691 , n68692 , n68693 , n68694 , n68695 , n68696 , n68697 , n68698 , n68699 , n68700 , n68701 , n68702 , n68703 , n68704 , n68705 , n68706 , n68707 , n68708 , n68709 , n68710 , n68711 , n68712 , n68713 , n68714 , n68715 , n68716 , n68717 , n68718 , n68719 , n68720 , n68721 , n68722 , n68723 , n68724 , n68725 , n68726 , n68727 , n68728 , n68729 , n68730 , n68731 , n68732 , n68733 , n68734 , n68735 , n68736 , n68737 , n68738 , n68739 , n68740 , n68741 , n68742 , n68743 , n68744 , n68745 , n68746 , n68747 , n68748 , n68749 , n68750 , n68751 , n68752 , n68753 , n68754 , n68755 , n68756 , n68757 , n68758 , n68759 , n68760 , n68761 , n68762 , n68763 , n68764 , n68765 , n68766 , n68767 , n68768 , n68769 , n68770 , n68771 , n68772 , n68773 , n68774 , n68775 , n68776 , n68777 , n68778 , n68779 , n68780 , n68781 , n68782 , n68783 , n68784 , n68785 , n68786 , n68787 , n68788 , n68789 , n68790 , n68791 , n68792 , n68793 , n68794 , n68795 , n68796 , n68797 , n68798 , n68799 , n68800 , n68801 , n68802 , n68803 , n68804 , n68805 , n68806 , n68807 , n68808 , n68809 , n68810 , n68811 , n68812 , n68813 , n68814 , n68815 , n68816 , n68817 , n68818 , n68819 , n68820 , n68821 , n68822 , n68823 , n68824 , n68825 , n68826 , n68827 , n68828 , n68829 , n68830 , n68831 , n68832 , n68833 , n68834 , n68835 , n68836 , n68837 , n68838 , n68839 , n68840 , n68841 , n68842 , n68843 , n68844 , n68845 , n68846 , n68847 , n68848 , n68849 , n68850 , n68851 , n68852 , n68853 , n68854 , n68855 , n68856 , n68857 , n68858 , n68859 , n68860 , n68861 , n68862 , n68863 , n68864 , n68865 , n68866 , n68867 , n68868 , n68869 , n68870 , n68871 , n68872 , n68873 , n68874 , n68875 , n68876 , n68877 , n68878 , n68879 , n68880 , n68881 , n68882 , n68883 , n68884 , n68885 , n68886 , n68887 , n68888 , n68889 , n68890 , n68891 , n68892 , n68893 , n68894 , n68895 , n68896 , n68897 , n68898 , n68899 , n68900 , n68901 , n68902 , n68903 , n68904 , n68905 , n68906 , n68907 , n68908 , n68909 , n68910 , n68911 , n68912 , n68913 , n68914 , n68915 , n68916 , n68917 , n68918 , n68919 , n68920 , n68921 , n68922 , n68923 , n68924 , n68925 , n68926 , n68927 , n68928 , n68929 , n68930 , n68931 , n68932 , n68933 , n68934 , n68935 , n68936 , n68937 , n68938 , n68939 , n68940 , n68941 , n68942 , n68943 , n68944 , n68945 , n68946 , n68947 , n68948 , n68949 , n68950 , n68951 , n68952 , n68953 , n68954 , n68955 , n68956 , n68957 , n68958 , n68959 , n68960 , n68961 , n68962 , n68963 , n68964 , n68965 , n68966 , n68967 , n68968 , n68969 , n68970 , n68971 , n68972 , n68973 , n68974 , n68975 , n68976 , n68977 , n68978 , n68979 , n68980 , n68981 , n68982 , n68983 , n68984 , n68985 , n68986 , n68987 , n68988 , n68989 , n68990 , n68991 , n68992 , n68993 , n68994 , n68995 , n68996 , n68997 , n68998 , n68999 , n69000 , n69001 , n69002 , n69003 , n69004 , n69005 , n69006 , n69007 , n69008 , n69009 , n69010 , n69011 , n69012 , n69013 , n69014 , n69015 , n69016 , n69017 , n69018 , n69019 , n69020 , n69021 , n69022 , n69023 , n69024 , n69025 , n69026 , n69027 , n69028 , n69029 , n69030 , n69031 , n69032 , n69033 , n69034 , n69035 , n69036 , n69037 , n69038 , n69039 , n69040 , n69041 , n69042 , n69043 , n69044 , n69045 , n69046 , n69047 , n69048 , n69049 , n69050 , n69051 , n69052 , n69053 , n69054 , n69055 , n69056 , n69057 , n69058 , n69059 , n69060 , n69061 , n69062 , n69063 , n69064 , n69065 , n69066 , n69067 , n69068 , n69069 , n69070 , n69071 , n69072 , n69073 , n69074 , n69075 , n69076 , n69077 , n69078 , n69079 , n69080 , n69081 , n69082 , n69083 , n69084 , n69085 , n69086 , n69087 , n69088 , n69089 , n69090 , n69091 , n69092 , n69093 , n69094 , n69095 , n69096 , n69097 , n69098 , n69099 , n69100 , n69101 , n69102 , n69103 , n69104 , n69105 , n69106 , n69107 , n69108 , n69109 , n69110 , n69111 , n69112 , n69113 , n69114 , n69115 , n69116 , n69117 , n69118 , n69119 , n69120 , n69121 , n69122 , n69123 , n69124 , n69125 , n69126 , n69127 , n69128 , n69129 , n69130 , n69131 , n69132 , n69133 , n69134 , n69135 , n69136 , n69137 , n69138 , n69139 , n69140 , n69141 , n69142 , n69143 , n69144 , n69145 , n69146 , n69147 , n69148 , n69149 , n69150 , n69151 , n69152 , n69153 , n69154 , n69155 , n69156 , n69157 , n69158 , n69159 , n69160 , n69161 , n69162 , n69163 , n69164 , n69165 , n69166 , n69167 , n69168 , n69169 , n69170 , n69171 , n69172 , n69173 , n69174 , n69175 , n69176 , n69177 , n69178 , n69179 , n69180 , n69181 , n69182 , n69183 , n69184 , n69185 , n69186 , n69187 , n69188 , n69189 , n69190 , n69191 , n69192 , n69193 , n69194 , n69195 , n69196 , n69197 , n69198 , n69199 , n69200 , n69201 , n69202 , n69203 , n69204 , n69205 , n69206 , n69207 , n69208 , n69209 , n69210 , n69211 , n69212 , n69213 , n69214 , n69215 , n69216 , n69217 , n69218 , n69219 , n69220 , n69221 , n69222 , n69223 , n69224 , n69225 , n69226 , n69227 , n69228 , n69229 , n69230 , n69231 , n69232 , n69233 , n69234 , n69235 , n69236 , n69237 , n69238 , n69239 , n69240 , n69241 , n69242 , n69243 , n69244 , n69245 , n69246 , n69247 , n69248 , n69249 , n69250 , n69251 , n69252 , n69253 , n69254 , n69255 , n69256 , n69257 , n69258 , n69259 , n69260 , n69261 , n69262 , n69263 , n69264 , n69265 , n69266 , n69267 , n69268 , n69269 , n69270 , n69271 , n69272 , n69273 , n69274 , n69275 , n69276 , n69277 , n69278 , n69279 , n69280 , n69281 , n69282 , n69283 , n69284 , n69285 , n69286 , n69287 , n69288 , n69289 , n69290 , n69291 , n69292 , n69293 , n69294 , n69295 , n69296 , n69297 , n69298 , n69299 , n69300 , n69301 , n69302 , n69303 , n69304 , n69305 , n69306 , n69307 , n69308 , n69309 , n69310 , n69311 , n69312 , n69313 , n69314 , n69315 , n69316 , n69317 , n69318 , n69319 , n69320 , n69321 , n69322 , n69323 , n69324 , n69325 , n69326 , n69327 , n69328 , n69329 , n69330 , n69331 , n69332 , n69333 , n69334 , n69335 , n69336 , n69337 , n69338 , n69339 , n69340 , n69341 , n69342 , n69343 , n69344 , n69345 , n69346 , n69347 , n69348 , n69349 , n69350 , n69351 , n69352 , n69353 , n69354 , n69355 , n69356 , n69357 , n69358 , n69359 , n69360 , n69361 , n69362 , n69363 , n69364 , n69365 , n69366 , n69367 , n69368 , n69369 , n69370 , n69371 , n69372 , n69373 , n69374 , n69375 , n69376 , n69377 , n69378 , n69379 , n69380 , n69381 , n69382 , n69383 , n69384 , n69385 , n69386 , n69387 , n69388 , n69389 , n69390 , n69391 , n69392 , n69393 , n69394 , n69395 , n69396 , n69397 , n69398 , n69399 , n69400 , n69401 , n69402 , n69403 , n69404 , n69405 , n69406 , n69407 , n69408 , n69409 , n69410 , n69411 , n69412 , n69413 , n69414 , n69415 , n69416 , n69417 , n69418 , n69419 , n69420 , n69421 , n69422 , n69423 , n69424 , n69425 , n69426 , n69427 , n69428 , n69429 , n69430 , n69431 , n69432 , n69433 , n69434 , n69435 , n69436 , n69437 , n69438 , n69439 , n69440 , n69441 , n69442 , n69443 , n69444 , n69445 , n69446 , n69447 , n69448 , n69449 , n69450 , n69451 , n69452 , n69453 , n69454 , n69455 , n69456 , n69457 , n69458 , n69459 , n69460 , n69461 , n69462 , n69463 , n69464 , n69465 , n69466 , n69467 , n69468 , n69469 , n69470 , n69471 , n69472 , n69473 , n69474 , n69475 , n69476 , n69477 , n69478 , n69479 , n69480 , n69481 , n69482 , n69483 , n69484 , n69485 , n69486 , n69487 , n69488 , n69489 , n69490 , n69491 , n69492 , n69493 , n69494 , n69495 , n69496 , n69497 , n69498 , n69499 , n69500 , n69501 , n69502 , n69503 , n69504 , n69505 , n69506 , n69507 , n69508 , n69509 , n69510 , n69511 , n69512 , n69513 , n69514 , n69515 , n69516 , n69517 , n69518 , n69519 , n69520 , n69521 , n69522 , n69523 , n69524 , n69525 , n69526 , n69527 , n69528 , n69529 , n69530 , n69531 , n69532 , n69533 , n69534 , n69535 , n69536 , n69537 , n69538 , n69539 , n69540 , n69541 , n69542 , n69543 , n69544 , n69545 , n69546 , n69547 , n69548 , n69549 , n69550 , n69551 , n69552 , n69553 , n69554 , n69555 , n69556 , n69557 , n69558 , n69559 , n69560 , n69561 , n69562 , n69563 , n69564 , n69565 , n69566 , n69567 , n69568 , n69569 , n69570 , n69571 , n69572 , n69573 , n69574 , n69575 , n69576 , n69577 , n69578 , n69579 , n69580 , n69581 , n69582 , n69583 , n69584 , n69585 , n69586 , n69587 , n69588 , n69589 , n69590 , n69591 , n69592 , n69593 , n69594 , n69595 , n69596 , n69597 , n69598 , n69599 , n69600 , n69601 , n69602 , n69603 , n69604 , n69605 , n69606 , n69607 , n69608 , n69609 , n69610 , n69611 , n69612 , n69613 , n69614 , n69615 , n69616 , n69617 , n69618 , n69619 , n69620 , n69621 , n69622 , n69623 , n69624 , n69625 , n69626 , n69627 , n69628 , n69629 , n69630 , n69631 , n69632 , n69633 , n69634 , n69635 , n69636 , n69637 , n69638 , n69639 , n69640 , n69641 , n69642 , n69643 , n69644 , n69645 , n69646 , n69647 , n69648 , n69649 , n69650 , n69651 , n69652 , n69653 , n69654 , n69655 , n69656 , n69657 , n69658 , n69659 , n69660 , n69661 , n69662 , n69663 , n69664 , n69665 , n69666 , n69667 , n69668 , n69669 , n69670 , n69671 , n69672 , n69673 , n69674 , n69675 , n69676 , n69677 , n69678 , n69679 , n69680 , n69681 , n69682 , n69683 , n69684 , n69685 , n69686 , n69687 , n69688 , n69689 , n69690 , n69691 , n69692 , n69693 , n69694 , n69695 , n69696 , n69697 , n69698 , n69699 , n69700 , n69701 , n69702 , n69703 , n69704 , n69705 , n69706 , n69707 , n69708 , n69709 , n69710 , n69711 , n69712 , n69713 , n69714 , n69715 , n69716 , n69717 , n69718 , n69719 , n69720 , n69721 , n69722 , n69723 , n69724 , n69725 , n69726 , n69727 , n69728 , n69729 , n69730 , n69731 , n69732 , n69733 , n69734 , n69735 , n69736 , n69737 , n69738 , n69739 , n69740 , n69741 , n69742 , n69743 , n69744 , n69745 , n69746 , n69747 , n69748 , n69749 , n69750 , n69751 , n69752 , n69753 , n69754 , n69755 , n69756 , n69757 , n69758 , n69759 , n69760 , n69761 , n69762 , n69763 , n69764 , n69765 , n69766 , n69767 , n69768 , n69769 , n69770 , n69771 , n69772 , n69773 , n69774 , n69775 , n69776 , n69777 , n69778 , n69779 , n69780 , n69781 , n69782 , n69783 , n69784 , n69785 , n69786 , n69787 , n69788 , n69789 , n69790 , n69791 , n69792 , n69793 , n69794 , n69795 , n69796 , n69797 , n69798 , n69799 , n69800 , n69801 , n69802 , n69803 , n69804 , n69805 , n69806 , n69807 , n69808 , n69809 , n69810 , n69811 , n69812 , n69813 , n69814 , n69815 , n69816 , n69817 , n69818 , n69819 , n69820 , n69821 , n69822 , n69823 , n69824 , n69825 , n69826 , n69827 , n69828 , n69829 , n69830 , n69831 , n69832 , n69833 , n69834 , n69835 , n69836 , n69837 , n69838 , n69839 , n69840 , n69841 , n69842 , n69843 , n69844 , n69845 , n69846 , n69847 , n69848 , n69849 , n69850 , n69851 , n69852 , n69853 , n69854 , n69855 , n69856 , n69857 , n69858 , n69859 , n69860 , n69861 , n69862 , n69863 , n69864 , n69865 , n69866 , n69867 , n69868 , n69869 , n69870 , n69871 , n69872 , n69873 , n69874 , n69875 , n69876 , n69877 , n69878 , n69879 , n69880 , n69881 , n69882 , n69883 , n69884 , n69885 , n69886 , n69887 , n69888 , n69889 , n69890 , n69891 , n69892 , n69893 , n69894 , n69895 , n69896 , n69897 , n69898 , n69899 , n69900 , n69901 , n69902 , n69903 , n69904 , n69905 , n69906 , n69907 , n69908 , n69909 , n69910 , n69911 , n69912 , n69913 , n69914 , n69915 , n69916 , n69917 , n69918 , n69919 , n69920 , n69921 , n69922 , n69923 , n69924 , n69925 , n69926 , n69927 , n69928 , n69929 , n69930 , n69931 , n69932 , n69933 , n69934 , n69935 , n69936 , n69937 , n69938 , n69939 , n69940 , n69941 , n69942 , n69943 , n69944 , n69945 , n69946 , n69947 , n69948 , n69949 , n69950 , n69951 , n69952 , n69953 , n69954 , n69955 , n69956 , n69957 , n69958 , n69959 , n69960 , n69961 , n69962 , n69963 , n69964 , n69965 , n69966 , n69967 , n69968 , n69969 , n69970 , n69971 , n69972 , n69973 , n69974 , n69975 , n69976 , n69977 , n69978 , n69979 , n69980 , n69981 , n69982 , n69983 , n69984 , n69985 , n69986 , n69987 , n69988 , n69989 , n69990 , n69991 , n69992 , n69993 , n69994 , n69995 , n69996 , n69997 , n69998 , n69999 , n70000 , n70001 , n70002 , n70003 , n70004 , n70005 , n70006 , n70007 , n70008 , n70009 , n70010 , n70011 , n70012 , n70013 , n70014 , n70015 , n70016 , n70017 , n70018 , n70019 , n70020 , n70021 , n70022 , n70023 , n70024 , n70025 , n70026 , n70027 , n70028 , n70029 , n70030 , n70031 , n70032 , n70033 , n70034 , n70035 , n70036 , n70037 , n70038 , n70039 , n70040 , n70041 , n70042 , n70043 , n70044 , n70045 , n70046 , n70047 , n70048 , n70049 , n70050 , n70051 , n70052 , n70053 , n70054 , n70055 , n70056 , n70057 , n70058 , n70059 , n70060 , n70061 , n70062 , n70063 , n70064 , n70065 , n70066 , n70067 , n70068 , n70069 , n70070 , n70071 , n70072 , n70073 , n70074 , n70075 , n70076 , n70077 , n70078 , n70079 , n70080 , n70081 , n70082 , n70083 , n70084 , n70085 , n70086 , n70087 , n70088 , n70089 , n70090 , n70091 , n70092 , n70093 , n70094 , n70095 , n70096 , n70097 , n70098 , n70099 , n70100 , n70101 , n70102 , n70103 , n70104 , n70105 , n70106 , n70107 , n70108 , n70109 , n70110 , n70111 , n70112 , n70113 , n70114 , n70115 , n70116 , n70117 , n70118 , n70119 , n70120 , n70121 , n70122 , n70123 , n70124 , n70125 , n70126 , n70127 , n70128 , n70129 , n70130 , n70131 , n70132 , n70133 , n70134 , n70135 , n70136 , n70137 , n70138 , n70139 , n70140 , n70141 , n70142 , n70143 , n70144 , n70145 , n70146 , n70147 , n70148 , n70149 , n70150 , n70151 , n70152 , n70153 , n70154 , n70155 , n70156 , n70157 , n70158 , n70159 , n70160 , n70161 , n70162 , n70163 , n70164 , n70165 , n70166 , n70167 , n70168 , n70169 , n70170 , n70171 , n70172 , n70173 , n70174 , n70175 , n70176 , n70177 , n70178 , n70179 , n70180 , n70181 , n70182 , n70183 , n70184 , n70185 , n70186 , n70187 , n70188 , n70189 , n70190 , n70191 , n70192 , n70193 , n70194 , n70195 , n70196 , n70197 , n70198 , n70199 , n70200 , n70201 , n70202 , n70203 , n70204 , n70205 , n70206 , n70207 , n70208 , n70209 , n70210 , n70211 , n70212 , n70213 , n70214 , n70215 , n70216 , n70217 , n70218 , n70219 , n70220 , n70221 , n70222 , n70223 , n70224 , n70225 , n70226 , n70227 , n70228 , n70229 , n70230 , n70231 , n70232 , n70233 , n70234 , n70235 , n70236 , n70237 , n70238 , n70239 , n70240 , n70241 , n70242 , n70243 , n70244 , n70245 , n70246 , n70247 , n70248 , n70249 , n70250 , n70251 , n70252 , n70253 , n70254 , n70255 , n70256 , n70257 , n70258 , n70259 , n70260 , n70261 , n70262 , n70263 , n70264 , n70265 , n70266 , n70267 , n70268 , n70269 , n70270 , n70271 , n70272 , n70273 , n70274 , n70275 , n70276 , n70277 , n70278 , n70279 , n70280 , n70281 , n70282 , n70283 , n70284 , n70285 , n70286 , n70287 , n70288 , n70289 , n70290 , n70291 , n70292 , n70293 , n70294 , n70295 , n70296 , n70297 , n70298 , n70299 , n70300 , n70301 , n70302 , n70303 , n70304 , n70305 , n70306 , n70307 , n70308 , n70309 , n70310 , n70311 , n70312 , n70313 , n70314 , n70315 , n70316 , n70317 , n70318 , n70319 , n70320 , n70321 , n70322 , n70323 , n70324 , n70325 , n70326 , n70327 , n70328 , n70329 , n70330 , n70331 , n70332 , n70333 , n70334 , n70335 , n70336 , n70337 , n70338 , n70339 , n70340 , n70341 , n70342 , n70343 , n70344 , n70345 , n70346 , n70347 , n70348 , n70349 , n70350 , n70351 , n70352 , n70353 , n70354 , n70355 , n70356 , n70357 , n70358 , n70359 , n70360 , n70361 , n70362 , n70363 , n70364 , n70365 , n70366 , n70367 , n70368 , n70369 , n70370 , n70371 , n70372 , n70373 , n70374 , n70375 , n70376 , n70377 , n70378 , n70379 , n70380 , n70381 , n70382 , n70383 , n70384 , n70385 , n70386 , n70387 , n70388 , n70389 , n70390 , n70391 , n70392 , n70393 , n70394 , n70395 , n70396 , n70397 , n70398 , n70399 , n70400 , n70401 , n70402 , n70403 , n70404 , n70405 , n70406 , n70407 , n70408 , n70409 , n70410 , n70411 , n70412 , n70413 , n70414 , n70415 , n70416 , n70417 , n70418 , n70419 , n70420 , n70421 , n70422 , n70423 , n70424 , n70425 , n70426 , n70427 , n70428 , n70429 , n70430 , n70431 , n70432 , n70433 , n70434 , n70435 , n70436 , n70437 , n70438 , n70439 , n70440 , n70441 , n70442 , n70443 , n70444 , n70445 , n70446 , n70447 , n70448 , n70449 , n70450 , n70451 , n70452 , n70453 , n70454 , n70455 , n70456 , n70457 , n70458 , n70459 , n70460 , n70461 , n70462 , n70463 , n70464 , n70465 , n70466 , n70467 , n70468 , n70469 , n70470 , n70471 , n70472 , n70473 , n70474 , n70475 , n70476 , n70477 , n70478 , n70479 , n70480 , n70481 , n70482 , n70483 , n70484 , n70485 , n70486 , n70487 , n70488 , n70489 , n70490 , n70491 , n70492 , n70493 , n70494 , n70495 , n70496 , n70497 , n70498 , n70499 , n70500 , n70501 , n70502 , n70503 , n70504 , n70505 , n70506 , n70507 , n70508 , n70509 , n70510 , n70511 , n70512 , n70513 , n70514 , n70515 , n70516 , n70517 , n70518 , n70519 , n70520 , n70521 , n70522 , n70523 , n70524 , n70525 , n70526 , n70527 , n70528 , n70529 , n70530 , n70531 , n70532 , n70533 , n70534 , n70535 , n70536 , n70537 , n70538 , n70539 , n70540 , n70541 , n70542 , n70543 , n70544 , n70545 , n70546 , n70547 , n70548 , n70549 , n70550 , n70551 , n70552 , n70553 , n70554 , n70555 , n70556 , n70557 , n70558 , n70559 , n70560 , n70561 , n70562 , n70563 , n70564 , n70565 , n70566 , n70567 , n70568 , n70569 , n70570 , n70571 , n70572 , n70573 , n70574 , n70575 , n70576 , n70577 , n70578 , n70579 , n70580 , n70581 , n70582 , n70583 , n70584 , n70585 , n70586 , n70587 , n70588 , n70589 , n70590 , n70591 , n70592 , n70593 , n70594 , n70595 , n70596 , n70597 , n70598 , n70599 , n70600 , n70601 , n70602 , n70603 , n70604 , n70605 , n70606 , n70607 , n70608 , n70609 , n70610 , n70611 , n70612 , n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , n70619 , n70620 , n70621 , n70622 , n70623 , n70624 , n70625 , n70626 , n70627 , n70628 , n70629 , n70630 , n70631 , n70632 , n70633 , n70634 , n70635 , n70636 , n70637 , n70638 , n70639 , n70640 , n70641 , n70642 , n70643 , n70644 , n70645 , n70646 , n70647 , n70648 , n70649 , n70650 , n70651 , n70652 , n70653 , n70654 , n70655 , n70656 , n70657 , n70658 , n70659 , n70660 , n70661 , n70662 , n70663 , n70664 , n70665 , n70666 , n70667 , n70668 , n70669 , n70670 , n70671 , n70672 , n70673 , n70674 , n70675 , n70676 , n70677 , n70678 , n70679 , n70680 , n70681 , n70682 , n70683 , n70684 , n70685 , n70686 , n70687 , n70688 , n70689 , n70690 , n70691 , n70692 , n70693 , n70694 , n70695 , n70696 , n70697 , n70698 , n70699 , n70700 , n70701 , n70702 , n70703 , n70704 , n70705 , n70706 , n70707 , n70708 , n70709 , n70710 , n70711 , n70712 , n70713 , n70714 , n70715 , n70716 , n70717 , n70718 , n70719 , n70720 , n70721 , n70722 , n70723 , n70724 , n70725 , n70726 , n70727 , n70728 , n70729 , n70730 , n70731 , n70732 , n70733 , n70734 , n70735 , n70736 , n70737 , n70738 , n70739 , n70740 , n70741 , n70742 , n70743 , n70744 , n70745 , n70746 , n70747 , n70748 , n70749 , n70750 , n70751 , n70752 , n70753 , n70754 , n70755 , n70756 , n70757 , n70758 , n70759 , n70760 , n70761 , n70762 , n70763 , n70764 , n70765 , n70766 , n70767 , n70768 , n70769 , n70770 , n70771 , n70772 , n70773 , n70774 , n70775 , n70776 , n70777 , n70778 , n70779 , n70780 , n70781 , n70782 , n70783 , n70784 , n70785 , n70786 , n70787 , n70788 , n70789 , n70790 , n70791 , n70792 , n70793 , n70794 , n70795 , n70796 , n70797 , n70798 , n70799 , n70800 , n70801 , n70802 , n70803 , n70804 , n70805 , n70806 , n70807 , n70808 , n70809 , n70810 , n70811 , n70812 , n70813 , n70814 , n70815 , n70816 , n70817 , n70818 , n70819 , n70820 , n70821 , n70822 , n70823 , n70824 , n70825 , n70826 , n70827 , n70828 , n70829 , n70830 , n70831 , n70832 , n70833 , n70834 , n70835 , n70836 , n70837 , n70838 , n70839 , n70840 , n70841 , n70842 , n70843 , n70844 , n70845 , n70846 , n70847 , n70848 , n70849 , n70850 , n70851 , n70852 , n70853 , n70854 , n70855 , n70856 , n70857 , n70858 , n70859 , n70860 , n70861 , n70862 , n70863 , n70864 , n70865 , n70866 , n70867 , n70868 , n70869 , n70870 , n70871 , n70872 , n70873 , n70874 , n70875 , n70876 , n70877 , n70878 , n70879 , n70880 , n70881 , n70882 , n70883 , n70884 , n70885 , n70886 , n70887 , n70888 , n70889 , n70890 , n70891 , n70892 , n70893 , n70894 , n70895 , n70896 , n70897 , n70898 , n70899 , n70900 , n70901 , n70902 , n70903 , n70904 , n70905 , n70906 , n70907 , n70908 , n70909 , n70910 , n70911 , n70912 , n70913 , n70914 , n70915 , n70916 , n70917 , n70918 , n70919 , n70920 , n70921 , n70922 , n70923 , n70924 , n70925 , n70926 , n70927 , n70928 , n70929 , n70930 , n70931 , n70932 , n70933 , n70934 , n70935 , n70936 , n70937 , n70938 , n70939 , n70940 , n70941 , n70942 , n70943 , n70944 , n70945 , n70946 , n70947 , n70948 , n70949 , n70950 , n70951 , n70952 , n70953 , n70954 , n70955 , n70956 , n70957 , n70958 , n70959 , n70960 , n70961 , n70962 , n70963 , n70964 , n70965 , n70966 , n70967 , n70968 , n70969 , n70970 , n70971 , n70972 , n70973 , n70974 , n70975 , n70976 , n70977 , n70978 , n70979 , n70980 , n70981 , n70982 , n70983 , n70984 , n70985 , n70986 , n70987 , n70988 , n70989 , n70990 , n70991 , n70992 , n70993 , n70994 , n70995 , n70996 , n70997 , n70998 , n70999 , n71000 , n71001 , n71002 , n71003 , n71004 , n71005 , n71006 , n71007 , n71008 , n71009 , n71010 , n71011 , n71012 , n71013 , n71014 , n71015 , n71016 , n71017 , n71018 , n71019 , n71020 , n71021 , n71022 , n71023 , n71024 , n71025 , n71026 , n71027 , n71028 , n71029 , n71030 , n71031 , n71032 , n71033 , n71034 , n71035 , n71036 , n71037 , n71038 , n71039 , n71040 , n71041 , n71042 , n71043 , n71044 , n71045 , n71046 , n71047 , n71048 , n71049 , n71050 , n71051 , n71052 , n71053 , n71054 , n71055 , n71056 , n71057 , n71058 , n71059 , n71060 , n71061 , n71062 , n71063 , n71064 , n71065 , n71066 , n71067 , n71068 , n71069 , n71070 , n71071 , n71072 , n71073 , n71074 , n71075 , n71076 , n71077 , n71078 , n71079 , n71080 , n71081 , n71082 , n71083 , n71084 , n71085 , n71086 , n71087 , n71088 , n71089 , n71090 , n71091 , n71092 , n71093 , n71094 , n71095 , n71096 , n71097 , n71098 , n71099 , n71100 , n71101 , n71102 , n71103 , n71104 , n71105 , n71106 , n71107 , n71108 , n71109 , n71110 , n71111 , n71112 , n71113 , n71114 , n71115 , n71116 , n71117 , n71118 , n71119 , n71120 , n71121 , n71122 , n71123 , n71124 , n71125 , n71126 , n71127 , n71128 , n71129 , n71130 , n71131 , n71132 , n71133 , n71134 , n71135 , n71136 , n71137 , n71138 , n71139 , n71140 , n71141 , n71142 , n71143 , n71144 , n71145 , n71146 , n71147 , n71148 , n71149 , n71150 , n71151 , n71152 , n71153 , n71154 , n71155 , n71156 , n71157 , n71158 , n71159 , n71160 , n71161 , n71162 , n71163 , n71164 , n71165 , n71166 , n71167 , n71168 , n71169 , n71170 , n71171 , n71172 , n71173 , n71174 , n71175 , n71176 , n71177 , n71178 , n71179 , n71180 , n71181 , n71182 , n71183 , n71184 , n71185 , n71186 , n71187 , n71188 , n71189 , n71190 , n71191 , n71192 , n71193 , n71194 , n71195 , n71196 , n71197 , n71198 , n71199 , n71200 , n71201 , n71202 , n71203 , n71204 , n71205 , n71206 , n71207 , n71208 , n71209 , n71210 , n71211 , n71212 , n71213 , n71214 , n71215 , n71216 , n71217 , n71218 , n71219 , n71220 , n71221 , n71222 , n71223 , n71224 , n71225 , n71226 , n71227 , n71228 , n71229 , n71230 , n71231 , n71232 , n71233 , n71234 , n71235 , n71236 , n71237 , n71238 , n71239 , n71240 , n71241 , n71242 , n71243 , n71244 , n71245 , n71246 , n71247 , n71248 , n71249 , n71250 , n71251 , n71252 , n71253 , n71254 , n71255 , n71256 , n71257 , n71258 , n71259 , n71260 , n71261 , n71262 , n71263 , n71264 , n71265 , n71266 , n71267 , n71268 , n71269 , n71270 , n71271 , n71272 , n71273 , n71274 , n71275 , n71276 , n71277 , n71278 , n71279 , n71280 , n71281 , n71282 , n71283 , n71284 , n71285 , n71286 , n71287 , n71288 , n71289 , n71290 , n71291 , n71292 , n71293 , n71294 , n71295 , n71296 , n71297 , n71298 , n71299 , n71300 , n71301 , n71302 , n71303 , n71304 , n71305 , n71306 , n71307 , n71308 , n71309 , n71310 , n71311 , n71312 , n71313 , n71314 , n71315 , n71316 , n71317 , n71318 , n71319 , n71320 , n71321 , n71322 , n71323 , n71324 , n71325 , n71326 , n71327 , n71328 , n71329 , n71330 , n71331 , n71332 , n71333 , n71334 , n71335 , n71336 , n71337 , n71338 , n71339 , n71340 , n71341 , n71342 , n71343 , n71344 , n71345 , n71346 , n71347 , n71348 , n71349 , n71350 , n71351 , n71352 , n71353 , n71354 , n71355 , n71356 , n71357 , n71358 , n71359 , n71360 , n71361 , n71362 , n71363 , n71364 , n71365 , n71366 , n71367 , n71368 , n71369 , n71370 , n71371 , n71372 , n71373 , n71374 , n71375 , n71376 , n71377 , n71378 , n71379 , n71380 , n71381 , n71382 , n71383 , n71384 , n71385 , n71386 , n71387 , n71388 , n71389 , n71390 , n71391 , n71392 , n71393 , n71394 , n71395 , n71396 , n71397 , n71398 , n71399 , n71400 , n71401 , n71402 , n71403 , n71404 , n71405 , n71406 , n71407 , n71408 , n71409 , n71410 , n71411 , n71412 , n71413 , n71414 , n71415 , n71416 , n71417 , n71418 , n71419 , n71420 , n71421 , n71422 , n71423 , n71424 , n71425 , n71426 , n71427 , n71428 , n71429 , n71430 , n71431 , n71432 , n71433 , n71434 , n71435 , n71436 , n71437 , n71438 , n71439 , n71440 , n71441 , n71442 , n71443 , n71444 , n71445 , n71446 , n71447 , n71448 , n71449 , n71450 , n71451 , n71452 , n71453 , n71454 , n71455 , n71456 , n71457 , n71458 , n71459 , n71460 , n71461 , n71462 , n71463 , n71464 , n71465 , n71466 , n71467 , n71468 , n71469 , n71470 , n71471 , n71472 , n71473 , n71474 , n71475 , n71476 , n71477 , n71478 , n71479 , n71480 , n71481 , n71482 , n71483 , n71484 , n71485 , n71486 , n71487 , n71488 , n71489 , n71490 , n71491 , n71492 , n71493 , n71494 , n71495 , n71496 , n71497 , n71498 , n71499 , n71500 , n71501 , n71502 , n71503 , n71504 , n71505 , n71506 , n71507 , n71508 , n71509 , n71510 , n71511 , n71512 , n71513 , n71514 , n71515 , n71516 , n71517 , n71518 , n71519 , n71520 , n71521 , n71522 , n71523 , n71524 , n71525 , n71526 , n71527 , n71528 , n71529 , n71530 , n71531 , n71532 , n71533 , n71534 , n71535 , n71536 , n71537 , n71538 , n71539 , n71540 , n71541 , n71542 , n71543 , n71544 , n71545 , n71546 , n71547 , n71548 , n71549 , n71550 , n71551 , n71552 , n71553 , n71554 , n71555 , n71556 , n71557 , n71558 , n71559 , n71560 , n71561 , n71562 , n71563 , n71564 , n71565 , n71566 , n71567 , n71568 , n71569 , n71570 , n71571 , n71572 , n71573 , n71574 , n71575 , n71576 , n71577 , n71578 , n71579 , n71580 , n71581 , n71582 , n71583 , n71584 , n71585 , n71586 , n71587 , n71588 , n71589 , n71590 , n71591 , n71592 , n71593 , n71594 , n71595 , n71596 , n71597 , n71598 , n71599 , n71600 , n71601 , n71602 , n71603 , n71604 , n71605 , n71606 , n71607 , n71608 , n71609 , n71610 , n71611 , n71612 , n71613 , n71614 , n71615 , n71616 , n71617 , n71618 , n71619 , n71620 , n71621 , n71622 , n71623 , n71624 , n71625 , n71626 , n71627 , n71628 , n71629 , n71630 , n71631 , n71632 , n71633 , n71634 , n71635 , n71636 , n71637 , n71638 , n71639 , n71640 , n71641 , n71642 , n71643 , n71644 , n71645 , n71646 , n71647 , n71648 , n71649 , n71650 , n71651 , n71652 , n71653 , n71654 , n71655 , n71656 , n71657 , n71658 , n71659 , n71660 , n71661 , n71662 , n71663 , n71664 , n71665 , n71666 , n71667 , n71668 , n71669 , n71670 , n71671 , n71672 , n71673 , n71674 , n71675 , n71676 , n71677 , n71678 , n71679 , n71680 , n71681 , n71682 , n71683 , n71684 , n71685 , n71686 , n71687 , n71688 , n71689 , n71690 , n71691 , n71692 , n71693 , n71694 , n71695 , n71696 , n71697 , n71698 , n71699 , n71700 , n71701 , n71702 , n71703 , n71704 , n71705 , n71706 , n71707 , n71708 , n71709 , n71710 , n71711 , n71712 , n71713 , n71714 , n71715 , n71716 , n71717 , n71718 , n71719 , n71720 , n71721 , n71722 , n71723 , n71724 , n71725 , n71726 , n71727 , n71728 , n71729 , n71730 , n71731 , n71732 , n71733 , n71734 , n71735 , n71736 , n71737 , n71738 , n71739 , n71740 , n71741 , n71742 , n71743 , n71744 , n71745 , n71746 , n71747 , n71748 , n71749 , n71750 , n71751 , n71752 , n71753 , n71754 , n71755 , n71756 , n71757 , n71758 , n71759 , n71760 , n71761 , n71762 , n71763 , n71764 , n71765 , n71766 , n71767 , n71768 , n71769 , n71770 , n71771 , n71772 , n71773 , n71774 , n71775 , n71776 , n71777 , n71778 , n71779 , n71780 , n71781 , n71782 , n71783 , n71784 , n71785 , n71786 , n71787 , n71788 , n71789 , n71790 , n71791 , n71792 , n71793 , n71794 , n71795 , n71796 , n71797 , n71798 , n71799 , n71800 , n71801 , n71802 , n71803 , n71804 , n71805 , n71806 , n71807 , n71808 , n71809 , n71810 , n71811 , n71812 , n71813 , n71814 , n71815 , n71816 , n71817 , n71818 , n71819 , n71820 , n71821 , n71822 , n71823 , n71824 , n71825 , n71826 , n71827 , n71828 , n71829 , n71830 , n71831 , n71832 , n71833 , n71834 , n71835 , n71836 , n71837 , n71838 , n71839 , n71840 , n71841 , n71842 , n71843 , n71844 , n71845 , n71846 , n71847 , n71848 , n71849 , n71850 , n71851 , n71852 , n71853 , n71854 , n71855 , n71856 , n71857 , n71858 , n71859 , n71860 , n71861 , n71862 , n71863 , n71864 , n71865 , n71866 , n71867 , n71868 , n71869 , n71870 , n71871 , n71872 , n71873 , n71874 , n71875 , n71876 , n71877 , n71878 , n71879 , n71880 , n71881 , n71882 , n71883 , n71884 , n71885 , n71886 , n71887 , n71888 , n71889 , n71890 , n71891 , n71892 , n71893 , n71894 , n71895 , n71896 , n71897 , n71898 , n71899 , n71900 , n71901 , n71902 , n71903 , n71904 , n71905 , n71906 , n71907 , n71908 , n71909 , n71910 , n71911 , n71912 , n71913 , n71914 , n71915 , n71916 , n71917 , n71918 , n71919 , n71920 , n71921 , n71922 , n71923 , n71924 , n71925 , n71926 , n71927 , n71928 , n71929 , n71930 , n71931 , n71932 , n71933 , n71934 , n71935 , n71936 , n71937 , n71938 , n71939 , n71940 , n71941 , n71942 , n71943 , n71944 , n71945 , n71946 , n71947 , n71948 , n71949 , n71950 , n71951 , n71952 , n71953 , n71954 , n71955 , n71956 , n71957 , n71958 , n71959 , n71960 , n71961 , n71962 , n71963 , n71964 , n71965 , n71966 , n71967 , n71968 , n71969 , n71970 , n71971 , n71972 , n71973 , n71974 , n71975 , n71976 , n71977 , n71978 , n71979 , n71980 , n71981 , n71982 , n71983 , n71984 , n71985 , n71986 , n71987 , n71988 , n71989 , n71990 , n71991 , n71992 , n71993 , n71994 , n71995 , n71996 , n71997 , n71998 , n71999 , n72000 , n72001 , n72002 , n72003 , n72004 , n72005 , n72006 , n72007 , n72008 , n72009 , n72010 , n72011 , n72012 , n72013 , n72014 , n72015 , n72016 , n72017 , n72018 , n72019 , n72020 , n72021 , n72022 , n72023 , n72024 , n72025 , n72026 , n72027 , n72028 , n72029 , n72030 , n72031 , n72032 , n72033 , n72034 , n72035 , n72036 , n72037 , n72038 , n72039 , n72040 , n72041 , n72042 , n72043 , n72044 , n72045 , n72046 , n72047 , n72048 , n72049 , n72050 , n72051 , n72052 , n72053 , n72054 , n72055 , n72056 , n72057 , n72058 , n72059 , n72060 , n72061 , n72062 , n72063 , n72064 , n72065 , n72066 , n72067 , n72068 , n72069 , n72070 , n72071 , n72072 , n72073 , n72074 , n72075 , n72076 , n72077 , n72078 , n72079 , n72080 , n72081 , n72082 , n72083 , n72084 , n72085 , n72086 , n72087 , n72088 , n72089 , n72090 , n72091 , n72092 , n72093 , n72094 , n72095 , n72096 , n72097 , n72098 , n72099 , n72100 , n72101 , n72102 , n72103 , n72104 , n72105 , n72106 , n72107 , n72108 , n72109 , n72110 , n72111 , n72112 , n72113 , n72114 , n72115 , n72116 , n72117 , n72118 , n72119 , n72120 , n72121 , n72122 , n72123 , n72124 , n72125 , n72126 , n72127 , n72128 , n72129 , n72130 , n72131 , n72132 , n72133 , n72134 , n72135 , n72136 , n72137 , n72138 , n72139 , n72140 , n72141 , n72142 , n72143 , n72144 , n72145 , n72146 , n72147 , n72148 , n72149 , n72150 , n72151 , n72152 , n72153 , n72154 , n72155 , n72156 , n72157 , n72158 , n72159 , n72160 , n72161 , n72162 , n72163 , n72164 , n72165 , n72166 , n72167 , n72168 , n72169 , n72170 , n72171 , n72172 , n72173 , n72174 , n72175 , n72176 , n72177 , n72178 , n72179 , n72180 , n72181 , n72182 , n72183 , n72184 , n72185 , n72186 , n72187 , n72188 , n72189 , n72190 , n72191 , n72192 , n72193 , n72194 , n72195 , n72196 , n72197 , n72198 , n72199 , n72200 , n72201 , n72202 , n72203 , n72204 , n72205 , n72206 , n72207 , n72208 , n72209 , n72210 , n72211 , n72212 , n72213 , n72214 , n72215 , n72216 , n72217 , n72218 , n72219 , n72220 , n72221 , n72222 , n72223 , n72224 , n72225 , n72226 , n72227 , n72228 , n72229 , n72230 , n72231 , n72232 , n72233 , n72234 , n72235 , n72236 , n72237 , n72238 , n72239 , n72240 , n72241 , n72242 , n72243 , n72244 , n72245 , n72246 , n72247 , n72248 , n72249 , n72250 , n72251 , n72252 , n72253 , n72254 , n72255 , n72256 , n72257 , n72258 , n72259 , n72260 , n72261 , n72262 , n72263 , n72264 , n72265 , n72266 , n72267 , n72268 , n72269 , n72270 , n72271 , n72272 , n72273 , n72274 , n72275 , n72276 , n72277 , n72278 , n72279 , n72280 , n72281 , n72282 , n72283 , n72284 , n72285 , n72286 , n72287 , n72288 , n72289 , n72290 , n72291 , n72292 , n72293 , n72294 , n72295 , n72296 , n72297 , n72298 , n72299 , n72300 , n72301 , n72302 , n72303 , n72304 , n72305 , n72306 , n72307 , n72308 , n72309 , n72310 , n72311 , n72312 , n72313 , n72314 , n72315 , n72316 , n72317 , n72318 , n72319 , n72320 , n72321 , n72322 , n72323 , n72324 , n72325 , n72326 , n72327 , n72328 , n72329 , n72330 , n72331 , n72332 , n72333 , n72334 , n72335 , n72336 , n72337 , n72338 , n72339 , n72340 , n72341 , n72342 , n72343 , n72344 , n72345 , n72346 , n72347 , n72348 , n72349 , n72350 , n72351 , n72352 , n72353 , n72354 , n72355 , n72356 , n72357 , n72358 , n72359 , n72360 , n72361 , n72362 , n72363 , n72364 , n72365 , n72366 , n72367 , n72368 , n72369 , n72370 , n72371 , n72372 , n72373 , n72374 , n72375 , n72376 , n72377 , n72378 , n72379 , n72380 , n72381 , n72382 , n72383 , n72384 , n72385 , n72386 , n72387 , n72388 , n72389 , n72390 , n72391 , n72392 , n72393 , n72394 , n72395 , n72396 , n72397 , n72398 , n72399 , n72400 , n72401 , n72402 , n72403 , n72404 , n72405 , n72406 , n72407 , n72408 , n72409 , n72410 , n72411 , n72412 , n72413 , n72414 , n72415 , n72416 , n72417 , n72418 , n72419 , n72420 , n72421 , n72422 , n72423 , n72424 , n72425 , n72426 , n72427 , n72428 , n72429 , n72430 , n72431 , n72432 , n72433 , n72434 , n72435 , n72436 , n72437 , n72438 , n72439 , n72440 , n72441 , n72442 , n72443 , n72444 , n72445 , n72446 , n72447 , n72448 , n72449 , n72450 , n72451 , n72452 , n72453 , n72454 , n72455 , n72456 , n72457 , n72458 , n72459 , n72460 , n72461 , n72462 , n72463 , n72464 , n72465 , n72466 , n72467 , n72468 , n72469 , n72470 , n72471 , n72472 , n72473 , n72474 , n72475 , n72476 , n72477 , n72478 , n72479 , n72480 , n72481 , n72482 , n72483 , n72484 , n72485 , n72486 , n72487 , n72488 , n72489 , n72490 , n72491 , n72492 , n72493 , n72494 , n72495 , n72496 , n72497 , n72498 , n72499 , n72500 , n72501 , n72502 , n72503 , n72504 , n72505 , n72506 , n72507 , n72508 , n72509 , n72510 , n72511 , n72512 , n72513 , n72514 , n72515 , n72516 , n72517 , n72518 , n72519 , n72520 , n72521 , n72522 , n72523 , n72524 , n72525 , n72526 , n72527 , n72528 , n72529 , n72530 , n72531 , n72532 , n72533 , n72534 , n72535 , n72536 , n72537 , n72538 , n72539 , n72540 , n72541 , n72542 , n72543 , n72544 , n72545 , n72546 , n72547 , n72548 , n72549 , n72550 , n72551 , n72552 , n72553 , n72554 , n72555 , n72556 , n72557 , n72558 , n72559 , n72560 , n72561 , n72562 , n72563 , n72564 , n72565 , n72566 , n72567 , n72568 , n72569 , n72570 , n72571 , n72572 , n72573 , n72574 , n72575 , n72576 , n72577 , n72578 , n72579 , n72580 , n72581 , n72582 , n72583 , n72584 , n72585 , n72586 , n72587 , n72588 , n72589 , n72590 , n72591 , n72592 , n72593 , n72594 , n72595 , n72596 , n72597 , n72598 , n72599 , n72600 , n72601 , n72602 , n72603 , n72604 , n72605 , n72606 , n72607 , n72608 , n72609 , n72610 , n72611 , n72612 , n72613 , n72614 , n72615 , n72616 , n72617 , n72618 , n72619 , n72620 , n72621 , n72622 , n72623 , n72624 , n72625 , n72626 , n72627 , n72628 , n72629 , n72630 , n72631 , n72632 , n72633 , n72634 , n72635 , n72636 , n72637 , n72638 , n72639 , n72640 , n72641 , n72642 , n72643 , n72644 , n72645 , n72646 , n72647 , n72648 , n72649 , n72650 , n72651 , n72652 , n72653 , n72654 , n72655 , n72656 , n72657 , n72658 , n72659 , n72660 , n72661 , n72662 , n72663 , n72664 , n72665 , n72666 , n72667 , n72668 , n72669 , n72670 , n72671 , n72672 , n72673 , n72674 , n72675 , n72676 , n72677 , n72678 , n72679 , n72680 , n72681 , n72682 , n72683 , n72684 , n72685 , n72686 , n72687 , n72688 , n72689 , n72690 , n72691 , n72692 , n72693 , n72694 , n72695 , n72696 , n72697 , n72698 , n72699 , n72700 , n72701 , n72702 , n72703 , n72704 , n72705 , n72706 , n72707 , n72708 , n72709 , n72710 , n72711 , n72712 , n72713 , n72714 , n72715 , n72716 , n72717 , n72718 , n72719 , n72720 , n72721 , n72722 , n72723 , n72724 , n72725 , n72726 , n72727 , n72728 , n72729 , n72730 , n72731 , n72732 , n72733 , n72734 , n72735 , n72736 , n72737 , n72738 , n72739 , n72740 , n72741 , n72742 , n72743 , n72744 , n72745 , n72746 , n72747 , n72748 , n72749 , n72750 , n72751 , n72752 , n72753 , n72754 , n72755 , n72756 , n72757 , n72758 , n72759 , n72760 , n72761 , n72762 , n72763 , n72764 , n72765 , n72766 , n72767 , n72768 , n72769 , n72770 , n72771 , n72772 , n72773 , n72774 , n72775 , n72776 , n72777 , n72778 , n72779 , n72780 , n72781 , n72782 , n72783 , n72784 , n72785 , n72786 , n72787 , n72788 , n72789 , n72790 , n72791 , n72792 , n72793 , n72794 , n72795 , n72796 , n72797 , n72798 , n72799 , n72800 , n72801 , n72802 , n72803 , n72804 , n72805 , n72806 , n72807 , n72808 , n72809 , n72810 , n72811 , n72812 , n72813 , n72814 , n72815 , n72816 , n72817 , n72818 , n72819 , n72820 , n72821 , n72822 , n72823 , n72824 , n72825 , n72826 , n72827 , n72828 , n72829 , n72830 , n72831 , n72832 , n72833 , n72834 , n72835 , n72836 , n72837 , n72838 , n72839 , n72840 , n72841 , n72842 , n72843 , n72844 , n72845 , n72846 , n72847 , n72848 , n72849 , n72850 , n72851 , n72852 , n72853 , n72854 , n72855 , n72856 , n72857 , n72858 , n72859 , n72860 , n72861 , n72862 , n72863 , n72864 , n72865 , n72866 , n72867 , n72868 , n72869 , n72870 , n72871 , n72872 , n72873 , n72874 , n72875 , n72876 , n72877 , n72878 , n72879 , n72880 , n72881 , n72882 , n72883 , n72884 , n72885 , n72886 , n72887 , n72888 , n72889 , n72890 , n72891 , n72892 , n72893 , n72894 , n72895 , n72896 , n72897 , n72898 , n72899 , n72900 , n72901 , n72902 , n72903 , n72904 , n72905 , n72906 , n72907 , n72908 , n72909 , n72910 , n72911 , n72912 , n72913 , n72914 , n72915 , n72916 , n72917 , n72918 , n72919 , n72920 , n72921 , n72922 , n72923 , n72924 , n72925 , n72926 , n72927 , n72928 , n72929 , n72930 , n72931 , n72932 , n72933 , n72934 , n72935 , n72936 , n72937 , n72938 , n72939 , n72940 , n72941 , n72942 , n72943 , n72944 , n72945 , n72946 , n72947 , n72948 , n72949 , n72950 , n72951 , n72952 , n72953 , n72954 , n72955 , n72956 , n72957 , n72958 , n72959 , n72960 , n72961 , n72962 , n72963 , n72964 , n72965 , n72966 , n72967 , n72968 , n72969 , n72970 , n72971 , n72972 , n72973 , n72974 , n72975 , n72976 , n72977 , n72978 , n72979 , n72980 , n72981 , n72982 , n72983 , n72984 , n72985 , n72986 , n72987 , n72988 , n72989 , n72990 , n72991 , n72992 , n72993 , n72994 , n72995 , n72996 , n72997 , n72998 , n72999 , n73000 , n73001 , n73002 , n73003 , n73004 , n73005 , n73006 , n73007 , n73008 , n73009 , n73010 , n73011 , n73012 , n73013 , n73014 , n73015 , n73016 , n73017 , n73018 , n73019 , n73020 , n73021 , n73022 , n73023 , n73024 , n73025 , n73026 , n73027 , n73028 , n73029 , n73030 , n73031 , n73032 , n73033 , n73034 , n73035 , n73036 , n73037 , n73038 , n73039 , n73040 , n73041 , n73042 , n73043 , n73044 , n73045 , n73046 , n73047 , n73048 , n73049 , n73050 , n73051 , n73052 , n73053 , n73054 , n73055 , n73056 , n73057 , n73058 , n73059 , n73060 , n73061 , n73062 , n73063 , n73064 , n73065 , n73066 , n73067 , n73068 , n73069 , n73070 , n73071 , n73072 , n73073 , n73074 , n73075 , n73076 , n73077 , n73078 , n73079 , n73080 , n73081 , n73082 , n73083 , n73084 , n73085 , n73086 , n73087 , n73088 , n73089 , n73090 , n73091 , n73092 , n73093 , n73094 , n73095 , n73096 , n73097 , n73098 , n73099 , n73100 , n73101 , n73102 , n73103 , n73104 , n73105 , n73106 , n73107 , n73108 , n73109 , n73110 , n73111 , n73112 , n73113 , n73114 , n73115 , n73116 , n73117 , n73118 , n73119 , n73120 , n73121 , n73122 , n73123 , n73124 , n73125 , n73126 , n73127 , n73128 , n73129 , n73130 , n73131 , n73132 , n73133 , n73134 , n73135 , n73136 , n73137 , n73138 , n73139 , n73140 , n73141 , n73142 , n73143 , n73144 , n73145 , n73146 , n73147 , n73148 , n73149 , n73150 , n73151 , n73152 , n73153 , n73154 , n73155 , n73156 , n73157 , n73158 , n73159 , n73160 , n73161 , n73162 , n73163 , n73164 , n73165 , n73166 , n73167 , n73168 , n73169 , n73170 , n73171 , n73172 , n73173 , n73174 , n73175 , n73176 , n73177 , n73178 , n73179 , n73180 , n73181 , n73182 , n73183 , n73184 , n73185 , n73186 , n73187 , n73188 , n73189 , n73190 , n73191 , n73192 , n73193 , n73194 , n73195 , n73196 , n73197 , n73198 , n73199 , n73200 , n73201 , n73202 , n73203 , n73204 , n73205 , n73206 , n73207 , n73208 , n73209 , n73210 , n73211 , n73212 , n73213 , n73214 , n73215 , n73216 , n73217 , n73218 , n73219 , n73220 , n73221 , n73222 , n73223 , n73224 , n73225 , n73226 , n73227 , n73228 , n73229 , n73230 , n73231 , n73232 , n73233 , n73234 , n73235 , n73236 , n73237 , n73238 , n73239 , n73240 , n73241 , n73242 , n73243 , n73244 , n73245 , n73246 , n73247 , n73248 , n73249 , n73250 , n73251 , n73252 , n73253 , n73254 , n73255 , n73256 , n73257 , n73258 , n73259 , n73260 , n73261 , n73262 , n73263 , n73264 , n73265 , n73266 , n73267 , n73268 , n73269 , n73270 , n73271 , n73272 , n73273 , n73274 , n73275 , n73276 , n73277 , n73278 , n73279 , n73280 , n73281 , n73282 , n73283 , n73284 , n73285 , n73286 , n73287 , n73288 , n73289 , n73290 , n73291 , n73292 , n73293 , n73294 , n73295 , n73296 , n73297 , n73298 , n73299 , n73300 , n73301 , n73302 , n73303 , n73304 , n73305 , n73306 , n73307 , n73308 , n73309 , n73310 , n73311 , n73312 , n73313 , n73314 , n73315 , n73316 , n73317 , n73318 , n73319 , n73320 , n73321 , n73322 , n73323 , n73324 , n73325 , n73326 , n73327 , n73328 , n73329 , n73330 , n73331 , n73332 , n73333 , n73334 , n73335 , n73336 , n73337 , n73338 , n73339 , n73340 , n73341 , n73342 , n73343 , n73344 , n73345 , n73346 , n73347 , n73348 , n73349 , n73350 , n73351 , n73352 , n73353 , n73354 , n73355 , n73356 , n73357 , n73358 , n73359 , n73360 , n73361 , n73362 , n73363 , n73364 , n73365 , n73366 , n73367 , n73368 , n73369 , n73370 , n73371 , n73372 , n73373 , n73374 , n73375 , n73376 , n73377 , n73378 , n73379 , n73380 , n73381 , n73382 , n73383 , n73384 , n73385 , n73386 , n73387 , n73388 , n73389 , n73390 , n73391 , n73392 , n73393 , n73394 , n73395 , n73396 , n73397 , n73398 , n73399 , n73400 , n73401 , n73402 , n73403 , n73404 , n73405 , n73406 , n73407 , n73408 , n73409 , n73410 , n73411 , n73412 , n73413 , n73414 , n73415 , n73416 , n73417 , n73418 , n73419 , n73420 , n73421 , n73422 , n73423 , n73424 , n73425 , n73426 , n73427 , n73428 , n73429 , n73430 , n73431 , n73432 , n73433 , n73434 , n73435 , n73436 , n73437 , n73438 , n73439 , n73440 , n73441 , n73442 , n73443 , n73444 , n73445 , n73446 , n73447 , n73448 , n73449 , n73450 , n73451 , n73452 , n73453 , n73454 , n73455 , n73456 , n73457 , n73458 , n73459 , n73460 , n73461 , n73462 , n73463 , n73464 , n73465 , n73466 , n73467 , n73468 , n73469 , n73470 , n73471 , n73472 , n73473 , n73474 , n73475 , n73476 , n73477 , n73478 , n73479 , n73480 , n73481 , n73482 , n73483 , n73484 , n73485 , n73486 , n73487 , n73488 , n73489 , n73490 , n73491 , n73492 , n73493 , n73494 , n73495 , n73496 , n73497 , n73498 , n73499 , n73500 , n73501 , n73502 , n73503 , n73504 , n73505 , n73506 , n73507 , n73508 , n73509 , n73510 , n73511 , n73512 , n73513 , n73514 , n73515 , n73516 , n73517 , n73518 , n73519 , n73520 , n73521 , n73522 , n73523 , n73524 , n73525 , n73526 , n73527 , n73528 , n73529 , n73530 , n73531 , n73532 , n73533 , n73534 , n73535 , n73536 , n73537 , n73538 , n73539 , n73540 , n73541 , n73542 , n73543 , n73544 , n73545 , n73546 , n73547 , n73548 , n73549 , n73550 , n73551 , n73552 , n73553 , n73554 , n73555 , n73556 , n73557 , n73558 , n73559 , n73560 , n73561 , n73562 , n73563 , n73564 , n73565 , n73566 , n73567 , n73568 , n73569 , n73570 , n73571 , n73572 , n73573 , n73574 , n73575 , n73576 , n73577 , n73578 , n73579 , n73580 , n73581 , n73582 , n73583 , n73584 , n73585 , n73586 , n73587 , n73588 , n73589 , n73590 , n73591 , n73592 , n73593 , n73594 , n73595 , n73596 , n73597 , n73598 , n73599 , n73600 , n73601 , n73602 , n73603 , n73604 , n73605 , n73606 , n73607 , n73608 , n73609 , n73610 , n73611 , n73612 , n73613 , n73614 , n73615 , n73616 , n73617 , n73618 , n73619 , n73620 , n73621 , n73622 , n73623 , n73624 , n73625 , n73626 , n73627 , n73628 , n73629 , n73630 , n73631 , n73632 , n73633 , n73634 , n73635 , n73636 , n73637 , n73638 , n73639 , n73640 , n73641 , n73642 , n73643 , n73644 , n73645 , n73646 , n73647 , n73648 , n73649 , n73650 , n73651 , n73652 , n73653 , n73654 , n73655 , n73656 , n73657 , n73658 , n73659 , n73660 , n73661 , n73662 , n73663 , n73664 , n73665 , n73666 , n73667 , n73668 , n73669 , n73670 , n73671 , n73672 , n73673 , n73674 , n73675 , n73676 , n73677 , n73678 , n73679 , n73680 , n73681 , n73682 , n73683 , n73684 , n73685 , n73686 , n73687 , n73688 , n73689 , n73690 , n73691 , n73692 , n73693 , n73694 , n73695 , n73696 , n73697 , n73698 , n73699 , n73700 , n73701 , n73702 , n73703 , n73704 , n73705 , n73706 , n73707 , n73708 , n73709 , n73710 , n73711 , n73712 , n73713 , n73714 , n73715 , n73716 , n73717 , n73718 , n73719 , n73720 , n73721 , n73722 , n73723 , n73724 , n73725 , n73726 , n73727 , n73728 , n73729 , n73730 , n73731 , n73732 , n73733 , n73734 , n73735 , n73736 , n73737 , n73738 , n73739 , n73740 , n73741 , n73742 , n73743 , n73744 , n73745 , n73746 , n73747 , n73748 , n73749 , n73750 , n73751 , n73752 , n73753 , n73754 , n73755 , n73756 , n73757 , n73758 , n73759 , n73760 , n73761 , n73762 , n73763 , n73764 , n73765 , n73766 , n73767 , n73768 , n73769 , n73770 , n73771 , n73772 , n73773 , n73774 , n73775 , n73776 , n73777 , n73778 , n73779 , n73780 , n73781 , n73782 , n73783 , n73784 , n73785 , n73786 , n73787 , n73788 , n73789 , n73790 , n73791 , n73792 , n73793 , n73794 , n73795 , n73796 , n73797 , n73798 , n73799 , n73800 , n73801 , n73802 , n73803 , n73804 , n73805 , n73806 , n73807 , n73808 , n73809 , n73810 , n73811 , n73812 , n73813 , n73814 , n73815 , n73816 , n73817 , n73818 , n73819 , n73820 , n73821 , n73822 , n73823 , n73824 , n73825 , n73826 , n73827 , n73828 , n73829 , n73830 , n73831 , n73832 , n73833 , n73834 , n73835 , n73836 , n73837 , n73838 , n73839 , n73840 , n73841 , n73842 , n73843 , n73844 , n73845 , n73846 , n73847 , n73848 , n73849 , n73850 , n73851 , n73852 , n73853 , n73854 , n73855 , n73856 , n73857 , n73858 , n73859 , n73860 , n73861 , n73862 , n73863 , n73864 , n73865 , n73866 , n73867 , n73868 , n73869 , n73870 , n73871 , n73872 , n73873 , n73874 , n73875 , n73876 , n73877 , n73878 , n73879 , n73880 , n73881 , n73882 , n73883 , n73884 , n73885 , n73886 , n73887 , n73888 , n73889 , n73890 , n73891 , n73892 , n73893 , n73894 , n73895 , n73896 , n73897 , n73898 , n73899 , n73900 , n73901 , n73902 , n73903 , n73904 , n73905 , n73906 , n73907 , n73908 , n73909 , n73910 , n73911 , n73912 , n73913 , n73914 , n73915 , n73916 , n73917 , n73918 , n73919 , n73920 , n73921 , n73922 , n73923 , n73924 , n73925 , n73926 , n73927 , n73928 , n73929 , n73930 , n73931 , n73932 , n73933 , n73934 , n73935 , n73936 , n73937 , n73938 , n73939 , n73940 , n73941 , n73942 , n73943 , n73944 , n73945 , n73946 , n73947 , n73948 , n73949 , n73950 , n73951 , n73952 , n73953 , n73954 , n73955 , n73956 , n73957 , n73958 , n73959 , n73960 , n73961 , n73962 , n73963 , n73964 , n73965 , n73966 , n73967 , n73968 , n73969 , n73970 , n73971 , n73972 , n73973 , n73974 , n73975 , n73976 , n73977 , n73978 , n73979 , n73980 , n73981 , n73982 , n73983 , n73984 , n73985 , n73986 , n73987 , n73988 , n73989 , n73990 , n73991 , n73992 , n73993 , n73994 , n73995 , n73996 , n73997 , n73998 , n73999 , n74000 , n74001 , n74002 , n74003 , n74004 , n74005 , n74006 , n74007 , n74008 , n74009 , n74010 , n74011 , n74012 , n74013 , n74014 , n74015 , n74016 , n74017 , n74018 , n74019 , n74020 , n74021 , n74022 , n74023 , n74024 , n74025 , n74026 , n74027 , n74028 , n74029 , n74030 , n74031 , n74032 , n74033 , n74034 , n74035 , n74036 , n74037 , n74038 , n74039 , n74040 , n74041 , n74042 , n74043 , n74044 , n74045 , n74046 , n74047 , n74048 , n74049 , n74050 , n74051 , n74052 , n74053 , n74054 , n74055 , n74056 , n74057 , n74058 , n74059 , n74060 , n74061 , n74062 , n74063 , n74064 , n74065 , n74066 , n74067 , n74068 , n74069 , n74070 , n74071 , n74072 , n74073 , n74074 , n74075 , n74076 , n74077 , n74078 , n74079 , n74080 , n74081 , n74082 , n74083 , n74084 , n74085 , n74086 , n74087 , n74088 , n74089 , n74090 , n74091 , n74092 , n74093 , n74094 , n74095 , n74096 , n74097 , n74098 , n74099 , n74100 , n74101 , n74102 , n74103 , n74104 , n74105 , n74106 , n74107 , n74108 , n74109 , n74110 , n74111 , n74112 , n74113 , n74114 , n74115 , n74116 , n74117 , n74118 , n74119 , n74120 , n74121 , n74122 , n74123 , n74124 , n74125 , n74126 , n74127 , n74128 , n74129 , n74130 , n74131 , n74132 , n74133 , n74134 , n74135 , n74136 , n74137 , n74138 , n74139 , n74140 , n74141 , n74142 , n74143 , n74144 , n74145 , n74146 , n74147 , n74148 , n74149 , n74150 , n74151 , n74152 , n74153 , n74154 , n74155 , n74156 , n74157 , n74158 , n74159 , n74160 , n74161 , n74162 , n74163 , n74164 , n74165 , n74166 , n74167 , n74168 , n74169 , n74170 , n74171 , n74172 , n74173 , n74174 , n74175 , n74176 , n74177 , n74178 , n74179 , n74180 , n74181 , n74182 , n74183 , n74184 , n74185 , n74186 , n74187 , n74188 , n74189 , n74190 , n74191 , n74192 , n74193 , n74194 , n74195 , n74196 , n74197 , n74198 , n74199 , n74200 , n74201 , n74202 , n74203 , n74204 , n74205 , n74206 , n74207 , n74208 , n74209 , n74210 , n74211 , n74212 , n74213 , n74214 , n74215 , n74216 , n74217 , n74218 , n74219 , n74220 , n74221 , n74222 , n74223 , n74224 , n74225 , n74226 , n74227 , n74228 , n74229 , n74230 , n74231 , n74232 , n74233 , n74234 , n74235 , n74236 , n74237 , n74238 , n74239 , n74240 , n74241 , n74242 , n74243 , n74244 , n74245 , n74246 , n74247 , n74248 , n74249 , n74250 , n74251 , n74252 , n74253 , n74254 , n74255 , n74256 , n74257 , n74258 , n74259 , n74260 , n74261 , n74262 , n74263 , n74264 , n74265 , n74266 , n74267 , n74268 , n74269 , n74270 , n74271 , n74272 , n74273 , n74274 , n74275 , n74276 , n74277 , n74278 , n74279 , n74280 , n74281 , n74282 , n74283 , n74284 , n74285 , n74286 , n74287 , n74288 , n74289 , n74290 , n74291 , n74292 , n74293 , n74294 , n74295 , n74296 , n74297 , n74298 , n74299 , n74300 , n74301 , n74302 , n74303 , n74304 , n74305 , n74306 , n74307 , n74308 , n74309 , n74310 , n74311 , n74312 , n74313 , n74314 , n74315 , n74316 , n74317 , n74318 , n74319 , n74320 , n74321 , n74322 , n74323 , n74324 , n74325 , n74326 , n74327 , n74328 , n74329 , n74330 , n74331 , n74332 , n74333 , n74334 , n74335 , n74336 , n74337 , n74338 , n74339 , n74340 , n74341 , n74342 , n74343 , n74344 , n74345 , n74346 , n74347 , n74348 , n74349 , n74350 , n74351 , n74352 , n74353 , n74354 , n74355 , n74356 , n74357 , n74358 , n74359 , n74360 , n74361 , n74362 , n74363 , n74364 , n74365 , n74366 , n74367 , n74368 , n74369 , n74370 , n74371 , n74372 , n74373 , n74374 , n74375 , n74376 , n74377 , n74378 , n74379 , n74380 , n74381 , n74382 , n74383 , n74384 , n74385 , n74386 , n74387 , n74388 , n74389 , n74390 , n74391 , n74392 , n74393 , n74394 , n74395 , n74396 , n74397 , n74398 , n74399 , n74400 , n74401 , n74402 , n74403 , n74404 , n74405 , n74406 , n74407 , n74408 , n74409 , n74410 , n74411 , n74412 , n74413 , n74414 , n74415 , n74416 , n74417 , n74418 , n74419 , n74420 , n74421 , n74422 , n74423 , n74424 , n74425 , n74426 , n74427 , n74428 , n74429 , n74430 , n74431 , n74432 , n74433 , n74434 , n74435 , n74436 , n74437 , n74438 , n74439 , n74440 , n74441 , n74442 , n74443 , n74444 , n74445 , n74446 , n74447 , n74448 , n74449 , n74450 , n74451 , n74452 , n74453 , n74454 , n74455 , n74456 , n74457 , n74458 , n74459 , n74460 , n74461 , n74462 , n74463 , n74464 , n74465 , n74466 , n74467 , n74468 , n74469 , n74470 , n74471 , n74472 , n74473 , n74474 , n74475 , n74476 , n74477 , n74478 , n74479 , n74480 , n74481 , n74482 , n74483 , n74484 , n74485 , n74486 , n74487 , n74488 , n74489 , n74490 , n74491 , n74492 , n74493 , n74494 , n74495 , n74496 , n74497 , n74498 , n74499 , n74500 , n74501 , n74502 , n74503 , n74504 , n74505 , n74506 , n74507 , n74508 , n74509 , n74510 , n74511 , n74512 , n74513 , n74514 , n74515 , n74516 , n74517 , n74518 , n74519 , n74520 , n74521 , n74522 , n74523 , n74524 , n74525 , n74526 , n74527 , n74528 , n74529 , n74530 , n74531 , n74532 , n74533 , n74534 , n74535 , n74536 , n74537 , n74538 , n74539 , n74540 , n74541 , n74542 , n74543 , n74544 , n74545 , n74546 , n74547 , n74548 , n74549 , n74550 , n74551 , n74552 , n74553 , n74554 , n74555 , n74556 , n74557 , n74558 , n74559 , n74560 , n74561 , n74562 , n74563 , n74564 , n74565 , n74566 , n74567 , n74568 , n74569 , n74570 , n74571 , n74572 , n74573 , n74574 , n74575 , n74576 , n74577 , n74578 , n74579 , n74580 , n74581 , n74582 , n74583 , n74584 , n74585 , n74586 , n74587 , n74588 , n74589 , n74590 , n74591 , n74592 , n74593 , n74594 , n74595 , n74596 , n74597 , n74598 , n74599 , n74600 , n74601 , n74602 , n74603 , n74604 , n74605 , n74606 , n74607 , n74608 , n74609 , n74610 , n74611 , n74612 , n74613 , n74614 , n74615 , n74616 , n74617 , n74618 , n74619 , n74620 , n74621 , n74622 , n74623 , n74624 , n74625 , n74626 , n74627 , n74628 , n74629 , n74630 , n74631 , n74632 , n74633 , n74634 , n74635 , n74636 , n74637 , n74638 , n74639 , n74640 , n74641 , n74642 , n74643 , n74644 , n74645 , n74646 , n74647 , n74648 , n74649 , n74650 , n74651 , n74652 , n74653 , n74654 , n74655 , n74656 , n74657 , n74658 , n74659 , n74660 , n74661 , n74662 , n74663 , n74664 , n74665 , n74666 , n74667 , n74668 , n74669 , n74670 , n74671 , n74672 , n74673 , n74674 , n74675 , n74676 , n74677 , n74678 , n74679 , n74680 , n74681 , n74682 , n74683 , n74684 , n74685 , n74686 , n74687 , n74688 , n74689 , n74690 , n74691 , n74692 , n74693 , n74694 , n74695 , n74696 , n74697 , n74698 , n74699 , n74700 , n74701 , n74702 , n74703 , n74704 , n74705 , n74706 , n74707 , n74708 , n74709 , n74710 , n74711 , n74712 , n74713 , n74714 , n74715 , n74716 , n74717 , n74718 , n74719 , n74720 , n74721 , n74722 , n74723 , n74724 , n74725 , n74726 , n74727 , n74728 , n74729 , n74730 , n74731 , n74732 , n74733 , n74734 , n74735 , n74736 , n74737 , n74738 , n74739 , n74740 , n74741 , n74742 , n74743 , n74744 , n74745 , n74746 , n74747 , n74748 , n74749 , n74750 , n74751 , n74752 , n74753 , n74754 , n74755 , n74756 , n74757 , n74758 , n74759 , n74760 , n74761 , n74762 , n74763 , n74764 , n74765 , n74766 , n74767 , n74768 , n74769 , n74770 , n74771 , n74772 , n74773 , n74774 , n74775 , n74776 , n74777 , n74778 , n74779 , n74780 , n74781 , n74782 , n74783 , n74784 , n74785 , n74786 , n74787 , n74788 , n74789 , n74790 , n74791 , n74792 , n74793 , n74794 , n74795 , n74796 , n74797 , n74798 , n74799 , n74800 , n74801 , n74802 , n74803 , n74804 , n74805 , n74806 , n74807 , n74808 , n74809 , n74810 , n74811 , n74812 , n74813 , n74814 , n74815 , n74816 , n74817 , n74818 , n74819 , n74820 , n74821 , n74822 , n74823 , n74824 , n74825 , n74826 , n74827 , n74828 , n74829 , n74830 , n74831 , n74832 , n74833 , n74834 , n74835 , n74836 , n74837 , n74838 , n74839 , n74840 , n74841 , n74842 , n74843 , n74844 , n74845 , n74846 , n74847 , n74848 , n74849 , n74850 , n74851 , n74852 , n74853 , n74854 , n74855 , n74856 , n74857 , n74858 , n74859 , n74860 , n74861 , n74862 , n74863 , n74864 , n74865 , n74866 , n74867 , n74868 , n74869 , n74870 , n74871 , n74872 , n74873 , n74874 , n74875 , n74876 , n74877 , n74878 , n74879 , n74880 , n74881 , n74882 , n74883 , n74884 , n74885 , n74886 , n74887 , n74888 , n74889 , n74890 , n74891 , n74892 , n74893 , n74894 , n74895 , n74896 , n74897 , n74898 , n74899 , n74900 , n74901 , n74902 , n74903 , n74904 , n74905 , n74906 , n74907 , n74908 , n74909 , n74910 , n74911 , n74912 , n74913 , n74914 , n74915 , n74916 , n74917 , n74918 , n74919 , n74920 , n74921 , n74922 , n74923 , n74924 , n74925 , n74926 , n74927 , n74928 , n74929 , n74930 , n74931 , n74932 , n74933 , n74934 , n74935 , n74936 , n74937 , n74938 , n74939 , n74940 , n74941 , n74942 , n74943 , n74944 , n74945 , n74946 , n74947 , n74948 , n74949 , n74950 , n74951 , n74952 , n74953 , n74954 , n74955 , n74956 , n74957 , n74958 , n74959 , n74960 , n74961 , n74962 , n74963 , n74964 , n74965 , n74966 , n74967 , n74968 , n74969 , n74970 , n74971 , n74972 , n74973 , n74974 , n74975 , n74976 , n74977 , n74978 , n74979 , n74980 , n74981 , n74982 , n74983 , n74984 , n74985 , n74986 , n74987 , n74988 , n74989 , n74990 , n74991 , n74992 , n74993 , n74994 , n74995 , n74996 , n74997 , n74998 , n74999 , n75000 , n75001 , n75002 , n75003 , n75004 , n75005 , n75006 , n75007 , n75008 , n75009 , n75010 , n75011 , n75012 , n75013 , n75014 , n75015 , n75016 , n75017 , n75018 , n75019 , n75020 , n75021 , n75022 , n75023 , n75024 , n75025 , n75026 , n75027 , n75028 , n75029 , n75030 , n75031 , n75032 , n75033 , n75034 , n75035 , n75036 , n75037 , n75038 , n75039 , n75040 , n75041 , n75042 , n75043 , n75044 , n75045 , n75046 , n75047 , n75048 , n75049 , n75050 , n75051 , n75052 , n75053 , n75054 , n75055 , n75056 , n75057 , n75058 , n75059 , n75060 , n75061 , n75062 , n75063 , n75064 , n75065 , n75066 , n75067 , n75068 , n75069 , n75070 , n75071 , n75072 , n75073 , n75074 , n75075 , n75076 , n75077 , n75078 , n75079 , n75080 , n75081 , n75082 , n75083 , n75084 , n75085 , n75086 , n75087 , n75088 , n75089 , n75090 , n75091 , n75092 , n75093 , n75094 , n75095 , n75096 , n75097 , n75098 , n75099 , n75100 , n75101 , n75102 , n75103 , n75104 , n75105 , n75106 , n75107 , n75108 , n75109 , n75110 , n75111 , n75112 , n75113 , n75114 , n75115 , n75116 , n75117 , n75118 , n75119 , n75120 , n75121 , n75122 , n75123 , n75124 , n75125 , n75126 , n75127 , n75128 , n75129 , n75130 , n75131 , n75132 , n75133 , n75134 , n75135 , n75136 , n75137 , n75138 , n75139 , n75140 , n75141 , n75142 , n75143 , n75144 , n75145 , n75146 , n75147 , n75148 , n75149 , n75150 , n75151 , n75152 , n75153 , n75154 , n75155 , n75156 , n75157 , n75158 , n75159 , n75160 , n75161 , n75162 , n75163 , n75164 , n75165 , n75166 , n75167 , n75168 , n75169 , n75170 , n75171 , n75172 , n75173 , n75174 , n75175 , n75176 , n75177 , n75178 , n75179 , n75180 , n75181 , n75182 , n75183 , n75184 , n75185 , n75186 , n75187 , n75188 , n75189 , n75190 , n75191 , n75192 , n75193 , n75194 , n75195 , n75196 , n75197 , n75198 , n75199 , n75200 , n75201 , n75202 , n75203 , n75204 , n75205 , n75206 , n75207 , n75208 , n75209 , n75210 , n75211 , n75212 , n75213 , n75214 , n75215 , n75216 , n75217 , n75218 , n75219 , n75220 , n75221 , n75222 , n75223 , n75224 , n75225 , n75226 , n75227 , n75228 , n75229 , n75230 , n75231 , n75232 , n75233 , n75234 , n75235 , n75236 , n75237 , n75238 , n75239 , n75240 , n75241 , n75242 , n75243 , n75244 , n75245 , n75246 , n75247 , n75248 , n75249 , n75250 , n75251 , n75252 , n75253 , n75254 , n75255 , n75256 , n75257 , n75258 , n75259 , n75260 , n75261 , n75262 , n75263 , n75264 , n75265 , n75266 , n75267 , n75268 , n75269 , n75270 , n75271 , n75272 , n75273 , n75274 , n75275 , n75276 , n75277 , n75278 , n75279 , n75280 , n75281 , n75282 , n75283 , n75284 , n75285 , n75286 , n75287 , n75288 , n75289 , n75290 , n75291 , n75292 , n75293 , n75294 , n75295 , n75296 , n75297 , n75298 , n75299 , n75300 , n75301 , n75302 , n75303 , n75304 , n75305 , n75306 , n75307 , n75308 , n75309 , n75310 , n75311 , n75312 , n75313 , n75314 , n75315 , n75316 , n75317 , n75318 , n75319 , n75320 , n75321 , n75322 , n75323 , n75324 , n75325 , n75326 , n75327 , n75328 , n75329 , n75330 , n75331 , n75332 , n75333 , n75334 , n75335 , n75336 , n75337 , n75338 , n75339 , n75340 , n75341 , n75342 , n75343 , n75344 , n75345 , n75346 , n75347 , n75348 , n75349 , n75350 , n75351 , n75352 , n75353 , n75354 , n75355 , n75356 , n75357 , n75358 , n75359 , n75360 , n75361 , n75362 , n75363 , n75364 , n75365 , n75366 , n75367 , n75368 , n75369 , n75370 , n75371 , n75372 , n75373 , n75374 , n75375 , n75376 , n75377 , n75378 , n75379 , n75380 , n75381 , n75382 , n75383 , n75384 , n75385 , n75386 , n75387 , n75388 , n75389 , n75390 , n75391 , n75392 , n75393 , n75394 , n75395 , n75396 , n75397 , n75398 , n75399 , n75400 , n75401 , n75402 , n75403 , n75404 , n75405 , n75406 , n75407 , n75408 , n75409 , n75410 , n75411 , n75412 , n75413 , n75414 , n75415 , n75416 , n75417 , n75418 , n75419 , n75420 , n75421 , n75422 , n75423 , n75424 , n75425 , n75426 , n75427 , n75428 , n75429 , n75430 , n75431 , n75432 , n75433 , n75434 , n75435 , n75436 , n75437 , n75438 , n75439 , n75440 , n75441 , n75442 , n75443 , n75444 , n75445 , n75446 , n75447 , n75448 , n75449 , n75450 , n75451 , n75452 , n75453 , n75454 , n75455 , n75456 , n75457 , n75458 , n75459 , n75460 , n75461 , n75462 , n75463 , n75464 , n75465 , n75466 , n75467 , n75468 , n75469 , n75470 , n75471 , n75472 , n75473 , n75474 , n75475 , n75476 , n75477 , n75478 , n75479 , n75480 , n75481 , n75482 , n75483 , n75484 , n75485 , n75486 , n75487 , n75488 , n75489 , n75490 , n75491 , n75492 , n75493 , n75494 , n75495 , n75496 , n75497 , n75498 , n75499 , n75500 , n75501 , n75502 , n75503 , n75504 , n75505 , n75506 , n75507 , n75508 , n75509 , n75510 , n75511 , n75512 , n75513 , n75514 , n75515 , n75516 , n75517 , n75518 , n75519 , n75520 , n75521 , n75522 , n75523 , n75524 , n75525 , n75526 , n75527 , n75528 , n75529 , n75530 , n75531 , n75532 , n75533 , n75534 , n75535 , n75536 , n75537 , n75538 , n75539 , n75540 , n75541 , n75542 , n75543 , n75544 , n75545 , n75546 , n75547 , n75548 , n75549 , n75550 , n75551 , n75552 , n75553 , n75554 , n75555 , n75556 , n75557 , n75558 , n75559 , n75560 , n75561 , n75562 , n75563 , n75564 , n75565 , n75566 , n75567 , n75568 , n75569 , n75570 , n75571 , n75572 , n75573 , n75574 , n75575 , n75576 , n75577 , n75578 , n75579 , n75580 , n75581 , n75582 , n75583 , n75584 , n75585 , n75586 , n75587 , n75588 , n75589 , n75590 , n75591 , n75592 , n75593 , n75594 , n75595 , n75596 , n75597 , n75598 , n75599 , n75600 , n75601 , n75602 , n75603 , n75604 , n75605 , n75606 , n75607 , n75608 , n75609 , n75610 , n75611 , n75612 , n75613 , n75614 , n75615 , n75616 , n75617 , n75618 , n75619 , n75620 , n75621 , n75622 , n75623 , n75624 , n75625 , n75626 , n75627 , n75628 , n75629 , n75630 , n75631 , n75632 , n75633 , n75634 , n75635 , n75636 , n75637 , n75638 , n75639 , n75640 , n75641 , n75642 , n75643 , n75644 , n75645 , n75646 , n75647 , n75648 , n75649 , n75650 , n75651 , n75652 , n75653 , n75654 , n75655 , n75656 , n75657 , n75658 , n75659 , n75660 , n75661 , n75662 , n75663 , n75664 , n75665 , n75666 , n75667 , n75668 , n75669 , n75670 , n75671 , n75672 , n75673 , n75674 , n75675 , n75676 , n75677 , n75678 , n75679 , n75680 , n75681 , n75682 , n75683 , n75684 , n75685 , n75686 , n75687 , n75688 , n75689 , n75690 , n75691 , n75692 , n75693 , n75694 , n75695 , n75696 , n75697 , n75698 , n75699 , n75700 , n75701 , n75702 , n75703 , n75704 , n75705 , n75706 , n75707 , n75708 , n75709 , n75710 , n75711 , n75712 , n75713 , n75714 , n75715 , n75716 , n75717 , n75718 , n75719 , n75720 , n75721 , n75722 , n75723 , n75724 , n75725 , n75726 , n75727 , n75728 , n75729 , n75730 , n75731 , n75732 , n75733 , n75734 , n75735 , n75736 , n75737 , n75738 , n75739 , n75740 , n75741 , n75742 , n75743 , n75744 , n75745 , n75746 , n75747 , n75748 , n75749 , n75750 , n75751 , n75752 , n75753 , n75754 , n75755 , n75756 , n75757 , n75758 , n75759 , n75760 , n75761 , n75762 , n75763 , n75764 , n75765 , n75766 , n75767 , n75768 , n75769 , n75770 , n75771 , n75772 , n75773 , n75774 , n75775 , n75776 , n75777 , n75778 , n75779 , n75780 , n75781 , n75782 , n75783 , n75784 , n75785 , n75786 , n75787 , n75788 , n75789 , n75790 , n75791 , n75792 , n75793 , n75794 , n75795 , n75796 , n75797 , n75798 , n75799 , n75800 , n75801 , n75802 , n75803 , n75804 , n75805 , n75806 , n75807 , n75808 , n75809 , n75810 , n75811 , n75812 , n75813 , n75814 , n75815 , n75816 , n75817 , n75818 , n75819 , n75820 , n75821 , n75822 , n75823 , n75824 , n75825 , n75826 , n75827 , n75828 , n75829 , n75830 , n75831 , n75832 , n75833 , n75834 , n75835 , n75836 , n75837 , n75838 , n75839 , n75840 , n75841 , n75842 , n75843 , n75844 , n75845 , n75846 , n75847 , n75848 , n75849 , n75850 , n75851 , n75852 , n75853 , n75854 , n75855 , n75856 , n75857 , n75858 , n75859 , n75860 , n75861 , n75862 , n75863 , n75864 , n75865 , n75866 , n75867 , n75868 , n75869 , n75870 , n75871 , n75872 , n75873 , n75874 , n75875 , n75876 , n75877 , n75878 , n75879 , n75880 , n75881 , n75882 , n75883 , n75884 , n75885 , n75886 , n75887 , n75888 , n75889 , n75890 , n75891 , n75892 , n75893 , n75894 , n75895 , n75896 , n75897 , n75898 , n75899 , n75900 , n75901 , n75902 , n75903 , n75904 , n75905 , n75906 , n75907 , n75908 , n75909 , n75910 , n75911 , n75912 , n75913 , n75914 , n75915 , n75916 , n75917 , n75918 , n75919 , n75920 , n75921 , n75922 , n75923 , n75924 , n75925 , n75926 , n75927 , n75928 , n75929 , n75930 , n75931 , n75932 , n75933 , n75934 , n75935 , n75936 , n75937 , n75938 , n75939 , n75940 , n75941 , n75942 , n75943 , n75944 , n75945 , n75946 , n75947 , n75948 , n75949 , n75950 , n75951 , n75952 , n75953 , n75954 , n75955 , n75956 , n75957 , n75958 , n75959 , n75960 , n75961 , n75962 , n75963 , n75964 , n75965 , n75966 , n75967 , n75968 , n75969 , n75970 , n75971 , n75972 , n75973 , n75974 , n75975 , n75976 , n75977 , n75978 , n75979 , n75980 , n75981 , n75982 , n75983 , n75984 , n75985 , n75986 , n75987 , n75988 , n75989 , n75990 , n75991 , n75992 , n75993 , n75994 , n75995 , n75996 , n75997 , n75998 , n75999 , n76000 , n76001 , n76002 , n76003 , n76004 , n76005 , n76006 , n76007 , n76008 , n76009 , n76010 , n76011 , n76012 , n76013 , n76014 , n76015 , n76016 , n76017 , n76018 , n76019 , n76020 , n76021 , n76022 , n76023 , n76024 , n76025 , n76026 , n76027 , n76028 , n76029 , n76030 , n76031 , n76032 , n76033 , n76034 , n76035 , n76036 , n76037 , n76038 , n76039 , n76040 , n76041 , n76042 , n76043 , n76044 , n76045 , n76046 , n76047 , n76048 , n76049 , n76050 , n76051 , n76052 , n76053 , n76054 , n76055 , n76056 , n76057 , n76058 , n76059 , n76060 , n76061 , n76062 , n76063 , n76064 , n76065 , n76066 , n76067 , n76068 , n76069 , n76070 , n76071 , n76072 , n76073 , n76074 , n76075 , n76076 , n76077 , n76078 , n76079 , n76080 , n76081 , n76082 , n76083 , n76084 , n76085 , n76086 , n76087 , n76088 , n76089 , n76090 , n76091 , n76092 , n76093 , n76094 , n76095 , n76096 , n76097 , n76098 , n76099 , n76100 , n76101 , n76102 , n76103 , n76104 , n76105 , n76106 , n76107 , n76108 , n76109 , n76110 , n76111 , n76112 , n76113 , n76114 , n76115 , n76116 , n76117 , n76118 , n76119 , n76120 , n76121 , n76122 , n76123 , n76124 , n76125 , n76126 , n76127 , n76128 , n76129 , n76130 , n76131 , n76132 , n76133 , n76134 , n76135 , n76136 , n76137 , n76138 , n76139 , n76140 , n76141 , n76142 , n76143 , n76144 , n76145 , n76146 , n76147 , n76148 , n76149 , n76150 , n76151 , n76152 , n76153 , n76154 , n76155 , n76156 , n76157 , n76158 , n76159 , n76160 , n76161 , n76162 , n76163 , n76164 , n76165 , n76166 , n76167 , n76168 , n76169 , n76170 , n76171 , n76172 , n76173 , n76174 , n76175 , n76176 , n76177 , n76178 , n76179 , n76180 , n76181 , n76182 , n76183 , n76184 , n76185 , n76186 , n76187 , n76188 , n76189 , n76190 , n76191 , n76192 , n76193 , n76194 , n76195 , n76196 , n76197 , n76198 , n76199 , n76200 , n76201 , n76202 , n76203 , n76204 , n76205 , n76206 , n76207 , n76208 , n76209 , n76210 , n76211 , n76212 , n76213 , n76214 , n76215 , n76216 , n76217 , n76218 , n76219 , n76220 , n76221 , n76222 , n76223 , n76224 , n76225 , n76226 , n76227 , n76228 , n76229 , n76230 , n76231 , n76232 , n76233 , n76234 , n76235 , n76236 , n76237 , n76238 , n76239 , n76240 , n76241 , n76242 , n76243 , n76244 , n76245 , n76246 , n76247 , n76248 , n76249 , n76250 , n76251 , n76252 , n76253 , n76254 , n76255 , n76256 , n76257 , n76258 , n76259 , n76260 , n76261 , n76262 , n76263 , n76264 , n76265 , n76266 , n76267 , n76268 , n76269 , n76270 , n76271 , n76272 , n76273 , n76274 , n76275 , n76276 , n76277 , n76278 , n76279 , n76280 , n76281 , n76282 , n76283 , n76284 , n76285 , n76286 , n76287 , n76288 , n76289 , n76290 , n76291 , n76292 , n76293 , n76294 , n76295 , n76296 , n76297 , n76298 , n76299 , n76300 , n76301 , n76302 , n76303 , n76304 , n76305 , n76306 , n76307 , n76308 , n76309 , n76310 , n76311 , n76312 , n76313 , n76314 , n76315 , n76316 , n76317 , n76318 , n76319 , n76320 , n76321 , n76322 , n76323 , n76324 , n76325 , n76326 , n76327 , n76328 , n76329 , n76330 , n76331 , n76332 , n76333 , n76334 , n76335 , n76336 , n76337 , n76338 , n76339 , n76340 , n76341 , n76342 , n76343 , n76344 , n76345 , n76346 , n76347 , n76348 , n76349 , n76350 , n76351 , n76352 , n76353 , n76354 , n76355 , n76356 , n76357 , n76358 , n76359 , n76360 , n76361 , n76362 , n76363 , n76364 , n76365 , n76366 , n76367 , n76368 , n76369 , n76370 , n76371 , n76372 , n76373 , n76374 , n76375 , n76376 , n76377 , n76378 , n76379 , n76380 , n76381 , n76382 , n76383 , n76384 , n76385 , n76386 , n76387 , n76388 , n76389 , n76390 , n76391 , n76392 , n76393 , n76394 , n76395 , n76396 , n76397 , n76398 , n76399 , n76400 , n76401 , n76402 , n76403 , n76404 , n76405 , n76406 , n76407 , n76408 , n76409 , n76410 , n76411 , n76412 , n76413 , n76414 , n76415 , n76416 , n76417 , n76418 , n76419 , n76420 , n76421 , n76422 , n76423 , n76424 , n76425 , n76426 , n76427 , n76428 , n76429 , n76430 , n76431 , n76432 , n76433 , n76434 , n76435 , n76436 , n76437 , n76438 , n76439 , n76440 , n76441 , n76442 , n76443 , n76444 , n76445 , n76446 , n76447 , n76448 , n76449 , n76450 , n76451 , n76452 , n76453 , n76454 , n76455 , n76456 , n76457 , n76458 , n76459 , n76460 , n76461 , n76462 , n76463 , n76464 , n76465 , n76466 , n76467 , n76468 , n76469 , n76470 , n76471 , n76472 , n76473 , n76474 , n76475 , n76476 , n76477 , n76478 , n76479 , n76480 , n76481 , n76482 , n76483 , n76484 , n76485 , n76486 , n76487 , n76488 , n76489 , n76490 , n76491 , n76492 , n76493 , n76494 , n76495 , n76496 , n76497 , n76498 , n76499 , n76500 , n76501 , n76502 , n76503 , n76504 , n76505 , n76506 , n76507 , n76508 , n76509 , n76510 , n76511 , n76512 , n76513 , n76514 , n76515 , n76516 , n76517 , n76518 , n76519 , n76520 , n76521 , n76522 , n76523 , n76524 , n76525 , n76526 , n76527 , n76528 , n76529 , n76530 , n76531 , n76532 , n76533 , n76534 , n76535 , n76536 , n76537 , n76538 , n76539 , n76540 , n76541 , n76542 , n76543 , n76544 , n76545 , n76546 , n76547 , n76548 , n76549 , n76550 , n76551 , n76552 , n76553 , n76554 , n76555 , n76556 , n76557 , n76558 , n76559 , n76560 , n76561 , n76562 , n76563 , n76564 , n76565 , n76566 , n76567 , n76568 , n76569 , n76570 , n76571 , n76572 , n76573 , n76574 , n76575 , n76576 , n76577 , n76578 , n76579 , n76580 , n76581 , n76582 , n76583 , n76584 , n76585 , n76586 , n76587 , n76588 , n76589 , n76590 , n76591 , n76592 , n76593 , n76594 , n76595 , n76596 , n76597 , n76598 , n76599 , n76600 , n76601 , n76602 , n76603 , n76604 , n76605 , n76606 , n76607 , n76608 , n76609 , n76610 , n76611 , n76612 , n76613 , n76614 , n76615 , n76616 , n76617 , n76618 , n76619 , n76620 , n76621 , n76622 , n76623 , n76624 , n76625 , n76626 , n76627 , n76628 , n76629 , n76630 , n76631 , n76632 , n76633 , n76634 , n76635 , n76636 , n76637 , n76638 , n76639 , n76640 , n76641 , n76642 , n76643 , n76644 , n76645 , n76646 , n76647 , n76648 , n76649 , n76650 , n76651 , n76652 , n76653 , n76654 , n76655 , n76656 , n76657 , n76658 , n76659 , n76660 , n76661 , n76662 , n76663 , n76664 , n76665 , n76666 , n76667 , n76668 , n76669 , n76670 , n76671 , n76672 , n76673 , n76674 , n76675 , n76676 , n76677 , n76678 , n76679 , n76680 , n76681 , n76682 , n76683 , n76684 , n76685 , n76686 , n76687 , n76688 , n76689 , n76690 , n76691 , n76692 , n76693 , n76694 , n76695 , n76696 , n76697 , n76698 , n76699 , n76700 , n76701 , n76702 , n76703 , n76704 , n76705 , n76706 , n76707 , n76708 , n76709 , n76710 , n76711 , n76712 , n76713 , n76714 , n76715 , n76716 , n76717 , n76718 , n76719 , n76720 , n76721 , n76722 , n76723 , n76724 , n76725 , n76726 , n76727 , n76728 , n76729 , n76730 , n76731 , n76732 , n76733 , n76734 , n76735 , n76736 , n76737 , n76738 , n76739 , n76740 , n76741 , n76742 , n76743 , n76744 , n76745 , n76746 , n76747 , n76748 , n76749 , n76750 , n76751 , n76752 , n76753 , n76754 , n76755 , n76756 , n76757 , n76758 , n76759 , n76760 , n76761 , n76762 , n76763 , n76764 , n76765 , n76766 , n76767 , n76768 , n76769 , n76770 , n76771 , n76772 , n76773 , n76774 , n76775 , n76776 , n76777 , n76778 , n76779 , n76780 , n76781 , n76782 , n76783 , n76784 , n76785 , n76786 , n76787 , n76788 , n76789 , n76790 , n76791 , n76792 , n76793 , n76794 , n76795 , n76796 , n76797 , n76798 , n76799 , n76800 , n76801 , n76802 , n76803 , n76804 , n76805 , n76806 , n76807 , n76808 , n76809 , n76810 , n76811 , n76812 , n76813 , n76814 , n76815 , n76816 , n76817 , n76818 , n76819 , n76820 , n76821 , n76822 , n76823 , n76824 , n76825 , n76826 , n76827 , n76828 , n76829 , n76830 , n76831 , n76832 , n76833 , n76834 , n76835 , n76836 , n76837 , n76838 , n76839 , n76840 , n76841 , n76842 , n76843 , n76844 , n76845 , n76846 , n76847 , n76848 , n76849 , n76850 , n76851 , n76852 , n76853 , n76854 , n76855 , n76856 , n76857 , n76858 , n76859 , n76860 , n76861 , n76862 , n76863 , n76864 , n76865 , n76866 , n76867 , n76868 , n76869 , n76870 , n76871 , n76872 , n76873 , n76874 , n76875 , n76876 , n76877 , n76878 , n76879 , n76880 , n76881 , n76882 , n76883 , n76884 , n76885 , n76886 , n76887 , n76888 , n76889 , n76890 , n76891 , n76892 , n76893 , n76894 , n76895 , n76896 , n76897 , n76898 , n76899 , n76900 , n76901 , n76902 , n76903 , n76904 , n76905 , n76906 , n76907 , n76908 , n76909 , n76910 , n76911 , n76912 , n76913 , n76914 , n76915 , n76916 , n76917 , n76918 , n76919 , n76920 , n76921 , n76922 , n76923 , n76924 , n76925 , n76926 , n76927 , n76928 , n76929 , n76930 , n76931 , n76932 , n76933 , n76934 , n76935 , n76936 , n76937 , n76938 , n76939 , n76940 , n76941 , n76942 , n76943 , n76944 , n76945 , n76946 , n76947 , n76948 , n76949 , n76950 , n76951 , n76952 , n76953 , n76954 , n76955 , n76956 , n76957 , n76958 , n76959 , n76960 , n76961 , n76962 , n76963 , n76964 , n76965 , n76966 , n76967 , n76968 , n76969 , n76970 , n76971 , n76972 , n76973 , n76974 , n76975 , n76976 , n76977 , n76978 , n76979 , n76980 , n76981 , n76982 , n76983 , n76984 , n76985 , n76986 , n76987 , n76988 , n76989 , n76990 , n76991 , n76992 , n76993 , n76994 , n76995 , n76996 , n76997 , n76998 , n76999 , n77000 , n77001 , n77002 , n77003 , n77004 , n77005 , n77006 , n77007 , n77008 , n77009 , n77010 , n77011 , n77012 , n77013 , n77014 , n77015 , n77016 , n77017 , n77018 , n77019 , n77020 , n77021 , n77022 , n77023 , n77024 , n77025 , n77026 , n77027 , n77028 , n77029 , n77030 , n77031 , n77032 , n77033 , n77034 , n77035 , n77036 , n77037 , n77038 , n77039 , n77040 , n77041 , n77042 , n77043 , n77044 , n77045 , n77046 , n77047 , n77048 , n77049 , n77050 , n77051 , n77052 , n77053 , n77054 , n77055 , n77056 , n77057 , n77058 , n77059 , n77060 , n77061 , n77062 , n77063 , n77064 , n77065 , n77066 , n77067 , n77068 , n77069 , n77070 , n77071 , n77072 , n77073 , n77074 , n77075 , n77076 , n77077 , n77078 , n77079 , n77080 , n77081 , n77082 , n77083 , n77084 , n77085 , n77086 , n77087 , n77088 , n77089 , n77090 , n77091 , n77092 , n77093 , n77094 , n77095 , n77096 , n77097 , n77098 , n77099 , n77100 , n77101 , n77102 , n77103 , n77104 , n77105 , n77106 , n77107 , n77108 , n77109 , n77110 , n77111 , n77112 , n77113 , n77114 , n77115 , n77116 , n77117 , n77118 , n77119 , n77120 , n77121 , n77122 , n77123 , n77124 , n77125 , n77126 , n77127 , n77128 , n77129 , n77130 , n77131 , n77132 , n77133 , n77134 , n77135 , n77136 , n77137 , n77138 , n77139 , n77140 , n77141 , n77142 , n77143 , n77144 , n77145 , n77146 , n77147 , n77148 , n77149 , n77150 , n77151 , n77152 , n77153 , n77154 , n77155 , n77156 , n77157 , n77158 , n77159 , n77160 , n77161 , n77162 , n77163 , n77164 , n77165 , n77166 , n77167 , n77168 , n77169 , n77170 , n77171 , n77172 , n77173 , n77174 , n77175 , n77176 , n77177 , n77178 , n77179 , n77180 , n77181 , n77182 , n77183 , n77184 , n77185 , n77186 , n77187 , n77188 , n77189 , n77190 , n77191 , n77192 , n77193 , n77194 , n77195 , n77196 , n77197 , n77198 , n77199 , n77200 , n77201 , n77202 , n77203 , n77204 , n77205 , n77206 , n77207 , n77208 , n77209 , n77210 , n77211 , n77212 , n77213 , n77214 , n77215 , n77216 , n77217 , n77218 , n77219 , n77220 , n77221 , n77222 , n77223 , n77224 , n77225 , n77226 , n77227 , n77228 , n77229 , n77230 , n77231 , n77232 , n77233 , n77234 , n77235 , n77236 , n77237 , n77238 , n77239 , n77240 , n77241 , n77242 , n77243 , n77244 , n77245 , n77246 , n77247 , n77248 , n77249 , n77250 , n77251 , n77252 , n77253 , n77254 , n77255 , n77256 , n77257 , n77258 , n77259 , n77260 , n77261 , n77262 , n77263 , n77264 , n77265 , n77266 , n77267 , n77268 , n77269 , n77270 , n77271 , n77272 , n77273 , n77274 , n77275 , n77276 , n77277 , n77278 , n77279 , n77280 , n77281 , n77282 , n77283 , n77284 , n77285 , n77286 , n77287 , n77288 , n77289 , n77290 , n77291 , n77292 , n77293 , n77294 , n77295 , n77296 , n77297 , n77298 , n77299 , n77300 , n77301 , n77302 , n77303 , n77304 , n77305 , n77306 , n77307 , n77308 , n77309 , n77310 , n77311 , n77312 , n77313 , n77314 , n77315 , n77316 , n77317 , n77318 , n77319 , n77320 , n77321 , n77322 , n77323 , n77324 , n77325 , n77326 , n77327 , n77328 , n77329 , n77330 , n77331 , n77332 , n77333 , n77334 , n77335 , n77336 , n77337 , n77338 , n77339 , n77340 , n77341 , n77342 , n77343 , n77344 , n77345 , n77346 , n77347 , n77348 , n77349 , n77350 , n77351 , n77352 , n77353 , n77354 , n77355 , n77356 , n77357 , n77358 , n77359 , n77360 , n77361 , n77362 , n77363 , n77364 , n77365 , n77366 , n77367 , n77368 , n77369 , n77370 , n77371 , n77372 , n77373 , n77374 , n77375 , n77376 , n77377 , n77378 , n77379 , n77380 , n77381 , n77382 , n77383 , n77384 , n77385 , n77386 , n77387 , n77388 , n77389 , n77390 , n77391 , n77392 , n77393 , n77394 , n77395 , n77396 , n77397 , n77398 , n77399 , n77400 , n77401 , n77402 , n77403 , n77404 , n77405 , n77406 , n77407 , n77408 , n77409 , n77410 , n77411 , n77412 , n77413 , n77414 , n77415 , n77416 , n77417 , n77418 , n77419 , n77420 , n77421 , n77422 , n77423 , n77424 , n77425 , n77426 , n77427 , n77428 , n77429 , n77430 , n77431 , n77432 , n77433 , n77434 , n77435 , n77436 , n77437 , n77438 , n77439 , n77440 , n77441 , n77442 , n77443 , n77444 , n77445 , n77446 , n77447 , n77448 , n77449 , n77450 , n77451 , n77452 , n77453 , n77454 , n77455 , n77456 , n77457 , n77458 , n77459 , n77460 , n77461 , n77462 , n77463 , n77464 , n77465 , n77466 , n77467 , n77468 , n77469 , n77470 , n77471 , n77472 , n77473 , n77474 , n77475 , n77476 , n77477 , n77478 , n77479 , n77480 , n77481 , n77482 , n77483 , n77484 , n77485 , n77486 , n77487 , n77488 , n77489 , n77490 , n77491 , n77492 , n77493 , n77494 , n77495 , n77496 , n77497 , n77498 , n77499 , n77500 , n77501 , n77502 , n77503 , n77504 , n77505 , n77506 , n77507 , n77508 , n77509 , n77510 , n77511 , n77512 , n77513 , n77514 , n77515 , n77516 , n77517 , n77518 , n77519 , n77520 , n77521 , n77522 , n77523 , n77524 , n77525 , n77526 , n77527 , n77528 , n77529 , n77530 , n77531 , n77532 , n77533 , n77534 , n77535 , n77536 , n77537 , n77538 , n77539 , n77540 , n77541 , n77542 , n77543 , n77544 , n77545 , n77546 , n77547 , n77548 , n77549 , n77550 , n77551 , n77552 , n77553 , n77554 , n77555 , n77556 , n77557 , n77558 , n77559 , n77560 , n77561 , n77562 , n77563 , n77564 , n77565 , n77566 , n77567 , n77568 , n77569 , n77570 , n77571 , n77572 , n77573 , n77574 , n77575 , n77576 , n77577 , n77578 , n77579 , n77580 , n77581 , n77582 , n77583 , n77584 , n77585 , n77586 , n77587 , n77588 , n77589 , n77590 , n77591 , n77592 , n77593 , n77594 , n77595 , n77596 , n77597 , n77598 , n77599 , n77600 , n77601 , n77602 , n77603 , n77604 , n77605 , n77606 , n77607 , n77608 , n77609 , n77610 , n77611 , n77612 , n77613 , n77614 , n77615 , n77616 , n77617 , n77618 , n77619 , n77620 , n77621 , n77622 , n77623 , n77624 , n77625 , n77626 , n77627 , n77628 , n77629 , n77630 , n77631 , n77632 , n77633 , n77634 , n77635 , n77636 , n77637 , n77638 , n77639 , n77640 , n77641 , n77642 , n77643 , n77644 , n77645 , n77646 , n77647 , n77648 , n77649 , n77650 , n77651 , n77652 , n77653 , n77654 , n77655 , n77656 , n77657 , n77658 , n77659 , n77660 , n77661 , n77662 , n77663 , n77664 , n77665 , n77666 , n77667 , n77668 , n77669 , n77670 , n77671 , n77672 , n77673 , n77674 , n77675 , n77676 , n77677 , n77678 , n77679 , n77680 , n77681 , n77682 , n77683 , n77684 , n77685 , n77686 , n77687 , n77688 , n77689 , n77690 , n77691 , n77692 , n77693 , n77694 , n77695 , n77696 , n77697 , n77698 , n77699 , n77700 , n77701 , n77702 , n77703 , n77704 , n77705 , n77706 , n77707 , n77708 , n77709 , n77710 , n77711 , n77712 , n77713 , n77714 , n77715 , n77716 , n77717 , n77718 , n77719 , n77720 , n77721 , n77722 , n77723 , n77724 , n77725 , n77726 , n77727 , n77728 , n77729 , n77730 , n77731 , n77732 , n77733 , n77734 , n77735 , n77736 , n77737 , n77738 , n77739 , n77740 , n77741 , n77742 , n77743 , n77744 , n77745 , n77746 , n77747 , n77748 , n77749 , n77750 , n77751 , n77752 , n77753 , n77754 , n77755 , n77756 , n77757 , n77758 , n77759 , n77760 , n77761 , n77762 , n77763 , n77764 , n77765 , n77766 , n77767 , n77768 , n77769 , n77770 , n77771 , n77772 , n77773 , n77774 , n77775 , n77776 , n77777 , n77778 , n77779 , n77780 , n77781 , n77782 , n77783 , n77784 , n77785 , n77786 , n77787 , n77788 , n77789 , n77790 , n77791 , n77792 , n77793 , n77794 , n77795 , n77796 , n77797 , n77798 , n77799 , n77800 , n77801 , n77802 , n77803 , n77804 , n77805 , n77806 , n77807 , n77808 , n77809 , n77810 , n77811 , n77812 , n77813 , n77814 , n77815 , n77816 , n77817 , n77818 , n77819 , n77820 , n77821 , n77822 , n77823 , n77824 , n77825 , n77826 , n77827 , n77828 , n77829 , n77830 , n77831 , n77832 , n77833 , n77834 , n77835 , n77836 , n77837 , n77838 , n77839 , n77840 , n77841 , n77842 , n77843 , n77844 , n77845 , n77846 , n77847 , n77848 , n77849 , n77850 , n77851 , n77852 , n77853 , n77854 , n77855 , n77856 , n77857 , n77858 , n77859 , n77860 , n77861 , n77862 , n77863 , n77864 , n77865 , n77866 , n77867 , n77868 , n77869 , n77870 , n77871 , n77872 , n77873 , n77874 , n77875 , n77876 , n77877 , n77878 , n77879 , n77880 , n77881 , n77882 , n77883 , n77884 , n77885 , n77886 , n77887 , n77888 , n77889 , n77890 , n77891 , n77892 , n77893 , n77894 , n77895 , n77896 , n77897 , n77898 , n77899 , n77900 , n77901 , n77902 , n77903 , n77904 , n77905 , n77906 , n77907 , n77908 , n77909 , n77910 , n77911 , n77912 , n77913 , n77914 , n77915 , n77916 , n77917 , n77918 , n77919 , n77920 , n77921 , n77922 , n77923 , n77924 , n77925 , n77926 , n77927 , n77928 , n77929 , n77930 , n77931 , n77932 , n77933 , n77934 , n77935 , n77936 , n77937 , n77938 , n77939 , n77940 , n77941 , n77942 , n77943 , n77944 , n77945 , n77946 , n77947 , n77948 , n77949 , n77950 , n77951 , n77952 , n77953 , n77954 , n77955 , n77956 , n77957 , n77958 , n77959 , n77960 , n77961 , n77962 , n77963 , n77964 , n77965 , n77966 , n77967 , n77968 , n77969 , n77970 , n77971 , n77972 , n77973 , n77974 , n77975 , n77976 , n77977 , n77978 , n77979 , n77980 , n77981 , n77982 , n77983 , n77984 , n77985 , n77986 , n77987 , n77988 , n77989 , n77990 , n77991 , n77992 , n77993 , n77994 , n77995 , n77996 , n77997 , n77998 , n77999 , n78000 , n78001 , n78002 , n78003 , n78004 , n78005 , n78006 , n78007 , n78008 , n78009 , n78010 , n78011 , n78012 , n78013 , n78014 , n78015 , n78016 , n78017 , n78018 , n78019 , n78020 , n78021 , n78022 , n78023 , n78024 , n78025 , n78026 , n78027 , n78028 , n78029 , n78030 , n78031 , n78032 , n78033 , n78034 , n78035 , n78036 , n78037 , n78038 , n78039 , n78040 , n78041 , n78042 , n78043 , n78044 , n78045 , n78046 , n78047 , n78048 , n78049 , n78050 , n78051 , n78052 , n78053 , n78054 , n78055 , n78056 , n78057 , n78058 , n78059 , n78060 , n78061 , n78062 , n78063 , n78064 , n78065 , n78066 , n78067 , n78068 , n78069 , n78070 , n78071 , n78072 , n78073 , n78074 , n78075 , n78076 , n78077 , n78078 , n78079 , n78080 , n78081 , n78082 , n78083 , n78084 , n78085 , n78086 , n78087 , n78088 , n78089 , n78090 , n78091 , n78092 , n78093 , n78094 , n78095 , n78096 , n78097 , n78098 , n78099 , n78100 , n78101 , n78102 , n78103 , n78104 , n78105 , n78106 , n78107 , n78108 , n78109 , n78110 , n78111 , n78112 , n78113 , n78114 , n78115 , n78116 , n78117 , n78118 , n78119 , n78120 , n78121 , n78122 , n78123 , n78124 , n78125 , n78126 , n78127 , n78128 , n78129 , n78130 , n78131 , n78132 , n78133 , n78134 , n78135 , n78136 , n78137 , n78138 , n78139 , n78140 , n78141 , n78142 , n78143 , n78144 , n78145 , n78146 , n78147 , n78148 , n78149 , n78150 , n78151 , n78152 , n78153 , n78154 , n78155 , n78156 , n78157 , n78158 , n78159 , n78160 , n78161 , n78162 , n78163 , n78164 , n78165 , n78166 , n78167 , n78168 , n78169 , n78170 , n78171 , n78172 , n78173 , n78174 , n78175 , n78176 , n78177 , n78178 , n78179 , n78180 , n78181 , n78182 , n78183 , n78184 , n78185 , n78186 , n78187 , n78188 , n78189 , n78190 , n78191 , n78192 , n78193 , n78194 , n78195 , n78196 , n78197 , n78198 , n78199 , n78200 , n78201 , n78202 , n78203 , n78204 , n78205 , n78206 , n78207 , n78208 , n78209 , n78210 , n78211 , n78212 , n78213 , n78214 , n78215 , n78216 , n78217 , n78218 , n78219 , n78220 , n78221 , n78222 , n78223 , n78224 , n78225 , n78226 , n78227 , n78228 , n78229 , n78230 , n78231 , n78232 , n78233 , n78234 , n78235 , n78236 , n78237 , n78238 ;
  assign n5832 = decrypt_pad & ~\u1_uk_K_r3_reg[3]/NET0131  ;
  assign n5833 = ~decrypt_pad & ~\u1_uk_K_r3_reg[12]/NET0131  ;
  assign n5834 = ~n5832 & ~n5833 ;
  assign n5835 = \u1_R3_reg[1]/NET0131  & ~n5834 ;
  assign n5836 = ~\u1_R3_reg[1]/NET0131  & n5834 ;
  assign n5837 = ~n5835 & ~n5836 ;
  assign n5826 = decrypt_pad & ~\u1_uk_K_r3_reg[39]/NET0131  ;
  assign n5827 = ~decrypt_pad & ~\u1_uk_K_r3_reg[48]/NET0131  ;
  assign n5828 = ~n5826 & ~n5827 ;
  assign n5829 = \u1_R3_reg[32]/NET0131  & ~n5828 ;
  assign n5830 = ~\u1_R3_reg[32]/NET0131  & n5828 ;
  assign n5831 = ~n5829 & ~n5830 ;
  assign n5845 = decrypt_pad & ~\u1_uk_K_r3_reg[33]/NET0131  ;
  assign n5846 = ~decrypt_pad & ~\u1_uk_K_r3_reg[10]/NET0131  ;
  assign n5847 = ~n5845 & ~n5846 ;
  assign n5848 = \u1_R3_reg[5]/NET0131  & ~n5847 ;
  assign n5849 = ~\u1_R3_reg[5]/NET0131  & n5847 ;
  assign n5850 = ~n5848 & ~n5849 ;
  assign n5855 = n5831 & ~n5850 ;
  assign n5856 = ~n5837 & n5855 ;
  assign n5857 = n5831 & n5837 ;
  assign n5858 = n5850 & n5857 ;
  assign n5859 = ~n5856 & ~n5858 ;
  assign n5838 = ~n5831 & n5837 ;
  assign n5839 = decrypt_pad & ~\u1_uk_K_r3_reg[18]/NET0131  ;
  assign n5840 = ~decrypt_pad & ~\u1_uk_K_r3_reg[27]/NET0131  ;
  assign n5841 = ~n5839 & ~n5840 ;
  assign n5842 = \u1_R3_reg[2]/NET0131  & ~n5841 ;
  assign n5843 = ~\u1_R3_reg[2]/NET0131  & n5841 ;
  assign n5844 = ~n5842 & ~n5843 ;
  assign n5851 = n5844 & n5850 ;
  assign n5852 = ~n5844 & ~n5850 ;
  assign n5853 = ~n5851 & ~n5852 ;
  assign n5854 = n5838 & n5853 ;
  assign n5860 = decrypt_pad & ~\u1_uk_K_r3_reg[27]/NET0131  ;
  assign n5861 = ~decrypt_pad & ~\u1_uk_K_r3_reg[4]/NET0131  ;
  assign n5862 = ~n5860 & ~n5861 ;
  assign n5863 = \u1_R3_reg[3]/NET0131  & ~n5862 ;
  assign n5864 = ~\u1_R3_reg[3]/NET0131  & n5862 ;
  assign n5865 = ~n5863 & ~n5864 ;
  assign n5866 = ~n5854 & n5865 ;
  assign n5867 = n5859 & n5866 ;
  assign n5869 = ~n5831 & n5850 ;
  assign n5870 = ~n5837 & ~n5855 ;
  assign n5871 = ~n5869 & n5870 ;
  assign n5868 = ~n5831 & n5852 ;
  assign n5872 = ~n5865 & ~n5868 ;
  assign n5873 = ~n5871 & n5872 ;
  assign n5874 = ~n5867 & ~n5873 ;
  assign n5875 = n5844 & ~n5850 ;
  assign n5876 = n5837 & n5875 ;
  assign n5877 = n5831 & n5876 ;
  assign n5878 = decrypt_pad & ~\u1_uk_K_r3_reg[5]/NET0131  ;
  assign n5879 = ~decrypt_pad & ~\u1_uk_K_r3_reg[39]/NET0131  ;
  assign n5880 = ~n5878 & ~n5879 ;
  assign n5881 = \u1_R3_reg[4]/NET0131  & ~n5880 ;
  assign n5882 = ~\u1_R3_reg[4]/NET0131  & n5880 ;
  assign n5883 = ~n5881 & ~n5882 ;
  assign n5884 = ~n5831 & ~n5837 ;
  assign n5885 = n5851 & n5884 ;
  assign n5886 = ~n5883 & ~n5885 ;
  assign n5887 = ~n5877 & n5886 ;
  assign n5888 = ~n5874 & n5887 ;
  assign n5892 = n5831 & n5844 ;
  assign n5893 = ~n5865 & ~n5892 ;
  assign n5894 = ~n5844 & n5884 ;
  assign n5895 = n5893 & ~n5894 ;
  assign n5898 = n5831 & n5850 ;
  assign n5899 = ~n5837 & ~n5844 ;
  assign n5900 = n5898 & n5899 ;
  assign n5896 = ~n5831 & n5844 ;
  assign n5897 = n5865 & ~n5896 ;
  assign n5901 = ~n5838 & n5897 ;
  assign n5902 = ~n5900 & n5901 ;
  assign n5903 = ~n5895 & ~n5902 ;
  assign n5889 = n5837 & n5852 ;
  assign n5890 = n5831 & n5889 ;
  assign n5891 = n5837 & n5851 ;
  assign n5904 = n5883 & ~n5891 ;
  assign n5905 = ~n5890 & n5904 ;
  assign n5906 = ~n5903 & n5905 ;
  assign n5907 = ~n5888 & ~n5906 ;
  assign n5908 = ~\u1_L3_reg[17]/NET0131  & n5907 ;
  assign n5909 = \u1_L3_reg[17]/NET0131  & ~n5907 ;
  assign n5910 = ~n5908 & ~n5909 ;
  assign n5941 = decrypt_pad & ~\u2_uk_K_r13_reg[7]/NET0131  ;
  assign n5942 = ~decrypt_pad & ~\u2_uk_K_r13_reg[45]/NET0131  ;
  assign n5943 = ~n5941 & ~n5942 ;
  assign n5944 = \u2_R13_reg[27]/P0001  & ~n5943 ;
  assign n5945 = ~\u2_R13_reg[27]/P0001  & n5943 ;
  assign n5946 = ~n5944 & ~n5945 ;
  assign n5917 = decrypt_pad & ~\u2_uk_K_r13_reg[9]/NET0131  ;
  assign n5918 = ~decrypt_pad & ~\u2_uk_K_r13_reg[43]/NET0131  ;
  assign n5919 = ~n5917 & ~n5918 ;
  assign n5920 = \u2_R13_reg[24]/NET0131  & ~n5919 ;
  assign n5921 = ~\u2_R13_reg[24]/NET0131  & n5919 ;
  assign n5922 = ~n5920 & ~n5921 ;
  assign n5911 = decrypt_pad & ~\u2_uk_K_r13_reg[29]/NET0131  ;
  assign n5912 = ~decrypt_pad & ~\u2_uk_K_r13_reg[8]/NET0131  ;
  assign n5913 = ~n5911 & ~n5912 ;
  assign n5914 = \u2_R13_reg[26]/NET0131  & ~n5913 ;
  assign n5915 = ~\u2_R13_reg[26]/NET0131  & n5913 ;
  assign n5916 = ~n5914 & ~n5915 ;
  assign n5924 = decrypt_pad & ~\u2_uk_K_r13_reg[44]/NET0131  ;
  assign n5925 = ~decrypt_pad & ~\u2_uk_K_r13_reg[23]/NET0131  ;
  assign n5926 = ~n5924 & ~n5925 ;
  assign n5927 = \u2_R13_reg[25]/NET0131  & ~n5926 ;
  assign n5928 = ~\u2_R13_reg[25]/NET0131  & n5926 ;
  assign n5929 = ~n5927 & ~n5928 ;
  assign n5931 = decrypt_pad & ~\u2_uk_K_r13_reg[45]/NET0131  ;
  assign n5932 = ~decrypt_pad & ~\u2_uk_K_r13_reg[51]/NET0131  ;
  assign n5933 = ~n5931 & ~n5932 ;
  assign n5934 = \u2_R13_reg[29]/NET0131  & ~n5933 ;
  assign n5935 = ~\u2_R13_reg[29]/NET0131  & n5933 ;
  assign n5936 = ~n5934 & ~n5935 ;
  assign n5954 = n5929 & n5936 ;
  assign n5955 = ~n5916 & n5954 ;
  assign n5956 = n5922 & n5955 ;
  assign n5948 = n5916 & n5922 ;
  assign n5957 = ~n5929 & n5948 ;
  assign n5958 = ~n5956 & ~n5957 ;
  assign n5959 = n5946 & ~n5958 ;
  assign n5947 = n5936 & ~n5946 ;
  assign n5949 = ~n5922 & n5929 ;
  assign n5950 = n5922 & ~n5929 ;
  assign n5951 = ~n5949 & ~n5950 ;
  assign n5952 = ~n5948 & ~n5951 ;
  assign n5953 = n5947 & n5952 ;
  assign n5938 = ~n5922 & n5936 ;
  assign n5939 = ~n5929 & n5938 ;
  assign n5940 = n5916 & n5939 ;
  assign n5923 = ~n5916 & ~n5922 ;
  assign n5930 = n5923 & ~n5929 ;
  assign n5937 = n5930 & ~n5936 ;
  assign n5960 = decrypt_pad & ~\u2_uk_K_r13_reg[49]/NET0131  ;
  assign n5961 = ~decrypt_pad & ~\u2_uk_K_r13_reg[28]/NET0131  ;
  assign n5962 = ~n5960 & ~n5961 ;
  assign n5963 = \u2_R13_reg[28]/NET0131  & ~n5962 ;
  assign n5964 = ~\u2_R13_reg[28]/NET0131  & n5962 ;
  assign n5965 = ~n5963 & ~n5964 ;
  assign n5966 = ~n5937 & n5965 ;
  assign n5967 = ~n5940 & n5966 ;
  assign n5968 = ~n5953 & n5967 ;
  assign n5969 = ~n5959 & n5968 ;
  assign n5980 = ~n5938 & ~n5949 ;
  assign n5977 = ~n5929 & ~n5936 ;
  assign n5978 = n5916 & ~n5922 ;
  assign n5979 = n5977 & ~n5978 ;
  assign n5976 = ~n5916 & n5936 ;
  assign n5981 = ~n5946 & ~n5976 ;
  assign n5982 = ~n5979 & n5981 ;
  assign n5983 = n5980 & n5982 ;
  assign n5972 = ~n5947 & n5950 ;
  assign n5973 = n5938 & ~n5946 ;
  assign n5974 = ~n5972 & ~n5973 ;
  assign n5975 = ~n5916 & ~n5974 ;
  assign n5970 = ~n5923 & ~n5948 ;
  assign n5971 = n5954 & ~n5970 ;
  assign n5984 = ~n5965 & ~n5971 ;
  assign n5985 = ~n5975 & n5984 ;
  assign n5986 = ~n5983 & n5985 ;
  assign n5987 = ~n5969 & ~n5986 ;
  assign n5990 = n5916 & n5949 ;
  assign n5991 = ~n5936 & n5990 ;
  assign n5992 = n5946 & ~n5979 ;
  assign n5993 = ~n5940 & n5992 ;
  assign n5994 = ~n5991 & n5993 ;
  assign n5988 = ~n5946 & n5970 ;
  assign n5989 = ~n5929 & ~n5946 ;
  assign n5995 = ~n5988 & ~n5989 ;
  assign n5996 = ~n5994 & n5995 ;
  assign n5997 = ~n5987 & ~n5996 ;
  assign n5998 = \u2_L13_reg[22]/NET0131  & n5997 ;
  assign n5999 = ~\u2_L13_reg[22]/NET0131  & ~n5997 ;
  assign n6000 = ~n5998 & ~n5999 ;
  assign n6001 = decrypt_pad & ~\u2_uk_K_r13_reg[20]/NET0131  ;
  assign n6002 = ~decrypt_pad & ~\u2_uk_K_r13_reg[24]/NET0131  ;
  assign n6003 = ~n6001 & ~n6002 ;
  assign n6004 = \u2_R13_reg[4]/NET0131  & ~n6003 ;
  assign n6005 = ~\u2_R13_reg[4]/NET0131  & n6003 ;
  assign n6006 = ~n6004 & ~n6005 ;
  assign n6007 = decrypt_pad & ~\u2_uk_K_r13_reg[10]/NET0131  ;
  assign n6008 = ~decrypt_pad & ~\u2_uk_K_r13_reg[46]/NET0131  ;
  assign n6009 = ~n6007 & ~n6008 ;
  assign n6010 = \u2_R13_reg[3]/NET0131  & ~n6009 ;
  assign n6011 = ~\u2_R13_reg[3]/NET0131  & n6009 ;
  assign n6012 = ~n6010 & ~n6011 ;
  assign n6013 = decrypt_pad & ~\u2_uk_K_r13_reg[18]/NET0131  ;
  assign n6014 = ~decrypt_pad & ~\u2_uk_K_r13_reg[54]/NET0131  ;
  assign n6015 = ~n6013 & ~n6014 ;
  assign n6016 = \u2_R13_reg[1]/NET0131  & ~n6015 ;
  assign n6017 = ~\u2_R13_reg[1]/NET0131  & n6015 ;
  assign n6018 = ~n6016 & ~n6017 ;
  assign n6020 = decrypt_pad & ~\u2_uk_K_r13_reg[48]/NET0131  ;
  assign n6021 = ~decrypt_pad & ~\u2_uk_K_r13_reg[27]/NET0131  ;
  assign n6022 = ~n6020 & ~n6021 ;
  assign n6023 = \u2_R13_reg[5]/NET0131  & ~n6022 ;
  assign n6024 = ~\u2_R13_reg[5]/NET0131  & n6022 ;
  assign n6025 = ~n6023 & ~n6024 ;
  assign n6043 = ~n6018 & n6025 ;
  assign n6026 = decrypt_pad & ~\u2_uk_K_r13_reg[54]/NET0131  ;
  assign n6027 = ~decrypt_pad & ~\u2_uk_K_r13_reg[33]/NET0131  ;
  assign n6028 = ~n6026 & ~n6027 ;
  assign n6029 = \u2_R13_reg[32]/NET0131  & ~n6028 ;
  assign n6030 = ~\u2_R13_reg[32]/NET0131  & n6028 ;
  assign n6031 = ~n6029 & ~n6030 ;
  assign n6032 = ~n6025 & ~n6031 ;
  assign n6035 = decrypt_pad & ~\u2_uk_K_r13_reg[33]/NET0131  ;
  assign n6036 = ~decrypt_pad & ~\u2_uk_K_r13_reg[12]/NET0131  ;
  assign n6037 = ~n6035 & ~n6036 ;
  assign n6038 = \u2_R13_reg[2]/NET0131  & ~n6037 ;
  assign n6039 = ~\u2_R13_reg[2]/NET0131  & n6037 ;
  assign n6040 = ~n6038 & ~n6039 ;
  assign n6073 = n6032 & n6040 ;
  assign n6074 = ~n6043 & ~n6073 ;
  assign n6075 = n6012 & ~n6074 ;
  assign n6064 = n6025 & ~n6031 ;
  assign n6070 = n6012 & ~n6040 ;
  assign n6082 = n6018 & ~n6070 ;
  assign n6083 = n6064 & ~n6082 ;
  assign n6071 = ~n6018 & n6031 ;
  assign n6046 = ~n6018 & n6040 ;
  assign n6076 = ~n6012 & n6031 ;
  assign n6077 = ~n6046 & ~n6076 ;
  assign n6078 = ~n6071 & ~n6077 ;
  assign n6079 = ~n6018 & ~n6025 ;
  assign n6080 = n6031 & ~n6040 ;
  assign n6081 = n6079 & n6080 ;
  assign n6084 = ~n6078 & ~n6081 ;
  assign n6085 = ~n6083 & n6084 ;
  assign n6086 = ~n6075 & n6085 ;
  assign n6087 = n6006 & ~n6086 ;
  assign n6044 = ~n6031 & ~n6040 ;
  assign n6045 = ~n6043 & n6044 ;
  assign n6047 = ~n6025 & n6046 ;
  assign n6048 = n6031 & n6047 ;
  assign n6049 = ~n6045 & ~n6048 ;
  assign n6050 = ~n6012 & ~n6049 ;
  assign n6019 = n6012 & n6018 ;
  assign n6033 = n6025 & n6031 ;
  assign n6034 = ~n6032 & ~n6033 ;
  assign n6041 = n6034 & n6040 ;
  assign n6042 = n6019 & n6041 ;
  assign n6051 = n6018 & ~n6025 ;
  assign n6052 = ~n6043 & ~n6051 ;
  assign n6053 = ~n6019 & n6052 ;
  assign n6054 = ~n6034 & ~n6040 ;
  assign n6055 = ~n6053 & n6054 ;
  assign n6056 = ~n6042 & ~n6055 ;
  assign n6057 = ~n6050 & n6056 ;
  assign n6058 = ~n6006 & ~n6057 ;
  assign n6061 = n6025 & n6040 ;
  assign n6062 = n6018 & n6061 ;
  assign n6063 = n6031 & n6062 ;
  assign n6065 = n6040 & ~n6064 ;
  assign n6066 = ~n6046 & ~n6051 ;
  assign n6067 = ~n6065 & ~n6066 ;
  assign n6068 = ~n6063 & ~n6067 ;
  assign n6069 = ~n6012 & ~n6068 ;
  assign n6059 = n6012 & n6032 ;
  assign n6060 = n6046 & n6059 ;
  assign n6072 = n6070 & n6071 ;
  assign n6088 = ~n6060 & ~n6072 ;
  assign n6089 = ~n6069 & n6088 ;
  assign n6090 = ~n6058 & n6089 ;
  assign n6091 = ~n6087 & n6090 ;
  assign n6092 = ~\u2_L13_reg[31]/NET0131  & ~n6091 ;
  assign n6093 = \u2_L13_reg[31]/NET0131  & n6091 ;
  assign n6094 = ~n6092 & ~n6093 ;
  assign n6101 = decrypt_pad & ~\u2_uk_K_r13_reg[16]/NET0131  ;
  assign n6102 = ~decrypt_pad & ~\u2_uk_K_r13_reg[50]/NET0131  ;
  assign n6103 = ~n6101 & ~n6102 ;
  assign n6104 = \u2_R13_reg[23]/NET0131  & ~n6103 ;
  assign n6105 = ~\u2_R13_reg[23]/NET0131  & n6103 ;
  assign n6106 = ~n6104 & ~n6105 ;
  assign n6107 = decrypt_pad & ~\u2_uk_K_r13_reg[31]/NET0131  ;
  assign n6108 = ~decrypt_pad & ~\u2_uk_K_r13_reg[37]/NET0131  ;
  assign n6109 = ~n6107 & ~n6108 ;
  assign n6110 = \u2_R13_reg[22]/NET0131  & ~n6109 ;
  assign n6111 = ~\u2_R13_reg[22]/NET0131  & n6109 ;
  assign n6112 = ~n6110 & ~n6111 ;
  assign n6114 = decrypt_pad & ~\u2_uk_K_r13_reg[21]/NET0131  ;
  assign n6115 = ~decrypt_pad & ~\u2_uk_K_r13_reg[0]/NET0131  ;
  assign n6116 = ~n6114 & ~n6115 ;
  assign n6117 = \u2_R13_reg[20]/NET0131  & ~n6116 ;
  assign n6118 = ~\u2_R13_reg[20]/NET0131  & n6116 ;
  assign n6119 = ~n6117 & ~n6118 ;
  assign n6133 = decrypt_pad & ~\u2_uk_K_r13_reg[37]/NET0131  ;
  assign n6134 = ~decrypt_pad & ~\u2_uk_K_r13_reg[16]/NET0131  ;
  assign n6135 = ~n6133 & ~n6134 ;
  assign n6136 = \u2_R13_reg[25]/NET0131  & ~n6135 ;
  assign n6137 = ~\u2_R13_reg[25]/NET0131  & n6135 ;
  assign n6138 = ~n6136 & ~n6137 ;
  assign n6139 = n6119 & ~n6138 ;
  assign n6121 = decrypt_pad & ~\u2_uk_K_r13_reg[36]/NET0131  ;
  assign n6122 = ~decrypt_pad & ~\u2_uk_K_r13_reg[15]/NET0131  ;
  assign n6123 = ~n6121 & ~n6122 ;
  assign n6124 = \u2_R13_reg[21]/NET0131  & ~n6123 ;
  assign n6125 = ~\u2_R13_reg[21]/NET0131  & n6123 ;
  assign n6126 = ~n6124 & ~n6125 ;
  assign n6148 = ~n6119 & ~n6126 ;
  assign n6176 = ~n6139 & ~n6148 ;
  assign n6177 = n6112 & n6176 ;
  assign n6178 = n6126 & n6138 ;
  assign n6179 = ~n6119 & n6178 ;
  assign n6145 = n6119 & n6138 ;
  assign n6146 = ~n6126 & n6145 ;
  assign n6180 = ~n6112 & ~n6146 ;
  assign n6181 = ~n6179 & n6180 ;
  assign n6182 = ~n6177 & ~n6181 ;
  assign n6183 = ~n6106 & ~n6182 ;
  assign n6095 = decrypt_pad & ~\u2_uk_K_r13_reg[42]/NET0131  ;
  assign n6096 = ~decrypt_pad & ~\u2_uk_K_r13_reg[21]/NET0131  ;
  assign n6097 = ~n6095 & ~n6096 ;
  assign n6098 = \u2_R13_reg[24]/NET0131  & ~n6097 ;
  assign n6099 = ~\u2_R13_reg[24]/NET0131  & n6097 ;
  assign n6100 = ~n6098 & ~n6099 ;
  assign n6127 = n6112 & ~n6119 ;
  assign n6128 = n6126 & n6127 ;
  assign n6173 = n6106 & ~n6128 ;
  assign n6170 = ~n6112 & ~n6126 ;
  assign n6171 = n6139 & n6170 ;
  assign n6172 = n6126 & n6145 ;
  assign n6174 = ~n6171 & ~n6172 ;
  assign n6175 = n6173 & n6174 ;
  assign n6184 = n6100 & ~n6175 ;
  assign n6185 = ~n6183 & n6184 ;
  assign n6129 = ~n6112 & n6126 ;
  assign n6151 = n6129 & ~n6138 ;
  assign n6152 = n6119 & n6151 ;
  assign n6147 = n6112 & n6146 ;
  assign n6149 = n6138 & n6148 ;
  assign n6150 = n6106 & n6149 ;
  assign n6155 = ~n6147 & ~n6150 ;
  assign n6156 = ~n6152 & n6155 ;
  assign n6130 = n6119 & n6129 ;
  assign n6131 = ~n6128 & ~n6130 ;
  assign n6132 = ~n6106 & ~n6131 ;
  assign n6142 = n6119 & ~n6126 ;
  assign n6143 = n6106 & n6112 ;
  assign n6144 = n6142 & n6143 ;
  assign n6113 = n6106 & ~n6112 ;
  assign n6120 = n6113 & ~n6119 ;
  assign n6140 = ~n6106 & ~n6112 ;
  assign n6141 = n6139 & n6140 ;
  assign n6153 = ~n6120 & ~n6141 ;
  assign n6154 = ~n6144 & n6153 ;
  assign n6157 = ~n6132 & n6154 ;
  assign n6158 = n6156 & n6157 ;
  assign n6159 = ~n6100 & ~n6158 ;
  assign n6164 = n6126 & n6139 ;
  assign n6165 = ~n6106 & n6164 ;
  assign n6166 = ~n6150 & ~n6165 ;
  assign n6167 = ~n6112 & ~n6166 ;
  assign n6160 = n6112 & n6145 ;
  assign n6161 = ~n6119 & n6151 ;
  assign n6162 = ~n6160 & ~n6161 ;
  assign n6163 = n6106 & ~n6162 ;
  assign n6168 = ~n6138 & n6148 ;
  assign n6169 = n6140 & n6168 ;
  assign n6186 = ~n6163 & ~n6169 ;
  assign n6187 = ~n6167 & n6186 ;
  assign n6188 = ~n6159 & n6187 ;
  assign n6189 = ~n6185 & n6188 ;
  assign n6190 = ~\u2_L13_reg[11]/NET0131  & n6189 ;
  assign n6191 = \u2_L13_reg[11]/NET0131  & ~n6189 ;
  assign n6192 = ~n6190 & ~n6191 ;
  assign n6193 = decrypt_pad & ~\u2_uk_K_r13_reg[8]/NET0131  ;
  assign n6194 = ~decrypt_pad & ~\u2_uk_K_r13_reg[42]/NET0131  ;
  assign n6195 = ~n6193 & ~n6194 ;
  assign n6196 = \u2_R13_reg[31]/P0001  & ~n6195 ;
  assign n6197 = ~\u2_R13_reg[31]/P0001  & n6195 ;
  assign n6198 = ~n6196 & ~n6197 ;
  assign n6199 = decrypt_pad & ~\u2_uk_K_r13_reg[51]/NET0131  ;
  assign n6200 = ~decrypt_pad & ~\u2_uk_K_r13_reg[30]/NET0131  ;
  assign n6201 = ~n6199 & ~n6200 ;
  assign n6202 = \u2_R13_reg[30]/NET0131  & ~n6201 ;
  assign n6203 = ~\u2_R13_reg[30]/NET0131  & n6201 ;
  assign n6204 = ~n6202 & ~n6203 ;
  assign n6205 = decrypt_pad & ~\u2_uk_K_r13_reg[50]/NET0131  ;
  assign n6206 = ~decrypt_pad & ~\u2_uk_K_r13_reg[29]/NET0131  ;
  assign n6207 = ~n6205 & ~n6206 ;
  assign n6208 = \u2_R13_reg[29]/NET0131  & ~n6207 ;
  assign n6209 = ~\u2_R13_reg[29]/NET0131  & n6207 ;
  assign n6210 = ~n6208 & ~n6209 ;
  assign n6211 = ~n6204 & ~n6210 ;
  assign n6212 = decrypt_pad & ~\u2_uk_K_r13_reg[23]/NET0131  ;
  assign n6213 = ~decrypt_pad & ~\u2_uk_K_r13_reg[2]/NET0131  ;
  assign n6214 = ~n6212 & ~n6213 ;
  assign n6215 = \u2_R13_reg[28]/NET0131  & ~n6214 ;
  assign n6216 = ~\u2_R13_reg[28]/NET0131  & n6214 ;
  assign n6217 = ~n6215 & ~n6216 ;
  assign n6218 = n6211 & ~n6217 ;
  assign n6219 = ~n6198 & ~n6218 ;
  assign n6220 = ~n6204 & n6217 ;
  assign n6221 = decrypt_pad & ~\u2_uk_K_r13_reg[35]/NET0131  ;
  assign n6222 = ~decrypt_pad & ~\u2_uk_K_r13_reg[14]/NET0131  ;
  assign n6223 = ~n6221 & ~n6222 ;
  assign n6224 = \u2_R13_reg[1]/NET0131  & ~n6223 ;
  assign n6225 = ~\u2_R13_reg[1]/NET0131  & n6223 ;
  assign n6226 = ~n6224 & ~n6225 ;
  assign n6227 = n6210 & ~n6226 ;
  assign n6228 = ~n6220 & ~n6227 ;
  assign n6229 = n6210 & n6217 ;
  assign n6230 = ~n6226 & n6229 ;
  assign n6231 = ~n6204 & n6230 ;
  assign n6232 = ~n6228 & ~n6231 ;
  assign n6233 = n6198 & ~n6232 ;
  assign n6234 = ~n6219 & ~n6233 ;
  assign n6235 = n6210 & n6226 ;
  assign n6236 = ~n6217 & n6235 ;
  assign n6237 = n6204 & n6236 ;
  assign n6238 = ~n6234 & ~n6237 ;
  assign n6239 = decrypt_pad & ~\u2_uk_K_r13_reg[14]/NET0131  ;
  assign n6240 = ~decrypt_pad & ~\u2_uk_K_r13_reg[52]/NET0131  ;
  assign n6241 = ~n6239 & ~n6240 ;
  assign n6242 = \u2_R13_reg[32]/NET0131  & ~n6241 ;
  assign n6243 = ~\u2_R13_reg[32]/NET0131  & n6241 ;
  assign n6244 = ~n6242 & ~n6243 ;
  assign n6245 = ~n6238 & n6244 ;
  assign n6246 = ~n6217 & ~n6226 ;
  assign n6247 = ~n6210 & n6246 ;
  assign n6248 = ~n6204 & n6247 ;
  assign n6256 = n6198 & ~n6248 ;
  assign n6249 = ~n6210 & ~n6217 ;
  assign n6250 = n6226 & n6249 ;
  assign n6251 = n6204 & n6250 ;
  assign n6252 = ~n6204 & n6210 ;
  assign n6253 = n6217 & ~n6226 ;
  assign n6254 = ~n6252 & ~n6253 ;
  assign n6255 = ~n6228 & n6254 ;
  assign n6257 = ~n6251 & ~n6255 ;
  assign n6258 = n6256 & n6257 ;
  assign n6259 = n6204 & n6217 ;
  assign n6260 = ~n6210 & n6259 ;
  assign n6261 = n6244 & n6260 ;
  assign n6262 = ~n6198 & ~n6231 ;
  assign n6263 = ~n6261 & n6262 ;
  assign n6264 = ~n6258 & ~n6263 ;
  assign n6265 = ~n6226 & n6260 ;
  assign n6266 = n6198 & ~n6250 ;
  assign n6267 = ~n6265 & n6266 ;
  assign n6268 = n6204 & ~n6217 ;
  assign n6269 = ~n6226 & n6268 ;
  assign n6270 = ~n6198 & ~n6235 ;
  assign n6271 = ~n6269 & n6270 ;
  assign n6272 = ~n6267 & ~n6271 ;
  assign n6273 = ~n6198 & n6220 ;
  assign n6274 = n6235 & n6259 ;
  assign n6275 = ~n6273 & ~n6274 ;
  assign n6276 = ~n6231 & n6275 ;
  assign n6277 = ~n6272 & n6276 ;
  assign n6278 = ~n6244 & ~n6277 ;
  assign n6279 = ~n6264 & ~n6278 ;
  assign n6280 = ~n6245 & n6279 ;
  assign n6281 = \u2_L13_reg[5]/NET0131  & ~n6280 ;
  assign n6282 = ~\u2_L13_reg[5]/NET0131  & n6280 ;
  assign n6283 = ~n6281 & ~n6282 ;
  assign n6284 = decrypt_pad & ~\u2_uk_K_r13_reg[47]/NET0131  ;
  assign n6285 = ~decrypt_pad & ~\u2_uk_K_r13_reg[26]/NET0131  ;
  assign n6286 = ~n6284 & ~n6285 ;
  assign n6287 = \u2_R13_reg[16]/NET0131  & ~n6286 ;
  assign n6288 = ~\u2_R13_reg[16]/NET0131  & n6286 ;
  assign n6289 = ~n6287 & ~n6288 ;
  assign n6305 = decrypt_pad & ~\u2_uk_K_r13_reg[6]/NET0131  ;
  assign n6306 = ~decrypt_pad & ~\u2_uk_K_r13_reg[10]/NET0131  ;
  assign n6307 = ~n6305 & ~n6306 ;
  assign n6308 = \u2_R13_reg[14]/NET0131  & ~n6307 ;
  assign n6309 = ~\u2_R13_reg[14]/NET0131  & n6307 ;
  assign n6310 = ~n6308 & ~n6309 ;
  assign n6319 = decrypt_pad & ~\u2_uk_K_r13_reg[39]/NET0131  ;
  assign n6320 = ~decrypt_pad & ~\u2_uk_K_r13_reg[18]/NET0131  ;
  assign n6321 = ~n6319 & ~n6320 ;
  assign n6322 = \u2_R13_reg[15]/NET0131  & ~n6321 ;
  assign n6323 = ~\u2_R13_reg[15]/NET0131  & n6321 ;
  assign n6324 = ~n6322 & ~n6323 ;
  assign n6290 = decrypt_pad & ~\u2_uk_K_r13_reg[11]/NET0131  ;
  assign n6291 = ~decrypt_pad & ~\u2_uk_K_r13_reg[47]/NET0131  ;
  assign n6292 = ~n6290 & ~n6291 ;
  assign n6293 = \u2_R13_reg[12]/NET0131  & ~n6292 ;
  assign n6294 = ~\u2_R13_reg[12]/NET0131  & n6292 ;
  assign n6295 = ~n6293 & ~n6294 ;
  assign n6311 = decrypt_pad & ~\u2_uk_K_r13_reg[27]/NET0131  ;
  assign n6312 = ~decrypt_pad & ~\u2_uk_K_r13_reg[6]/NET0131  ;
  assign n6313 = ~n6311 & ~n6312 ;
  assign n6314 = \u2_R13_reg[17]/NET0131  & ~n6313 ;
  assign n6315 = ~\u2_R13_reg[17]/NET0131  & n6313 ;
  assign n6316 = ~n6314 & ~n6315 ;
  assign n6326 = ~n6295 & n6316 ;
  assign n6355 = n6324 & n6326 ;
  assign n6296 = decrypt_pad & ~\u2_uk_K_r13_reg[5]/NET0131  ;
  assign n6297 = ~decrypt_pad & ~\u2_uk_K_r13_reg[41]/NET0131  ;
  assign n6298 = ~n6296 & ~n6297 ;
  assign n6299 = \u2_R13_reg[13]/NET0131  & ~n6298 ;
  assign n6300 = ~\u2_R13_reg[13]/NET0131  & n6298 ;
  assign n6301 = ~n6299 & ~n6300 ;
  assign n6352 = ~n6301 & ~n6316 ;
  assign n6356 = ~n6301 & n6324 ;
  assign n6357 = n6295 & ~n6356 ;
  assign n6358 = ~n6352 & n6357 ;
  assign n6359 = ~n6355 & ~n6358 ;
  assign n6360 = ~n6310 & ~n6359 ;
  assign n6334 = ~n6310 & n6316 ;
  assign n6335 = n6295 & ~n6334 ;
  assign n6364 = n6335 & n6356 ;
  assign n6353 = ~n6295 & n6352 ;
  assign n6354 = ~n6324 & n6353 ;
  assign n6302 = ~n6295 & ~n6301 ;
  assign n6342 = ~n6310 & ~n6316 ;
  assign n6343 = n6302 & n6342 ;
  assign n6346 = ~n6295 & n6310 ;
  assign n6361 = n6301 & ~n6316 ;
  assign n6362 = n6346 & n6361 ;
  assign n6363 = ~n6343 & ~n6362 ;
  assign n6365 = ~n6354 & n6363 ;
  assign n6366 = ~n6364 & n6365 ;
  assign n6367 = ~n6360 & n6366 ;
  assign n6368 = ~n6289 & ~n6367 ;
  assign n6303 = n6295 & n6301 ;
  assign n6304 = ~n6302 & ~n6303 ;
  assign n6317 = n6310 & n6316 ;
  assign n6318 = ~n6304 & n6317 ;
  assign n6325 = ~n6318 & n6324 ;
  assign n6327 = n6301 & ~n6310 ;
  assign n6328 = n6326 & n6327 ;
  assign n6329 = n6295 & ~n6316 ;
  assign n6330 = ~n6327 & n6329 ;
  assign n6331 = ~n6328 & ~n6330 ;
  assign n6332 = ~n6318 & n6331 ;
  assign n6333 = ~n6325 & ~n6332 ;
  assign n6336 = n6301 & n6316 ;
  assign n6337 = ~n6302 & n6324 ;
  assign n6338 = ~n6336 & n6337 ;
  assign n6339 = ~n6335 & n6338 ;
  assign n6340 = ~n6333 & ~n6339 ;
  assign n6341 = n6289 & ~n6340 ;
  assign n6344 = ~n6318 & ~n6343 ;
  assign n6345 = ~n6324 & ~n6344 ;
  assign n6347 = n6295 & ~n6310 ;
  assign n6348 = ~n6346 & ~n6347 ;
  assign n6349 = n6301 & n6324 ;
  assign n6350 = ~n6334 & n6349 ;
  assign n6351 = ~n6348 & n6350 ;
  assign n6369 = ~n6345 & ~n6351 ;
  assign n6370 = ~n6341 & n6369 ;
  assign n6371 = ~n6368 & n6370 ;
  assign n6372 = \u2_L13_reg[10]/NET0131  & n6371 ;
  assign n6373 = ~\u2_L13_reg[10]/NET0131  & ~n6371 ;
  assign n6374 = ~n6372 & ~n6373 ;
  assign n6379 = n5922 & n5929 ;
  assign n6380 = ~n5937 & ~n6379 ;
  assign n6381 = n5946 & ~n6380 ;
  assign n6375 = n5940 & ~n5946 ;
  assign n6376 = n5916 & ~n5936 ;
  assign n6377 = ~n5976 & ~n6376 ;
  assign n6378 = ~n5951 & ~n6377 ;
  assign n6382 = n5965 & ~n6378 ;
  assign n6383 = ~n6375 & n6382 ;
  assign n6384 = ~n6381 & n6383 ;
  assign n6388 = ~n5939 & n5946 ;
  assign n6389 = ~n5954 & ~n5977 ;
  assign n6390 = ~n5946 & ~n5948 ;
  assign n6391 = n6389 & n6390 ;
  assign n6392 = ~n6388 & ~n6391 ;
  assign n6385 = n5952 & n6377 ;
  assign n6386 = n5936 & n5957 ;
  assign n6387 = n5977 & n5978 ;
  assign n6393 = ~n5965 & ~n6387 ;
  assign n6394 = ~n6386 & n6393 ;
  assign n6395 = ~n6385 & n6394 ;
  assign n6396 = ~n6392 & n6395 ;
  assign n6397 = ~n6384 & ~n6396 ;
  assign n6398 = \u2_L13_reg[12]/NET0131  & n6397 ;
  assign n6399 = ~\u2_L13_reg[12]/NET0131  & ~n6397 ;
  assign n6400 = ~n6398 & ~n6399 ;
  assign n6461 = decrypt_pad & ~\u2_uk_K_r13_reg[30]/NET0131  ;
  assign n6462 = ~decrypt_pad & ~\u2_uk_K_r13_reg[9]/NET0131  ;
  assign n6463 = ~n6461 & ~n6462 ;
  assign n6464 = \u2_R13_reg[20]/NET0131  & ~n6463 ;
  assign n6465 = ~\u2_R13_reg[20]/NET0131  & n6463 ;
  assign n6466 = ~n6464 & ~n6465 ;
  assign n6433 = decrypt_pad & ~\u2_uk_K_r13_reg[15]/NET0131  ;
  assign n6434 = ~decrypt_pad & ~\u2_uk_K_r13_reg[49]/NET0131  ;
  assign n6435 = ~n6433 & ~n6434 ;
  assign n6436 = \u2_R13_reg[19]/NET0131  & ~n6435 ;
  assign n6437 = ~\u2_R13_reg[19]/NET0131  & n6435 ;
  assign n6438 = ~n6436 & ~n6437 ;
  assign n6421 = decrypt_pad & ~\u2_uk_K_r13_reg[28]/NET0131  ;
  assign n6422 = ~decrypt_pad & ~\u2_uk_K_r13_reg[7]/NET0131  ;
  assign n6423 = ~n6421 & ~n6422 ;
  assign n6424 = \u2_R13_reg[18]/NET0131  & ~n6423 ;
  assign n6425 = ~\u2_R13_reg[18]/NET0131  & n6423 ;
  assign n6426 = ~n6424 & ~n6425 ;
  assign n6401 = decrypt_pad & ~\u2_uk_K_r13_reg[38]/NET0131  ;
  assign n6402 = ~decrypt_pad & ~\u2_uk_K_r13_reg[44]/NET0131  ;
  assign n6403 = ~n6401 & ~n6402 ;
  assign n6404 = \u2_R13_reg[17]/NET0131  & ~n6403 ;
  assign n6405 = ~\u2_R13_reg[17]/NET0131  & n6403 ;
  assign n6406 = ~n6404 & ~n6405 ;
  assign n6407 = decrypt_pad & ~\u2_uk_K_r13_reg[43]/NET0131  ;
  assign n6408 = ~decrypt_pad & ~\u2_uk_K_r13_reg[22]/NET0131  ;
  assign n6409 = ~n6407 & ~n6408 ;
  assign n6410 = \u2_R13_reg[16]/NET0131  & ~n6409 ;
  assign n6411 = ~\u2_R13_reg[16]/NET0131  & n6409 ;
  assign n6412 = ~n6410 & ~n6411 ;
  assign n6413 = n6406 & n6412 ;
  assign n6414 = decrypt_pad & ~\u2_uk_K_r13_reg[0]/NET0131  ;
  assign n6415 = ~decrypt_pad & ~\u2_uk_K_r13_reg[38]/NET0131  ;
  assign n6416 = ~n6414 & ~n6415 ;
  assign n6417 = \u2_R13_reg[21]/NET0131  & ~n6416 ;
  assign n6418 = ~\u2_R13_reg[21]/NET0131  & n6416 ;
  assign n6419 = ~n6417 & ~n6418 ;
  assign n6451 = n6413 & n6419 ;
  assign n6486 = ~n6426 & n6451 ;
  assign n6440 = ~n6406 & n6412 ;
  assign n6468 = ~n6419 & ~n6426 ;
  assign n6487 = n6440 & n6468 ;
  assign n6445 = ~n6412 & n6419 ;
  assign n6473 = ~n6406 & n6445 ;
  assign n6475 = n6406 & n6426 ;
  assign n6481 = ~n6419 & n6475 ;
  assign n6488 = ~n6473 & ~n6481 ;
  assign n6489 = ~n6487 & n6488 ;
  assign n6490 = ~n6486 & n6489 ;
  assign n6491 = ~n6438 & ~n6490 ;
  assign n6441 = n6419 & n6440 ;
  assign n6479 = n6426 & n6441 ;
  assign n6427 = n6406 & ~n6426 ;
  assign n6428 = ~n6412 & n6427 ;
  assign n6429 = n6412 & n6426 ;
  assign n6430 = n6419 & ~n6429 ;
  assign n6431 = ~n6428 & n6430 ;
  assign n6480 = ~n6419 & n6428 ;
  assign n6454 = n6412 & ~n6419 ;
  assign n6482 = n6438 & ~n6454 ;
  assign n6483 = ~n6481 & n6482 ;
  assign n6484 = ~n6480 & ~n6483 ;
  assign n6485 = ~n6431 & ~n6484 ;
  assign n6492 = ~n6479 & ~n6485 ;
  assign n6493 = ~n6491 & n6492 ;
  assign n6494 = ~n6466 & ~n6493 ;
  assign n6420 = n6413 & ~n6419 ;
  assign n6432 = ~n6420 & ~n6431 ;
  assign n6439 = ~n6432 & n6438 ;
  assign n6444 = ~n6426 & ~n6438 ;
  assign n6446 = n6406 & n6445 ;
  assign n6447 = ~n6412 & ~n6419 ;
  assign n6448 = ~n6406 & n6447 ;
  assign n6449 = ~n6446 & ~n6448 ;
  assign n6450 = n6444 & ~n6449 ;
  assign n6442 = ~n6420 & ~n6441 ;
  assign n6443 = ~n6426 & ~n6442 ;
  assign n6452 = n6426 & ~n6438 ;
  assign n6453 = n6451 & n6452 ;
  assign n6455 = ~n6406 & n6426 ;
  assign n6456 = n6454 & n6455 ;
  assign n6457 = ~n6453 & ~n6456 ;
  assign n6458 = ~n6443 & n6457 ;
  assign n6459 = ~n6450 & n6458 ;
  assign n6460 = ~n6439 & n6459 ;
  assign n6467 = ~n6460 & n6466 ;
  assign n6469 = n6413 & n6468 ;
  assign n6470 = n6426 & n6448 ;
  assign n6471 = ~n6469 & ~n6470 ;
  assign n6472 = n6438 & ~n6471 ;
  assign n6474 = n6426 & n6473 ;
  assign n6476 = n6447 & n6475 ;
  assign n6477 = ~n6474 & ~n6476 ;
  assign n6478 = ~n6438 & ~n6477 ;
  assign n6495 = ~n6472 & ~n6478 ;
  assign n6496 = ~n6467 & n6495 ;
  assign n6497 = ~n6494 & n6496 ;
  assign n6498 = ~\u2_L13_reg[14]/NET0131  & ~n6497 ;
  assign n6499 = \u2_L13_reg[14]/NET0131  & n6497 ;
  assign n6500 = ~n6498 & ~n6499 ;
  assign n6504 = n6018 & ~n6044 ;
  assign n6505 = ~n6012 & ~n6034 ;
  assign n6506 = ~n6504 & n6505 ;
  assign n6501 = n6031 & n6052 ;
  assign n6502 = n6012 & n6501 ;
  assign n6503 = n6041 & ~n6052 ;
  assign n6507 = ~n6502 & ~n6503 ;
  assign n6508 = ~n6506 & n6507 ;
  assign n6509 = ~n6006 & ~n6508 ;
  assign n6510 = ~n6040 & n6064 ;
  assign n6511 = ~n6073 & ~n6510 ;
  assign n6512 = n6019 & ~n6511 ;
  assign n6514 = ~n6018 & ~n6040 ;
  assign n6515 = ~n6031 & ~n6514 ;
  assign n6516 = n6033 & n6514 ;
  assign n6517 = ~n6515 & ~n6516 ;
  assign n6518 = n6012 & ~n6517 ;
  assign n6519 = ~n6012 & ~n6080 ;
  assign n6520 = ~n6515 & n6519 ;
  assign n6513 = n6051 & n6080 ;
  assign n6521 = ~n6062 & ~n6513 ;
  assign n6522 = ~n6520 & n6521 ;
  assign n6523 = ~n6518 & n6522 ;
  assign n6524 = n6006 & ~n6523 ;
  assign n6525 = ~n6512 & ~n6524 ;
  assign n6526 = ~n6509 & n6525 ;
  assign n6527 = ~\u2_L13_reg[17]/NET0131  & ~n6526 ;
  assign n6528 = \u2_L13_reg[17]/NET0131  & n6526 ;
  assign n6529 = ~n6527 & ~n6528 ;
  assign n6530 = n6325 & ~n6362 ;
  assign n6531 = n6310 & ~n6316 ;
  assign n6532 = ~n6335 & ~n6531 ;
  assign n6533 = n6289 & n6301 ;
  assign n6534 = n6532 & n6533 ;
  assign n6535 = ~n6304 & n6531 ;
  assign n6536 = ~n6324 & ~n6535 ;
  assign n6537 = ~n6534 & n6536 ;
  assign n6538 = ~n6530 & ~n6537 ;
  assign n6539 = ~n6289 & ~n6328 ;
  assign n6543 = n6303 & n6317 ;
  assign n6546 = n6539 & ~n6543 ;
  assign n6540 = ~n6316 & n6324 ;
  assign n6541 = ~n6303 & n6540 ;
  assign n6542 = n6348 & n6541 ;
  assign n6544 = ~n6336 & ~n6531 ;
  assign n6545 = n6357 & n6544 ;
  assign n6547 = ~n6542 & ~n6545 ;
  assign n6548 = n6546 & n6547 ;
  assign n6551 = ~n6316 & ~n6347 ;
  assign n6552 = n6356 & ~n6551 ;
  assign n6549 = n6303 & n6531 ;
  assign n6550 = n6289 & ~n6549 ;
  assign n6553 = ~n6301 & n6346 ;
  assign n6554 = n6550 & ~n6553 ;
  assign n6555 = ~n6552 & n6554 ;
  assign n6556 = ~n6548 & ~n6555 ;
  assign n6557 = ~n6538 & ~n6556 ;
  assign n6558 = ~\u2_L13_reg[1]/NET0131  & ~n6557 ;
  assign n6559 = \u2_L13_reg[1]/NET0131  & n6557 ;
  assign n6560 = ~n6558 & ~n6559 ;
  assign n6565 = ~n6226 & ~n6259 ;
  assign n6563 = n6210 & n6220 ;
  assign n6564 = n6204 & ~n6210 ;
  assign n6566 = ~n6563 & ~n6564 ;
  assign n6567 = ~n6565 & n6566 ;
  assign n6568 = n6198 & ~n6567 ;
  assign n6569 = n6226 & n6260 ;
  assign n6570 = n6220 & ~n6226 ;
  assign n6571 = ~n6198 & ~n6570 ;
  assign n6572 = ~n6569 & n6571 ;
  assign n6573 = ~n6568 & ~n6572 ;
  assign n6574 = ~n6230 & ~n6247 ;
  assign n6575 = n6204 & ~n6574 ;
  assign n6576 = n6211 & n6226 ;
  assign n6577 = ~n6217 & n6576 ;
  assign n6578 = n6244 & ~n6577 ;
  assign n6579 = ~n6575 & n6578 ;
  assign n6580 = ~n6573 & n6579 ;
  assign n6583 = ~n6198 & n6210 ;
  assign n6584 = n6246 & n6583 ;
  assign n6590 = ~n6244 & ~n6584 ;
  assign n6591 = ~n6248 & n6590 ;
  assign n6587 = ~n6198 & n6226 ;
  assign n6588 = ~n6210 & ~n6587 ;
  assign n6589 = n6268 & ~n6588 ;
  assign n6592 = ~n6265 & ~n6589 ;
  assign n6593 = n6591 & n6592 ;
  assign n6581 = ~n6230 & ~n6260 ;
  assign n6582 = n6198 & ~n6581 ;
  assign n6585 = ~n6273 & ~n6563 ;
  assign n6586 = n6226 & ~n6585 ;
  assign n6594 = ~n6582 & ~n6586 ;
  assign n6595 = n6593 & n6594 ;
  assign n6596 = ~n6580 & ~n6595 ;
  assign n6561 = n6198 & n6218 ;
  assign n6562 = n6235 & n6273 ;
  assign n6597 = ~n6561 & ~n6562 ;
  assign n6598 = ~n6596 & n6597 ;
  assign n6599 = ~\u2_L13_reg[21]/NET0131  & ~n6598 ;
  assign n6600 = \u2_L13_reg[21]/NET0131  & n6598 ;
  assign n6601 = ~n6599 & ~n6600 ;
  assign n6608 = ~n6327 & ~n6336 ;
  assign n6609 = ~n6356 & n6608 ;
  assign n6610 = ~n6295 & ~n6334 ;
  assign n6611 = ~n6609 & n6610 ;
  assign n6602 = n6295 & n6316 ;
  assign n6603 = ~n6301 & n6316 ;
  assign n6604 = ~n6310 & n6603 ;
  assign n6605 = ~n6602 & ~n6604 ;
  assign n6606 = ~n6324 & ~n6347 ;
  assign n6607 = ~n6605 & n6606 ;
  assign n6612 = n6550 & ~n6607 ;
  assign n6613 = ~n6611 & n6612 ;
  assign n6614 = n6349 & ~n6532 ;
  assign n6615 = ~n6301 & n6347 ;
  assign n6616 = n6539 & ~n6615 ;
  assign n6617 = ~n6614 & n6616 ;
  assign n6618 = ~n6613 & ~n6617 ;
  assign n6624 = ~n6352 & ~n6553 ;
  assign n6625 = ~n6289 & ~n6624 ;
  assign n6620 = ~n6303 & n6316 ;
  assign n6619 = n6303 & ~n6316 ;
  assign n6621 = ~n6302 & ~n6310 ;
  assign n6622 = ~n6619 & n6621 ;
  assign n6623 = ~n6620 & n6622 ;
  assign n6626 = ~n6324 & ~n6623 ;
  assign n6627 = ~n6625 & n6626 ;
  assign n6628 = n6347 & n6603 ;
  assign n6629 = n6324 & ~n6328 ;
  assign n6630 = ~n6628 & n6629 ;
  assign n6631 = ~n6627 & ~n6630 ;
  assign n6632 = ~n6618 & ~n6631 ;
  assign n6633 = \u2_L13_reg[26]/NET0131  & n6632 ;
  assign n6634 = ~\u2_L13_reg[26]/NET0131  & ~n6632 ;
  assign n6635 = ~n6633 & ~n6634 ;
  assign n6638 = ~n6419 & ~n6427 ;
  assign n6639 = ~n6429 & n6638 ;
  assign n6637 = ~n6406 & ~n6412 ;
  assign n6640 = ~n6451 & ~n6637 ;
  assign n6641 = ~n6639 & n6640 ;
  assign n6642 = n6438 & ~n6641 ;
  assign n6643 = ~n6428 & ~n6441 ;
  assign n6644 = ~n6438 & ~n6643 ;
  assign n6636 = n6419 & n6427 ;
  assign n6645 = n6420 & n6426 ;
  assign n6646 = ~n6636 & ~n6645 ;
  assign n6647 = ~n6644 & n6646 ;
  assign n6648 = ~n6642 & n6647 ;
  assign n6649 = n6466 & ~n6648 ;
  assign n6658 = ~n6454 & ~n6475 ;
  assign n6659 = ~n6413 & ~n6438 ;
  assign n6660 = ~n6658 & n6659 ;
  assign n6656 = ~n6419 & n6438 ;
  assign n6657 = n6427 & n6656 ;
  assign n6654 = n6444 & n6637 ;
  assign n6655 = n6445 & n6475 ;
  assign n6661 = ~n6654 & ~n6655 ;
  assign n6662 = ~n6657 & n6661 ;
  assign n6663 = ~n6660 & n6662 ;
  assign n6664 = ~n6466 & ~n6663 ;
  assign n6650 = ~n6470 & ~n6645 ;
  assign n6651 = ~n6426 & n6473 ;
  assign n6652 = n6650 & ~n6651 ;
  assign n6653 = n6438 & ~n6652 ;
  assign n6665 = n6440 & n6452 ;
  assign n6666 = ~n6486 & ~n6665 ;
  assign n6667 = ~n6653 & n6666 ;
  assign n6668 = ~n6664 & n6667 ;
  assign n6669 = ~n6649 & n6668 ;
  assign n6670 = ~\u2_L13_reg[25]/NET0131  & ~n6669 ;
  assign n6671 = \u2_L13_reg[25]/NET0131  & n6669 ;
  assign n6672 = ~n6670 & ~n6671 ;
  assign n6696 = ~n6126 & n6139 ;
  assign n6697 = ~n6172 & ~n6696 ;
  assign n6698 = ~n6128 & ~n6170 ;
  assign n6699 = ~n6138 & ~n6698 ;
  assign n6700 = n6697 & ~n6699 ;
  assign n6701 = n6106 & ~n6700 ;
  assign n6673 = n6112 & n6164 ;
  assign n6693 = ~n6112 & n6176 ;
  assign n6694 = ~n6673 & ~n6693 ;
  assign n6695 = ~n6106 & ~n6694 ;
  assign n6702 = n6112 & n6149 ;
  assign n6703 = ~n6695 & ~n6702 ;
  assign n6704 = ~n6701 & n6703 ;
  assign n6705 = ~n6100 & ~n6704 ;
  assign n6674 = ~n6112 & ~n6119 ;
  assign n6675 = n6126 & n6674 ;
  assign n6676 = ~n6179 & ~n6675 ;
  assign n6677 = ~n6673 & n6676 ;
  assign n6678 = n6106 & ~n6677 ;
  assign n6679 = ~n6119 & ~n6138 ;
  assign n6683 = n6112 & n6679 ;
  assign n6684 = n6138 & n6674 ;
  assign n6685 = ~n6683 & ~n6684 ;
  assign n6686 = ~n6126 & ~n6685 ;
  assign n6680 = ~n6129 & n6679 ;
  assign n6681 = ~n6160 & ~n6680 ;
  assign n6682 = ~n6106 & ~n6681 ;
  assign n6687 = ~n6141 & ~n6147 ;
  assign n6688 = ~n6682 & n6687 ;
  assign n6689 = ~n6686 & n6688 ;
  assign n6690 = ~n6678 & n6689 ;
  assign n6691 = n6100 & ~n6690 ;
  assign n6692 = n6113 & n6178 ;
  assign n6706 = ~n6171 & ~n6692 ;
  assign n6707 = ~n6691 & n6706 ;
  assign n6708 = ~n6705 & n6707 ;
  assign n6709 = \u2_L13_reg[29]/NET0131  & ~n6708 ;
  assign n6710 = ~\u2_L13_reg[29]/NET0131  & n6708 ;
  assign n6711 = ~n6709 & ~n6710 ;
  assign n6718 = decrypt_pad & ~\u2_uk_K_r13_reg[13]/NET0131  ;
  assign n6719 = ~decrypt_pad & ~\u2_uk_K_r13_reg[17]/NET0131  ;
  assign n6720 = ~n6718 & ~n6719 ;
  assign n6721 = \u2_R13_reg[5]/NET0131  & ~n6720 ;
  assign n6722 = ~\u2_R13_reg[5]/NET0131  & n6720 ;
  assign n6723 = ~n6721 & ~n6722 ;
  assign n6725 = decrypt_pad & ~\u2_uk_K_r13_reg[34]/NET0131  ;
  assign n6726 = ~decrypt_pad & ~\u2_uk_K_r13_reg[13]/NET0131  ;
  assign n6727 = ~n6725 & ~n6726 ;
  assign n6728 = \u2_R13_reg[4]/NET0131  & ~n6727 ;
  assign n6729 = ~\u2_R13_reg[4]/NET0131  & n6727 ;
  assign n6730 = ~n6728 & ~n6729 ;
  assign n6732 = decrypt_pad & ~\u2_uk_K_r13_reg[26]/NET0131  ;
  assign n6733 = ~decrypt_pad & ~\u2_uk_K_r13_reg[5]/NET0131  ;
  assign n6734 = ~n6732 & ~n6733 ;
  assign n6735 = \u2_R13_reg[9]/NET0131  & ~n6734 ;
  assign n6736 = ~\u2_R13_reg[9]/NET0131  & n6734 ;
  assign n6737 = ~n6735 & ~n6736 ;
  assign n6739 = n6730 & ~n6737 ;
  assign n6740 = ~n6723 & ~n6739 ;
  assign n6741 = n6723 & n6730 ;
  assign n6742 = ~n6737 & n6741 ;
  assign n6743 = ~n6740 & ~n6742 ;
  assign n6744 = ~n6730 & n6737 ;
  assign n6712 = decrypt_pad & ~\u2_uk_K_r13_reg[4]/NET0131  ;
  assign n6713 = ~decrypt_pad & ~\u2_uk_K_r13_reg[40]/NET0131  ;
  assign n6714 = ~n6712 & ~n6713 ;
  assign n6715 = \u2_R13_reg[6]/NET0131  & ~n6714 ;
  assign n6716 = ~\u2_R13_reg[6]/NET0131  & n6714 ;
  assign n6717 = ~n6715 & ~n6716 ;
  assign n6745 = ~n6717 & ~n6730 ;
  assign n6746 = ~n6744 & ~n6745 ;
  assign n6747 = n6743 & n6746 ;
  assign n6748 = decrypt_pad & ~\u2_uk_K_r13_reg[55]/NET0131  ;
  assign n6749 = ~decrypt_pad & ~\u2_uk_K_r13_reg[34]/NET0131  ;
  assign n6750 = ~n6748 & ~n6749 ;
  assign n6751 = \u2_R13_reg[7]/NET0131  & ~n6750 ;
  assign n6752 = ~\u2_R13_reg[7]/NET0131  & n6750 ;
  assign n6753 = ~n6751 & ~n6752 ;
  assign n6754 = ~n6747 & n6753 ;
  assign n6755 = ~n6723 & n6737 ;
  assign n6756 = ~n6746 & ~n6755 ;
  assign n6757 = n6717 & n6742 ;
  assign n6724 = n6717 & ~n6723 ;
  assign n6731 = n6724 & ~n6730 ;
  assign n6758 = ~n6731 & ~n6753 ;
  assign n6759 = ~n6757 & n6758 ;
  assign n6760 = ~n6756 & n6759 ;
  assign n6761 = ~n6754 & ~n6760 ;
  assign n6762 = n6730 & n6755 ;
  assign n6763 = ~n6753 & ~n6762 ;
  assign n6764 = ~n6717 & n6730 ;
  assign n6765 = ~n6763 & n6764 ;
  assign n6738 = n6731 & n6737 ;
  assign n6766 = decrypt_pad & ~\u2_uk_K_r13_reg[46]/NET0131  ;
  assign n6767 = ~decrypt_pad & ~\u2_uk_K_r13_reg[25]/P0001  ;
  assign n6768 = ~n6766 & ~n6767 ;
  assign n6769 = \u2_R13_reg[8]/NET0131  & ~n6768 ;
  assign n6770 = ~\u2_R13_reg[8]/NET0131  & n6768 ;
  assign n6771 = ~n6769 & ~n6770 ;
  assign n6772 = ~n6738 & n6771 ;
  assign n6773 = ~n6765 & n6772 ;
  assign n6774 = ~n6761 & n6773 ;
  assign n6778 = n6753 & ~n6756 ;
  assign n6779 = n6730 & ~n6755 ;
  assign n6780 = ~n6724 & n6779 ;
  assign n6781 = ~n6730 & n6755 ;
  assign n6782 = ~n6780 & ~n6781 ;
  assign n6783 = n6759 & n6782 ;
  assign n6784 = ~n6778 & ~n6783 ;
  assign n6775 = n6717 & ~n6744 ;
  assign n6776 = n6740 & n6775 ;
  assign n6777 = ~n6757 & ~n6771 ;
  assign n6785 = ~n6776 & n6777 ;
  assign n6786 = ~n6784 & n6785 ;
  assign n6787 = ~n6774 & ~n6786 ;
  assign n6788 = ~\u2_L13_reg[28]/NET0131  & n6787 ;
  assign n6789 = \u2_L13_reg[28]/NET0131  & ~n6787 ;
  assign n6790 = ~n6788 & ~n6789 ;
  assign n6791 = n6717 & n6753 ;
  assign n6792 = n6762 & n6791 ;
  assign n6793 = n6717 & n6730 ;
  assign n6794 = ~n6755 & ~n6793 ;
  assign n6795 = n6763 & ~n6794 ;
  assign n6805 = ~n6792 & ~n6795 ;
  assign n6796 = n6723 & ~n6737 ;
  assign n6797 = ~n6781 & ~n6796 ;
  assign n6798 = ~n6717 & ~n6797 ;
  assign n6799 = n6717 & n6744 ;
  assign n6800 = n6723 & n6799 ;
  assign n6801 = ~n6717 & ~n6723 ;
  assign n6802 = n6737 & ~n6753 ;
  assign n6803 = n6801 & n6802 ;
  assign n6804 = ~n6800 & ~n6803 ;
  assign n6806 = ~n6798 & n6804 ;
  assign n6807 = n6805 & n6806 ;
  assign n6808 = ~n6771 & ~n6807 ;
  assign n6814 = ~n6723 & ~n6737 ;
  assign n6815 = ~n6775 & ~n6814 ;
  assign n6816 = ~n6779 & ~n6815 ;
  assign n6809 = ~n6717 & n6723 ;
  assign n6812 = n6730 & n6809 ;
  assign n6813 = n6737 & n6812 ;
  assign n6817 = ~n6737 & n6801 ;
  assign n6818 = n6730 & n6817 ;
  assign n6819 = ~n6813 & ~n6818 ;
  assign n6820 = ~n6816 & n6819 ;
  assign n6821 = n6771 & ~n6820 ;
  assign n6810 = ~n6724 & ~n6809 ;
  assign n6811 = n6744 & n6810 ;
  assign n6822 = ~n6753 & ~n6811 ;
  assign n6823 = ~n6821 & n6822 ;
  assign n6825 = n6717 & ~n6741 ;
  assign n6826 = ~n6740 & n6771 ;
  assign n6827 = ~n6825 & n6826 ;
  assign n6824 = n6731 & ~n6737 ;
  assign n6828 = n6753 & ~n6812 ;
  assign n6829 = ~n6824 & n6828 ;
  assign n6830 = ~n6827 & n6829 ;
  assign n6831 = ~n6823 & ~n6830 ;
  assign n6832 = ~n6808 & ~n6831 ;
  assign n6833 = \u2_L13_reg[2]/NET0131  & n6832 ;
  assign n6834 = ~\u2_L13_reg[2]/NET0131  & ~n6832 ;
  assign n6835 = ~n6833 & ~n6834 ;
  assign n6840 = ~n6164 & ~n6684 ;
  assign n6841 = ~n6147 & n6840 ;
  assign n6842 = n6106 & ~n6841 ;
  assign n6836 = n6126 & n6679 ;
  assign n6837 = ~n6702 & ~n6836 ;
  assign n6838 = ~n6106 & ~n6837 ;
  assign n6839 = n6140 & n6145 ;
  assign n6843 = ~n6171 & ~n6839 ;
  assign n6844 = ~n6838 & n6843 ;
  assign n6845 = ~n6842 & n6844 ;
  assign n6846 = ~n6100 & ~n6845 ;
  assign n6854 = ~n6151 & ~n6674 ;
  assign n6855 = ~n6106 & ~n6854 ;
  assign n6856 = n6112 & n6178 ;
  assign n6857 = n6113 & n6145 ;
  assign n6858 = ~n6856 & ~n6857 ;
  assign n6859 = ~n6161 & n6858 ;
  assign n6860 = ~n6855 & n6859 ;
  assign n6861 = n6100 & ~n6860 ;
  assign n6847 = ~n6168 & ~n6179 ;
  assign n6848 = ~n6164 & n6847 ;
  assign n6849 = n6143 & ~n6848 ;
  assign n6850 = n6112 & n6697 ;
  assign n6851 = ~n6112 & ~n6679 ;
  assign n6852 = ~n6106 & ~n6851 ;
  assign n6853 = ~n6850 & n6852 ;
  assign n6862 = ~n6849 & ~n6853 ;
  assign n6863 = ~n6861 & n6862 ;
  assign n6864 = ~n6846 & n6863 ;
  assign n6865 = ~\u2_L13_reg[4]/NET0131  & ~n6864 ;
  assign n6866 = \u2_L13_reg[4]/NET0131  & n6864 ;
  assign n6867 = ~n6865 & ~n6866 ;
  assign n6869 = n6724 & ~n6737 ;
  assign n6870 = n6763 & ~n6869 ;
  assign n6871 = n6753 & ~n6799 ;
  assign n6872 = ~n6817 & n6871 ;
  assign n6873 = ~n6870 & ~n6872 ;
  assign n6868 = n6745 & n6796 ;
  assign n6874 = n6771 & ~n6868 ;
  assign n6875 = n6804 & n6874 ;
  assign n6876 = ~n6873 & n6875 ;
  assign n6878 = n6744 & ~n6810 ;
  assign n6877 = ~n6730 & n6796 ;
  assign n6879 = ~n6753 & ~n6771 ;
  assign n6880 = ~n6877 & n6879 ;
  assign n6881 = ~n6818 & n6880 ;
  assign n6882 = ~n6878 & n6881 ;
  assign n6883 = ~n6876 & ~n6882 ;
  assign n6884 = ~n6757 & ~n6813 ;
  assign n6885 = ~n6883 & n6884 ;
  assign n6888 = ~n6717 & ~n6743 ;
  assign n6886 = n6775 & ~n6796 ;
  assign n6887 = n6744 & n6809 ;
  assign n6889 = n6753 & ~n6771 ;
  assign n6890 = ~n6887 & n6889 ;
  assign n6891 = ~n6886 & n6890 ;
  assign n6892 = ~n6888 & n6891 ;
  assign n6893 = ~n6885 & ~n6892 ;
  assign n6894 = ~\u2_L13_reg[13]/NET0131  & ~n6893 ;
  assign n6895 = \u2_L13_reg[13]/NET0131  & n6893 ;
  assign n6896 = ~n6894 & ~n6895 ;
  assign n6899 = n6119 & ~n6129 ;
  assign n6900 = ~n6836 & ~n6899 ;
  assign n6901 = n6106 & ~n6900 ;
  assign n6898 = ~n6106 & ~n6847 ;
  assign n6897 = n6112 & n6172 ;
  assign n6902 = ~n6100 & ~n6897 ;
  assign n6903 = ~n6898 & n6902 ;
  assign n6904 = ~n6901 & n6903 ;
  assign n6907 = n6112 & n6179 ;
  assign n6908 = ~n6106 & n6142 ;
  assign n6909 = n6100 & ~n6151 ;
  assign n6910 = ~n6908 & n6909 ;
  assign n6911 = ~n6907 & n6910 ;
  assign n6905 = ~n6130 & ~n6149 ;
  assign n6906 = n6106 & ~n6905 ;
  assign n6912 = ~n6686 & ~n6906 ;
  assign n6913 = n6911 & n6912 ;
  assign n6914 = ~n6904 & ~n6913 ;
  assign n6915 = n6140 & n6146 ;
  assign n6916 = ~n6167 & ~n6915 ;
  assign n6917 = ~n6914 & n6916 ;
  assign n6918 = \u2_L13_reg[19]/P0001  & n6917 ;
  assign n6919 = ~\u2_L13_reg[19]/P0001  & ~n6917 ;
  assign n6920 = ~n6918 & ~n6919 ;
  assign n6921 = n6076 & ~n6514 ;
  assign n6922 = ~n6059 & ~n6079 ;
  assign n6923 = ~n6921 & n6922 ;
  assign n6924 = ~n6047 & ~n6923 ;
  assign n6925 = ~n6012 & ~n6018 ;
  assign n6926 = n6061 & ~n6071 ;
  assign n6927 = ~n6925 & n6926 ;
  assign n6928 = ~n6924 & ~n6927 ;
  assign n6929 = ~n6006 & ~n6928 ;
  assign n6941 = n6019 & ~n6080 ;
  assign n6942 = n6034 & n6941 ;
  assign n6943 = ~n6060 & ~n6516 ;
  assign n6944 = ~n6942 & n6943 ;
  assign n6945 = n6006 & ~n6944 ;
  assign n6937 = ~n6031 & ~n6052 ;
  assign n6938 = ~n6048 & ~n6937 ;
  assign n6939 = n6006 & ~n6012 ;
  assign n6940 = ~n6938 & n6939 ;
  assign n6930 = n6064 & n6514 ;
  assign n6931 = ~n6513 & ~n6930 ;
  assign n6932 = ~n6063 & n6931 ;
  assign n6933 = ~n6012 & ~n6932 ;
  assign n6934 = n6018 & n6032 ;
  assign n6935 = ~n6071 & ~n6934 ;
  assign n6936 = n6070 & ~n6935 ;
  assign n6946 = ~n6933 & ~n6936 ;
  assign n6947 = ~n6940 & n6946 ;
  assign n6948 = ~n6945 & n6947 ;
  assign n6949 = ~n6929 & n6948 ;
  assign n6950 = ~\u2_L13_reg[23]/P0001  & n6949 ;
  assign n6951 = \u2_L13_reg[23]/P0001  & ~n6949 ;
  assign n6952 = ~n6950 & ~n6951 ;
  assign n6966 = n6246 & n6252 ;
  assign n6965 = n6217 & n6235 ;
  assign n6967 = n6198 & ~n6965 ;
  assign n6968 = ~n6966 & n6967 ;
  assign n6969 = ~n6230 & ~n6236 ;
  assign n6970 = n6219 & n6969 ;
  assign n6971 = ~n6968 & ~n6970 ;
  assign n6972 = ~n6237 & ~n6576 ;
  assign n6973 = ~n6265 & n6972 ;
  assign n6974 = ~n6971 & n6973 ;
  assign n6975 = n6244 & ~n6974 ;
  assign n6959 = n6227 & ~n6259 ;
  assign n6960 = ~n6244 & ~n6959 ;
  assign n6961 = ~n6564 & ~n6960 ;
  assign n6962 = n6226 & ~n6252 ;
  assign n6963 = n6198 & ~n6962 ;
  assign n6964 = ~n6961 & n6963 ;
  assign n6953 = ~n6231 & ~n6255 ;
  assign n6954 = ~n6198 & ~n6953 ;
  assign n6955 = n6259 & n6587 ;
  assign n6956 = ~n6584 & ~n6955 ;
  assign n6957 = ~n6251 & n6956 ;
  assign n6958 = ~n6244 & ~n6957 ;
  assign n6976 = ~n6954 & ~n6958 ;
  assign n6977 = ~n6964 & n6976 ;
  assign n6978 = ~n6975 & n6977 ;
  assign n6979 = \u2_L13_reg[27]/NET0131  & n6978 ;
  assign n6980 = ~\u2_L13_reg[27]/NET0131  & ~n6978 ;
  assign n6981 = ~n6979 & ~n6980 ;
  assign n6982 = n6376 & n6379 ;
  assign n6983 = ~n5946 & ~n6386 ;
  assign n6984 = n5922 & ~n5936 ;
  assign n6985 = ~n5938 & ~n6984 ;
  assign n6986 = n5929 & ~n6985 ;
  assign n6987 = ~n5916 & ~n6985 ;
  assign n6988 = ~n5949 & ~n6987 ;
  assign n6989 = ~n6986 & ~n6988 ;
  assign n6990 = n6983 & ~n6989 ;
  assign n6991 = n5922 & ~n6376 ;
  assign n6992 = n5980 & ~n6991 ;
  assign n6993 = n5946 & ~n5955 ;
  assign n6994 = ~n6992 & n6993 ;
  assign n6995 = ~n6990 & ~n6994 ;
  assign n6996 = ~n6982 & ~n6995 ;
  assign n6997 = n5965 & ~n6996 ;
  assign n7000 = ~n5916 & n5950 ;
  assign n7001 = ~n5946 & ~n6389 ;
  assign n7002 = ~n7000 & n7001 ;
  assign n6998 = ~n5955 & ~n5989 ;
  assign n6999 = n6991 & n6998 ;
  assign n7003 = ~n5991 & ~n6999 ;
  assign n7004 = ~n7002 & n7003 ;
  assign n7005 = ~n5965 & ~n7004 ;
  assign n7006 = ~n5946 & n5965 ;
  assign n7007 = n5940 & ~n7006 ;
  assign n7008 = ~n5956 & ~n5990 ;
  assign n7009 = ~n5946 & ~n7008 ;
  assign n7010 = ~n7007 & ~n7009 ;
  assign n7011 = ~n7005 & n7010 ;
  assign n7012 = ~n6997 & n7011 ;
  assign n7013 = \u2_L13_reg[32]/NET0131  & n7012 ;
  assign n7014 = ~\u2_L13_reg[32]/NET0131  & ~n7012 ;
  assign n7015 = ~n7013 & ~n7014 ;
  assign n7016 = decrypt_pad & ~\u2_uk_K_r13_reg[24]/NET0131  ;
  assign n7017 = ~decrypt_pad & ~\u2_uk_K_r13_reg[3]/NET0131  ;
  assign n7018 = ~n7016 & ~n7017 ;
  assign n7019 = \u2_R13_reg[12]/NET0131  & ~n7018 ;
  assign n7020 = ~\u2_R13_reg[12]/NET0131  & n7018 ;
  assign n7021 = ~n7019 & ~n7020 ;
  assign n7028 = decrypt_pad & ~\u2_uk_K_r13_reg[41]/NET0131  ;
  assign n7029 = ~decrypt_pad & ~\u2_uk_K_r13_reg[20]/NET0131  ;
  assign n7030 = ~n7028 & ~n7029 ;
  assign n7031 = \u2_R13_reg[11]/NET0131  & ~n7030 ;
  assign n7032 = ~\u2_R13_reg[11]/NET0131  & n7030 ;
  assign n7033 = ~n7031 & ~n7032 ;
  assign n7044 = decrypt_pad & ~\u2_uk_K_r13_reg[32]/NET0131  ;
  assign n7045 = ~decrypt_pad & ~\u2_uk_K_r13_reg[11]/NET0131  ;
  assign n7046 = ~n7044 & ~n7045 ;
  assign n7047 = \u2_R13_reg[9]/NET0131  & ~n7046 ;
  assign n7048 = ~\u2_R13_reg[9]/NET0131  & n7046 ;
  assign n7049 = ~n7047 & ~n7048 ;
  assign n7050 = decrypt_pad & ~\u2_uk_K_r13_reg[40]/NET0131  ;
  assign n7051 = ~decrypt_pad & ~\u2_uk_K_r13_reg[19]/NET0131  ;
  assign n7052 = ~n7050 & ~n7051 ;
  assign n7053 = \u2_R13_reg[10]/NET0131  & ~n7052 ;
  assign n7054 = ~\u2_R13_reg[10]/NET0131  & n7052 ;
  assign n7055 = ~n7053 & ~n7054 ;
  assign n7022 = decrypt_pad & ~\u2_uk_K_r13_reg[3]/NET0131  ;
  assign n7023 = ~decrypt_pad & ~\u2_uk_K_r13_reg[39]/NET0131  ;
  assign n7024 = ~n7022 & ~n7023 ;
  assign n7025 = \u2_R13_reg[8]/NET0131  & ~n7024 ;
  assign n7026 = ~\u2_R13_reg[8]/NET0131  & n7024 ;
  assign n7027 = ~n7025 & ~n7026 ;
  assign n7035 = decrypt_pad & ~\u2_uk_K_r13_reg[12]/NET0131  ;
  assign n7036 = ~decrypt_pad & ~\u2_uk_K_r13_reg[48]/NET0131  ;
  assign n7037 = ~n7035 & ~n7036 ;
  assign n7038 = \u2_R13_reg[13]/NET0131  & ~n7037 ;
  assign n7039 = ~\u2_R13_reg[13]/NET0131  & n7037 ;
  assign n7040 = ~n7038 & ~n7039 ;
  assign n7062 = ~n7027 & n7040 ;
  assign n7063 = n7055 & n7062 ;
  assign n7064 = n7049 & n7063 ;
  assign n7065 = ~n7033 & n7064 ;
  assign n7059 = n7049 & n7055 ;
  assign n7041 = ~n7027 & ~n7040 ;
  assign n7042 = n7027 & n7040 ;
  assign n7043 = ~n7041 & ~n7042 ;
  assign n7056 = ~n7049 & ~n7055 ;
  assign n7060 = ~n7043 & ~n7056 ;
  assign n7061 = ~n7059 & n7060 ;
  assign n7034 = ~n7027 & n7033 ;
  assign n7057 = ~n7034 & n7056 ;
  assign n7058 = n7043 & n7057 ;
  assign n7066 = ~n7027 & n7049 ;
  assign n7067 = n7033 & ~n7055 ;
  assign n7068 = n7066 & n7067 ;
  assign n7069 = ~n7040 & n7049 ;
  assign n7070 = n7027 & n7055 ;
  assign n7071 = n7069 & n7070 ;
  assign n7072 = ~n7068 & ~n7071 ;
  assign n7073 = ~n7058 & n7072 ;
  assign n7074 = ~n7061 & n7073 ;
  assign n7075 = ~n7065 & n7074 ;
  assign n7076 = ~n7021 & ~n7075 ;
  assign n7077 = n7021 & n7055 ;
  assign n7078 = ~n7027 & n7069 ;
  assign n7079 = n7077 & n7078 ;
  assign n7080 = n7040 & ~n7049 ;
  assign n7081 = n7027 & n7069 ;
  assign n7082 = ~n7063 & ~n7081 ;
  assign n7083 = ~n7080 & n7082 ;
  assign n7084 = n7021 & n7033 ;
  assign n7085 = ~n7083 & n7084 ;
  assign n7100 = ~n7079 & ~n7085 ;
  assign n7086 = n7055 & n7080 ;
  assign n7087 = n7041 & ~n7055 ;
  assign n7088 = ~n7049 & n7087 ;
  assign n7089 = ~n7086 & ~n7088 ;
  assign n7090 = n7033 & ~n7089 ;
  assign n7091 = n7021 & ~n7033 ;
  assign n7096 = n7042 & n7049 ;
  assign n7092 = n7049 & ~n7055 ;
  assign n7093 = n7040 & n7092 ;
  assign n7094 = n7027 & ~n7049 ;
  assign n7095 = ~n7040 & n7094 ;
  assign n7097 = ~n7093 & ~n7095 ;
  assign n7098 = ~n7096 & n7097 ;
  assign n7099 = n7091 & ~n7098 ;
  assign n7101 = ~n7090 & ~n7099 ;
  assign n7102 = n7100 & n7101 ;
  assign n7103 = ~n7076 & n7102 ;
  assign n7104 = ~\u2_L13_reg[6]/NET0131  & ~n7103 ;
  assign n7105 = \u2_L13_reg[6]/NET0131  & n7103 ;
  assign n7106 = ~n7104 & ~n7105 ;
  assign n7107 = n5946 & ~n5965 ;
  assign n7108 = n5916 & n6986 ;
  assign n7109 = n5916 & ~n5950 ;
  assign n7110 = n6985 & ~n7109 ;
  assign n7111 = ~n7108 & ~n7110 ;
  assign n7112 = n7107 & ~n7111 ;
  assign n7113 = ~n5916 & ~n5977 ;
  assign n7114 = n6985 & n7113 ;
  assign n7115 = ~n7006 & ~n7107 ;
  assign n7116 = ~n6386 & n7115 ;
  assign n7117 = ~n7114 & n7116 ;
  assign n7118 = ~n7108 & n7117 ;
  assign n7119 = ~n7112 & ~n7118 ;
  assign n7120 = ~n6387 & ~n7119 ;
  assign n7121 = ~n5949 & ~n6984 ;
  assign n7122 = n5916 & ~n7121 ;
  assign n7123 = ~n5930 & n5965 ;
  assign n7124 = ~n6986 & n7123 ;
  assign n7125 = ~n7122 & n7124 ;
  assign n7126 = n6983 & n7125 ;
  assign n7127 = ~n7120 & ~n7126 ;
  assign n7128 = \u2_L13_reg[7]/NET0131  & ~n7127 ;
  assign n7129 = ~\u2_L13_reg[7]/NET0131  & n7127 ;
  assign n7130 = ~n7128 & ~n7129 ;
  assign n7145 = ~n6426 & n6445 ;
  assign n7146 = ~n6441 & ~n6446 ;
  assign n7147 = ~n7145 & n7146 ;
  assign n7148 = ~n6438 & ~n7147 ;
  assign n7143 = ~n6451 & ~n6487 ;
  assign n7144 = n6438 & ~n7143 ;
  assign n7149 = ~n6428 & n6650 ;
  assign n7150 = ~n7144 & n7149 ;
  assign n7151 = ~n7148 & n7150 ;
  assign n7152 = ~n6466 & ~n7151 ;
  assign n7136 = ~n6426 & n6448 ;
  assign n7137 = ~n6441 & ~n7136 ;
  assign n7138 = n6438 & ~n7137 ;
  assign n7139 = n6412 & n6444 ;
  assign n7140 = n6477 & ~n7139 ;
  assign n7141 = ~n7138 & n7140 ;
  assign n7142 = n6466 & ~n7141 ;
  assign n7131 = ~n6419 & n6665 ;
  assign n7132 = ~n6427 & ~n6455 ;
  assign n7133 = n6445 & ~n7132 ;
  assign n7134 = ~n6481 & ~n7133 ;
  assign n7135 = n6438 & ~n7134 ;
  assign n7153 = ~n7131 & ~n7135 ;
  assign n7154 = ~n7142 & n7153 ;
  assign n7155 = ~n7152 & n7154 ;
  assign n7156 = ~\u2_L13_reg[8]/NET0131  & ~n7155 ;
  assign n7157 = \u2_L13_reg[8]/NET0131  & n7155 ;
  assign n7158 = ~n7156 & ~n7157 ;
  assign n7167 = n7033 & n7078 ;
  assign n7165 = n7040 & ~n7066 ;
  assign n7166 = ~n7094 & n7165 ;
  assign n7168 = ~n7095 & ~n7166 ;
  assign n7169 = ~n7167 & n7168 ;
  assign n7170 = ~n7055 & ~n7169 ;
  assign n7159 = n7041 & n7055 ;
  assign n7171 = n7027 & ~n7055 ;
  assign n7172 = ~n7040 & n7171 ;
  assign n7173 = ~n7159 & ~n7172 ;
  assign n7174 = ~n7033 & ~n7173 ;
  assign n7175 = n7021 & ~n7064 ;
  assign n7176 = ~n7174 & n7175 ;
  assign n7177 = ~n7170 & n7176 ;
  assign n7178 = n7040 & n7094 ;
  assign n7179 = n7033 & ~n7178 ;
  assign n7180 = ~n7042 & n7049 ;
  assign n7181 = ~n7041 & n7180 ;
  assign n7182 = n7179 & ~n7181 ;
  assign n7183 = ~n7033 & ~n7087 ;
  assign n7184 = ~n7166 & n7183 ;
  assign n7185 = ~n7182 & ~n7184 ;
  assign n7186 = ~n7021 & ~n7088 ;
  assign n7187 = ~n7185 & n7186 ;
  assign n7188 = ~n7177 & ~n7187 ;
  assign n7160 = ~n7049 & n7159 ;
  assign n7161 = ~n7071 & ~n7160 ;
  assign n7162 = n7033 & ~n7161 ;
  assign n7163 = ~n7033 & n7055 ;
  assign n7164 = n7094 & n7163 ;
  assign n7189 = ~n7162 & ~n7164 ;
  assign n7190 = ~n7188 & n7189 ;
  assign n7191 = ~\u2_L13_reg[16]/NET0131  & ~n7190 ;
  assign n7192 = \u2_L13_reg[16]/NET0131  & n7190 ;
  assign n7193 = ~n7191 & ~n7192 ;
  assign n7204 = ~n7043 & n7056 ;
  assign n7205 = n7082 & ~n7204 ;
  assign n7206 = ~n7033 & ~n7205 ;
  assign n7207 = ~n7021 & ~n7206 ;
  assign n7210 = ~n7033 & n7060 ;
  assign n7214 = n7021 & ~n7058 ;
  assign n7208 = ~n7049 & ~n7062 ;
  assign n7209 = n7067 & n7208 ;
  assign n7211 = n7033 & n7055 ;
  assign n7212 = ~n7041 & n7211 ;
  assign n7213 = ~n7094 & n7212 ;
  assign n7215 = ~n7209 & ~n7213 ;
  assign n7216 = n7214 & n7215 ;
  assign n7217 = ~n7210 & n7216 ;
  assign n7218 = ~n7207 & ~n7217 ;
  assign n7195 = ~n7055 & n7062 ;
  assign n7196 = ~n7159 & ~n7195 ;
  assign n7197 = n7055 & n7094 ;
  assign n7198 = ~n7078 & ~n7197 ;
  assign n7199 = n7196 & n7198 ;
  assign n7200 = n7033 & ~n7199 ;
  assign n7201 = n7055 & n7095 ;
  assign n7202 = ~n7200 & ~n7201 ;
  assign n7203 = ~n7021 & ~n7202 ;
  assign n7220 = n7034 & n7093 ;
  assign n7194 = n7067 & n7095 ;
  assign n7219 = n7096 & n7163 ;
  assign n7221 = ~n7194 & ~n7219 ;
  assign n7222 = ~n7220 & n7221 ;
  assign n7223 = ~n7203 & n7222 ;
  assign n7224 = ~n7218 & n7223 ;
  assign n7225 = ~\u2_L13_reg[24]/NET0131  & ~n7224 ;
  assign n7226 = \u2_L13_reg[24]/NET0131  & n7224 ;
  assign n7227 = ~n7225 & ~n7226 ;
  assign n7228 = ~n7069 & n7070 ;
  assign n7229 = ~n7040 & n7092 ;
  assign n7230 = ~n7228 & ~n7229 ;
  assign n7231 = n7033 & ~n7230 ;
  assign n7235 = ~n7027 & n7086 ;
  assign n7232 = ~n7066 & ~n7171 ;
  assign n7233 = ~n7033 & ~n7069 ;
  assign n7234 = ~n7232 & n7233 ;
  assign n7236 = ~n7204 & ~n7234 ;
  assign n7237 = ~n7235 & n7236 ;
  assign n7238 = ~n7231 & n7237 ;
  assign n7239 = ~n7021 & ~n7238 ;
  assign n7240 = n7033 & ~n7196 ;
  assign n7241 = ~n7194 & ~n7240 ;
  assign n7242 = n7021 & ~n7241 ;
  assign n7246 = n7055 & ~n7233 ;
  assign n7247 = ~n7179 & n7246 ;
  assign n7243 = ~n7070 & ~n7078 ;
  assign n7244 = n7091 & ~n7243 ;
  assign n7245 = n7077 & n7180 ;
  assign n7248 = ~n7244 & ~n7245 ;
  assign n7249 = ~n7247 & n7248 ;
  assign n7250 = ~n7242 & n7249 ;
  assign n7251 = ~n7239 & n7250 ;
  assign n7252 = \u2_L13_reg[30]/NET0131  & ~n7251 ;
  assign n7253 = ~\u2_L13_reg[30]/NET0131  & n7251 ;
  assign n7254 = ~n7252 & ~n7253 ;
  assign n7257 = n6438 & ~n6455 ;
  assign n7258 = n6419 & ~n6426 ;
  assign n7259 = ~n6454 & ~n7258 ;
  assign n7260 = ~n6441 & ~n7259 ;
  assign n7261 = ~n7257 & ~n7260 ;
  assign n7255 = ~n6420 & ~n7145 ;
  assign n7256 = n6438 & ~n7255 ;
  assign n7262 = ~n6466 & ~n7256 ;
  assign n7263 = ~n7261 & n7262 ;
  assign n7264 = n6412 & ~n7258 ;
  assign n7265 = n6438 & ~n6445 ;
  assign n7266 = ~n6637 & n7265 ;
  assign n7267 = ~n7264 & n7266 ;
  assign n7268 = ~n6438 & n6446 ;
  assign n7269 = ~n6456 & n6466 ;
  assign n7270 = ~n6486 & n7269 ;
  assign n7271 = ~n7268 & n7270 ;
  assign n7272 = ~n7267 & n7271 ;
  assign n7273 = ~n7263 & ~n7272 ;
  assign n7274 = ~n6438 & ~n6469 ;
  assign n7275 = ~n6479 & n7274 ;
  assign n7276 = ~n7136 & n7275 ;
  assign n7277 = n6438 & ~n6487 ;
  assign n7278 = ~n6474 & n7277 ;
  assign n7279 = ~n7276 & ~n7278 ;
  assign n7280 = ~n7273 & ~n7279 ;
  assign n7281 = ~\u2_L13_reg[3]/NET0131  & ~n7280 ;
  assign n7282 = \u2_L13_reg[3]/NET0131  & n7280 ;
  assign n7283 = ~n7281 & ~n7282 ;
  assign n7299 = ~n6501 & ~n6937 ;
  assign n7300 = n6040 & ~n7299 ;
  assign n7287 = ~n6033 & n6052 ;
  assign n7298 = n6070 & n7287 ;
  assign n7301 = ~n6513 & ~n7298 ;
  assign n7302 = ~n7300 & n7301 ;
  assign n7303 = n6006 & ~n7302 ;
  assign n7288 = ~n6012 & n7287 ;
  assign n7284 = n6018 & n6080 ;
  assign n7285 = n6012 & ~n6052 ;
  assign n7286 = ~n7284 & n7285 ;
  assign n7289 = ~n6034 & n6046 ;
  assign n7290 = n6025 & n7284 ;
  assign n7291 = ~n7289 & ~n7290 ;
  assign n7292 = ~n7286 & n7291 ;
  assign n7293 = ~n7288 & n7292 ;
  assign n7294 = ~n6006 & ~n7293 ;
  assign n7295 = ~n6031 & n6062 ;
  assign n7296 = ~n7290 & ~n7295 ;
  assign n7297 = ~n6012 & ~n7296 ;
  assign n7304 = ~n7294 & ~n7297 ;
  assign n7305 = ~n7303 & n7304 ;
  assign n7306 = ~\u2_L13_reg[9]/NET0131  & ~n7305 ;
  assign n7307 = \u2_L13_reg[9]/NET0131  & n7305 ;
  assign n7308 = ~n7306 & ~n7307 ;
  assign n7315 = n6753 & ~n6797 ;
  assign n7311 = n6717 & n6737 ;
  assign n7312 = n6730 & ~n6753 ;
  assign n7313 = ~n6796 & n7312 ;
  assign n7314 = ~n7311 & n7313 ;
  assign n7316 = n6771 & ~n6824 ;
  assign n7317 = ~n7314 & n7316 ;
  assign n7318 = ~n7315 & n7317 ;
  assign n7309 = n6723 & ~n6753 ;
  assign n7321 = n6730 & n6737 ;
  assign n7322 = ~n6801 & n7321 ;
  assign n7323 = ~n7309 & n7322 ;
  assign n7319 = ~n6730 & ~n6791 ;
  assign n7320 = n6810 & n7319 ;
  assign n7324 = ~n6817 & ~n7320 ;
  assign n7325 = ~n7323 & n7324 ;
  assign n7326 = n6777 & n7325 ;
  assign n7327 = ~n7318 & ~n7326 ;
  assign n7310 = n6744 & n7309 ;
  assign n7328 = n6730 & n7311 ;
  assign n7329 = ~n6868 & ~n7328 ;
  assign n7330 = n6753 & ~n7329 ;
  assign n7331 = ~n7310 & ~n7330 ;
  assign n7332 = ~n7327 & n7331 ;
  assign n7333 = ~\u2_L13_reg[18]/P0001  & ~n7332 ;
  assign n7334 = \u2_L13_reg[18]/P0001  & n7332 ;
  assign n7335 = ~n7333 & ~n7334 ;
  assign n7378 = decrypt_pad & ~\u2_uk_K_r12_reg[34]/NET0131  ;
  assign n7379 = ~decrypt_pad & ~\u2_uk_K_r12_reg[10]/P0001  ;
  assign n7380 = ~n7378 & ~n7379 ;
  assign n7381 = \u2_R12_reg[4]/NET0131  & ~n7380 ;
  assign n7382 = ~\u2_R12_reg[4]/NET0131  & n7380 ;
  assign n7383 = ~n7381 & ~n7382 ;
  assign n7355 = decrypt_pad & ~\u2_uk_K_r12_reg[32]/NET0131  ;
  assign n7356 = ~decrypt_pad & ~\u2_uk_K_r12_reg[40]/NET0131  ;
  assign n7357 = ~n7355 & ~n7356 ;
  assign n7358 = \u2_R12_reg[1]/NET0131  & ~n7357 ;
  assign n7359 = ~\u2_R12_reg[1]/NET0131  & n7357 ;
  assign n7360 = ~n7358 & ~n7359 ;
  assign n7336 = decrypt_pad & ~\u2_uk_K_r12_reg[24]/NET0131  ;
  assign n7337 = ~decrypt_pad & ~\u2_uk_K_r12_reg[32]/NET0131  ;
  assign n7338 = ~n7336 & ~n7337 ;
  assign n7339 = \u2_R12_reg[3]/NET0131  & ~n7338 ;
  assign n7340 = ~\u2_R12_reg[3]/NET0131  & n7338 ;
  assign n7341 = ~n7339 & ~n7340 ;
  assign n7342 = decrypt_pad & ~\u2_uk_K_r12_reg[47]/NET0131  ;
  assign n7343 = ~decrypt_pad & ~\u2_uk_K_r12_reg[55]/NET0131  ;
  assign n7344 = ~n7342 & ~n7343 ;
  assign n7345 = \u2_R12_reg[2]/NET0131  & ~n7344 ;
  assign n7346 = ~\u2_R12_reg[2]/NET0131  & n7344 ;
  assign n7347 = ~n7345 & ~n7346 ;
  assign n7348 = decrypt_pad & ~\u2_uk_K_r12_reg[5]/NET0131  ;
  assign n7349 = ~decrypt_pad & ~\u2_uk_K_r12_reg[13]/NET0131  ;
  assign n7350 = ~n7348 & ~n7349 ;
  assign n7351 = \u2_R12_reg[5]/NET0131  & ~n7350 ;
  assign n7352 = ~\u2_R12_reg[5]/NET0131  & n7350 ;
  assign n7353 = ~n7351 & ~n7352 ;
  assign n7362 = decrypt_pad & ~\u2_uk_K_r12_reg[11]/NET0131  ;
  assign n7363 = ~decrypt_pad & ~\u2_uk_K_r12_reg[19]/NET0131  ;
  assign n7364 = ~n7362 & ~n7363 ;
  assign n7365 = \u2_R12_reg[32]/NET0131  & ~n7364 ;
  assign n7366 = ~\u2_R12_reg[32]/NET0131  & n7364 ;
  assign n7367 = ~n7365 & ~n7366 ;
  assign n7368 = n7353 & ~n7367 ;
  assign n7369 = n7347 & n7368 ;
  assign n7417 = n7341 & n7369 ;
  assign n7354 = ~n7347 & ~n7353 ;
  assign n7418 = n7354 & ~n7367 ;
  assign n7419 = ~n7417 & ~n7418 ;
  assign n7420 = n7360 & ~n7419 ;
  assign n7385 = n7347 & n7360 ;
  assign n7412 = ~n7353 & n7385 ;
  assign n7413 = n7367 & n7412 ;
  assign n7410 = ~n7347 & n7367 ;
  assign n7414 = n7353 & n7410 ;
  assign n7415 = ~n7413 & ~n7414 ;
  assign n7416 = n7341 & ~n7415 ;
  assign n7374 = n7353 & ~n7360 ;
  assign n7421 = n7374 & n7410 ;
  assign n7422 = ~n7416 & ~n7421 ;
  assign n7423 = ~n7420 & n7422 ;
  assign n7424 = ~n7383 & ~n7423 ;
  assign n7397 = ~n7353 & ~n7367 ;
  assign n7398 = n7347 & n7397 ;
  assign n7399 = ~n7374 & ~n7398 ;
  assign n7400 = n7341 & ~n7399 ;
  assign n7392 = ~n7341 & n7360 ;
  assign n7393 = ~n7347 & ~n7360 ;
  assign n7394 = ~n7353 & n7393 ;
  assign n7395 = ~n7392 & ~n7394 ;
  assign n7396 = n7367 & ~n7395 ;
  assign n7401 = n7341 & ~n7347 ;
  assign n7402 = n7360 & ~n7401 ;
  assign n7403 = ~n7354 & ~n7367 ;
  assign n7404 = ~n7402 & n7403 ;
  assign n7405 = ~n7396 & ~n7404 ;
  assign n7406 = ~n7400 & n7405 ;
  assign n7407 = n7383 & ~n7406 ;
  assign n7371 = ~n7353 & ~n7360 ;
  assign n7372 = n7367 & n7371 ;
  assign n7373 = n7347 & n7372 ;
  assign n7375 = ~n7347 & ~n7367 ;
  assign n7376 = ~n7374 & n7375 ;
  assign n7377 = ~n7373 & ~n7376 ;
  assign n7384 = ~n7377 & ~n7383 ;
  assign n7370 = ~n7360 & n7369 ;
  assign n7361 = n7354 & n7360 ;
  assign n7386 = n7353 & n7367 ;
  assign n7387 = n7385 & n7386 ;
  assign n7388 = ~n7361 & ~n7387 ;
  assign n7389 = ~n7370 & n7388 ;
  assign n7390 = ~n7384 & n7389 ;
  assign n7391 = ~n7341 & ~n7390 ;
  assign n7408 = n7341 & ~n7360 ;
  assign n7409 = n7398 & n7408 ;
  assign n7411 = n7408 & n7410 ;
  assign n7425 = ~n7409 & ~n7411 ;
  assign n7426 = ~n7391 & n7425 ;
  assign n7427 = ~n7407 & n7426 ;
  assign n7428 = ~n7424 & n7427 ;
  assign n7429 = ~\u2_L12_reg[31]/NET0131  & ~n7428 ;
  assign n7430 = \u2_L12_reg[31]/NET0131  & n7428 ;
  assign n7431 = ~n7429 & ~n7430 ;
  assign n7438 = decrypt_pad & ~\u2_uk_K_r12_reg[30]/NET0131  ;
  assign n7439 = ~decrypt_pad & ~\u2_uk_K_r12_reg[36]/NET0131  ;
  assign n7440 = ~n7438 & ~n7439 ;
  assign n7441 = \u2_R12_reg[23]/NET0131  & ~n7440 ;
  assign n7442 = ~\u2_R12_reg[23]/NET0131  & n7440 ;
  assign n7443 = ~n7441 & ~n7442 ;
  assign n7444 = decrypt_pad & ~\u2_uk_K_r12_reg[45]/NET0131  ;
  assign n7445 = ~decrypt_pad & ~\u2_uk_K_r12_reg[23]/NET0131  ;
  assign n7446 = ~n7444 & ~n7445 ;
  assign n7447 = \u2_R12_reg[22]/NET0131  & ~n7446 ;
  assign n7448 = ~\u2_R12_reg[22]/NET0131  & n7446 ;
  assign n7449 = ~n7447 & ~n7448 ;
  assign n7451 = decrypt_pad & ~\u2_uk_K_r12_reg[35]/NET0131  ;
  assign n7452 = ~decrypt_pad & ~\u2_uk_K_r12_reg[45]/NET0131  ;
  assign n7453 = ~n7451 & ~n7452 ;
  assign n7454 = \u2_R12_reg[20]/NET0131  & ~n7453 ;
  assign n7455 = ~\u2_R12_reg[20]/NET0131  & n7453 ;
  assign n7456 = ~n7454 & ~n7455 ;
  assign n7470 = decrypt_pad & ~\u2_uk_K_r12_reg[51]/NET0131  ;
  assign n7471 = ~decrypt_pad & ~\u2_uk_K_r12_reg[2]/NET0131  ;
  assign n7472 = ~n7470 & ~n7471 ;
  assign n7473 = \u2_R12_reg[25]/NET0131  & ~n7472 ;
  assign n7474 = ~\u2_R12_reg[25]/NET0131  & n7472 ;
  assign n7475 = ~n7473 & ~n7474 ;
  assign n7476 = n7456 & ~n7475 ;
  assign n7458 = decrypt_pad & ~\u2_uk_K_r12_reg[50]/NET0131  ;
  assign n7459 = ~decrypt_pad & ~\u2_uk_K_r12_reg[1]/NET0131  ;
  assign n7460 = ~n7458 & ~n7459 ;
  assign n7461 = \u2_R12_reg[21]/NET0131  & ~n7460 ;
  assign n7462 = ~\u2_R12_reg[21]/NET0131  & n7460 ;
  assign n7463 = ~n7461 & ~n7462 ;
  assign n7485 = ~n7456 & ~n7463 ;
  assign n7513 = ~n7476 & ~n7485 ;
  assign n7514 = n7449 & n7513 ;
  assign n7515 = n7463 & n7475 ;
  assign n7516 = ~n7456 & n7515 ;
  assign n7482 = n7456 & n7475 ;
  assign n7483 = ~n7463 & n7482 ;
  assign n7517 = ~n7449 & ~n7483 ;
  assign n7518 = ~n7516 & n7517 ;
  assign n7519 = ~n7514 & ~n7518 ;
  assign n7520 = ~n7443 & ~n7519 ;
  assign n7432 = decrypt_pad & ~\u2_uk_K_r12_reg[1]/NET0131  ;
  assign n7433 = ~decrypt_pad & ~\u2_uk_K_r12_reg[7]/P0001  ;
  assign n7434 = ~n7432 & ~n7433 ;
  assign n7435 = \u2_R12_reg[24]/NET0131  & ~n7434 ;
  assign n7436 = ~\u2_R12_reg[24]/NET0131  & n7434 ;
  assign n7437 = ~n7435 & ~n7436 ;
  assign n7464 = n7449 & ~n7456 ;
  assign n7465 = n7463 & n7464 ;
  assign n7510 = n7443 & ~n7465 ;
  assign n7507 = ~n7449 & ~n7463 ;
  assign n7508 = n7476 & n7507 ;
  assign n7509 = n7463 & n7482 ;
  assign n7511 = ~n7508 & ~n7509 ;
  assign n7512 = n7510 & n7511 ;
  assign n7521 = n7437 & ~n7512 ;
  assign n7522 = ~n7520 & n7521 ;
  assign n7466 = ~n7449 & n7463 ;
  assign n7488 = n7466 & ~n7475 ;
  assign n7489 = n7456 & n7488 ;
  assign n7484 = n7449 & n7483 ;
  assign n7486 = n7475 & n7485 ;
  assign n7487 = n7443 & n7486 ;
  assign n7492 = ~n7484 & ~n7487 ;
  assign n7493 = ~n7489 & n7492 ;
  assign n7467 = n7456 & n7466 ;
  assign n7468 = ~n7465 & ~n7467 ;
  assign n7469 = ~n7443 & ~n7468 ;
  assign n7479 = n7456 & ~n7463 ;
  assign n7480 = n7443 & n7449 ;
  assign n7481 = n7479 & n7480 ;
  assign n7450 = n7443 & ~n7449 ;
  assign n7457 = n7450 & ~n7456 ;
  assign n7477 = ~n7443 & ~n7449 ;
  assign n7478 = n7476 & n7477 ;
  assign n7490 = ~n7457 & ~n7478 ;
  assign n7491 = ~n7481 & n7490 ;
  assign n7494 = ~n7469 & n7491 ;
  assign n7495 = n7493 & n7494 ;
  assign n7496 = ~n7437 & ~n7495 ;
  assign n7501 = n7463 & n7476 ;
  assign n7502 = ~n7443 & n7501 ;
  assign n7503 = ~n7487 & ~n7502 ;
  assign n7504 = ~n7449 & ~n7503 ;
  assign n7497 = n7449 & n7482 ;
  assign n7498 = ~n7456 & n7488 ;
  assign n7499 = ~n7497 & ~n7498 ;
  assign n7500 = n7443 & ~n7499 ;
  assign n7505 = ~n7475 & n7485 ;
  assign n7506 = n7477 & n7505 ;
  assign n7523 = ~n7500 & ~n7506 ;
  assign n7524 = ~n7504 & n7523 ;
  assign n7525 = ~n7496 & n7524 ;
  assign n7526 = ~n7522 & n7525 ;
  assign n7527 = \u2_L12_reg[11]/NET0131  & ~n7526 ;
  assign n7528 = ~\u2_L12_reg[11]/NET0131  & n7526 ;
  assign n7529 = ~n7527 & ~n7528 ;
  assign n7530 = decrypt_pad & ~\u2_uk_K_r12_reg[8]/NET0131  ;
  assign n7531 = ~decrypt_pad & ~\u2_uk_K_r12_reg[14]/NET0131  ;
  assign n7532 = ~n7530 & ~n7531 ;
  assign n7533 = \u2_R12_reg[28]/NET0131  & ~n7532 ;
  assign n7534 = ~\u2_R12_reg[28]/NET0131  & n7532 ;
  assign n7535 = ~n7533 & ~n7534 ;
  assign n7536 = decrypt_pad & ~\u2_uk_K_r12_reg[21]/NET0131  ;
  assign n7537 = ~decrypt_pad & ~\u2_uk_K_r12_reg[31]/NET0131  ;
  assign n7538 = ~n7536 & ~n7537 ;
  assign n7539 = \u2_R12_reg[27]/NET0131  & ~n7538 ;
  assign n7540 = ~\u2_R12_reg[27]/NET0131  & n7538 ;
  assign n7541 = ~n7539 & ~n7540 ;
  assign n7549 = decrypt_pad & ~\u2_uk_K_r12_reg[43]/NET0131  ;
  assign n7550 = ~decrypt_pad & ~\u2_uk_K_r12_reg[49]/NET0131  ;
  assign n7551 = ~n7549 & ~n7550 ;
  assign n7552 = \u2_R12_reg[26]/NET0131  & ~n7551 ;
  assign n7553 = ~\u2_R12_reg[26]/NET0131  & n7551 ;
  assign n7554 = ~n7552 & ~n7553 ;
  assign n7562 = decrypt_pad & ~\u2_uk_K_r12_reg[23]/NET0131  ;
  assign n7563 = ~decrypt_pad & ~\u2_uk_K_r12_reg[29]/NET0131  ;
  assign n7564 = ~n7562 & ~n7563 ;
  assign n7565 = \u2_R12_reg[24]/NET0131  & ~n7564 ;
  assign n7566 = ~\u2_R12_reg[24]/NET0131  & n7564 ;
  assign n7567 = ~n7565 & ~n7566 ;
  assign n7542 = decrypt_pad & ~\u2_uk_K_r12_reg[0]/NET0131  ;
  assign n7543 = ~decrypt_pad & ~\u2_uk_K_r12_reg[37]/NET0131  ;
  assign n7544 = ~n7542 & ~n7543 ;
  assign n7545 = \u2_R12_reg[29]/NET0131  & ~n7544 ;
  assign n7546 = ~\u2_R12_reg[29]/NET0131  & n7544 ;
  assign n7547 = ~n7545 & ~n7546 ;
  assign n7555 = decrypt_pad & ~\u2_uk_K_r12_reg[31]/NET0131  ;
  assign n7556 = ~decrypt_pad & ~\u2_uk_K_r12_reg[9]/NET0131  ;
  assign n7557 = ~n7555 & ~n7556 ;
  assign n7558 = \u2_R12_reg[25]/NET0131  & ~n7557 ;
  assign n7559 = ~\u2_R12_reg[25]/NET0131  & n7557 ;
  assign n7560 = ~n7558 & ~n7559 ;
  assign n7572 = ~n7547 & ~n7560 ;
  assign n7573 = ~n7567 & n7572 ;
  assign n7592 = n7554 & n7573 ;
  assign n7588 = n7554 & n7567 ;
  assign n7593 = n7547 & n7588 ;
  assign n7594 = ~n7547 & n7567 ;
  assign n7595 = n7560 & n7594 ;
  assign n7596 = ~n7593 & ~n7595 ;
  assign n7597 = ~n7592 & n7596 ;
  assign n7598 = ~n7541 & ~n7597 ;
  assign n7548 = ~n7541 & n7547 ;
  assign n7561 = ~n7554 & ~n7560 ;
  assign n7568 = n7561 & n7567 ;
  assign n7602 = ~n7548 & n7568 ;
  assign n7587 = ~n7554 & ~n7567 ;
  assign n7599 = n7547 & n7560 ;
  assign n7600 = ~n7548 & ~n7599 ;
  assign n7601 = n7587 & ~n7600 ;
  assign n7603 = n7588 & n7599 ;
  assign n7604 = ~n7601 & ~n7603 ;
  assign n7605 = ~n7602 & n7604 ;
  assign n7606 = ~n7598 & n7605 ;
  assign n7607 = ~n7535 & ~n7606 ;
  assign n7576 = n7554 & ~n7560 ;
  assign n7578 = ~n7554 & n7560 ;
  assign n7579 = n7547 & n7578 ;
  assign n7580 = ~n7576 & ~n7579 ;
  assign n7581 = n7541 & n7567 ;
  assign n7582 = ~n7580 & n7581 ;
  assign n7569 = n7560 & ~n7567 ;
  assign n7570 = ~n7568 & ~n7569 ;
  assign n7571 = n7548 & ~n7570 ;
  assign n7574 = ~n7554 & n7573 ;
  assign n7575 = n7547 & ~n7567 ;
  assign n7577 = n7575 & n7576 ;
  assign n7583 = ~n7574 & ~n7577 ;
  assign n7584 = ~n7571 & n7583 ;
  assign n7585 = ~n7582 & n7584 ;
  assign n7586 = n7535 & ~n7585 ;
  assign n7589 = ~n7587 & ~n7588 ;
  assign n7590 = ~n7541 & n7560 ;
  assign n7591 = ~n7589 & n7590 ;
  assign n7608 = ~n7547 & n7554 ;
  assign n7609 = n7569 & n7608 ;
  assign n7612 = ~n7577 & ~n7609 ;
  assign n7610 = n7567 & n7572 ;
  assign n7611 = ~n7554 & n7572 ;
  assign n7613 = ~n7610 & ~n7611 ;
  assign n7614 = n7612 & n7613 ;
  assign n7615 = n7541 & ~n7614 ;
  assign n7616 = ~n7591 & ~n7615 ;
  assign n7617 = ~n7586 & n7616 ;
  assign n7618 = ~n7607 & n7617 ;
  assign n7619 = ~\u2_L12_reg[22]/NET0131  & ~n7618 ;
  assign n7620 = \u2_L12_reg[22]/NET0131  & n7618 ;
  assign n7621 = ~n7619 & ~n7620 ;
  assign n7649 = decrypt_pad & ~\u2_uk_K_r12_reg[20]/NET0131  ;
  assign n7650 = ~decrypt_pad & ~\u2_uk_K_r12_reg[53]/NET0131  ;
  assign n7651 = ~n7649 & ~n7650 ;
  assign n7652 = \u2_R12_reg[14]/NET0131  & ~n7651 ;
  assign n7653 = ~\u2_R12_reg[14]/NET0131  & n7651 ;
  assign n7654 = ~n7652 & ~n7653 ;
  assign n7622 = decrypt_pad & ~\u2_uk_K_r12_reg[19]/NET0131  ;
  assign n7623 = ~decrypt_pad & ~\u2_uk_K_r12_reg[27]/NET0131  ;
  assign n7624 = ~n7622 & ~n7623 ;
  assign n7625 = \u2_R12_reg[13]/NET0131  & ~n7624 ;
  assign n7626 = ~\u2_R12_reg[13]/NET0131  & n7624 ;
  assign n7627 = ~n7625 & ~n7626 ;
  assign n7635 = decrypt_pad & ~\u2_uk_K_r12_reg[25]/NET0131  ;
  assign n7636 = ~decrypt_pad & ~\u2_uk_K_r12_reg[33]/NET0131  ;
  assign n7637 = ~n7635 & ~n7636 ;
  assign n7638 = \u2_R12_reg[12]/NET0131  & ~n7637 ;
  assign n7639 = ~\u2_R12_reg[12]/NET0131  & n7637 ;
  assign n7640 = ~n7638 & ~n7639 ;
  assign n7641 = decrypt_pad & ~\u2_uk_K_r12_reg[41]/NET0131  ;
  assign n7642 = ~decrypt_pad & ~\u2_uk_K_r12_reg[17]/NET0131  ;
  assign n7643 = ~n7641 & ~n7642 ;
  assign n7644 = \u2_R12_reg[17]/NET0131  & ~n7643 ;
  assign n7645 = ~\u2_R12_reg[17]/NET0131  & n7643 ;
  assign n7646 = ~n7644 & ~n7645 ;
  assign n7678 = n7640 & n7646 ;
  assign n7679 = n7627 & n7678 ;
  assign n7628 = decrypt_pad & ~\u2_uk_K_r12_reg[53]/NET0131  ;
  assign n7629 = ~decrypt_pad & ~\u2_uk_K_r12_reg[4]/NET0131  ;
  assign n7630 = ~n7628 & ~n7629 ;
  assign n7631 = \u2_R12_reg[15]/NET0131  & ~n7630 ;
  assign n7632 = ~\u2_R12_reg[15]/NET0131  & n7630 ;
  assign n7633 = ~n7631 & ~n7632 ;
  assign n7660 = ~n7627 & ~n7646 ;
  assign n7680 = ~n7640 & n7660 ;
  assign n7681 = ~n7633 & n7680 ;
  assign n7682 = ~n7679 & ~n7681 ;
  assign n7683 = n7654 & ~n7682 ;
  assign n7634 = n7627 & n7633 ;
  assign n7647 = n7640 & ~n7646 ;
  assign n7648 = n7634 & n7647 ;
  assign n7656 = ~n7640 & n7646 ;
  assign n7657 = n7627 & n7656 ;
  assign n7658 = ~n7654 & n7657 ;
  assign n7686 = ~n7648 & ~n7658 ;
  assign n7684 = n7633 & n7656 ;
  assign n7685 = ~n7627 & n7684 ;
  assign n7667 = ~n7633 & ~n7654 ;
  assign n7668 = n7627 & ~n7640 ;
  assign n7669 = ~n7627 & n7640 ;
  assign n7670 = ~n7668 & ~n7669 ;
  assign n7671 = n7667 & ~n7670 ;
  assign n7672 = decrypt_pad & ~\u2_uk_K_r12_reg[4]/NET0131  ;
  assign n7673 = ~decrypt_pad & ~\u2_uk_K_r12_reg[12]/NET0131  ;
  assign n7674 = ~n7672 & ~n7673 ;
  assign n7675 = \u2_R12_reg[16]/NET0131  & ~n7674 ;
  assign n7676 = ~\u2_R12_reg[16]/NET0131  & n7674 ;
  assign n7677 = ~n7675 & ~n7676 ;
  assign n7687 = ~n7671 & n7677 ;
  assign n7688 = ~n7685 & n7687 ;
  assign n7689 = n7686 & n7688 ;
  assign n7690 = ~n7683 & n7689 ;
  assign n7702 = ~n7627 & n7678 ;
  assign n7703 = ~n7654 & n7702 ;
  assign n7692 = n7633 & n7680 ;
  assign n7693 = n7634 & n7654 ;
  assign n7694 = ~n7640 & n7693 ;
  assign n7705 = ~n7692 & ~n7694 ;
  assign n7706 = ~n7703 & n7705 ;
  assign n7661 = ~n7640 & ~n7654 ;
  assign n7662 = n7660 & n7661 ;
  assign n7699 = ~n7646 & n7668 ;
  assign n7700 = n7654 & n7699 ;
  assign n7701 = ~n7662 & ~n7700 ;
  assign n7695 = n7647 & n7654 ;
  assign n7696 = ~n7627 & n7646 ;
  assign n7697 = ~n7695 & ~n7696 ;
  assign n7698 = ~n7633 & ~n7697 ;
  assign n7691 = n7633 & n7679 ;
  assign n7704 = ~n7677 & ~n7691 ;
  assign n7707 = ~n7698 & n7704 ;
  assign n7708 = n7701 & n7707 ;
  assign n7709 = n7706 & n7708 ;
  assign n7710 = ~n7690 & ~n7709 ;
  assign n7663 = ~n7627 & n7654 ;
  assign n7664 = n7647 & n7663 ;
  assign n7665 = ~n7662 & ~n7664 ;
  assign n7666 = n7633 & ~n7665 ;
  assign n7655 = n7648 & ~n7654 ;
  assign n7659 = ~n7633 & n7658 ;
  assign n7711 = ~n7655 & ~n7659 ;
  assign n7712 = ~n7666 & n7711 ;
  assign n7713 = ~n7710 & n7712 ;
  assign n7714 = ~\u2_L12_reg[20]/NET0131  & ~n7713 ;
  assign n7715 = \u2_L12_reg[20]/NET0131  & n7713 ;
  assign n7716 = ~n7714 & ~n7715 ;
  assign n7721 = n7361 & n7367 ;
  assign n7722 = n7383 & ~n7721 ;
  assign n7717 = ~n7367 & ~n7393 ;
  assign n7718 = ~n7421 & ~n7717 ;
  assign n7719 = n7341 & ~n7718 ;
  assign n7720 = n7353 & n7385 ;
  assign n7723 = ~n7341 & ~n7410 ;
  assign n7724 = ~n7717 & n7723 ;
  assign n7725 = ~n7720 & ~n7724 ;
  assign n7726 = ~n7719 & n7725 ;
  assign n7727 = n7722 & n7726 ;
  assign n7732 = ~n7347 & n7368 ;
  assign n7733 = ~n7398 & ~n7732 ;
  assign n7734 = n7360 & ~n7733 ;
  assign n7735 = n7360 & n7386 ;
  assign n7736 = ~n7372 & ~n7735 ;
  assign n7737 = ~n7734 & n7736 ;
  assign n7738 = n7341 & ~n7737 ;
  assign n7728 = ~n7386 & ~n7397 ;
  assign n7729 = ~n7360 & ~n7728 ;
  assign n7730 = ~n7418 & ~n7729 ;
  assign n7731 = ~n7341 & ~n7730 ;
  assign n7739 = ~n7370 & ~n7383 ;
  assign n7740 = ~n7413 & n7739 ;
  assign n7741 = ~n7731 & n7740 ;
  assign n7742 = ~n7738 & n7741 ;
  assign n7743 = ~n7727 & ~n7742 ;
  assign n7744 = ~\u2_L12_reg[17]/NET0131  & n7743 ;
  assign n7745 = \u2_L12_reg[17]/NET0131  & ~n7743 ;
  assign n7746 = ~n7744 & ~n7745 ;
  assign n7770 = ~n7463 & n7476 ;
  assign n7771 = ~n7509 & ~n7770 ;
  assign n7772 = ~n7465 & ~n7507 ;
  assign n7773 = ~n7475 & ~n7772 ;
  assign n7774 = n7771 & ~n7773 ;
  assign n7775 = n7443 & ~n7774 ;
  assign n7747 = n7449 & n7501 ;
  assign n7767 = ~n7449 & n7513 ;
  assign n7768 = ~n7747 & ~n7767 ;
  assign n7769 = ~n7443 & ~n7768 ;
  assign n7776 = n7449 & n7486 ;
  assign n7777 = ~n7769 & ~n7776 ;
  assign n7778 = ~n7775 & n7777 ;
  assign n7779 = ~n7437 & ~n7778 ;
  assign n7748 = ~n7449 & ~n7456 ;
  assign n7749 = n7463 & n7748 ;
  assign n7750 = ~n7516 & ~n7749 ;
  assign n7751 = ~n7747 & n7750 ;
  assign n7752 = n7443 & ~n7751 ;
  assign n7753 = ~n7456 & ~n7475 ;
  assign n7757 = n7449 & n7753 ;
  assign n7758 = n7475 & n7748 ;
  assign n7759 = ~n7757 & ~n7758 ;
  assign n7760 = ~n7463 & ~n7759 ;
  assign n7754 = ~n7466 & n7753 ;
  assign n7755 = ~n7497 & ~n7754 ;
  assign n7756 = ~n7443 & ~n7755 ;
  assign n7761 = ~n7478 & ~n7484 ;
  assign n7762 = ~n7756 & n7761 ;
  assign n7763 = ~n7760 & n7762 ;
  assign n7764 = ~n7752 & n7763 ;
  assign n7765 = n7437 & ~n7764 ;
  assign n7766 = n7450 & n7515 ;
  assign n7780 = ~n7508 & ~n7766 ;
  assign n7781 = ~n7765 & n7780 ;
  assign n7782 = ~n7779 & n7781 ;
  assign n7783 = \u2_L12_reg[29]/NET0131  & ~n7782 ;
  assign n7784 = ~\u2_L12_reg[29]/NET0131  & n7782 ;
  assign n7785 = ~n7783 & ~n7784 ;
  assign n7804 = decrypt_pad & ~\u2_uk_K_r12_reg[18]/NET0131  ;
  assign n7805 = ~decrypt_pad & ~\u2_uk_K_r12_reg[26]/NET0131  ;
  assign n7806 = ~n7804 & ~n7805 ;
  assign n7807 = \u2_R12_reg[6]/NET0131  & ~n7806 ;
  assign n7808 = ~\u2_R12_reg[6]/NET0131  & n7806 ;
  assign n7809 = ~n7807 & ~n7808 ;
  assign n7792 = decrypt_pad & ~\u2_uk_K_r12_reg[40]/NET0131  ;
  assign n7793 = ~decrypt_pad & ~\u2_uk_K_r12_reg[48]/NET0131  ;
  assign n7794 = ~n7792 & ~n7793 ;
  assign n7795 = \u2_R12_reg[9]/NET0131  & ~n7794 ;
  assign n7796 = ~\u2_R12_reg[9]/NET0131  & n7794 ;
  assign n7797 = ~n7795 & ~n7796 ;
  assign n7798 = decrypt_pad & ~\u2_uk_K_r12_reg[27]/NET0131  ;
  assign n7799 = ~decrypt_pad & ~\u2_uk_K_r12_reg[3]/NET0131  ;
  assign n7800 = ~n7798 & ~n7799 ;
  assign n7801 = \u2_R12_reg[5]/NET0131  & ~n7800 ;
  assign n7802 = ~\u2_R12_reg[5]/NET0131  & n7800 ;
  assign n7803 = ~n7801 & ~n7802 ;
  assign n7823 = ~n7797 & n7803 ;
  assign n7811 = decrypt_pad & ~\u2_uk_K_r12_reg[48]/NET0131  ;
  assign n7812 = ~decrypt_pad & ~\u2_uk_K_r12_reg[24]/NET0131  ;
  assign n7813 = ~n7811 & ~n7812 ;
  assign n7814 = \u2_R12_reg[4]/NET0131  & ~n7813 ;
  assign n7815 = ~\u2_R12_reg[4]/NET0131  & n7813 ;
  assign n7816 = ~n7814 & ~n7815 ;
  assign n7824 = n7797 & ~n7803 ;
  assign n7825 = ~n7816 & n7824 ;
  assign n7826 = ~n7823 & ~n7825 ;
  assign n7827 = ~n7809 & ~n7826 ;
  assign n7786 = decrypt_pad & ~\u2_uk_K_r12_reg[12]/NET0131  ;
  assign n7787 = ~decrypt_pad & ~\u2_uk_K_r12_reg[20]/NET0131  ;
  assign n7788 = ~n7786 & ~n7787 ;
  assign n7789 = \u2_R12_reg[7]/NET0131  & ~n7788 ;
  assign n7790 = ~\u2_R12_reg[7]/NET0131  & n7788 ;
  assign n7791 = ~n7789 & ~n7790 ;
  assign n7836 = n7809 & n7816 ;
  assign n7837 = n7791 & n7836 ;
  assign n7838 = n7824 & n7837 ;
  assign n7842 = decrypt_pad & ~\u2_uk_K_r12_reg[3]/NET0131  ;
  assign n7843 = ~decrypt_pad & ~\u2_uk_K_r12_reg[11]/NET0131  ;
  assign n7844 = ~n7842 & ~n7843 ;
  assign n7845 = \u2_R12_reg[8]/NET0131  & ~n7844 ;
  assign n7846 = ~\u2_R12_reg[8]/NET0131  & n7844 ;
  assign n7847 = ~n7845 & ~n7846 ;
  assign n7848 = ~n7838 & ~n7847 ;
  assign n7849 = ~n7827 & n7848 ;
  assign n7830 = n7797 & ~n7816 ;
  assign n7831 = n7803 & n7830 ;
  assign n7832 = n7809 & ~n7831 ;
  assign n7828 = ~n7791 & ~n7803 ;
  assign n7829 = ~n7809 & ~n7828 ;
  assign n7833 = ~n7797 & ~n7809 ;
  assign n7834 = ~n7829 & ~n7833 ;
  assign n7835 = ~n7832 & n7834 ;
  assign n7839 = ~n7824 & n7836 ;
  assign n7840 = ~n7825 & ~n7839 ;
  assign n7841 = ~n7791 & ~n7840 ;
  assign n7850 = ~n7835 & ~n7841 ;
  assign n7851 = n7849 & n7850 ;
  assign n7859 = ~n7809 & n7816 ;
  assign n7860 = n7797 & n7859 ;
  assign n7861 = n7809 & ~n7816 ;
  assign n7862 = n7791 & ~n7861 ;
  assign n7863 = ~n7860 & ~n7862 ;
  assign n7864 = n7803 & ~n7863 ;
  assign n7810 = ~n7803 & n7809 ;
  assign n7855 = n7797 & ~n7810 ;
  assign n7853 = ~n7791 & n7809 ;
  assign n7854 = ~n7828 & ~n7853 ;
  assign n7852 = ~n7797 & n7816 ;
  assign n7856 = ~n7830 & ~n7852 ;
  assign n7857 = ~n7854 & n7856 ;
  assign n7858 = ~n7855 & n7857 ;
  assign n7865 = ~n7803 & n7833 ;
  assign n7866 = n7816 & n7865 ;
  assign n7867 = n7847 & ~n7866 ;
  assign n7868 = ~n7858 & n7867 ;
  assign n7869 = ~n7864 & n7868 ;
  assign n7870 = ~n7851 & ~n7869 ;
  assign n7817 = n7810 & ~n7816 ;
  assign n7818 = ~n7797 & n7817 ;
  assign n7819 = n7803 & n7816 ;
  assign n7820 = ~n7809 & n7819 ;
  assign n7821 = ~n7818 & ~n7820 ;
  assign n7822 = n7791 & ~n7821 ;
  assign n7871 = ~n7810 & ~n7816 ;
  assign n7872 = n7797 & ~n7854 ;
  assign n7873 = n7871 & n7872 ;
  assign n7874 = ~n7822 & ~n7873 ;
  assign n7875 = ~n7870 & n7874 ;
  assign n7876 = \u2_L12_reg[2]/NET0131  & n7875 ;
  assign n7877 = ~\u2_L12_reg[2]/NET0131  & ~n7875 ;
  assign n7878 = ~n7876 & ~n7877 ;
  assign n7932 = decrypt_pad & ~\u2_uk_K_r12_reg[28]/NET0131  ;
  assign n7933 = ~decrypt_pad & ~\u2_uk_K_r12_reg[38]/NET0131  ;
  assign n7934 = ~n7932 & ~n7933 ;
  assign n7935 = \u2_R12_reg[32]/NET0131  & ~n7934 ;
  assign n7936 = ~\u2_R12_reg[32]/NET0131  & n7934 ;
  assign n7937 = ~n7935 & ~n7936 ;
  assign n7899 = decrypt_pad & ~\u2_uk_K_r12_reg[22]/NET0131  ;
  assign n7900 = ~decrypt_pad & ~\u2_uk_K_r12_reg[28]/NET0131  ;
  assign n7901 = ~n7899 & ~n7900 ;
  assign n7902 = \u2_R12_reg[31]/P0001  & ~n7901 ;
  assign n7903 = ~\u2_R12_reg[31]/P0001  & n7901 ;
  assign n7904 = ~n7902 & ~n7903 ;
  assign n7879 = decrypt_pad & ~\u2_uk_K_r12_reg[38]/NET0131  ;
  assign n7880 = ~decrypt_pad & ~\u2_uk_K_r12_reg[16]/NET0131  ;
  assign n7881 = ~n7879 & ~n7880 ;
  assign n7882 = \u2_R12_reg[30]/NET0131  & ~n7881 ;
  assign n7883 = ~\u2_R12_reg[30]/NET0131  & n7881 ;
  assign n7884 = ~n7882 & ~n7883 ;
  assign n7885 = decrypt_pad & ~\u2_uk_K_r12_reg[9]/NET0131  ;
  assign n7886 = ~decrypt_pad & ~\u2_uk_K_r12_reg[15]/NET0131  ;
  assign n7887 = ~n7885 & ~n7886 ;
  assign n7888 = \u2_R12_reg[29]/NET0131  & ~n7887 ;
  assign n7889 = ~\u2_R12_reg[29]/NET0131  & n7887 ;
  assign n7890 = ~n7888 & ~n7889 ;
  assign n7907 = decrypt_pad & ~\u2_uk_K_r12_reg[37]/NET0131  ;
  assign n7908 = ~decrypt_pad & ~\u2_uk_K_r12_reg[43]/NET0131  ;
  assign n7909 = ~n7907 & ~n7908 ;
  assign n7910 = \u2_R12_reg[28]/NET0131  & ~n7909 ;
  assign n7911 = ~\u2_R12_reg[28]/NET0131  & n7909 ;
  assign n7912 = ~n7910 & ~n7911 ;
  assign n7914 = ~n7890 & n7912 ;
  assign n7892 = decrypt_pad & ~\u2_uk_K_r12_reg[49]/NET0131  ;
  assign n7893 = ~decrypt_pad & ~\u2_uk_K_r12_reg[0]/NET0131  ;
  assign n7894 = ~n7892 & ~n7893 ;
  assign n7895 = \u2_R12_reg[1]/NET0131  & ~n7894 ;
  assign n7896 = ~\u2_R12_reg[1]/NET0131  & n7894 ;
  assign n7897 = ~n7895 & ~n7896 ;
  assign n7956 = n7897 & n7912 ;
  assign n7957 = ~n7914 & ~n7956 ;
  assign n7958 = ~n7884 & ~n7957 ;
  assign n7942 = ~n7897 & ~n7912 ;
  assign n7955 = n7890 & n7942 ;
  assign n7891 = n7884 & n7890 ;
  assign n7959 = n7891 & ~n7897 ;
  assign n7960 = ~n7955 & ~n7959 ;
  assign n7961 = ~n7958 & n7960 ;
  assign n7962 = n7904 & ~n7961 ;
  assign n7944 = ~n7884 & ~n7890 ;
  assign n7963 = ~n7912 & n7944 ;
  assign n7964 = ~n7904 & n7963 ;
  assign n7965 = n7891 & ~n7912 ;
  assign n7966 = n7897 & n7965 ;
  assign n7967 = ~n7964 & ~n7966 ;
  assign n7968 = ~n7962 & n7967 ;
  assign n7969 = n7937 & ~n7968 ;
  assign n7915 = n7884 & n7914 ;
  assign n7916 = ~n7897 & n7915 ;
  assign n7917 = n7897 & ~n7912 ;
  assign n7918 = ~n7890 & n7917 ;
  assign n7919 = ~n7916 & ~n7918 ;
  assign n7920 = n7904 & ~n7919 ;
  assign n7898 = n7891 & n7897 ;
  assign n7905 = ~n7884 & ~n7904 ;
  assign n7906 = ~n7898 & ~n7905 ;
  assign n7913 = ~n7906 & n7912 ;
  assign n7923 = ~n7897 & n7912 ;
  assign n7924 = ~n7904 & ~n7923 ;
  assign n7921 = ~n7884 & ~n7897 ;
  assign n7922 = ~n7890 & n7897 ;
  assign n7925 = ~n7921 & ~n7922 ;
  assign n7926 = n7924 & n7925 ;
  assign n7927 = n7890 & n7923 ;
  assign n7928 = ~n7884 & n7927 ;
  assign n7929 = ~n7926 & ~n7928 ;
  assign n7930 = ~n7913 & n7929 ;
  assign n7931 = ~n7920 & n7930 ;
  assign n7938 = ~n7931 & ~n7937 ;
  assign n7943 = n7891 & n7942 ;
  assign n7945 = n7897 & n7944 ;
  assign n7946 = n7912 & n7945 ;
  assign n7947 = ~n7943 & ~n7946 ;
  assign n7948 = n7884 & n7918 ;
  assign n7949 = ~n7890 & n7942 ;
  assign n7950 = ~n7884 & n7949 ;
  assign n7951 = ~n7948 & ~n7950 ;
  assign n7952 = n7947 & n7951 ;
  assign n7953 = n7904 & ~n7952 ;
  assign n7939 = n7884 & ~n7904 ;
  assign n7940 = n7914 & n7937 ;
  assign n7941 = n7939 & n7940 ;
  assign n7954 = ~n7904 & n7928 ;
  assign n7970 = ~n7941 & ~n7954 ;
  assign n7971 = ~n7953 & n7970 ;
  assign n7972 = ~n7938 & n7971 ;
  assign n7973 = ~n7969 & n7972 ;
  assign n7974 = \u2_L12_reg[5]/NET0131  & ~n7973 ;
  assign n7975 = ~\u2_L12_reg[5]/NET0131  & n7973 ;
  assign n7976 = ~n7974 & ~n7975 ;
  assign n7981 = ~n7501 & ~n7758 ;
  assign n7982 = ~n7484 & n7981 ;
  assign n7983 = n7443 & ~n7982 ;
  assign n7977 = n7463 & n7753 ;
  assign n7978 = ~n7776 & ~n7977 ;
  assign n7979 = ~n7443 & ~n7978 ;
  assign n7980 = n7477 & n7482 ;
  assign n7984 = ~n7508 & ~n7980 ;
  assign n7985 = ~n7979 & n7984 ;
  assign n7986 = ~n7983 & n7985 ;
  assign n7987 = ~n7437 & ~n7986 ;
  assign n7995 = ~n7488 & ~n7748 ;
  assign n7996 = ~n7443 & ~n7995 ;
  assign n7997 = n7449 & n7515 ;
  assign n7998 = n7450 & n7482 ;
  assign n7999 = ~n7997 & ~n7998 ;
  assign n8000 = ~n7498 & n7999 ;
  assign n8001 = ~n7996 & n8000 ;
  assign n8002 = n7437 & ~n8001 ;
  assign n7988 = ~n7505 & ~n7516 ;
  assign n7989 = ~n7501 & n7988 ;
  assign n7990 = n7480 & ~n7989 ;
  assign n7991 = n7449 & n7771 ;
  assign n7992 = ~n7449 & ~n7753 ;
  assign n7993 = ~n7443 & ~n7992 ;
  assign n7994 = ~n7991 & n7993 ;
  assign n8003 = ~n7990 & ~n7994 ;
  assign n8004 = ~n8002 & n8003 ;
  assign n8005 = ~n7987 & n8004 ;
  assign n8006 = ~\u2_L12_reg[4]/NET0131  & ~n8005 ;
  assign n8007 = \u2_L12_reg[4]/NET0131  & n8005 ;
  assign n8008 = ~n8006 & ~n8007 ;
  assign n8027 = n7627 & ~n7654 ;
  assign n8028 = n7647 & ~n8027 ;
  assign n8029 = ~n7658 & ~n8028 ;
  assign n8030 = ~n7633 & ~n8029 ;
  assign n8022 = n7654 & n7679 ;
  assign n8023 = n7656 & n7663 ;
  assign n8024 = ~n8022 & ~n8023 ;
  assign n8025 = ~n7699 & ~n7703 ;
  assign n8026 = n7633 & ~n8025 ;
  assign n8031 = n8024 & ~n8026 ;
  assign n8032 = ~n8030 & n8031 ;
  assign n8033 = n7677 & ~n8032 ;
  assign n8009 = n7640 & ~n7654 ;
  assign n8010 = n7627 & n8009 ;
  assign n8011 = n7667 & n7678 ;
  assign n8016 = ~n8010 & ~n8011 ;
  assign n8017 = ~n7681 & n8016 ;
  assign n8012 = n7646 & ~n7654 ;
  assign n8013 = n7633 & n7669 ;
  assign n8014 = ~n8012 & n8013 ;
  assign n8015 = ~n7654 & n7684 ;
  assign n8018 = ~n8014 & ~n8015 ;
  assign n8019 = n8017 & n8018 ;
  assign n8020 = n7701 & n8019 ;
  assign n8021 = ~n7677 & ~n8020 ;
  assign n8034 = ~n7662 & n8024 ;
  assign n8035 = ~n7633 & ~n8034 ;
  assign n8036 = ~n7655 & ~n7694 ;
  assign n8037 = ~n8035 & n8036 ;
  assign n8038 = ~n8021 & n8037 ;
  assign n8039 = ~n8033 & n8038 ;
  assign n8040 = ~\u2_L12_reg[10]/NET0131  & ~n8039 ;
  assign n8041 = \u2_L12_reg[10]/NET0131  & n8039 ;
  assign n8042 = ~n8040 & ~n8041 ;
  assign n8051 = ~n7567 & ~n7578 ;
  assign n8052 = ~n7541 & ~n7560 ;
  assign n8053 = n7547 & ~n8052 ;
  assign n8054 = n8051 & n8053 ;
  assign n8043 = ~n7575 & ~n7594 ;
  assign n8044 = n7576 & n8043 ;
  assign n8055 = ~n7535 & ~n8044 ;
  assign n8056 = ~n8054 & n8055 ;
  assign n8045 = ~n7572 & ~n7599 ;
  assign n8046 = ~n7588 & n8045 ;
  assign n8047 = ~n7541 & ~n8046 ;
  assign n8048 = ~n7547 & n7569 ;
  assign n8049 = ~n7610 & ~n8048 ;
  assign n8050 = ~n7554 & ~n8049 ;
  assign n8057 = ~n8047 & ~n8050 ;
  assign n8058 = n8056 & n8057 ;
  assign n8060 = n7560 & n7567 ;
  assign n8061 = ~n7574 & ~n8060 ;
  assign n8062 = n7541 & ~n8061 ;
  assign n8059 = n7554 & ~n8049 ;
  assign n8064 = n7554 & ~n8052 ;
  assign n8065 = ~n7561 & n7575 ;
  assign n8066 = ~n8064 & n8065 ;
  assign n8063 = n7547 & n7568 ;
  assign n8067 = n7535 & ~n8063 ;
  assign n8068 = ~n8066 & n8067 ;
  assign n8069 = ~n8059 & n8068 ;
  assign n8070 = ~n8062 & n8069 ;
  assign n8071 = ~n8058 & ~n8070 ;
  assign n8072 = \u2_L12_reg[12]/NET0131  & n8071 ;
  assign n8073 = ~\u2_L12_reg[12]/NET0131  & ~n8071 ;
  assign n8074 = ~n8072 & ~n8073 ;
  assign n8075 = ~n7797 & n7859 ;
  assign n8076 = ~n7823 & ~n8075 ;
  assign n8077 = ~n7819 & ~n8076 ;
  assign n8078 = n7797 & n7817 ;
  assign n8079 = ~n8077 & ~n8078 ;
  assign n8080 = ~n7847 & ~n8079 ;
  assign n8081 = n7823 & n7836 ;
  assign n8082 = n7797 & n7820 ;
  assign n8083 = ~n8081 & ~n8082 ;
  assign n8084 = ~n8080 & n8083 ;
  assign n8085 = ~n7791 & ~n8084 ;
  assign n8086 = ~n7803 & ~n7830 ;
  assign n8087 = ~n7852 & n8086 ;
  assign n8088 = n7803 & n8075 ;
  assign n8089 = ~n8087 & ~n8088 ;
  assign n8090 = n7791 & ~n8089 ;
  assign n8092 = n7829 & n7830 ;
  assign n8091 = ~n7823 & n7837 ;
  assign n8093 = ~n7847 & ~n8091 ;
  assign n8094 = ~n8092 & n8093 ;
  assign n8095 = ~n8090 & n8094 ;
  assign n8096 = ~n7833 & n8086 ;
  assign n8097 = ~n7791 & ~n8096 ;
  assign n8098 = n7797 & n7861 ;
  assign n8099 = n7791 & ~n7865 ;
  assign n8100 = ~n8098 & n8099 ;
  assign n8101 = ~n8097 & ~n8100 ;
  assign n8102 = ~n7816 & n7833 ;
  assign n8103 = n7803 & n8102 ;
  assign n8104 = n7847 & ~n8103 ;
  assign n8105 = ~n7835 & n8104 ;
  assign n8106 = n8083 & n8105 ;
  assign n8107 = ~n8101 & n8106 ;
  assign n8108 = ~n8095 & ~n8107 ;
  assign n8109 = ~n8085 & ~n8108 ;
  assign n8110 = ~\u2_L12_reg[13]/NET0131  & n8109 ;
  assign n8111 = \u2_L12_reg[13]/NET0131  & ~n8109 ;
  assign n8112 = ~n8110 & ~n8111 ;
  assign n8113 = ~n7912 & ~n7921 ;
  assign n8114 = n7890 & ~n8113 ;
  assign n8115 = ~n7918 & ~n8114 ;
  assign n8116 = n7904 & ~n8115 ;
  assign n8117 = n7923 & n7944 ;
  assign n8118 = ~n8116 & ~n8117 ;
  assign n8119 = ~n7937 & ~n8118 ;
  assign n8135 = n7922 & n7939 ;
  assign n8125 = ~n7884 & n7890 ;
  assign n8134 = n7912 & n8125 ;
  assign n8136 = ~n7943 & ~n8134 ;
  assign n8137 = ~n8135 & n8136 ;
  assign n8132 = n7904 & n7949 ;
  assign n8133 = n7897 & n7915 ;
  assign n8138 = ~n8132 & ~n8133 ;
  assign n8139 = n8137 & n8138 ;
  assign n8140 = n7937 & ~n8139 ;
  assign n8120 = ~n7884 & n7937 ;
  assign n8121 = ~n7914 & ~n7943 ;
  assign n8122 = ~n8120 & ~n8121 ;
  assign n8123 = ~n7950 & ~n8122 ;
  assign n8124 = ~n7904 & ~n8123 ;
  assign n8128 = ~n7904 & ~n8125 ;
  assign n8126 = n7904 & n8125 ;
  assign n8127 = n7884 & ~n7890 ;
  assign n8129 = n7917 & ~n8127 ;
  assign n8130 = ~n8126 & n8129 ;
  assign n8131 = ~n8128 & n8130 ;
  assign n8141 = ~n8124 & ~n8131 ;
  assign n8142 = ~n8140 & n8141 ;
  assign n8143 = ~n8119 & n8142 ;
  assign n8144 = ~\u2_L12_reg[15]/NET0131  & ~n8143 ;
  assign n8145 = \u2_L12_reg[15]/NET0131  & n8143 ;
  assign n8146 = ~n8144 & ~n8145 ;
  assign n8147 = decrypt_pad & ~\u2_uk_K_r12_reg[44]/P0001  ;
  assign n8148 = ~decrypt_pad & ~\u2_uk_K_r12_reg[50]/NET0131  ;
  assign n8149 = ~n8147 & ~n8148 ;
  assign n8150 = \u2_R12_reg[20]/NET0131  & ~n8149 ;
  assign n8151 = ~\u2_R12_reg[20]/NET0131  & n8149 ;
  assign n8152 = ~n8150 & ~n8151 ;
  assign n8180 = decrypt_pad & ~\u2_uk_K_r12_reg[29]/NET0131  ;
  assign n8181 = ~decrypt_pad & ~\u2_uk_K_r12_reg[35]/NET0131  ;
  assign n8182 = ~n8180 & ~n8181 ;
  assign n8183 = \u2_R12_reg[19]/NET0131  & ~n8182 ;
  assign n8184 = ~\u2_R12_reg[19]/NET0131  & n8182 ;
  assign n8185 = ~n8183 & ~n8184 ;
  assign n8153 = decrypt_pad & ~\u2_uk_K_r12_reg[52]/NET0131  ;
  assign n8154 = ~decrypt_pad & ~\u2_uk_K_r12_reg[30]/NET0131  ;
  assign n8155 = ~n8153 & ~n8154 ;
  assign n8156 = \u2_R12_reg[17]/NET0131  & ~n8155 ;
  assign n8157 = ~\u2_R12_reg[17]/NET0131  & n8155 ;
  assign n8158 = ~n8156 & ~n8157 ;
  assign n8166 = decrypt_pad & ~\u2_uk_K_r12_reg[2]/NET0131  ;
  assign n8167 = ~decrypt_pad & ~\u2_uk_K_r12_reg[8]/NET0131  ;
  assign n8168 = ~n8166 & ~n8167 ;
  assign n8169 = \u2_R12_reg[16]/NET0131  & ~n8168 ;
  assign n8170 = ~\u2_R12_reg[16]/NET0131  & n8168 ;
  assign n8171 = ~n8169 & ~n8170 ;
  assign n8173 = decrypt_pad & ~\u2_uk_K_r12_reg[14]/NET0131  ;
  assign n8174 = ~decrypt_pad & ~\u2_uk_K_r12_reg[51]/NET0131  ;
  assign n8175 = ~n8173 & ~n8174 ;
  assign n8176 = \u2_R12_reg[21]/NET0131  & ~n8175 ;
  assign n8177 = ~\u2_R12_reg[21]/NET0131  & n8175 ;
  assign n8178 = ~n8176 & ~n8177 ;
  assign n8188 = ~n8171 & n8178 ;
  assign n8189 = ~n8158 & n8188 ;
  assign n8186 = n8158 & ~n8178 ;
  assign n8213 = n8171 & n8186 ;
  assign n8226 = ~n8189 & ~n8213 ;
  assign n8159 = decrypt_pad & ~\u2_uk_K_r12_reg[42]/NET0131  ;
  assign n8160 = ~decrypt_pad & ~\u2_uk_K_r12_reg[52]/NET0131  ;
  assign n8161 = ~n8159 & ~n8160 ;
  assign n8162 = \u2_R12_reg[18]/NET0131  & ~n8161 ;
  assign n8163 = ~\u2_R12_reg[18]/NET0131  & n8161 ;
  assign n8164 = ~n8162 & ~n8163 ;
  assign n8193 = n8171 & n8178 ;
  assign n8224 = ~n8164 & n8193 ;
  assign n8225 = n8164 & n8188 ;
  assign n8227 = ~n8224 & ~n8225 ;
  assign n8228 = n8226 & n8227 ;
  assign n8229 = n8185 & ~n8228 ;
  assign n8215 = ~n8164 & ~n8185 ;
  assign n8200 = ~n8171 & ~n8178 ;
  assign n8201 = ~n8158 & n8200 ;
  assign n8216 = n8158 & n8188 ;
  assign n8217 = ~n8201 & ~n8216 ;
  assign n8218 = n8215 & ~n8217 ;
  assign n8219 = n8158 & ~n8185 ;
  assign n8220 = n8164 & ~n8219 ;
  assign n8165 = n8158 & ~n8164 ;
  assign n8221 = ~n8165 & n8193 ;
  assign n8222 = ~n8220 & n8221 ;
  assign n8214 = ~n8164 & n8213 ;
  assign n8190 = n8171 & ~n8178 ;
  assign n8207 = ~n8158 & n8164 ;
  assign n8223 = n8190 & n8207 ;
  assign n8230 = ~n8214 & ~n8223 ;
  assign n8231 = ~n8222 & n8230 ;
  assign n8232 = ~n8218 & n8231 ;
  assign n8233 = ~n8229 & n8232 ;
  assign n8234 = n8152 & ~n8233 ;
  assign n8194 = n8158 & n8193 ;
  assign n8195 = ~n8164 & n8194 ;
  assign n8191 = ~n8158 & ~n8164 ;
  assign n8192 = n8190 & n8191 ;
  assign n8187 = n8164 & n8186 ;
  assign n8196 = ~n8187 & ~n8189 ;
  assign n8197 = ~n8192 & n8196 ;
  assign n8198 = ~n8195 & n8197 ;
  assign n8199 = ~n8185 & ~n8198 ;
  assign n8202 = n8164 & n8178 ;
  assign n8203 = n8171 & n8202 ;
  assign n8172 = n8165 & ~n8171 ;
  assign n8204 = ~n8172 & ~n8201 ;
  assign n8205 = ~n8203 & n8204 ;
  assign n8206 = n8185 & ~n8205 ;
  assign n8179 = n8172 & ~n8178 ;
  assign n8208 = n8193 & n8207 ;
  assign n8209 = ~n8179 & ~n8208 ;
  assign n8210 = ~n8206 & n8209 ;
  assign n8211 = ~n8199 & n8210 ;
  assign n8212 = ~n8152 & ~n8211 ;
  assign n8235 = ~n8171 & n8186 ;
  assign n8236 = ~n8189 & ~n8235 ;
  assign n8237 = n8164 & ~n8236 ;
  assign n8238 = ~n8185 & n8237 ;
  assign n8239 = n8164 & n8201 ;
  assign n8240 = ~n8214 & ~n8239 ;
  assign n8241 = n8185 & ~n8240 ;
  assign n8242 = ~n8238 & ~n8241 ;
  assign n8243 = ~n8212 & n8242 ;
  assign n8244 = ~n8234 & n8243 ;
  assign n8245 = ~\u2_L12_reg[14]/NET0131  & ~n8244 ;
  assign n8246 = \u2_L12_reg[14]/NET0131  & n8244 ;
  assign n8247 = ~n8245 & ~n8246 ;
  assign n8250 = n7456 & ~n7466 ;
  assign n8251 = ~n7977 & ~n8250 ;
  assign n8252 = n7443 & ~n8251 ;
  assign n8249 = ~n7443 & ~n7988 ;
  assign n8248 = n7449 & n7509 ;
  assign n8253 = ~n7437 & ~n8248 ;
  assign n8254 = ~n8249 & n8253 ;
  assign n8255 = ~n8252 & n8254 ;
  assign n8258 = n7449 & n7516 ;
  assign n8259 = ~n7443 & n7479 ;
  assign n8260 = n7437 & ~n7488 ;
  assign n8261 = ~n8259 & n8260 ;
  assign n8262 = ~n8258 & n8261 ;
  assign n8256 = ~n7467 & ~n7486 ;
  assign n8257 = n7443 & ~n8256 ;
  assign n8263 = ~n7760 & ~n8257 ;
  assign n8264 = n8262 & n8263 ;
  assign n8265 = ~n8255 & ~n8264 ;
  assign n8266 = n7477 & n7483 ;
  assign n8267 = ~n7504 & ~n8266 ;
  assign n8268 = ~n8265 & n8267 ;
  assign n8269 = ~\u2_L12_reg[19]/NET0131  & ~n8268 ;
  assign n8270 = \u2_L12_reg[19]/NET0131  & n8268 ;
  assign n8271 = ~n8269 & ~n8270 ;
  assign n8272 = ~n7654 & n7669 ;
  assign n8273 = ~n7696 & ~n8272 ;
  assign n8274 = n7677 & ~n8273 ;
  assign n8275 = n7633 & ~n7700 ;
  assign n8276 = n8024 & n8275 ;
  assign n8277 = ~n8274 & n8276 ;
  assign n8279 = n7654 & n7680 ;
  assign n8278 = n7627 & n7695 ;
  assign n8280 = ~n7633 & ~n8278 ;
  assign n8281 = ~n8279 & n8280 ;
  assign n8282 = ~n8277 & ~n8281 ;
  assign n8283 = n7647 & ~n7654 ;
  assign n8284 = ~n7633 & ~n7702 ;
  assign n8285 = ~n8283 & n8284 ;
  assign n8286 = ~n7646 & n7661 ;
  assign n8287 = n7633 & ~n7664 ;
  assign n8288 = ~n8286 & n8287 ;
  assign n8289 = ~n8285 & ~n8288 ;
  assign n8290 = ~n7647 & ~n7656 ;
  assign n8291 = n8027 & ~n8290 ;
  assign n8292 = ~n7677 & ~n8022 ;
  assign n8293 = ~n8291 & n8292 ;
  assign n8294 = ~n8289 & n8293 ;
  assign n8296 = ~n7647 & n8027 ;
  assign n8297 = ~n7657 & ~n8296 ;
  assign n8298 = ~n7633 & ~n8297 ;
  assign n8295 = ~n7640 & n7663 ;
  assign n8299 = n7677 & ~n8295 ;
  assign n8300 = ~n8278 & n8299 ;
  assign n8301 = ~n8298 & n8300 ;
  assign n8302 = ~n8294 & ~n8301 ;
  assign n8303 = ~n8282 & ~n8302 ;
  assign n8304 = ~\u2_L12_reg[1]/NET0131  & ~n8303 ;
  assign n8305 = \u2_L12_reg[1]/NET0131  & n8303 ;
  assign n8306 = ~n8304 & ~n8305 ;
  assign n8312 = ~n7924 & ~n7939 ;
  assign n8313 = ~n8133 & ~n8312 ;
  assign n8316 = n7904 & ~n7945 ;
  assign n8314 = n7890 & n7917 ;
  assign n8315 = n7891 & n7912 ;
  assign n8317 = ~n8314 & ~n8315 ;
  assign n8318 = n8316 & n8317 ;
  assign n8319 = ~n8313 & ~n8318 ;
  assign n8310 = ~n7927 & ~n7949 ;
  assign n8311 = n7884 & ~n8310 ;
  assign n8320 = n7897 & n7963 ;
  assign n8321 = n7937 & ~n8320 ;
  assign n8322 = ~n8311 & n8321 ;
  assign n8323 = ~n8319 & n8322 ;
  assign n8332 = ~n7916 & ~n7950 ;
  assign n8327 = n7897 & n8134 ;
  assign n8328 = ~n7904 & n7955 ;
  assign n8333 = ~n8327 & ~n8328 ;
  assign n8334 = n8332 & n8333 ;
  assign n8325 = ~n7915 & ~n7927 ;
  assign n8326 = n7904 & ~n8325 ;
  assign n8329 = ~n7937 & ~n7965 ;
  assign n8308 = n7905 & n7956 ;
  assign n8324 = n7917 & n7939 ;
  assign n8330 = ~n8308 & ~n8324 ;
  assign n8331 = n8329 & n8330 ;
  assign n8335 = ~n8326 & n8331 ;
  assign n8336 = n8334 & n8335 ;
  assign n8337 = ~n8323 & ~n8336 ;
  assign n8307 = n7904 & n7963 ;
  assign n8309 = n7890 & n8308 ;
  assign n8338 = ~n8307 & ~n8309 ;
  assign n8339 = ~n8337 & n8338 ;
  assign n8340 = ~\u2_L12_reg[21]/NET0131  & ~n8339 ;
  assign n8341 = \u2_L12_reg[21]/NET0131  & n8339 ;
  assign n8342 = ~n8340 & ~n8341 ;
  assign n8344 = n7360 & n7397 ;
  assign n8363 = ~n7360 & n7368 ;
  assign n8364 = ~n8344 & ~n8363 ;
  assign n8365 = ~n7373 & n8364 ;
  assign n8366 = n7383 & ~n8365 ;
  assign n8367 = n7368 & n7393 ;
  assign n8368 = ~n7721 & ~n8367 ;
  assign n8369 = ~n8366 & n8368 ;
  assign n8370 = ~n7341 & ~n8369 ;
  assign n8357 = n7360 & n7368 ;
  assign n8358 = ~n7413 & ~n8357 ;
  assign n8359 = n7341 & ~n8358 ;
  assign n8360 = ~n7409 & ~n7421 ;
  assign n8361 = ~n8359 & n8360 ;
  assign n8362 = n7383 & ~n8361 ;
  assign n8345 = ~n7369 & ~n8344 ;
  assign n8346 = n7341 & ~n8345 ;
  assign n8349 = ~n7394 & ~n7720 ;
  assign n8343 = n7367 & n7392 ;
  assign n8347 = ~n7341 & n7347 ;
  assign n8348 = n7386 & n8347 ;
  assign n8350 = ~n8343 & ~n8348 ;
  assign n8351 = n8349 & n8350 ;
  assign n8352 = ~n8346 & n8351 ;
  assign n8353 = ~n7383 & ~n8352 ;
  assign n8354 = n7341 & n7418 ;
  assign n8355 = ~n8348 & ~n8354 ;
  assign n8356 = n7360 & ~n8355 ;
  assign n8371 = ~n7411 & ~n8356 ;
  assign n8372 = ~n8353 & n8371 ;
  assign n8373 = ~n8362 & n8372 ;
  assign n8374 = ~n8370 & n8373 ;
  assign n8375 = \u2_L12_reg[23]/NET0131  & ~n8374 ;
  assign n8376 = ~\u2_L12_reg[23]/NET0131  & n8374 ;
  assign n8377 = ~n8375 & ~n8376 ;
  assign n8384 = n8164 & ~n8171 ;
  assign n8394 = n8158 & ~n8384 ;
  assign n8395 = ~n8185 & ~n8394 ;
  assign n8397 = ~n8225 & ~n8395 ;
  assign n8398 = n8158 & ~n8397 ;
  assign n8396 = n8190 & n8395 ;
  assign n8400 = n8185 & ~n8186 ;
  assign n8383 = ~n8158 & ~n8171 ;
  assign n8399 = ~n8185 & ~n8383 ;
  assign n8401 = ~n8164 & ~n8399 ;
  assign n8402 = ~n8400 & n8401 ;
  assign n8403 = ~n8396 & ~n8402 ;
  assign n8404 = ~n8398 & n8403 ;
  assign n8405 = ~n8152 & ~n8404 ;
  assign n8380 = ~n8158 & n8193 ;
  assign n8381 = ~n8185 & ~n8380 ;
  assign n8382 = ~n8172 & n8381 ;
  assign n8385 = ~n8191 & ~n8384 ;
  assign n8386 = ~n8178 & ~n8385 ;
  assign n8387 = n8185 & ~n8383 ;
  assign n8388 = ~n8194 & n8387 ;
  assign n8389 = ~n8386 & n8388 ;
  assign n8390 = ~n8382 & ~n8389 ;
  assign n8378 = n8165 & n8178 ;
  assign n8379 = n8171 & n8187 ;
  assign n8391 = ~n8378 & ~n8379 ;
  assign n8392 = ~n8390 & n8391 ;
  assign n8393 = n8152 & ~n8392 ;
  assign n8408 = ~n8239 & ~n8379 ;
  assign n8409 = n8188 & n8191 ;
  assign n8410 = n8408 & ~n8409 ;
  assign n8411 = n8185 & ~n8410 ;
  assign n8406 = n8171 & ~n8185 ;
  assign n8407 = n8207 & n8406 ;
  assign n8412 = ~n8195 & ~n8407 ;
  assign n8413 = ~n8411 & n8412 ;
  assign n8414 = ~n8393 & n8413 ;
  assign n8415 = ~n8405 & n8414 ;
  assign n8416 = ~\u2_L12_reg[25]/NET0131  & ~n8415 ;
  assign n8417 = \u2_L12_reg[25]/NET0131  & n8415 ;
  assign n8418 = ~n8416 & ~n8417 ;
  assign n8428 = ~n7695 & ~n8286 ;
  assign n8429 = n7627 & ~n8428 ;
  assign n8436 = n7677 & ~n7692 ;
  assign n8437 = ~n8429 & n8436 ;
  assign n8430 = ~n7657 & ~n7684 ;
  assign n8431 = n7654 & ~n8430 ;
  assign n8432 = ~n7627 & n8012 ;
  assign n8433 = ~n7678 & ~n8432 ;
  assign n8434 = ~n7633 & ~n8009 ;
  assign n8435 = ~n8433 & n8434 ;
  assign n8438 = ~n8431 & ~n8435 ;
  assign n8439 = n8437 & n8438 ;
  assign n8440 = ~n7656 & n7693 ;
  assign n8441 = ~n7677 & ~n8272 ;
  assign n8442 = ~n8440 & n8441 ;
  assign n8443 = n7686 & n8442 ;
  assign n8444 = ~n8439 & ~n8443 ;
  assign n8419 = ~n7646 & ~n7670 ;
  assign n8420 = ~n7679 & ~n8419 ;
  assign n8421 = ~n7654 & ~n8420 ;
  assign n8422 = ~n7660 & ~n8295 ;
  assign n8423 = ~n7677 & ~n8422 ;
  assign n8424 = ~n8421 & ~n8423 ;
  assign n8425 = ~n7633 & ~n8424 ;
  assign n8426 = n7633 & n8012 ;
  assign n8427 = ~n7670 & n8426 ;
  assign n8445 = ~n8425 & ~n8427 ;
  assign n8446 = ~n8444 & n8445 ;
  assign n8447 = ~\u2_L12_reg[26]/NET0131  & ~n8446 ;
  assign n8448 = \u2_L12_reg[26]/NET0131  & n8446 ;
  assign n8449 = ~n8447 & ~n8448 ;
  assign n8453 = ~n7823 & ~n7824 ;
  assign n8454 = n7816 & n8453 ;
  assign n8452 = n7823 & n7861 ;
  assign n8455 = n7791 & ~n7859 ;
  assign n8456 = ~n8452 & n8455 ;
  assign n8457 = ~n8454 & n8456 ;
  assign n8459 = ~n7791 & ~n7817 ;
  assign n8458 = ~n7831 & ~n8102 ;
  assign n8460 = ~n8081 & n8458 ;
  assign n8461 = n8459 & n8460 ;
  assign n8462 = ~n8457 & ~n8461 ;
  assign n8450 = ~n7859 & ~n7861 ;
  assign n8451 = n7824 & ~n8450 ;
  assign n8463 = n7847 & ~n8451 ;
  assign n8464 = ~n8462 & n8463 ;
  assign n8465 = n7791 & n8458 ;
  assign n8466 = ~n7819 & ~n7825 ;
  assign n8467 = ~n8075 & n8466 ;
  assign n8468 = n8459 & n8467 ;
  assign n8469 = ~n8465 & ~n8468 ;
  assign n8470 = n7809 & n8087 ;
  assign n8471 = ~n7847 & ~n8081 ;
  assign n8472 = ~n8470 & n8471 ;
  assign n8473 = ~n8469 & n8472 ;
  assign n8474 = ~n8464 & ~n8473 ;
  assign n8475 = ~\u2_L12_reg[28]/NET0131  & n8474 ;
  assign n8476 = \u2_L12_reg[28]/NET0131  & ~n8474 ;
  assign n8477 = ~n8475 & ~n8476 ;
  assign n8478 = ~n8185 & ~n8223 ;
  assign n8479 = n8172 & n8178 ;
  assign n8480 = n8188 & n8207 ;
  assign n8481 = n8185 & ~n8187 ;
  assign n8482 = ~n8480 & n8481 ;
  assign n8483 = ~n8479 & n8482 ;
  assign n8484 = ~n8478 & ~n8483 ;
  assign n8486 = ~n8164 & n8201 ;
  assign n8487 = ~n8380 & ~n8486 ;
  assign n8488 = n8185 & ~n8487 ;
  assign n8485 = n8171 & n8215 ;
  assign n8489 = n8152 & ~n8485 ;
  assign n8490 = ~n8237 & n8489 ;
  assign n8491 = ~n8488 & n8490 ;
  assign n8492 = n8188 & ~n8207 ;
  assign n8493 = n8381 & ~n8492 ;
  assign n8494 = n8185 & ~n8192 ;
  assign n8495 = ~n8194 & n8494 ;
  assign n8496 = ~n8493 & ~n8495 ;
  assign n8497 = ~n8152 & ~n8172 ;
  assign n8498 = n8408 & n8497 ;
  assign n8499 = ~n8496 & n8498 ;
  assign n8500 = ~n8491 & ~n8499 ;
  assign n8501 = ~n8484 & ~n8500 ;
  assign n8502 = ~\u2_L12_reg[8]/NET0131  & ~n8501 ;
  assign n8503 = \u2_L12_reg[8]/NET0131  & n8501 ;
  assign n8504 = ~n8502 & ~n8503 ;
  assign n8505 = ~n7927 & ~n7963 ;
  assign n8506 = ~n8314 & n8505 ;
  assign n8507 = ~n7904 & ~n8506 ;
  assign n8508 = n7904 & ~n7923 ;
  assign n8509 = n8114 & n8508 ;
  assign n8510 = ~n7916 & ~n7945 ;
  assign n8511 = ~n7966 & n8510 ;
  assign n8512 = ~n8509 & n8511 ;
  assign n8513 = ~n8507 & n8512 ;
  assign n8514 = n7937 & ~n8513 ;
  assign n8518 = n7904 & ~n7965 ;
  assign n8516 = ~n7897 & n8125 ;
  assign n8517 = n7897 & ~n8125 ;
  assign n8519 = ~n8516 & ~n8517 ;
  assign n8520 = n8518 & n8519 ;
  assign n8515 = n7939 & n7956 ;
  assign n8521 = ~n7948 & ~n8515 ;
  assign n8522 = ~n8328 & n8521 ;
  assign n8523 = ~n8520 & n8522 ;
  assign n8524 = ~n7937 & ~n8523 ;
  assign n8527 = ~n7904 & ~n7947 ;
  assign n8525 = ~n7897 & n7904 ;
  assign n8526 = n8127 & n8525 ;
  assign n8528 = ~n7954 & ~n8526 ;
  assign n8529 = ~n8527 & n8528 ;
  assign n8530 = ~n8524 & n8529 ;
  assign n8531 = ~n8514 & n8530 ;
  assign n8532 = \u2_L12_reg[27]/NET0131  & n8531 ;
  assign n8533 = ~\u2_L12_reg[27]/NET0131  & ~n8531 ;
  assign n8534 = ~n8532 & ~n8533 ;
  assign n8540 = ~n7560 & n7593 ;
  assign n8539 = n7561 & ~n8043 ;
  assign n8541 = ~n8048 & ~n8539 ;
  assign n8542 = ~n8540 & n8541 ;
  assign n8543 = ~n7541 & ~n8542 ;
  assign n8535 = n7567 & ~n8052 ;
  assign n8536 = n7608 & n8535 ;
  assign n8537 = ~n7573 & ~n7579 ;
  assign n8538 = n7541 & ~n8537 ;
  assign n8544 = ~n8536 & ~n8538 ;
  assign n8545 = ~n8543 & n8544 ;
  assign n8546 = n7535 & ~n8545 ;
  assign n8553 = ~n7541 & ~n7568 ;
  assign n8554 = ~n8045 & n8553 ;
  assign n8551 = ~n7579 & ~n7608 ;
  assign n8552 = n8535 & n8551 ;
  assign n8555 = ~n7609 & ~n8552 ;
  assign n8556 = ~n8554 & n8555 ;
  assign n8557 = ~n7535 & ~n8556 ;
  assign n8547 = n7590 & ~n7594 ;
  assign n8548 = n7589 & n8547 ;
  assign n8549 = n7535 & ~n7541 ;
  assign n8550 = n7577 & ~n8549 ;
  assign n8558 = ~n8548 & ~n8550 ;
  assign n8559 = ~n8557 & n8558 ;
  assign n8560 = ~n8546 & n8559 ;
  assign n8561 = \u2_L12_reg[32]/NET0131  & n8560 ;
  assign n8562 = ~\u2_L12_reg[32]/NET0131  & ~n8560 ;
  assign n8563 = ~n8561 & ~n8562 ;
  assign n8565 = ~n8224 & ~n8235 ;
  assign n8566 = n8185 & ~n8565 ;
  assign n8564 = ~n8185 & n8216 ;
  assign n8567 = ~n8195 & ~n8223 ;
  assign n8568 = ~n8564 & n8567 ;
  assign n8569 = ~n8566 & n8568 ;
  assign n8570 = n8152 & ~n8569 ;
  assign n8572 = ~n8164 & n8188 ;
  assign n8571 = ~n8190 & n8207 ;
  assign n8573 = ~n8213 & ~n8571 ;
  assign n8574 = ~n8572 & n8573 ;
  assign n8575 = ~n8152 & ~n8574 ;
  assign n8576 = ~n8480 & n8494 ;
  assign n8577 = ~n8575 & n8576 ;
  assign n8578 = n8152 & ~n8208 ;
  assign n8579 = ~n8200 & ~n8202 ;
  assign n8580 = ~n8380 & n8579 ;
  assign n8581 = ~n8578 & ~n8580 ;
  assign n8582 = ~n8185 & ~n8214 ;
  assign n8583 = ~n8486 & n8582 ;
  assign n8584 = ~n8581 & n8583 ;
  assign n8585 = ~n8577 & ~n8584 ;
  assign n8586 = ~n8570 & ~n8585 ;
  assign n8587 = ~\u2_L12_reg[3]/NET0131  & ~n8586 ;
  assign n8588 = \u2_L12_reg[3]/NET0131  & n8586 ;
  assign n8589 = ~n8587 & ~n8588 ;
  assign n8623 = decrypt_pad & ~\u2_uk_K_r12_reg[13]/NET0131  ;
  assign n8624 = ~decrypt_pad & ~\u2_uk_K_r12_reg[46]/NET0131  ;
  assign n8625 = ~n8623 & ~n8624 ;
  assign n8626 = \u2_R12_reg[12]/NET0131  & ~n8625 ;
  assign n8627 = ~\u2_R12_reg[12]/NET0131  & n8625 ;
  assign n8628 = ~n8626 & ~n8627 ;
  assign n8590 = decrypt_pad & ~\u2_uk_K_r12_reg[26]/NET0131  ;
  assign n8591 = ~decrypt_pad & ~\u2_uk_K_r12_reg[34]/NET0131  ;
  assign n8592 = ~n8590 & ~n8591 ;
  assign n8593 = \u2_R12_reg[13]/NET0131  & ~n8592 ;
  assign n8594 = ~\u2_R12_reg[13]/NET0131  & n8592 ;
  assign n8595 = ~n8593 & ~n8594 ;
  assign n8603 = decrypt_pad & ~\u2_uk_K_r12_reg[17]/NET0131  ;
  assign n8604 = ~decrypt_pad & ~\u2_uk_K_r12_reg[25]/NET0131  ;
  assign n8605 = ~n8603 & ~n8604 ;
  assign n8606 = \u2_R12_reg[8]/NET0131  & ~n8605 ;
  assign n8607 = ~\u2_R12_reg[8]/NET0131  & n8605 ;
  assign n8608 = ~n8606 & ~n8607 ;
  assign n8610 = ~n8595 & ~n8608 ;
  assign n8611 = n8595 & n8608 ;
  assign n8612 = ~n8610 & ~n8611 ;
  assign n8596 = decrypt_pad & ~\u2_uk_K_r12_reg[46]/NET0131  ;
  assign n8597 = ~decrypt_pad & ~\u2_uk_K_r12_reg[54]/NET0131  ;
  assign n8598 = ~n8596 & ~n8597 ;
  assign n8599 = \u2_R12_reg[9]/NET0131  & ~n8598 ;
  assign n8600 = ~\u2_R12_reg[9]/NET0131  & n8598 ;
  assign n8601 = ~n8599 & ~n8600 ;
  assign n8613 = decrypt_pad & ~\u2_uk_K_r12_reg[54]/NET0131  ;
  assign n8614 = ~decrypt_pad & ~\u2_uk_K_r12_reg[5]/NET0131  ;
  assign n8615 = ~n8613 & ~n8614 ;
  assign n8616 = \u2_R12_reg[10]/NET0131  & ~n8615 ;
  assign n8617 = ~\u2_R12_reg[10]/NET0131  & n8615 ;
  assign n8618 = ~n8616 & ~n8617 ;
  assign n8664 = ~n8601 & n8618 ;
  assign n8665 = ~n8612 & n8664 ;
  assign n8653 = n8595 & ~n8608 ;
  assign n8654 = n8601 & n8653 ;
  assign n8635 = decrypt_pad & ~\u2_uk_K_r12_reg[55]/NET0131  ;
  assign n8636 = ~decrypt_pad & ~\u2_uk_K_r12_reg[6]/NET0131  ;
  assign n8637 = ~n8635 & ~n8636 ;
  assign n8638 = \u2_R12_reg[11]/NET0131  & ~n8637 ;
  assign n8639 = ~\u2_R12_reg[11]/NET0131  & n8637 ;
  assign n8640 = ~n8638 & ~n8639 ;
  assign n8655 = n8618 & ~n8640 ;
  assign n8656 = n8654 & n8655 ;
  assign n8661 = ~n8595 & n8601 ;
  assign n8662 = n8618 & n8661 ;
  assign n8663 = n8608 & n8662 ;
  assign n8666 = ~n8656 & ~n8663 ;
  assign n8667 = ~n8665 & n8666 ;
  assign n8646 = n8601 & ~n8618 ;
  assign n8657 = n8595 & n8640 ;
  assign n8658 = n8612 & ~n8657 ;
  assign n8659 = n8646 & ~n8658 ;
  assign n8630 = ~n8601 & ~n8618 ;
  assign n8660 = n8630 & n8658 ;
  assign n8668 = ~n8659 & ~n8660 ;
  assign n8669 = n8667 & n8668 ;
  assign n8670 = ~n8628 & ~n8669 ;
  assign n8602 = n8595 & ~n8601 ;
  assign n8609 = ~n8601 & n8608 ;
  assign n8619 = ~n8608 & ~n8618 ;
  assign n8620 = ~n8609 & ~n8619 ;
  assign n8621 = n8612 & n8620 ;
  assign n8622 = ~n8602 & ~n8621 ;
  assign n8629 = ~n8622 & n8628 ;
  assign n8631 = n8610 & n8630 ;
  assign n8632 = n8602 & n8618 ;
  assign n8633 = ~n8631 & ~n8632 ;
  assign n8634 = ~n8629 & n8633 ;
  assign n8641 = ~n8634 & n8640 ;
  assign n8642 = n8618 & n8628 ;
  assign n8643 = n8601 & n8610 ;
  assign n8644 = n8642 & n8643 ;
  assign n8645 = n8628 & ~n8640 ;
  assign n8647 = n8595 & n8646 ;
  assign n8648 = ~n8595 & n8609 ;
  assign n8649 = n8601 & n8611 ;
  assign n8650 = ~n8648 & ~n8649 ;
  assign n8651 = ~n8647 & n8650 ;
  assign n8652 = n8645 & ~n8651 ;
  assign n8671 = ~n8644 & ~n8652 ;
  assign n8672 = ~n8641 & n8671 ;
  assign n8673 = ~n8670 & n8672 ;
  assign n8674 = ~\u2_L12_reg[6]/NET0131  & ~n8673 ;
  assign n8675 = \u2_L12_reg[6]/NET0131  & n8673 ;
  assign n8676 = ~n8674 & ~n8675 ;
  assign n8679 = n7554 & n8043 ;
  assign n8677 = n7554 & n7560 ;
  assign n8678 = ~n8043 & ~n8677 ;
  assign n8680 = ~n7611 & ~n8678 ;
  assign n8681 = ~n8679 & n8680 ;
  assign n8682 = ~n7535 & n7541 ;
  assign n8683 = ~n8549 & ~n8682 ;
  assign n8684 = ~n7592 & n8683 ;
  assign n8685 = ~n8681 & n8684 ;
  assign n8688 = ~n7576 & n8051 ;
  assign n8687 = n7560 & ~n8043 ;
  assign n8686 = n7567 & n7608 ;
  assign n8689 = n8549 & ~n8686 ;
  assign n8690 = ~n8687 & n8689 ;
  assign n8691 = ~n8688 & n8690 ;
  assign n8692 = ~n8685 & ~n8691 ;
  assign n8693 = ~n8540 & ~n8692 ;
  assign n8694 = n7547 & ~n7560 ;
  assign n8695 = n8679 & ~n8694 ;
  assign n8696 = ~n8678 & n8682 ;
  assign n8697 = ~n8695 & n8696 ;
  assign n8698 = ~n8693 & ~n8697 ;
  assign n8699 = ~\u2_L12_reg[7]/NET0131  & n8698 ;
  assign n8700 = \u2_L12_reg[7]/NET0131  & ~n8698 ;
  assign n8701 = ~n8699 & ~n8700 ;
  assign n8702 = ~n7369 & ~n7414 ;
  assign n8703 = n7392 & ~n8702 ;
  assign n8706 = n7736 & n8364 ;
  assign n8707 = n7347 & ~n8706 ;
  assign n8704 = ~n7371 & ~n8357 ;
  assign n8705 = n7401 & ~n8704 ;
  assign n8708 = n7722 & ~n8705 ;
  assign n8709 = ~n8707 & n8708 ;
  assign n8710 = ~n7374 & ~n7412 ;
  assign n8711 = ~n8344 & n8710 ;
  assign n8712 = n7341 & ~n8711 ;
  assign n8715 = ~n7341 & ~n8704 ;
  assign n8714 = n7347 & n7729 ;
  assign n8713 = ~n7347 & n7735 ;
  assign n8716 = ~n7383 & ~n8713 ;
  assign n8717 = ~n8714 & n8716 ;
  assign n8718 = ~n8715 & n8717 ;
  assign n8719 = ~n8712 & n8718 ;
  assign n8720 = ~n8709 & ~n8719 ;
  assign n8721 = ~n8703 & ~n8720 ;
  assign n8722 = ~\u2_L12_reg[9]/NET0131  & ~n8721 ;
  assign n8723 = \u2_L12_reg[9]/NET0131  & n8721 ;
  assign n8724 = ~n8722 & ~n8723 ;
  assign n8725 = n8618 & ~n8654 ;
  assign n8727 = n8640 & n8643 ;
  assign n8726 = n8602 & ~n8608 ;
  assign n8728 = ~n8618 & ~n8726 ;
  assign n8729 = n8650 & n8728 ;
  assign n8730 = ~n8727 & n8729 ;
  assign n8731 = ~n8725 & ~n8730 ;
  assign n8732 = n8610 & n8618 ;
  assign n8733 = ~n8601 & n8732 ;
  assign n8734 = n8640 & ~n8663 ;
  assign n8735 = ~n8733 & n8734 ;
  assign n8736 = n8608 & n8618 ;
  assign n8737 = ~n8595 & ~n8619 ;
  assign n8738 = ~n8736 & n8737 ;
  assign n8739 = ~n8735 & n8738 ;
  assign n8740 = ~n8731 & ~n8739 ;
  assign n8741 = n8628 & ~n8740 ;
  assign n8742 = ~n8601 & n8736 ;
  assign n8743 = ~n8640 & ~n8742 ;
  assign n8744 = ~n8735 & ~n8743 ;
  assign n8749 = n8610 & ~n8618 ;
  assign n8750 = ~n8649 & ~n8726 ;
  assign n8751 = ~n8749 & n8750 ;
  assign n8752 = ~n8640 & ~n8751 ;
  assign n8746 = ~n8610 & n8640 ;
  assign n8745 = ~n8601 & ~n8611 ;
  assign n8747 = ~n8649 & ~n8745 ;
  assign n8748 = n8746 & n8747 ;
  assign n8753 = ~n8631 & ~n8748 ;
  assign n8754 = ~n8752 & n8753 ;
  assign n8755 = ~n8628 & ~n8754 ;
  assign n8756 = ~n8744 & ~n8755 ;
  assign n8757 = ~n8741 & n8756 ;
  assign n8758 = ~\u2_L12_reg[16]/NET0131  & ~n8757 ;
  assign n8759 = \u2_L12_reg[16]/NET0131  & n8757 ;
  assign n8760 = ~n8758 & ~n8759 ;
  assign n8765 = n7791 & ~n7826 ;
  assign n8762 = ~n7803 & n7852 ;
  assign n8763 = ~n7860 & ~n8762 ;
  assign n8764 = ~n7791 & ~n8763 ;
  assign n8766 = ~n7818 & ~n8764 ;
  assign n8767 = ~n8765 & n8766 ;
  assign n8768 = n7847 & ~n8767 ;
  assign n8775 = n7803 & ~n7853 ;
  assign n8776 = n7871 & ~n8775 ;
  assign n8774 = n7836 & ~n8453 ;
  assign n8772 = n7791 & n7797 ;
  assign n8773 = n7819 & n8772 ;
  assign n8777 = ~n7865 & ~n8773 ;
  assign n8778 = ~n8774 & n8777 ;
  assign n8779 = ~n8776 & n8778 ;
  assign n8780 = ~n7847 & ~n8779 ;
  assign n8761 = ~n7791 & n7831 ;
  assign n8769 = n7797 & n7836 ;
  assign n8770 = ~n8103 & ~n8769 ;
  assign n8771 = n7791 & ~n8770 ;
  assign n8781 = ~n8761 & ~n8771 ;
  assign n8782 = ~n8780 & n8781 ;
  assign n8783 = ~n8768 & n8782 ;
  assign n8784 = ~\u2_L12_reg[18]/P0001  & ~n8783 ;
  assign n8785 = \u2_L12_reg[18]/P0001  & n8783 ;
  assign n8786 = ~n8784 & ~n8785 ;
  assign n8796 = ~n8618 & n8640 ;
  assign n8807 = ~n8601 & ~n8653 ;
  assign n8808 = n8796 & n8807 ;
  assign n8803 = ~n8630 & ~n8640 ;
  assign n8804 = ~n8612 & n8803 ;
  assign n8805 = ~n8609 & n8618 ;
  assign n8806 = n8746 & n8805 ;
  assign n8809 = ~n8804 & ~n8806 ;
  assign n8810 = ~n8808 & n8809 ;
  assign n8811 = ~n8660 & n8810 ;
  assign n8812 = n8628 & ~n8811 ;
  assign n8787 = n8595 & n8619 ;
  assign n8788 = ~n8732 & ~n8787 ;
  assign n8789 = ~n8643 & ~n8742 ;
  assign n8790 = n8788 & n8789 ;
  assign n8791 = n8640 & ~n8790 ;
  assign n8792 = ~n8595 & n8742 ;
  assign n8793 = ~n8791 & ~n8792 ;
  assign n8794 = ~n8628 & ~n8793 ;
  assign n8799 = ~n8612 & n8630 ;
  assign n8800 = ~n8621 & ~n8799 ;
  assign n8801 = ~n8628 & ~n8640 ;
  assign n8802 = ~n8800 & n8801 ;
  assign n8795 = n8649 & n8655 ;
  assign n8797 = ~n8648 & ~n8654 ;
  assign n8798 = n8796 & ~n8797 ;
  assign n8813 = ~n8795 & ~n8798 ;
  assign n8814 = ~n8802 & n8813 ;
  assign n8815 = ~n8794 & n8814 ;
  assign n8816 = ~n8812 & n8815 ;
  assign n8817 = ~\u2_L12_reg[24]/NET0131  & ~n8816 ;
  assign n8818 = \u2_L12_reg[24]/NET0131  & n8816 ;
  assign n8819 = ~n8817 & ~n8818 ;
  assign n8821 = ~n8618 & n8648 ;
  assign n8822 = n8788 & ~n8821 ;
  assign n8823 = n8628 & ~n8822 ;
  assign n8824 = ~n8661 & ~n8736 ;
  assign n8825 = ~n8628 & ~n8662 ;
  assign n8826 = ~n8824 & n8825 ;
  assign n8827 = ~n8823 & ~n8826 ;
  assign n8828 = n8640 & ~n8827 ;
  assign n8832 = n8618 & n8726 ;
  assign n8829 = ~n8601 & ~n8608 ;
  assign n8830 = ~n8640 & ~n8829 ;
  assign n8831 = n8824 & n8830 ;
  assign n8833 = ~n8799 & ~n8831 ;
  assign n8834 = ~n8832 & n8833 ;
  assign n8835 = ~n8628 & ~n8834 ;
  assign n8836 = ~n8643 & ~n8736 ;
  assign n8837 = n8645 & ~n8836 ;
  assign n8839 = n8601 & ~n8611 ;
  assign n8840 = n8642 & n8839 ;
  assign n8820 = n8655 & n8661 ;
  assign n8838 = n8657 & n8742 ;
  assign n8841 = ~n8820 & ~n8838 ;
  assign n8842 = ~n8840 & n8841 ;
  assign n8843 = ~n8837 & n8842 ;
  assign n8844 = ~n8835 & n8843 ;
  assign n8845 = ~n8828 & n8844 ;
  assign n8846 = \u2_L12_reg[30]/NET0131  & ~n8845 ;
  assign n8847 = ~\u2_L12_reg[30]/NET0131  & n8845 ;
  assign n8848 = ~n8846 & ~n8847 ;
  assign n8855 = decrypt_pad & ~\u2_uk_K_r11_reg[2]/NET0131  ;
  assign n8856 = ~decrypt_pad & ~\u2_uk_K_r11_reg[35]/NET0131  ;
  assign n8857 = ~n8855 & ~n8856 ;
  assign n8858 = \u2_R11_reg[26]/NET0131  & ~n8857 ;
  assign n8859 = ~\u2_R11_reg[26]/NET0131  & n8857 ;
  assign n8860 = ~n8858 & ~n8859 ;
  assign n8849 = decrypt_pad & ~\u2_uk_K_r11_reg[37]/NET0131  ;
  assign n8850 = ~decrypt_pad & ~\u2_uk_K_r11_reg[15]/NET0131  ;
  assign n8851 = ~n8849 & ~n8850 ;
  assign n8852 = \u2_R11_reg[24]/NET0131  & ~n8851 ;
  assign n8853 = ~\u2_R11_reg[24]/NET0131  & n8851 ;
  assign n8854 = ~n8852 & ~n8853 ;
  assign n8879 = decrypt_pad & ~\u2_uk_K_r11_reg[14]/NET0131  ;
  assign n8880 = ~decrypt_pad & ~\u2_uk_K_r11_reg[23]/NET0131  ;
  assign n8881 = ~n8879 & ~n8880 ;
  assign n8882 = \u2_R11_reg[29]/NET0131  & ~n8881 ;
  assign n8883 = ~\u2_R11_reg[29]/NET0131  & n8881 ;
  assign n8884 = ~n8882 & ~n8883 ;
  assign n8890 = ~n8854 & ~n8884 ;
  assign n8891 = n8860 & n8890 ;
  assign n8864 = decrypt_pad & ~\u2_uk_K_r11_reg[35]/NET0131  ;
  assign n8865 = ~decrypt_pad & ~\u2_uk_K_r11_reg[44]/NET0131  ;
  assign n8866 = ~n8864 & ~n8865 ;
  assign n8867 = \u2_R11_reg[27]/NET0131  & ~n8866 ;
  assign n8868 = ~\u2_R11_reg[27]/NET0131  & n8866 ;
  assign n8869 = ~n8867 & ~n8868 ;
  assign n8908 = n8854 & n8869 ;
  assign n8909 = ~n8891 & ~n8908 ;
  assign n8870 = decrypt_pad & ~\u2_uk_K_r11_reg[45]/NET0131  ;
  assign n8871 = ~decrypt_pad & ~\u2_uk_K_r11_reg[50]/NET0131  ;
  assign n8872 = ~n8870 & ~n8871 ;
  assign n8873 = \u2_R11_reg[25]/NET0131  & ~n8872 ;
  assign n8874 = ~\u2_R11_reg[25]/NET0131  & n8872 ;
  assign n8875 = ~n8873 & ~n8874 ;
  assign n8910 = n8860 & n8869 ;
  assign n8911 = ~n8875 & ~n8910 ;
  assign n8912 = ~n8909 & n8911 ;
  assign n8861 = ~n8854 & ~n8860 ;
  assign n8862 = n8854 & n8860 ;
  assign n8863 = ~n8861 & ~n8862 ;
  assign n8878 = n8869 & ~n8875 ;
  assign n8913 = ~n8878 & n8884 ;
  assign n8914 = ~n8863 & n8913 ;
  assign n8885 = ~n8860 & ~n8884 ;
  assign n8898 = n8860 & n8875 ;
  assign n8899 = ~n8885 & ~n8898 ;
  assign n8900 = n8854 & ~n8869 ;
  assign n8901 = ~n8899 & n8900 ;
  assign n8902 = decrypt_pad & ~\u2_uk_K_r11_reg[22]/NET0131  ;
  assign n8903 = ~decrypt_pad & ~\u2_uk_K_r11_reg[0]/NET0131  ;
  assign n8904 = ~n8902 & ~n8903 ;
  assign n8905 = \u2_R11_reg[28]/NET0131  & ~n8904 ;
  assign n8906 = ~\u2_R11_reg[28]/NET0131  & n8904 ;
  assign n8907 = ~n8905 & ~n8906 ;
  assign n8915 = ~n8901 & ~n8907 ;
  assign n8916 = ~n8914 & n8915 ;
  assign n8917 = ~n8912 & n8916 ;
  assign n8918 = ~n8860 & ~n8875 ;
  assign n8919 = n8854 & n8884 ;
  assign n8920 = n8918 & n8919 ;
  assign n8887 = ~n8854 & n8884 ;
  assign n8921 = n8875 & n8887 ;
  assign n8922 = ~n8920 & ~n8921 ;
  assign n8923 = ~n8869 & ~n8922 ;
  assign n8924 = ~n8898 & ~n8918 ;
  assign n8925 = ~n8885 & n8908 ;
  assign n8926 = n8924 & n8925 ;
  assign n8894 = ~n8875 & ~n8884 ;
  assign n8927 = n8861 & n8894 ;
  assign n8888 = n8860 & ~n8875 ;
  assign n8889 = n8887 & n8888 ;
  assign n8928 = ~n8889 & n8907 ;
  assign n8929 = ~n8927 & n8928 ;
  assign n8930 = ~n8926 & n8929 ;
  assign n8931 = ~n8923 & n8930 ;
  assign n8932 = ~n8917 & ~n8931 ;
  assign n8892 = n8875 & n8891 ;
  assign n8893 = ~n8889 & ~n8892 ;
  assign n8895 = n8854 & n8894 ;
  assign n8896 = n8893 & ~n8895 ;
  assign n8897 = n8869 & ~n8896 ;
  assign n8876 = ~n8869 & n8875 ;
  assign n8877 = ~n8863 & n8876 ;
  assign n8886 = n8878 & n8885 ;
  assign n8933 = ~n8877 & ~n8886 ;
  assign n8934 = ~n8897 & n8933 ;
  assign n8935 = ~n8932 & n8934 ;
  assign n8936 = ~\u2_L11_reg[22]/NET0131  & ~n8935 ;
  assign n8937 = \u2_L11_reg[22]/NET0131  & n8935 ;
  assign n8938 = ~n8936 & ~n8937 ;
  assign n8939 = decrypt_pad & ~\u2_uk_K_r11_reg[13]/NET0131  ;
  assign n8940 = ~decrypt_pad & ~\u2_uk_K_r11_reg[18]/NET0131  ;
  assign n8941 = ~n8939 & ~n8940 ;
  assign n8942 = \u2_R11_reg[3]/NET0131  & ~n8941 ;
  assign n8943 = ~\u2_R11_reg[3]/NET0131  & n8941 ;
  assign n8944 = ~n8942 & ~n8943 ;
  assign n8983 = decrypt_pad & ~\u2_uk_K_r11_reg[48]/NET0131  ;
  assign n8984 = ~decrypt_pad & ~\u2_uk_K_r11_reg[53]/P0001  ;
  assign n8985 = ~n8983 & ~n8984 ;
  assign n8986 = \u2_R11_reg[4]/NET0131  & ~n8985 ;
  assign n8987 = ~\u2_R11_reg[4]/NET0131  & n8985 ;
  assign n8988 = ~n8986 & ~n8987 ;
  assign n8958 = decrypt_pad & ~\u2_uk_K_r11_reg[4]/NET0131  ;
  assign n8959 = ~decrypt_pad & ~\u2_uk_K_r11_reg[41]/NET0131  ;
  assign n8960 = ~n8958 & ~n8959 ;
  assign n8961 = \u2_R11_reg[2]/NET0131  & ~n8960 ;
  assign n8962 = ~\u2_R11_reg[2]/NET0131  & n8960 ;
  assign n8963 = ~n8961 & ~n8962 ;
  assign n8952 = decrypt_pad & ~\u2_uk_K_r11_reg[19]/NET0131  ;
  assign n8953 = ~decrypt_pad & ~\u2_uk_K_r11_reg[24]/NET0131  ;
  assign n8954 = ~n8952 & ~n8953 ;
  assign n8955 = \u2_R11_reg[5]/NET0131  & ~n8954 ;
  assign n8956 = ~\u2_R11_reg[5]/NET0131  & n8954 ;
  assign n8957 = ~n8955 & ~n8956 ;
  assign n8945 = decrypt_pad & ~\u2_uk_K_r11_reg[46]/NET0131  ;
  assign n8946 = ~decrypt_pad & ~\u2_uk_K_r11_reg[26]/NET0131  ;
  assign n8947 = ~n8945 & ~n8946 ;
  assign n8948 = \u2_R11_reg[1]/NET0131  & ~n8947 ;
  assign n8949 = ~\u2_R11_reg[1]/NET0131  & n8947 ;
  assign n8950 = ~n8948 & ~n8949 ;
  assign n8967 = decrypt_pad & ~\u2_uk_K_r11_reg[25]/NET0131  ;
  assign n8968 = ~decrypt_pad & ~\u2_uk_K_r11_reg[5]/NET0131  ;
  assign n8969 = ~n8967 & ~n8968 ;
  assign n8970 = \u2_R11_reg[32]/NET0131  & ~n8969 ;
  assign n8971 = ~\u2_R11_reg[32]/NET0131  & n8969 ;
  assign n8972 = ~n8970 & ~n8971 ;
  assign n9014 = ~n8950 & n8972 ;
  assign n9015 = ~n8957 & n9014 ;
  assign n9016 = n8963 & n9015 ;
  assign n8978 = ~n8950 & n8957 ;
  assign n8995 = ~n8963 & ~n8972 ;
  assign n9017 = ~n8978 & n8995 ;
  assign n9018 = ~n9016 & ~n9017 ;
  assign n9019 = ~n8988 & ~n9018 ;
  assign n8993 = n8957 & ~n8972 ;
  assign n9020 = ~n8950 & n8993 ;
  assign n9021 = n8963 & n9020 ;
  assign n8999 = n8950 & n8963 ;
  assign n9012 = n8957 & n8999 ;
  assign n9013 = n8972 & n9012 ;
  assign n8964 = ~n8957 & ~n8963 ;
  assign n9022 = n8950 & n8964 ;
  assign n9023 = ~n9013 & ~n9022 ;
  assign n9024 = ~n9021 & n9023 ;
  assign n9025 = ~n9019 & n9024 ;
  assign n9026 = ~n8944 & ~n9025 ;
  assign n8979 = ~n8957 & ~n8972 ;
  assign n8980 = n8963 & n8979 ;
  assign n8981 = ~n8978 & ~n8980 ;
  assign n8982 = n8944 & ~n8981 ;
  assign n8951 = ~n8944 & n8950 ;
  assign n8965 = ~n8950 & n8964 ;
  assign n8966 = ~n8951 & ~n8965 ;
  assign n8973 = ~n8966 & n8972 ;
  assign n8974 = n8944 & ~n8963 ;
  assign n8975 = n8950 & ~n8974 ;
  assign n8976 = ~n8964 & ~n8972 ;
  assign n8977 = ~n8975 & n8976 ;
  assign n8989 = ~n8977 & n8988 ;
  assign n8990 = ~n8973 & n8989 ;
  assign n8991 = ~n8982 & n8990 ;
  assign n9000 = ~n8957 & n8999 ;
  assign n9001 = n8972 & n9000 ;
  assign n9002 = n8957 & n8972 ;
  assign n9003 = ~n8963 & n9002 ;
  assign n9004 = ~n9001 & ~n9003 ;
  assign n9005 = n8944 & ~n9004 ;
  assign n8992 = n8944 & n8963 ;
  assign n8994 = n8992 & n8993 ;
  assign n8996 = ~n8957 & n8995 ;
  assign n8997 = ~n8994 & ~n8996 ;
  assign n8998 = n8950 & ~n8997 ;
  assign n9006 = ~n8963 & n8972 ;
  assign n9007 = n8978 & n9006 ;
  assign n9008 = ~n8988 & ~n9007 ;
  assign n9009 = ~n8998 & n9008 ;
  assign n9010 = ~n9005 & n9009 ;
  assign n9011 = ~n8991 & ~n9010 ;
  assign n9027 = n8974 & n9014 ;
  assign n9028 = ~n8950 & n8979 ;
  assign n9029 = n8992 & n9028 ;
  assign n9030 = ~n9027 & ~n9029 ;
  assign n9031 = ~n9011 & n9030 ;
  assign n9032 = ~n9026 & n9031 ;
  assign n9033 = ~\u2_L11_reg[31]/NET0131  & ~n9032 ;
  assign n9034 = \u2_L11_reg[31]/NET0131  & n9032 ;
  assign n9035 = ~n9033 & ~n9034 ;
  assign n9042 = decrypt_pad & ~\u2_uk_K_r11_reg[44]/NET0131  ;
  assign n9043 = ~decrypt_pad & ~\u2_uk_K_r11_reg[22]/NET0131  ;
  assign n9044 = ~n9042 & ~n9043 ;
  assign n9045 = \u2_R11_reg[23]/NET0131  & ~n9044 ;
  assign n9046 = ~\u2_R11_reg[23]/NET0131  & n9044 ;
  assign n9047 = ~n9045 & ~n9046 ;
  assign n9048 = decrypt_pad & ~\u2_uk_K_r11_reg[0]/NET0131  ;
  assign n9049 = ~decrypt_pad & ~\u2_uk_K_r11_reg[9]/NET0131  ;
  assign n9050 = ~n9048 & ~n9049 ;
  assign n9051 = \u2_R11_reg[22]/NET0131  & ~n9050 ;
  assign n9052 = ~\u2_R11_reg[22]/NET0131  & n9050 ;
  assign n9053 = ~n9051 & ~n9052 ;
  assign n9055 = decrypt_pad & ~\u2_uk_K_r11_reg[49]/NET0131  ;
  assign n9056 = ~decrypt_pad & ~\u2_uk_K_r11_reg[31]/NET0131  ;
  assign n9057 = ~n9055 & ~n9056 ;
  assign n9058 = \u2_R11_reg[20]/NET0131  & ~n9057 ;
  assign n9059 = ~\u2_R11_reg[20]/NET0131  & n9057 ;
  assign n9060 = ~n9058 & ~n9059 ;
  assign n9062 = decrypt_pad & ~\u2_uk_K_r11_reg[9]/NET0131  ;
  assign n9063 = ~decrypt_pad & ~\u2_uk_K_r11_reg[42]/NET0131  ;
  assign n9064 = ~n9062 & ~n9063 ;
  assign n9065 = \u2_R11_reg[21]/NET0131  & ~n9064 ;
  assign n9066 = ~\u2_R11_reg[21]/NET0131  & n9064 ;
  assign n9067 = ~n9065 & ~n9066 ;
  assign n9068 = ~n9060 & n9067 ;
  assign n9074 = decrypt_pad & ~\u2_uk_K_r11_reg[38]/NET0131  ;
  assign n9075 = ~decrypt_pad & ~\u2_uk_K_r11_reg[43]/NET0131  ;
  assign n9076 = ~n9074 & ~n9075 ;
  assign n9077 = \u2_R11_reg[25]/NET0131  & ~n9076 ;
  assign n9078 = ~\u2_R11_reg[25]/NET0131  & n9076 ;
  assign n9079 = ~n9077 & ~n9078 ;
  assign n9105 = n9060 & n9079 ;
  assign n9117 = ~n9068 & ~n9105 ;
  assign n9118 = n9053 & ~n9117 ;
  assign n9119 = n9067 & n9079 ;
  assign n9120 = ~n9060 & n9119 ;
  assign n9083 = n9060 & ~n9067 ;
  assign n9090 = n9079 & n9083 ;
  assign n9121 = ~n9053 & ~n9090 ;
  assign n9122 = ~n9120 & n9121 ;
  assign n9123 = ~n9118 & ~n9122 ;
  assign n9124 = ~n9047 & ~n9123 ;
  assign n9036 = decrypt_pad & ~\u2_uk_K_r11_reg[15]/NET0131  ;
  assign n9037 = ~decrypt_pad & ~\u2_uk_K_r11_reg[52]/NET0131  ;
  assign n9038 = ~n9036 & ~n9037 ;
  assign n9039 = \u2_R11_reg[24]/NET0131  & ~n9038 ;
  assign n9040 = ~\u2_R11_reg[24]/NET0131  & n9038 ;
  assign n9041 = ~n9039 & ~n9040 ;
  assign n9080 = n9060 & ~n9079 ;
  assign n9111 = ~n9067 & n9080 ;
  assign n9112 = ~n9053 & n9111 ;
  assign n9113 = n9067 & n9105 ;
  assign n9069 = n9053 & n9068 ;
  assign n9114 = n9047 & ~n9069 ;
  assign n9115 = ~n9113 & n9114 ;
  assign n9116 = ~n9112 & n9115 ;
  assign n9125 = n9041 & ~n9116 ;
  assign n9126 = ~n9124 & n9125 ;
  assign n9091 = n9053 & n9090 ;
  assign n9070 = ~n9053 & n9067 ;
  assign n9071 = n9060 & n9070 ;
  assign n9086 = n9071 & ~n9079 ;
  assign n9087 = ~n9060 & n9079 ;
  assign n9088 = ~n9067 & n9087 ;
  assign n9089 = n9047 & n9088 ;
  assign n9094 = ~n9086 & ~n9089 ;
  assign n9095 = ~n9091 & n9094 ;
  assign n9072 = ~n9069 & ~n9071 ;
  assign n9073 = ~n9047 & ~n9072 ;
  assign n9084 = n9047 & n9053 ;
  assign n9085 = n9083 & n9084 ;
  assign n9054 = n9047 & ~n9053 ;
  assign n9061 = n9054 & ~n9060 ;
  assign n9081 = ~n9047 & ~n9053 ;
  assign n9082 = n9080 & n9081 ;
  assign n9092 = ~n9061 & ~n9082 ;
  assign n9093 = ~n9085 & n9092 ;
  assign n9096 = ~n9073 & n9093 ;
  assign n9097 = n9095 & n9096 ;
  assign n9098 = ~n9041 & ~n9097 ;
  assign n9099 = n9067 & n9080 ;
  assign n9100 = ~n9060 & ~n9079 ;
  assign n9101 = ~n9067 & n9100 ;
  assign n9102 = ~n9099 & ~n9101 ;
  assign n9103 = n9081 & ~n9102 ;
  assign n9104 = ~n9053 & ~n9100 ;
  assign n9106 = ~n9070 & ~n9105 ;
  assign n9107 = ~n9104 & ~n9106 ;
  assign n9108 = ~n9053 & n9088 ;
  assign n9109 = ~n9107 & ~n9108 ;
  assign n9110 = n9047 & ~n9109 ;
  assign n9127 = ~n9103 & ~n9110 ;
  assign n9128 = ~n9098 & n9127 ;
  assign n9129 = ~n9126 & n9128 ;
  assign n9130 = \u2_L11_reg[11]/NET0131  & ~n9129 ;
  assign n9131 = ~\u2_L11_reg[11]/NET0131  & n9129 ;
  assign n9132 = ~n9130 & ~n9131 ;
  assign n9133 = decrypt_pad & ~\u2_uk_K_r11_reg[34]/NET0131  ;
  assign n9134 = ~decrypt_pad & ~\u2_uk_K_r11_reg[39]/NET0131  ;
  assign n9135 = ~n9133 & ~n9134 ;
  assign n9136 = \u2_R11_reg[14]/NET0131  & ~n9135 ;
  assign n9137 = ~\u2_R11_reg[14]/NET0131  & n9135 ;
  assign n9138 = ~n9136 & ~n9137 ;
  assign n9139 = decrypt_pad & ~\u2_uk_K_r11_reg[10]/NET0131  ;
  assign n9140 = ~decrypt_pad & ~\u2_uk_K_r11_reg[47]/NET0131  ;
  assign n9141 = ~n9139 & ~n9140 ;
  assign n9142 = \u2_R11_reg[15]/NET0131  & ~n9141 ;
  assign n9143 = ~\u2_R11_reg[15]/NET0131  & n9141 ;
  assign n9144 = ~n9142 & ~n9143 ;
  assign n9145 = n9138 & n9144 ;
  assign n9146 = decrypt_pad & ~\u2_uk_K_r11_reg[33]/NET0131  ;
  assign n9147 = ~decrypt_pad & ~\u2_uk_K_r11_reg[13]/NET0131  ;
  assign n9148 = ~n9146 & ~n9147 ;
  assign n9149 = \u2_R11_reg[13]/NET0131  & ~n9148 ;
  assign n9150 = ~\u2_R11_reg[13]/NET0131  & n9148 ;
  assign n9151 = ~n9149 & ~n9150 ;
  assign n9152 = n9145 & n9151 ;
  assign n9153 = decrypt_pad & ~\u2_uk_K_r11_reg[39]/NET0131  ;
  assign n9154 = ~decrypt_pad & ~\u2_uk_K_r11_reg[19]/NET0131  ;
  assign n9155 = ~n9153 & ~n9154 ;
  assign n9156 = \u2_R11_reg[12]/NET0131  & ~n9155 ;
  assign n9157 = ~\u2_R11_reg[12]/NET0131  & n9155 ;
  assign n9158 = ~n9156 & ~n9157 ;
  assign n9159 = n9152 & ~n9158 ;
  assign n9171 = decrypt_pad & ~\u2_uk_K_r11_reg[18]/NET0131  ;
  assign n9172 = ~decrypt_pad & ~\u2_uk_K_r11_reg[55]/NET0131  ;
  assign n9173 = ~n9171 & ~n9172 ;
  assign n9174 = \u2_R11_reg[16]/NET0131  & ~n9173 ;
  assign n9175 = ~\u2_R11_reg[16]/NET0131  & n9173 ;
  assign n9176 = ~n9174 & ~n9175 ;
  assign n9160 = decrypt_pad & ~\u2_uk_K_r11_reg[55]/NET0131  ;
  assign n9161 = ~decrypt_pad & ~\u2_uk_K_r11_reg[3]/NET0131  ;
  assign n9162 = ~n9160 & ~n9161 ;
  assign n9163 = \u2_R11_reg[17]/NET0131  & ~n9162 ;
  assign n9164 = ~\u2_R11_reg[17]/NET0131  & n9162 ;
  assign n9165 = ~n9163 & ~n9164 ;
  assign n9180 = ~n9151 & ~n9165 ;
  assign n9181 = ~n9138 & ~n9158 ;
  assign n9182 = n9180 & n9181 ;
  assign n9191 = ~n9176 & ~n9182 ;
  assign n9192 = ~n9159 & n9191 ;
  assign n9177 = n9151 & ~n9158 ;
  assign n9178 = ~n9165 & n9177 ;
  assign n9179 = n9138 & n9178 ;
  assign n9188 = ~n9151 & n9158 ;
  assign n9189 = ~n9138 & n9188 ;
  assign n9190 = n9165 & n9189 ;
  assign n9193 = ~n9179 & ~n9190 ;
  assign n9194 = n9192 & n9193 ;
  assign n9166 = n9158 & ~n9165 ;
  assign n9167 = n9138 & n9166 ;
  assign n9168 = ~n9151 & n9165 ;
  assign n9169 = ~n9167 & ~n9168 ;
  assign n9170 = ~n9144 & ~n9169 ;
  assign n9183 = ~n9158 & n9180 ;
  assign n9184 = n9158 & n9165 ;
  assign n9185 = n9151 & n9184 ;
  assign n9186 = ~n9183 & ~n9185 ;
  assign n9187 = n9144 & ~n9186 ;
  assign n9195 = ~n9170 & ~n9187 ;
  assign n9196 = n9194 & n9195 ;
  assign n9202 = ~n9177 & ~n9188 ;
  assign n9203 = ~n9138 & ~n9202 ;
  assign n9204 = n9138 & ~n9151 ;
  assign n9205 = ~n9158 & n9204 ;
  assign n9206 = ~n9165 & n9205 ;
  assign n9207 = ~n9203 & ~n9206 ;
  assign n9208 = ~n9144 & ~n9207 ;
  assign n9199 = ~n9158 & n9165 ;
  assign n9209 = n9151 & n9199 ;
  assign n9210 = ~n9138 & n9209 ;
  assign n9211 = n9138 & n9185 ;
  assign n9212 = ~n9210 & ~n9211 ;
  assign n9200 = n9144 & n9199 ;
  assign n9201 = ~n9151 & n9200 ;
  assign n9197 = n9151 & n9166 ;
  assign n9198 = n9144 & n9197 ;
  assign n9213 = n9176 & ~n9198 ;
  assign n9214 = ~n9201 & n9213 ;
  assign n9215 = n9212 & n9214 ;
  assign n9216 = ~n9208 & n9215 ;
  assign n9217 = ~n9196 & ~n9216 ;
  assign n9224 = ~n9138 & n9198 ;
  assign n9218 = ~n9138 & ~n9144 ;
  assign n9219 = n9165 & n9218 ;
  assign n9220 = n9177 & n9219 ;
  assign n9221 = n9166 & n9204 ;
  assign n9222 = ~n9182 & ~n9221 ;
  assign n9223 = n9144 & ~n9222 ;
  assign n9225 = ~n9220 & ~n9223 ;
  assign n9226 = ~n9224 & n9225 ;
  assign n9227 = ~n9217 & n9226 ;
  assign n9228 = ~\u2_L11_reg[20]/NET0131  & ~n9227 ;
  assign n9229 = \u2_L11_reg[20]/NET0131  & n9227 ;
  assign n9230 = ~n9228 & ~n9229 ;
  assign n9284 = decrypt_pad & ~\u2_uk_K_r11_reg[42]/NET0131  ;
  assign n9285 = ~decrypt_pad & ~\u2_uk_K_r11_reg[51]/NET0131  ;
  assign n9286 = ~n9284 & ~n9285 ;
  assign n9287 = \u2_R11_reg[32]/NET0131  & ~n9286 ;
  assign n9288 = ~\u2_R11_reg[32]/NET0131  & n9286 ;
  assign n9289 = ~n9287 & ~n9288 ;
  assign n9261 = decrypt_pad & ~\u2_uk_K_r11_reg[36]/NET0131  ;
  assign n9262 = ~decrypt_pad & ~\u2_uk_K_r11_reg[14]/NET0131  ;
  assign n9263 = ~n9261 & ~n9262 ;
  assign n9264 = \u2_R11_reg[31]/P0001  & ~n9263 ;
  assign n9265 = ~\u2_R11_reg[31]/P0001  & n9263 ;
  assign n9266 = ~n9264 & ~n9265 ;
  assign n9237 = decrypt_pad & ~\u2_uk_K_r11_reg[23]/NET0131  ;
  assign n9238 = ~decrypt_pad & ~\u2_uk_K_r11_reg[1]/NET0131  ;
  assign n9239 = ~n9237 & ~n9238 ;
  assign n9240 = \u2_R11_reg[29]/NET0131  & ~n9239 ;
  assign n9241 = ~\u2_R11_reg[29]/NET0131  & n9239 ;
  assign n9242 = ~n9240 & ~n9241 ;
  assign n9244 = decrypt_pad & ~\u2_uk_K_r11_reg[52]/NET0131  ;
  assign n9245 = ~decrypt_pad & ~\u2_uk_K_r11_reg[2]/NET0131  ;
  assign n9246 = ~n9244 & ~n9245 ;
  assign n9247 = \u2_R11_reg[30]/NET0131  & ~n9246 ;
  assign n9248 = ~\u2_R11_reg[30]/NET0131  & n9246 ;
  assign n9249 = ~n9247 & ~n9248 ;
  assign n9251 = decrypt_pad & ~\u2_uk_K_r11_reg[51]/NET0131  ;
  assign n9252 = ~decrypt_pad & ~\u2_uk_K_r11_reg[29]/NET0131  ;
  assign n9253 = ~n9251 & ~n9252 ;
  assign n9254 = \u2_R11_reg[28]/NET0131  & ~n9253 ;
  assign n9255 = ~\u2_R11_reg[28]/NET0131  & n9253 ;
  assign n9256 = ~n9254 & ~n9255 ;
  assign n9291 = ~n9249 & ~n9256 ;
  assign n9292 = ~n9242 & n9291 ;
  assign n9293 = ~n9266 & ~n9292 ;
  assign n9231 = decrypt_pad & ~\u2_uk_K_r11_reg[8]/NET0131  ;
  assign n9232 = ~decrypt_pad & ~\u2_uk_K_r11_reg[45]/NET0131  ;
  assign n9233 = ~n9231 & ~n9232 ;
  assign n9234 = \u2_R11_reg[1]/NET0131  & ~n9233 ;
  assign n9235 = ~\u2_R11_reg[1]/NET0131  & n9233 ;
  assign n9236 = ~n9234 & ~n9235 ;
  assign n9271 = ~n9249 & n9256 ;
  assign n9272 = ~n9236 & n9271 ;
  assign n9273 = n9242 & n9272 ;
  assign n9294 = ~n9236 & n9242 ;
  assign n9295 = ~n9271 & ~n9294 ;
  assign n9296 = ~n9273 & ~n9295 ;
  assign n9297 = n9266 & ~n9296 ;
  assign n9298 = ~n9293 & ~n9297 ;
  assign n9258 = n9236 & ~n9256 ;
  assign n9299 = n9242 & n9258 ;
  assign n9300 = n9249 & n9299 ;
  assign n9301 = ~n9298 & ~n9300 ;
  assign n9302 = n9289 & ~n9301 ;
  assign n9243 = ~n9236 & ~n9242 ;
  assign n9250 = n9243 & n9249 ;
  assign n9257 = n9250 & n9256 ;
  assign n9259 = ~n9242 & n9258 ;
  assign n9260 = ~n9257 & ~n9259 ;
  assign n9267 = ~n9260 & n9266 ;
  assign n9268 = n9242 & n9256 ;
  assign n9269 = n9249 & n9268 ;
  assign n9270 = n9236 & n9269 ;
  assign n9274 = ~n9266 & n9271 ;
  assign n9280 = ~n9270 & ~n9274 ;
  assign n9276 = n9249 & ~n9256 ;
  assign n9277 = ~n9236 & ~n9276 ;
  assign n9275 = n9236 & ~n9242 ;
  assign n9278 = ~n9266 & ~n9275 ;
  assign n9279 = ~n9277 & n9278 ;
  assign n9281 = ~n9273 & ~n9279 ;
  assign n9282 = n9280 & n9281 ;
  assign n9283 = ~n9267 & n9282 ;
  assign n9290 = ~n9283 & ~n9289 ;
  assign n9304 = n9276 & n9294 ;
  assign n9305 = ~n9236 & n9291 ;
  assign n9306 = ~n9242 & n9305 ;
  assign n9307 = ~n9304 & ~n9306 ;
  assign n9303 = n9249 & n9259 ;
  assign n9308 = n9271 & n9275 ;
  assign n9309 = ~n9303 & ~n9308 ;
  assign n9310 = n9307 & n9309 ;
  assign n9311 = n9266 & ~n9310 ;
  assign n9312 = n9274 & n9294 ;
  assign n9314 = ~n9242 & n9256 ;
  assign n9313 = n9249 & ~n9266 ;
  assign n9315 = n9289 & n9313 ;
  assign n9316 = n9314 & n9315 ;
  assign n9317 = ~n9312 & ~n9316 ;
  assign n9318 = ~n9311 & n9317 ;
  assign n9319 = ~n9290 & n9318 ;
  assign n9320 = ~n9302 & n9319 ;
  assign n9321 = \u2_L11_reg[5]/NET0131  & ~n9320 ;
  assign n9322 = ~\u2_L11_reg[5]/NET0131  & n9320 ;
  assign n9323 = ~n9321 & ~n9322 ;
  assign n9329 = ~n9138 & n9151 ;
  assign n9341 = n9166 & ~n9329 ;
  assign n9342 = ~n9210 & ~n9341 ;
  assign n9343 = ~n9144 & ~n9342 ;
  assign n9337 = n9199 & n9204 ;
  assign n9338 = ~n9211 & ~n9337 ;
  assign n9339 = ~n9178 & ~n9190 ;
  assign n9340 = n9144 & ~n9339 ;
  assign n9344 = n9338 & ~n9340 ;
  assign n9345 = ~n9343 & n9344 ;
  assign n9346 = n9176 & ~n9345 ;
  assign n9327 = ~n9180 & ~n9204 ;
  assign n9328 = n9144 & ~n9327 ;
  assign n9330 = ~n9219 & ~n9329 ;
  assign n9331 = ~n9328 & n9330 ;
  assign n9332 = n9158 & ~n9331 ;
  assign n9326 = ~n9145 & n9183 ;
  assign n9324 = ~n9138 & n9144 ;
  assign n9325 = n9199 & n9324 ;
  assign n9333 = ~n9179 & ~n9325 ;
  assign n9334 = ~n9326 & n9333 ;
  assign n9335 = ~n9332 & n9334 ;
  assign n9336 = ~n9176 & ~n9335 ;
  assign n9347 = ~n9182 & n9338 ;
  assign n9348 = ~n9144 & ~n9347 ;
  assign n9349 = ~n9159 & ~n9224 ;
  assign n9350 = ~n9348 & n9349 ;
  assign n9351 = ~n9336 & n9350 ;
  assign n9352 = ~n9346 & n9351 ;
  assign n9353 = ~\u2_L11_reg[10]/NET0131  & ~n9352 ;
  assign n9354 = \u2_L11_reg[10]/NET0131  & n9352 ;
  assign n9355 = ~n9353 & ~n9354 ;
  assign n9356 = ~n8869 & n8889 ;
  assign n9364 = n8907 & ~n8920 ;
  assign n9365 = ~n8892 & n9364 ;
  assign n9366 = ~n9356 & n9365 ;
  assign n9357 = n8854 & n8875 ;
  assign n9358 = ~n8927 & ~n9357 ;
  assign n9359 = n8869 & ~n9358 ;
  assign n9360 = n8860 & ~n8884 ;
  assign n9361 = n8854 & n9360 ;
  assign n9362 = ~n8921 & ~n9361 ;
  assign n9363 = ~n8898 & ~n9362 ;
  assign n9367 = ~n9359 & ~n9363 ;
  assign n9368 = n9366 & n9367 ;
  assign n9374 = n8875 & n8890 ;
  assign n9375 = ~n8895 & ~n9374 ;
  assign n9376 = ~n8860 & ~n9375 ;
  assign n9369 = ~n8890 & ~n8919 ;
  assign n9370 = n8888 & ~n9369 ;
  assign n9371 = n8860 & n8900 ;
  assign n9380 = ~n8907 & ~n9371 ;
  assign n9381 = ~n9370 & n9380 ;
  assign n9372 = ~n8878 & ~n8898 ;
  assign n9373 = n8887 & ~n9372 ;
  assign n9377 = n8875 & n8884 ;
  assign n9378 = ~n8894 & ~n9377 ;
  assign n9379 = ~n8869 & ~n9378 ;
  assign n9382 = ~n9373 & ~n9379 ;
  assign n9383 = n9381 & n9382 ;
  assign n9384 = ~n9376 & n9383 ;
  assign n9385 = ~n9368 & ~n9384 ;
  assign n9386 = \u2_L11_reg[12]/NET0131  & n9385 ;
  assign n9387 = ~\u2_L11_reg[12]/NET0131  & ~n9385 ;
  assign n9388 = ~n9386 & ~n9387 ;
  assign n9389 = decrypt_pad & ~\u2_uk_K_r11_reg[43]/NET0131  ;
  assign n9390 = ~decrypt_pad & ~\u2_uk_K_r11_reg[21]/NET0131  ;
  assign n9391 = ~n9389 & ~n9390 ;
  assign n9392 = \u2_R11_reg[19]/NET0131  & ~n9391 ;
  assign n9393 = ~\u2_R11_reg[19]/NET0131  & n9391 ;
  assign n9394 = ~n9392 & ~n9393 ;
  assign n9395 = decrypt_pad & ~\u2_uk_K_r11_reg[1]/NET0131  ;
  assign n9396 = ~decrypt_pad & ~\u2_uk_K_r11_reg[38]/NET0131  ;
  assign n9397 = ~n9395 & ~n9396 ;
  assign n9398 = \u2_R11_reg[18]/NET0131  & ~n9397 ;
  assign n9399 = ~\u2_R11_reg[18]/NET0131  & n9397 ;
  assign n9400 = ~n9398 & ~n9399 ;
  assign n9401 = decrypt_pad & ~\u2_uk_K_r11_reg[7]/NET0131  ;
  assign n9402 = ~decrypt_pad & ~\u2_uk_K_r11_reg[16]/NET0131  ;
  assign n9403 = ~n9401 & ~n9402 ;
  assign n9404 = \u2_R11_reg[17]/NET0131  & ~n9403 ;
  assign n9405 = ~\u2_R11_reg[17]/NET0131  & n9403 ;
  assign n9406 = ~n9404 & ~n9405 ;
  assign n9408 = decrypt_pad & ~\u2_uk_K_r11_reg[16]/NET0131  ;
  assign n9409 = ~decrypt_pad & ~\u2_uk_K_r11_reg[49]/NET0131  ;
  assign n9410 = ~n9408 & ~n9409 ;
  assign n9411 = \u2_R11_reg[16]/NET0131  & ~n9410 ;
  assign n9412 = ~\u2_R11_reg[16]/NET0131  & n9410 ;
  assign n9413 = ~n9411 & ~n9412 ;
  assign n9414 = decrypt_pad & ~\u2_uk_K_r11_reg[28]/NET0131  ;
  assign n9415 = ~decrypt_pad & ~\u2_uk_K_r11_reg[37]/NET0131  ;
  assign n9416 = ~n9414 & ~n9415 ;
  assign n9417 = \u2_R11_reg[21]/NET0131  & ~n9416 ;
  assign n9418 = ~\u2_R11_reg[21]/NET0131  & n9416 ;
  assign n9419 = ~n9417 & ~n9418 ;
  assign n9424 = n9413 & ~n9419 ;
  assign n9425 = ~n9406 & n9424 ;
  assign n9426 = ~n9400 & n9425 ;
  assign n9427 = ~n9413 & n9419 ;
  assign n9428 = ~n9406 & n9427 ;
  assign n9407 = ~n9400 & n9406 ;
  assign n9420 = n9413 & n9419 ;
  assign n9421 = n9407 & n9420 ;
  assign n9422 = n9406 & ~n9419 ;
  assign n9423 = n9400 & n9422 ;
  assign n9429 = ~n9421 & ~n9423 ;
  assign n9430 = ~n9428 & n9429 ;
  assign n9431 = ~n9426 & n9430 ;
  assign n9432 = ~n9394 & ~n9431 ;
  assign n9437 = n9400 & n9413 ;
  assign n9438 = n9419 & n9437 ;
  assign n9433 = ~n9413 & ~n9419 ;
  assign n9435 = ~n9406 & n9433 ;
  assign n9436 = n9407 & ~n9413 ;
  assign n9439 = ~n9435 & ~n9436 ;
  assign n9440 = ~n9438 & n9439 ;
  assign n9441 = n9394 & ~n9440 ;
  assign n9434 = n9407 & n9433 ;
  assign n9442 = n9400 & ~n9406 ;
  assign n9443 = n9420 & n9442 ;
  assign n9444 = ~n9434 & ~n9443 ;
  assign n9445 = ~n9441 & n9444 ;
  assign n9446 = ~n9432 & n9445 ;
  assign n9447 = decrypt_pad & ~\u2_uk_K_r11_reg[31]/NET0131  ;
  assign n9448 = ~decrypt_pad & ~\u2_uk_K_r11_reg[36]/NET0131  ;
  assign n9449 = ~n9447 & ~n9448 ;
  assign n9450 = \u2_R11_reg[20]/NET0131  & ~n9449 ;
  assign n9451 = ~\u2_R11_reg[20]/NET0131  & n9449 ;
  assign n9452 = ~n9450 & ~n9451 ;
  assign n9453 = ~n9446 & ~n9452 ;
  assign n9456 = ~n9400 & n9420 ;
  assign n9460 = ~n9428 & ~n9456 ;
  assign n9457 = n9413 & n9422 ;
  assign n9458 = n9400 & n9419 ;
  assign n9459 = ~n9413 & n9458 ;
  assign n9461 = ~n9457 & ~n9459 ;
  assign n9462 = n9460 & n9461 ;
  assign n9463 = n9394 & ~n9462 ;
  assign n9464 = ~n9394 & ~n9400 ;
  assign n9465 = n9406 & n9427 ;
  assign n9466 = ~n9435 & ~n9465 ;
  assign n9467 = n9464 & ~n9466 ;
  assign n9454 = ~n9407 & ~n9442 ;
  assign n9455 = n9424 & ~n9454 ;
  assign n9468 = n9394 & n9400 ;
  assign n9469 = n9420 & ~n9468 ;
  assign n9470 = n9454 & n9469 ;
  assign n9471 = ~n9455 & ~n9470 ;
  assign n9472 = ~n9467 & n9471 ;
  assign n9473 = ~n9463 & n9472 ;
  assign n9474 = n9452 & ~n9473 ;
  assign n9475 = n9406 & n9433 ;
  assign n9476 = ~n9428 & ~n9475 ;
  assign n9477 = n9400 & ~n9476 ;
  assign n9478 = ~n9394 & n9477 ;
  assign n9479 = ~n9400 & n9457 ;
  assign n9480 = n9400 & n9435 ;
  assign n9481 = ~n9479 & ~n9480 ;
  assign n9482 = n9394 & ~n9481 ;
  assign n9483 = ~n9478 & ~n9482 ;
  assign n9484 = ~n9474 & n9483 ;
  assign n9485 = ~n9453 & n9484 ;
  assign n9486 = ~\u2_L11_reg[14]/NET0131  & ~n9485 ;
  assign n9487 = \u2_L11_reg[14]/NET0131  & n9485 ;
  assign n9488 = ~n9486 & ~n9487 ;
  assign n9489 = n9242 & ~n9249 ;
  assign n9490 = ~n9236 & n9489 ;
  assign n9491 = ~n9259 & ~n9268 ;
  assign n9492 = ~n9490 & n9491 ;
  assign n9493 = n9266 & ~n9492 ;
  assign n9494 = n9243 & n9271 ;
  assign n9495 = ~n9493 & ~n9494 ;
  assign n9496 = ~n9289 & ~n9495 ;
  assign n9502 = n9275 & n9313 ;
  assign n9501 = ~n9249 & n9268 ;
  assign n9503 = ~n9304 & ~n9501 ;
  assign n9504 = ~n9502 & n9503 ;
  assign n9497 = n9249 & n9314 ;
  assign n9498 = n9236 & n9497 ;
  assign n9499 = n9243 & ~n9256 ;
  assign n9500 = n9266 & n9499 ;
  assign n9505 = ~n9498 & ~n9500 ;
  assign n9506 = n9504 & n9505 ;
  assign n9507 = n9289 & ~n9506 ;
  assign n9510 = ~n9266 & ~n9497 ;
  assign n9508 = n9258 & n9489 ;
  assign n9509 = ~n9289 & n9314 ;
  assign n9511 = ~n9508 & ~n9509 ;
  assign n9512 = n9510 & n9511 ;
  assign n9513 = n9307 & n9512 ;
  assign n9514 = n9275 & n9291 ;
  assign n9515 = n9266 & ~n9514 ;
  assign n9516 = ~n9300 & n9515 ;
  assign n9517 = ~n9513 & ~n9516 ;
  assign n9518 = ~n9507 & ~n9517 ;
  assign n9519 = ~n9496 & n9518 ;
  assign n9520 = ~\u2_L11_reg[15]/NET0131  & ~n9519 ;
  assign n9521 = \u2_L11_reg[15]/NET0131  & n9519 ;
  assign n9522 = ~n9520 & ~n9521 ;
  assign n9539 = ~n8950 & ~n8963 ;
  assign n9540 = ~n8972 & ~n9539 ;
  assign n9541 = ~n9007 & ~n9540 ;
  assign n9542 = n8944 & ~n9541 ;
  assign n9543 = ~n8944 & ~n9006 ;
  assign n9544 = ~n9540 & n9543 ;
  assign n9538 = n8972 & n9022 ;
  assign n9545 = ~n9012 & ~n9538 ;
  assign n9546 = ~n9544 & n9545 ;
  assign n9547 = ~n9542 & n9546 ;
  assign n9548 = n8988 & ~n9547 ;
  assign n9523 = n8957 & n8995 ;
  assign n9524 = ~n8980 & ~n9523 ;
  assign n9525 = n8944 & n8950 ;
  assign n9526 = ~n9524 & n9525 ;
  assign n9527 = ~n8979 & ~n9002 ;
  assign n9528 = ~n8950 & ~n9527 ;
  assign n9529 = ~n8996 & ~n9528 ;
  assign n9530 = ~n8944 & ~n9529 ;
  assign n9531 = n8950 & n9002 ;
  assign n9532 = ~n9015 & ~n9531 ;
  assign n9533 = n8944 & ~n9532 ;
  assign n9534 = ~n9001 & ~n9021 ;
  assign n9535 = ~n9533 & n9534 ;
  assign n9536 = ~n9530 & n9535 ;
  assign n9537 = ~n8988 & ~n9536 ;
  assign n9549 = ~n9526 & ~n9537 ;
  assign n9550 = ~n9548 & n9549 ;
  assign n9551 = ~\u2_L11_reg[17]/NET0131  & ~n9550 ;
  assign n9552 = \u2_L11_reg[17]/NET0131  & n9550 ;
  assign n9553 = ~n9551 & ~n9552 ;
  assign n9554 = ~n9168 & ~n9189 ;
  assign n9555 = n9176 & ~n9554 ;
  assign n9556 = n9144 & ~n9179 ;
  assign n9557 = n9338 & n9556 ;
  assign n9558 = ~n9555 & n9557 ;
  assign n9559 = n9138 & n9197 ;
  assign n9560 = ~n9144 & ~n9206 ;
  assign n9561 = ~n9559 & n9560 ;
  assign n9562 = ~n9558 & ~n9561 ;
  assign n9564 = ~n9138 & n9166 ;
  assign n9563 = n9158 & n9168 ;
  assign n9565 = ~n9144 & ~n9563 ;
  assign n9566 = ~n9564 & n9565 ;
  assign n9567 = ~n9165 & n9181 ;
  assign n9568 = n9144 & ~n9221 ;
  assign n9569 = ~n9567 & n9568 ;
  assign n9570 = ~n9566 & ~n9569 ;
  assign n9571 = n9151 & n9564 ;
  assign n9572 = ~n9176 & ~n9571 ;
  assign n9573 = n9212 & n9572 ;
  assign n9574 = ~n9570 & n9573 ;
  assign n9575 = ~n9166 & n9329 ;
  assign n9576 = ~n9209 & ~n9575 ;
  assign n9577 = ~n9144 & ~n9576 ;
  assign n9578 = n9176 & ~n9205 ;
  assign n9579 = ~n9559 & n9578 ;
  assign n9580 = ~n9577 & n9579 ;
  assign n9581 = ~n9574 & ~n9580 ;
  assign n9582 = ~n9562 & ~n9581 ;
  assign n9583 = ~\u2_L11_reg[1]/NET0131  & ~n9582 ;
  assign n9584 = \u2_L11_reg[1]/NET0131  & n9582 ;
  assign n9585 = ~n9583 & ~n9584 ;
  assign n9586 = ~n9266 & ~n9272 ;
  assign n9587 = ~n9498 & n9586 ;
  assign n9589 = n9266 & ~n9269 ;
  assign n9588 = ~n9249 & n9275 ;
  assign n9590 = ~n9299 & ~n9588 ;
  assign n9591 = n9589 & n9590 ;
  assign n9592 = ~n9587 & ~n9591 ;
  assign n9593 = n9256 & n9294 ;
  assign n9594 = ~n9499 & ~n9593 ;
  assign n9595 = n9249 & ~n9594 ;
  assign n9596 = n9289 & ~n9514 ;
  assign n9597 = ~n9595 & n9596 ;
  assign n9598 = ~n9592 & n9597 ;
  assign n9599 = n9258 & n9313 ;
  assign n9607 = ~n9289 & ~n9599 ;
  assign n9602 = ~n9256 & ~n9266 ;
  assign n9603 = n9294 & n9602 ;
  assign n9604 = n9242 & n9276 ;
  assign n9608 = ~n9603 & ~n9604 ;
  assign n9609 = n9607 & n9608 ;
  assign n9610 = ~n9257 & ~n9306 ;
  assign n9611 = n9609 & n9610 ;
  assign n9600 = ~n9497 & ~n9593 ;
  assign n9601 = n9266 & ~n9600 ;
  assign n9605 = ~n9274 & ~n9501 ;
  assign n9606 = n9236 & ~n9605 ;
  assign n9612 = ~n9601 & ~n9606 ;
  assign n9613 = n9611 & n9612 ;
  assign n9614 = ~n9598 & ~n9613 ;
  assign n9615 = n9266 & n9292 ;
  assign n9616 = n9236 & n9256 ;
  assign n9617 = ~n9266 & n9489 ;
  assign n9618 = n9616 & n9617 ;
  assign n9619 = ~n9615 & ~n9618 ;
  assign n9620 = ~n9614 & n9619 ;
  assign n9621 = ~\u2_L11_reg[21]/NET0131  & ~n9620 ;
  assign n9622 = \u2_L11_reg[21]/NET0131  & n9620 ;
  assign n9623 = ~n9621 & ~n9622 ;
  assign n9630 = decrypt_pad & ~\u2_uk_K_r11_reg[41]/NET0131  ;
  assign n9631 = ~decrypt_pad & ~\u2_uk_K_r11_reg[46]/NET0131  ;
  assign n9632 = ~n9630 & ~n9631 ;
  assign n9633 = \u2_R11_reg[5]/NET0131  & ~n9632 ;
  assign n9634 = ~\u2_R11_reg[5]/NET0131  & n9632 ;
  assign n9635 = ~n9633 & ~n9634 ;
  assign n9637 = decrypt_pad & ~\u2_uk_K_r11_reg[5]/NET0131  ;
  assign n9638 = ~decrypt_pad & ~\u2_uk_K_r11_reg[10]/NET0131  ;
  assign n9639 = ~n9637 & ~n9638 ;
  assign n9640 = \u2_R11_reg[4]/NET0131  & ~n9639 ;
  assign n9641 = ~\u2_R11_reg[4]/NET0131  & n9639 ;
  assign n9642 = ~n9640 & ~n9641 ;
  assign n9644 = decrypt_pad & ~\u2_uk_K_r11_reg[54]/NET0131  ;
  assign n9645 = ~decrypt_pad & ~\u2_uk_K_r11_reg[34]/NET0131  ;
  assign n9646 = ~n9644 & ~n9645 ;
  assign n9647 = \u2_R11_reg[9]/NET0131  & ~n9646 ;
  assign n9648 = ~\u2_R11_reg[9]/NET0131  & n9646 ;
  assign n9649 = ~n9647 & ~n9648 ;
  assign n9651 = n9642 & ~n9649 ;
  assign n9652 = ~n9635 & ~n9651 ;
  assign n9653 = n9635 & n9642 ;
  assign n9654 = ~n9649 & n9653 ;
  assign n9655 = ~n9652 & ~n9654 ;
  assign n9656 = ~n9642 & n9649 ;
  assign n9624 = decrypt_pad & ~\u2_uk_K_r11_reg[32]/NET0131  ;
  assign n9625 = ~decrypt_pad & ~\u2_uk_K_r11_reg[12]/NET0131  ;
  assign n9626 = ~n9624 & ~n9625 ;
  assign n9627 = \u2_R11_reg[6]/NET0131  & ~n9626 ;
  assign n9628 = ~\u2_R11_reg[6]/NET0131  & n9626 ;
  assign n9629 = ~n9627 & ~n9628 ;
  assign n9657 = ~n9629 & ~n9642 ;
  assign n9658 = ~n9656 & ~n9657 ;
  assign n9659 = n9655 & n9658 ;
  assign n9660 = decrypt_pad & ~\u2_uk_K_r11_reg[26]/NET0131  ;
  assign n9661 = ~decrypt_pad & ~\u2_uk_K_r11_reg[6]/NET0131  ;
  assign n9662 = ~n9660 & ~n9661 ;
  assign n9663 = \u2_R11_reg[7]/NET0131  & ~n9662 ;
  assign n9664 = ~\u2_R11_reg[7]/NET0131  & n9662 ;
  assign n9665 = ~n9663 & ~n9664 ;
  assign n9666 = ~n9659 & n9665 ;
  assign n9667 = ~n9635 & n9649 ;
  assign n9668 = ~n9658 & ~n9667 ;
  assign n9669 = n9629 & n9654 ;
  assign n9636 = n9629 & ~n9635 ;
  assign n9643 = n9636 & ~n9642 ;
  assign n9670 = ~n9643 & ~n9665 ;
  assign n9671 = ~n9669 & n9670 ;
  assign n9672 = ~n9668 & n9671 ;
  assign n9673 = ~n9666 & ~n9672 ;
  assign n9674 = n9642 & n9667 ;
  assign n9675 = ~n9665 & ~n9674 ;
  assign n9676 = ~n9629 & n9642 ;
  assign n9677 = ~n9675 & n9676 ;
  assign n9650 = n9643 & n9649 ;
  assign n9678 = decrypt_pad & ~\u2_uk_K_r11_reg[17]/NET0131  ;
  assign n9679 = ~decrypt_pad & ~\u2_uk_K_r11_reg[54]/NET0131  ;
  assign n9680 = ~n9678 & ~n9679 ;
  assign n9681 = \u2_R11_reg[8]/NET0131  & ~n9680 ;
  assign n9682 = ~\u2_R11_reg[8]/NET0131  & n9680 ;
  assign n9683 = ~n9681 & ~n9682 ;
  assign n9684 = ~n9650 & n9683 ;
  assign n9685 = ~n9677 & n9684 ;
  assign n9686 = ~n9673 & n9685 ;
  assign n9690 = n9665 & ~n9668 ;
  assign n9691 = n9642 & ~n9667 ;
  assign n9692 = ~n9636 & n9691 ;
  assign n9693 = ~n9642 & n9667 ;
  assign n9694 = ~n9692 & ~n9693 ;
  assign n9695 = n9671 & n9694 ;
  assign n9696 = ~n9690 & ~n9695 ;
  assign n9687 = n9629 & ~n9656 ;
  assign n9688 = n9652 & n9687 ;
  assign n9689 = ~n9669 & ~n9683 ;
  assign n9697 = ~n9688 & n9689 ;
  assign n9698 = ~n9696 & n9697 ;
  assign n9699 = ~n9686 & ~n9698 ;
  assign n9700 = ~\u2_L11_reg[28]/NET0131  & n9699 ;
  assign n9701 = \u2_L11_reg[28]/NET0131  & ~n9699 ;
  assign n9702 = ~n9700 & ~n9701 ;
  assign n9703 = ~n9111 & ~n9113 ;
  assign n9704 = ~n9053 & ~n9079 ;
  assign n9705 = n9067 & n9100 ;
  assign n9706 = ~n9704 & ~n9705 ;
  assign n9707 = ~n9070 & ~n9706 ;
  assign n9708 = n9703 & ~n9707 ;
  assign n9709 = n9047 & ~n9708 ;
  assign n9710 = n9053 & n9088 ;
  assign n9711 = ~n9709 & ~n9710 ;
  assign n9712 = ~n9041 & ~n9711 ;
  assign n9713 = n9053 & n9099 ;
  assign n9714 = ~n9053 & ~n9060 ;
  assign n9715 = n9067 & n9714 ;
  assign n9716 = ~n9120 & ~n9715 ;
  assign n9717 = ~n9713 & n9716 ;
  assign n9718 = n9047 & ~n9717 ;
  assign n9722 = n9053 & ~n9100 ;
  assign n9723 = ~n9105 & n9722 ;
  assign n9719 = ~n9067 & ~n9704 ;
  assign n9720 = n9047 & ~n9719 ;
  assign n9721 = ~n9053 & ~n9117 ;
  assign n9724 = ~n9720 & ~n9721 ;
  assign n9725 = ~n9723 & n9724 ;
  assign n9726 = ~n9718 & ~n9725 ;
  assign n9727 = n9041 & ~n9726 ;
  assign n9729 = ~n9713 & ~n9721 ;
  assign n9730 = ~n9041 & ~n9047 ;
  assign n9731 = ~n9729 & n9730 ;
  assign n9728 = n9054 & n9119 ;
  assign n9732 = ~n9112 & ~n9728 ;
  assign n9733 = ~n9731 & n9732 ;
  assign n9734 = ~n9727 & n9733 ;
  assign n9735 = ~n9712 & n9734 ;
  assign n9736 = \u2_L11_reg[29]/NET0131  & ~n9735 ;
  assign n9737 = ~\u2_L11_reg[29]/NET0131  & n9735 ;
  assign n9738 = ~n9736 & ~n9737 ;
  assign n9739 = n9629 & n9665 ;
  assign n9740 = n9674 & n9739 ;
  assign n9741 = n9629 & n9642 ;
  assign n9742 = ~n9667 & ~n9741 ;
  assign n9743 = n9675 & ~n9742 ;
  assign n9753 = ~n9740 & ~n9743 ;
  assign n9744 = n9635 & ~n9649 ;
  assign n9745 = ~n9693 & ~n9744 ;
  assign n9746 = ~n9629 & ~n9745 ;
  assign n9747 = n9629 & n9656 ;
  assign n9748 = n9635 & n9747 ;
  assign n9749 = ~n9629 & ~n9635 ;
  assign n9750 = n9649 & ~n9665 ;
  assign n9751 = n9749 & n9750 ;
  assign n9752 = ~n9748 & ~n9751 ;
  assign n9754 = ~n9746 & n9752 ;
  assign n9755 = n9753 & n9754 ;
  assign n9756 = ~n9683 & ~n9755 ;
  assign n9762 = ~n9635 & ~n9649 ;
  assign n9763 = ~n9687 & ~n9762 ;
  assign n9764 = ~n9691 & ~n9763 ;
  assign n9757 = ~n9629 & n9635 ;
  assign n9760 = n9642 & n9757 ;
  assign n9761 = n9649 & n9760 ;
  assign n9765 = ~n9649 & n9749 ;
  assign n9766 = n9642 & n9765 ;
  assign n9767 = ~n9761 & ~n9766 ;
  assign n9768 = ~n9764 & n9767 ;
  assign n9769 = n9683 & ~n9768 ;
  assign n9758 = ~n9636 & ~n9757 ;
  assign n9759 = n9656 & n9758 ;
  assign n9770 = ~n9665 & ~n9759 ;
  assign n9771 = ~n9769 & n9770 ;
  assign n9773 = n9629 & ~n9653 ;
  assign n9774 = ~n9652 & n9683 ;
  assign n9775 = ~n9773 & n9774 ;
  assign n9772 = n9643 & ~n9649 ;
  assign n9776 = n9665 & ~n9760 ;
  assign n9777 = ~n9772 & n9776 ;
  assign n9778 = ~n9775 & n9777 ;
  assign n9779 = ~n9771 & ~n9778 ;
  assign n9780 = ~n9756 & ~n9779 ;
  assign n9781 = \u2_L11_reg[2]/NET0131  & n9780 ;
  assign n9782 = ~\u2_L11_reg[2]/NET0131  & ~n9780 ;
  assign n9783 = ~n9781 & ~n9782 ;
  assign n9790 = ~n9197 & ~n9200 ;
  assign n9791 = ~n9209 & n9790 ;
  assign n9792 = n9138 & ~n9791 ;
  assign n9785 = n9138 & n9184 ;
  assign n9786 = n9168 & n9181 ;
  assign n9787 = ~n9785 & ~n9786 ;
  assign n9788 = ~n9144 & ~n9787 ;
  assign n9784 = ~n9138 & n9178 ;
  assign n9789 = n9144 & n9183 ;
  assign n9793 = ~n9784 & ~n9789 ;
  assign n9794 = ~n9788 & n9793 ;
  assign n9795 = ~n9792 & n9794 ;
  assign n9796 = n9176 & ~n9795 ;
  assign n9806 = ~n9189 & ~n9198 ;
  assign n9805 = n9152 & ~n9199 ;
  assign n9807 = ~n9210 & ~n9805 ;
  assign n9808 = n9806 & n9807 ;
  assign n9809 = ~n9176 & ~n9808 ;
  assign n9797 = ~n9165 & ~n9202 ;
  assign n9798 = ~n9185 & ~n9797 ;
  assign n9799 = n9218 & ~n9798 ;
  assign n9800 = n9165 & n9324 ;
  assign n9801 = ~n9202 & n9800 ;
  assign n9802 = ~n9180 & ~n9205 ;
  assign n9803 = ~n9144 & ~n9176 ;
  assign n9804 = ~n9802 & n9803 ;
  assign n9810 = ~n9801 & ~n9804 ;
  assign n9811 = ~n9799 & n9810 ;
  assign n9812 = ~n9809 & n9811 ;
  assign n9813 = ~n9796 & n9812 ;
  assign n9814 = ~\u2_L11_reg[26]/NET0131  & ~n9813 ;
  assign n9815 = \u2_L11_reg[26]/NET0131  & n9813 ;
  assign n9816 = ~n9814 & ~n9815 ;
  assign n9823 = ~n9407 & ~n9419 ;
  assign n9824 = ~n9437 & n9823 ;
  assign n9821 = n9406 & n9420 ;
  assign n9822 = ~n9406 & ~n9413 ;
  assign n9825 = ~n9821 & ~n9822 ;
  assign n9826 = ~n9824 & n9825 ;
  assign n9827 = n9394 & ~n9826 ;
  assign n9818 = ~n9406 & n9420 ;
  assign n9819 = ~n9436 & ~n9818 ;
  assign n9820 = ~n9394 & ~n9819 ;
  assign n9817 = n9407 & n9419 ;
  assign n9828 = n9422 & n9437 ;
  assign n9829 = ~n9817 & ~n9828 ;
  assign n9830 = ~n9820 & n9829 ;
  assign n9831 = ~n9827 & n9830 ;
  assign n9832 = n9452 & ~n9831 ;
  assign n9845 = n9394 & ~n9422 ;
  assign n9844 = ~n9394 & ~n9822 ;
  assign n9846 = ~n9400 & ~n9844 ;
  assign n9847 = ~n9845 & n9846 ;
  assign n9839 = ~n9394 & n9425 ;
  assign n9840 = n9394 & ~n9419 ;
  assign n9841 = n9400 & n9406 ;
  assign n9842 = ~n9413 & n9841 ;
  assign n9843 = ~n9840 & n9842 ;
  assign n9848 = ~n9839 & ~n9843 ;
  assign n9849 = ~n9847 & n9848 ;
  assign n9850 = ~n9452 & ~n9849 ;
  assign n9833 = ~n9480 & ~n9828 ;
  assign n9834 = ~n9400 & n9428 ;
  assign n9835 = n9833 & ~n9834 ;
  assign n9836 = n9394 & ~n9835 ;
  assign n9837 = ~n9394 & n9413 ;
  assign n9838 = n9442 & n9837 ;
  assign n9851 = ~n9421 & ~n9838 ;
  assign n9852 = ~n9836 & n9851 ;
  assign n9853 = ~n9850 & n9852 ;
  assign n9854 = ~n9832 & n9853 ;
  assign n9855 = ~\u2_L11_reg[25]/NET0131  & ~n9854 ;
  assign n9856 = \u2_L11_reg[25]/NET0131  & n9854 ;
  assign n9857 = ~n9855 & ~n9856 ;
  assign n9877 = ~n9053 & n9087 ;
  assign n9878 = ~n9099 & ~n9877 ;
  assign n9879 = ~n9091 & n9878 ;
  assign n9880 = n9047 & ~n9879 ;
  assign n9874 = ~n9705 & ~n9710 ;
  assign n9875 = ~n9047 & ~n9874 ;
  assign n9876 = n9081 & n9105 ;
  assign n9881 = ~n9112 & ~n9876 ;
  assign n9882 = ~n9875 & n9881 ;
  assign n9883 = ~n9880 & n9882 ;
  assign n9884 = ~n9041 & ~n9883 ;
  assign n9861 = n9047 & n9105 ;
  assign n9862 = ~n9705 & ~n9861 ;
  assign n9863 = ~n9053 & ~n9862 ;
  assign n9858 = n9070 & ~n9079 ;
  assign n9859 = ~n9714 & ~n9858 ;
  assign n9860 = ~n9047 & ~n9859 ;
  assign n9864 = n9053 & n9119 ;
  assign n9865 = ~n9860 & ~n9864 ;
  assign n9866 = ~n9863 & n9865 ;
  assign n9867 = n9041 & ~n9866 ;
  assign n9868 = ~n9101 & ~n9120 ;
  assign n9869 = ~n9099 & n9868 ;
  assign n9870 = n9084 & ~n9869 ;
  assign n9871 = n9053 & n9703 ;
  assign n9872 = ~n9047 & ~n9104 ;
  assign n9873 = ~n9871 & n9872 ;
  assign n9885 = ~n9870 & ~n9873 ;
  assign n9886 = ~n9867 & n9885 ;
  assign n9887 = ~n9884 & n9886 ;
  assign n9888 = ~\u2_L11_reg[4]/NET0131  & ~n9887 ;
  assign n9889 = \u2_L11_reg[4]/NET0131  & n9887 ;
  assign n9890 = ~n9888 & ~n9889 ;
  assign n9892 = n9636 & ~n9649 ;
  assign n9893 = n9675 & ~n9892 ;
  assign n9894 = n9665 & ~n9747 ;
  assign n9895 = ~n9765 & n9894 ;
  assign n9896 = ~n9893 & ~n9895 ;
  assign n9891 = n9657 & n9744 ;
  assign n9897 = n9683 & ~n9891 ;
  assign n9898 = n9752 & n9897 ;
  assign n9899 = ~n9896 & n9898 ;
  assign n9901 = n9656 & ~n9758 ;
  assign n9900 = ~n9642 & n9744 ;
  assign n9902 = ~n9665 & ~n9683 ;
  assign n9903 = ~n9900 & n9902 ;
  assign n9904 = ~n9766 & n9903 ;
  assign n9905 = ~n9901 & n9904 ;
  assign n9906 = ~n9899 & ~n9905 ;
  assign n9907 = ~n9669 & ~n9761 ;
  assign n9908 = ~n9906 & n9907 ;
  assign n9911 = ~n9629 & ~n9655 ;
  assign n9909 = n9687 & ~n9744 ;
  assign n9910 = n9656 & n9757 ;
  assign n9912 = n9665 & ~n9683 ;
  assign n9913 = ~n9910 & n9912 ;
  assign n9914 = ~n9909 & n9913 ;
  assign n9915 = ~n9911 & n9914 ;
  assign n9916 = ~n9908 & ~n9915 ;
  assign n9917 = ~\u2_L11_reg[13]/NET0131  & ~n9916 ;
  assign n9918 = \u2_L11_reg[13]/NET0131  & n9916 ;
  assign n9919 = ~n9917 & ~n9918 ;
  assign n9920 = ~n9090 & ~n9099 ;
  assign n9921 = n9081 & ~n9920 ;
  assign n9922 = ~n9047 & n9083 ;
  assign n9926 = n9041 & ~n9858 ;
  assign n9927 = ~n9922 & n9926 ;
  assign n9928 = ~n9108 & n9927 ;
  assign n9923 = ~n9071 & ~n9088 ;
  assign n9924 = n9047 & ~n9923 ;
  assign n9925 = n9053 & ~n9868 ;
  assign n9929 = ~n9924 & ~n9925 ;
  assign n9930 = n9928 & n9929 ;
  assign n9931 = ~n9047 & n9868 ;
  assign n9932 = n9060 & ~n9070 ;
  assign n9933 = n9047 & ~n9705 ;
  assign n9934 = ~n9932 & n9933 ;
  assign n9935 = ~n9108 & n9934 ;
  assign n9936 = ~n9931 & ~n9935 ;
  assign n9937 = n9053 & n9113 ;
  assign n9938 = ~n9041 & ~n9937 ;
  assign n9939 = ~n9936 & n9938 ;
  assign n9940 = ~n9930 & ~n9939 ;
  assign n9941 = ~n9921 & ~n9940 ;
  assign n9942 = ~\u2_L11_reg[19]/NET0131  & ~n9941 ;
  assign n9943 = \u2_L11_reg[19]/NET0131  & n9941 ;
  assign n9944 = ~n9942 & ~n9943 ;
  assign n9953 = ~n9006 & n9525 ;
  assign n9954 = n9527 & n9953 ;
  assign n9955 = n8988 & ~n9007 ;
  assign n9956 = ~n9029 & n9955 ;
  assign n9957 = ~n9954 & n9956 ;
  assign n9959 = ~n8944 & n8963 ;
  assign n9960 = n8957 & n9959 ;
  assign n9961 = ~n8951 & ~n9960 ;
  assign n9962 = n8972 & ~n9961 ;
  assign n9963 = ~n8965 & ~n8988 ;
  assign n9958 = n8979 & n9525 ;
  assign n9964 = ~n8994 & ~n9012 ;
  assign n9965 = ~n9958 & n9964 ;
  assign n9966 = n9963 & n9965 ;
  assign n9967 = ~n9962 & n9966 ;
  assign n9968 = ~n9957 & ~n9967 ;
  assign n9945 = n8950 & n8979 ;
  assign n9946 = ~n9020 & ~n9945 ;
  assign n9947 = ~n9016 & n9946 ;
  assign n9948 = n8988 & ~n9947 ;
  assign n9949 = ~n8950 & n9523 ;
  assign n9950 = ~n9538 & ~n9949 ;
  assign n9951 = ~n9948 & n9950 ;
  assign n9952 = ~n8944 & ~n9951 ;
  assign n9969 = n9531 & n9959 ;
  assign n9970 = ~n9014 & ~n9945 ;
  assign n9971 = n8974 & ~n9970 ;
  assign n9972 = ~n9969 & ~n9971 ;
  assign n9973 = ~n9952 & n9972 ;
  assign n9974 = ~n9968 & n9973 ;
  assign n9975 = \u2_L11_reg[23]/NET0131  & ~n9974 ;
  assign n9976 = ~\u2_L11_reg[23]/NET0131  & n9974 ;
  assign n9977 = ~n9975 & ~n9976 ;
  assign n9990 = ~n9305 & ~n9616 ;
  assign n9991 = n9242 & ~n9990 ;
  assign n9992 = n9266 & ~n9991 ;
  assign n9993 = ~n9299 & ~n9593 ;
  assign n9994 = n9293 & n9993 ;
  assign n9995 = ~n9992 & ~n9994 ;
  assign n9996 = ~n9257 & ~n9588 ;
  assign n9997 = ~n9300 & n9996 ;
  assign n9998 = ~n9995 & n9997 ;
  assign n9999 = n9289 & ~n9998 ;
  assign n9980 = n9266 & ~n9490 ;
  assign n9979 = n9236 & ~n9489 ;
  assign n9981 = ~n9604 & ~n9979 ;
  assign n9982 = n9980 & n9981 ;
  assign n9978 = n9313 & n9616 ;
  assign n9983 = ~n9603 & ~n9978 ;
  assign n9984 = ~n9303 & n9983 ;
  assign n9985 = ~n9982 & n9984 ;
  assign n9986 = ~n9289 & ~n9985 ;
  assign n9987 = ~n9304 & ~n9308 ;
  assign n9988 = ~n9266 & ~n9987 ;
  assign n9989 = n9250 & n9266 ;
  assign n10000 = ~n9312 & ~n9989 ;
  assign n10001 = ~n9988 & n10000 ;
  assign n10002 = ~n9986 & n10001 ;
  assign n10003 = ~n9999 & n10002 ;
  assign n10004 = ~\u2_L11_reg[27]/NET0131  & ~n10003 ;
  assign n10005 = \u2_L11_reg[27]/NET0131  & n10003 ;
  assign n10006 = ~n10004 & ~n10005 ;
  assign n10012 = n8869 & ~n9361 ;
  assign n10010 = ~n8854 & n8894 ;
  assign n10011 = ~n8860 & n9377 ;
  assign n10013 = ~n10010 & ~n10011 ;
  assign n10014 = n10012 & n10013 ;
  assign n10015 = n8918 & n9369 ;
  assign n10016 = n8888 & n8919 ;
  assign n10017 = ~n8869 & ~n9374 ;
  assign n10018 = ~n10016 & n10017 ;
  assign n10019 = ~n10015 & n10018 ;
  assign n10020 = ~n10014 & ~n10019 ;
  assign n10021 = n9357 & n9360 ;
  assign n10022 = n8907 & ~n10021 ;
  assign n10023 = ~n10020 & n10022 ;
  assign n10027 = n8854 & ~n9377 ;
  assign n10028 = n8869 & ~n9360 ;
  assign n10029 = n10027 & n10028 ;
  assign n10030 = n8862 & n9377 ;
  assign n10024 = n8885 & n9357 ;
  assign n10031 = ~n8907 & ~n10024 ;
  assign n10032 = ~n10030 & n10031 ;
  assign n10033 = ~n10029 & n10032 ;
  assign n10025 = n8854 & n8885 ;
  assign n10026 = n9379 & ~n10025 ;
  assign n10034 = n8893 & ~n10026 ;
  assign n10035 = n10033 & n10034 ;
  assign n10036 = ~n10023 & ~n10035 ;
  assign n10007 = n8876 & ~n8885 ;
  assign n10008 = n8863 & n10007 ;
  assign n10009 = n8869 & n8889 ;
  assign n10037 = ~n10008 & ~n10009 ;
  assign n10038 = ~n10036 & n10037 ;
  assign n10039 = \u2_L11_reg[32]/NET0131  & n10038 ;
  assign n10040 = ~\u2_L11_reg[32]/NET0131  & ~n10038 ;
  assign n10041 = ~n10039 & ~n10040 ;
  assign n10075 = decrypt_pad & ~\u2_uk_K_r11_reg[27]/NET0131  ;
  assign n10076 = ~decrypt_pad & ~\u2_uk_K_r11_reg[32]/NET0131  ;
  assign n10077 = ~n10075 & ~n10076 ;
  assign n10078 = \u2_R11_reg[12]/NET0131  & ~n10077 ;
  assign n10079 = ~\u2_R11_reg[12]/NET0131  & n10077 ;
  assign n10080 = ~n10078 & ~n10079 ;
  assign n10042 = decrypt_pad & ~\u2_uk_K_r11_reg[40]/NET0131  ;
  assign n10043 = ~decrypt_pad & ~\u2_uk_K_r11_reg[20]/NET0131  ;
  assign n10044 = ~n10042 & ~n10043 ;
  assign n10045 = \u2_R11_reg[13]/NET0131  & ~n10044 ;
  assign n10046 = ~\u2_R11_reg[13]/NET0131  & n10044 ;
  assign n10047 = ~n10045 & ~n10046 ;
  assign n10055 = decrypt_pad & ~\u2_uk_K_r11_reg[6]/NET0131  ;
  assign n10056 = ~decrypt_pad & ~\u2_uk_K_r11_reg[11]/NET0131  ;
  assign n10057 = ~n10055 & ~n10056 ;
  assign n10058 = \u2_R11_reg[8]/NET0131  & ~n10057 ;
  assign n10059 = ~\u2_R11_reg[8]/NET0131  & n10057 ;
  assign n10060 = ~n10058 & ~n10059 ;
  assign n10062 = ~n10047 & ~n10060 ;
  assign n10063 = n10047 & n10060 ;
  assign n10064 = ~n10062 & ~n10063 ;
  assign n10048 = decrypt_pad & ~\u2_uk_K_r11_reg[3]/NET0131  ;
  assign n10049 = ~decrypt_pad & ~\u2_uk_K_r11_reg[40]/NET0131  ;
  assign n10050 = ~n10048 & ~n10049 ;
  assign n10051 = \u2_R11_reg[9]/NET0131  & ~n10050 ;
  assign n10052 = ~\u2_R11_reg[9]/NET0131  & n10050 ;
  assign n10053 = ~n10051 & ~n10052 ;
  assign n10065 = decrypt_pad & ~\u2_uk_K_r11_reg[11]/NET0131  ;
  assign n10066 = ~decrypt_pad & ~\u2_uk_K_r11_reg[48]/NET0131  ;
  assign n10067 = ~n10065 & ~n10066 ;
  assign n10068 = \u2_R11_reg[10]/NET0131  & ~n10067 ;
  assign n10069 = ~\u2_R11_reg[10]/NET0131  & n10067 ;
  assign n10070 = ~n10068 & ~n10069 ;
  assign n10116 = ~n10053 & n10070 ;
  assign n10117 = ~n10064 & n10116 ;
  assign n10105 = n10047 & ~n10060 ;
  assign n10106 = n10053 & n10105 ;
  assign n10087 = decrypt_pad & ~\u2_uk_K_r11_reg[12]/NET0131  ;
  assign n10088 = ~decrypt_pad & ~\u2_uk_K_r11_reg[17]/NET0131  ;
  assign n10089 = ~n10087 & ~n10088 ;
  assign n10090 = \u2_R11_reg[11]/NET0131  & ~n10089 ;
  assign n10091 = ~\u2_R11_reg[11]/NET0131  & n10089 ;
  assign n10092 = ~n10090 & ~n10091 ;
  assign n10107 = n10070 & ~n10092 ;
  assign n10108 = n10106 & n10107 ;
  assign n10113 = ~n10047 & n10053 ;
  assign n10114 = n10070 & n10113 ;
  assign n10115 = n10060 & n10114 ;
  assign n10118 = ~n10108 & ~n10115 ;
  assign n10119 = ~n10117 & n10118 ;
  assign n10098 = n10053 & ~n10070 ;
  assign n10109 = n10047 & n10092 ;
  assign n10110 = n10064 & ~n10109 ;
  assign n10111 = n10098 & ~n10110 ;
  assign n10082 = ~n10053 & ~n10070 ;
  assign n10112 = n10082 & n10110 ;
  assign n10120 = ~n10111 & ~n10112 ;
  assign n10121 = n10119 & n10120 ;
  assign n10122 = ~n10080 & ~n10121 ;
  assign n10054 = n10047 & ~n10053 ;
  assign n10061 = ~n10053 & n10060 ;
  assign n10071 = ~n10060 & ~n10070 ;
  assign n10072 = ~n10061 & ~n10071 ;
  assign n10073 = n10064 & n10072 ;
  assign n10074 = ~n10054 & ~n10073 ;
  assign n10081 = ~n10074 & n10080 ;
  assign n10083 = n10062 & n10082 ;
  assign n10084 = n10054 & n10070 ;
  assign n10085 = ~n10083 & ~n10084 ;
  assign n10086 = ~n10081 & n10085 ;
  assign n10093 = ~n10086 & n10092 ;
  assign n10094 = n10070 & n10080 ;
  assign n10095 = n10053 & n10062 ;
  assign n10096 = n10094 & n10095 ;
  assign n10097 = n10080 & ~n10092 ;
  assign n10099 = n10047 & n10098 ;
  assign n10100 = ~n10047 & n10061 ;
  assign n10101 = n10053 & n10063 ;
  assign n10102 = ~n10100 & ~n10101 ;
  assign n10103 = ~n10099 & n10102 ;
  assign n10104 = n10097 & ~n10103 ;
  assign n10123 = ~n10096 & ~n10104 ;
  assign n10124 = ~n10093 & n10123 ;
  assign n10125 = ~n10122 & n10124 ;
  assign n10126 = ~\u2_L11_reg[6]/NET0131  & ~n10125 ;
  assign n10127 = \u2_L11_reg[6]/NET0131  & n10125 ;
  assign n10128 = ~n10126 & ~n10127 ;
  assign n10136 = ~n8898 & n9369 ;
  assign n10140 = ~n8860 & ~n8894 ;
  assign n10141 = ~n9369 & ~n10140 ;
  assign n10142 = ~n10136 & ~n10141 ;
  assign n10129 = ~n8869 & n8907 ;
  assign n10135 = n8869 & ~n8907 ;
  assign n10143 = ~n10129 & ~n10135 ;
  assign n10144 = ~n9370 & n10143 ;
  assign n10145 = ~n10142 & n10144 ;
  assign n10131 = ~n8918 & n10027 ;
  assign n10130 = ~n8854 & ~n8924 ;
  assign n10132 = ~n8921 & n10129 ;
  assign n10133 = ~n10130 & n10132 ;
  assign n10134 = ~n10131 & n10133 ;
  assign n10137 = ~n8891 & n10135 ;
  assign n10138 = ~n10030 & n10137 ;
  assign n10139 = ~n10136 & n10138 ;
  assign n10146 = ~n10134 & ~n10139 ;
  assign n10147 = ~n10145 & n10146 ;
  assign n10148 = ~\u2_L11_reg[7]/NET0131  & n10147 ;
  assign n10149 = \u2_L11_reg[7]/NET0131  & ~n10147 ;
  assign n10150 = ~n10148 & ~n10149 ;
  assign n10165 = ~n9400 & n9435 ;
  assign n10166 = ~n9818 & ~n10165 ;
  assign n10167 = n9394 & ~n10166 ;
  assign n10168 = n9413 & n9464 ;
  assign n10169 = ~n9477 & ~n10168 ;
  assign n10170 = ~n10167 & n10169 ;
  assign n10171 = n9452 & ~n10170 ;
  assign n10151 = n9394 & n9821 ;
  assign n10156 = ~n9436 & ~n10151 ;
  assign n10157 = n9833 & n10156 ;
  assign n10152 = n9427 & ~n9442 ;
  assign n10153 = ~n9818 & ~n10152 ;
  assign n10154 = ~n9394 & ~n10153 ;
  assign n10155 = n9394 & n9426 ;
  assign n10158 = ~n10154 & ~n10155 ;
  assign n10159 = n10157 & n10158 ;
  assign n10160 = ~n9452 & ~n10159 ;
  assign n10161 = n9427 & ~n9454 ;
  assign n10162 = ~n9423 & ~n10161 ;
  assign n10163 = n9394 & ~n10162 ;
  assign n10164 = ~n9419 & n9838 ;
  assign n10172 = ~n10163 & ~n10164 ;
  assign n10173 = ~n10160 & n10172 ;
  assign n10174 = ~n10171 & n10173 ;
  assign n10175 = ~\u2_L11_reg[8]/NET0131  & ~n10174 ;
  assign n10176 = \u2_L11_reg[8]/NET0131  & n10174 ;
  assign n10177 = ~n10175 & ~n10176 ;
  assign n10178 = n10070 & ~n10106 ;
  assign n10180 = n10092 & n10095 ;
  assign n10179 = n10054 & ~n10060 ;
  assign n10181 = ~n10070 & ~n10179 ;
  assign n10182 = n10102 & n10181 ;
  assign n10183 = ~n10180 & n10182 ;
  assign n10184 = ~n10178 & ~n10183 ;
  assign n10185 = n10062 & n10070 ;
  assign n10186 = ~n10053 & n10185 ;
  assign n10187 = n10092 & ~n10115 ;
  assign n10188 = ~n10186 & n10187 ;
  assign n10189 = n10060 & n10070 ;
  assign n10190 = ~n10047 & ~n10071 ;
  assign n10191 = ~n10189 & n10190 ;
  assign n10192 = ~n10188 & n10191 ;
  assign n10193 = ~n10184 & ~n10192 ;
  assign n10194 = n10080 & ~n10193 ;
  assign n10195 = ~n10053 & n10189 ;
  assign n10196 = ~n10092 & ~n10195 ;
  assign n10197 = ~n10188 & ~n10196 ;
  assign n10202 = n10062 & ~n10070 ;
  assign n10203 = ~n10101 & ~n10179 ;
  assign n10204 = ~n10202 & n10203 ;
  assign n10205 = ~n10092 & ~n10204 ;
  assign n10199 = ~n10062 & n10092 ;
  assign n10198 = ~n10053 & ~n10063 ;
  assign n10200 = ~n10101 & ~n10198 ;
  assign n10201 = n10199 & n10200 ;
  assign n10206 = ~n10083 & ~n10201 ;
  assign n10207 = ~n10205 & n10206 ;
  assign n10208 = ~n10080 & ~n10207 ;
  assign n10209 = ~n10197 & ~n10208 ;
  assign n10210 = ~n10194 & n10209 ;
  assign n10211 = ~\u2_L11_reg[16]/NET0131  & ~n10210 ;
  assign n10212 = \u2_L11_reg[16]/NET0131  & n10210 ;
  assign n10213 = ~n10211 & ~n10212 ;
  assign n10223 = ~n10070 & n10092 ;
  assign n10234 = ~n10053 & ~n10105 ;
  assign n10235 = n10223 & n10234 ;
  assign n10230 = ~n10082 & ~n10092 ;
  assign n10231 = ~n10064 & n10230 ;
  assign n10232 = ~n10061 & n10070 ;
  assign n10233 = n10199 & n10232 ;
  assign n10236 = ~n10231 & ~n10233 ;
  assign n10237 = ~n10235 & n10236 ;
  assign n10238 = ~n10112 & n10237 ;
  assign n10239 = n10080 & ~n10238 ;
  assign n10214 = n10047 & n10071 ;
  assign n10215 = ~n10185 & ~n10214 ;
  assign n10216 = ~n10095 & ~n10195 ;
  assign n10217 = n10215 & n10216 ;
  assign n10218 = n10092 & ~n10217 ;
  assign n10219 = ~n10047 & n10195 ;
  assign n10220 = ~n10218 & ~n10219 ;
  assign n10221 = ~n10080 & ~n10220 ;
  assign n10226 = ~n10064 & n10082 ;
  assign n10227 = ~n10073 & ~n10226 ;
  assign n10228 = ~n10080 & ~n10092 ;
  assign n10229 = ~n10227 & n10228 ;
  assign n10222 = n10101 & n10107 ;
  assign n10224 = ~n10100 & ~n10106 ;
  assign n10225 = n10223 & ~n10224 ;
  assign n10240 = ~n10222 & ~n10225 ;
  assign n10241 = ~n10229 & n10240 ;
  assign n10242 = ~n10221 & n10241 ;
  assign n10243 = ~n10239 & n10242 ;
  assign n10244 = ~\u2_L11_reg[24]/NET0131  & ~n10243 ;
  assign n10245 = \u2_L11_reg[24]/NET0131  & n10243 ;
  assign n10246 = ~n10244 & ~n10245 ;
  assign n10248 = ~n10070 & n10100 ;
  assign n10249 = n10215 & ~n10248 ;
  assign n10250 = n10080 & ~n10249 ;
  assign n10251 = ~n10113 & ~n10189 ;
  assign n10252 = ~n10080 & ~n10114 ;
  assign n10253 = ~n10251 & n10252 ;
  assign n10254 = ~n10250 & ~n10253 ;
  assign n10255 = n10092 & ~n10254 ;
  assign n10259 = n10070 & n10179 ;
  assign n10256 = ~n10053 & ~n10060 ;
  assign n10257 = ~n10092 & ~n10256 ;
  assign n10258 = n10251 & n10257 ;
  assign n10260 = ~n10226 & ~n10258 ;
  assign n10261 = ~n10259 & n10260 ;
  assign n10262 = ~n10080 & ~n10261 ;
  assign n10263 = ~n10095 & ~n10189 ;
  assign n10264 = n10097 & ~n10263 ;
  assign n10266 = n10053 & ~n10063 ;
  assign n10267 = n10094 & n10266 ;
  assign n10247 = n10107 & n10113 ;
  assign n10265 = n10109 & n10195 ;
  assign n10268 = ~n10247 & ~n10265 ;
  assign n10269 = ~n10267 & n10268 ;
  assign n10270 = ~n10264 & n10269 ;
  assign n10271 = ~n10262 & n10270 ;
  assign n10272 = ~n10255 & n10271 ;
  assign n10273 = \u2_L11_reg[30]/NET0131  & ~n10272 ;
  assign n10274 = ~\u2_L11_reg[30]/NET0131  & n10272 ;
  assign n10275 = ~n10273 & ~n10274 ;
  assign n10288 = ~n9456 & ~n9475 ;
  assign n10289 = n9394 & ~n10288 ;
  assign n10290 = ~n9394 & n9465 ;
  assign n10287 = n9400 & n9425 ;
  assign n10291 = ~n9421 & ~n10287 ;
  assign n10292 = ~n10290 & n10291 ;
  assign n10293 = ~n10289 & n10292 ;
  assign n10294 = n9452 & ~n10293 ;
  assign n10281 = ~n9433 & ~n9458 ;
  assign n10282 = ~n9818 & n10281 ;
  assign n10283 = ~n9394 & ~n10282 ;
  assign n10277 = ~n9424 & n9442 ;
  assign n10278 = ~n9400 & n9427 ;
  assign n10279 = ~n9457 & ~n10278 ;
  assign n10280 = n9394 & ~n10279 ;
  assign n10284 = ~n10277 & ~n10280 ;
  assign n10285 = ~n10283 & n10284 ;
  assign n10286 = ~n9452 & ~n10285 ;
  assign n10295 = ~n9443 & ~n9479 ;
  assign n10296 = ~n10165 & n10295 ;
  assign n10297 = ~n9394 & ~n10296 ;
  assign n10276 = n9428 & n9468 ;
  assign n10298 = ~n10155 & ~n10276 ;
  assign n10299 = ~n10297 & n10298 ;
  assign n10300 = ~n10286 & n10299 ;
  assign n10301 = ~n10294 & n10300 ;
  assign n10302 = ~\u2_L11_reg[3]/NET0131  & ~n10301 ;
  assign n10303 = \u2_L11_reg[3]/NET0131  & n10301 ;
  assign n10304 = ~n10302 & ~n10303 ;
  assign n10310 = ~n8978 & ~n9000 ;
  assign n10311 = ~n9945 & n10310 ;
  assign n10312 = n8944 & ~n10311 ;
  assign n10305 = n8950 & ~n8993 ;
  assign n10306 = ~n8978 & ~n10305 ;
  assign n10307 = ~n8944 & n10306 ;
  assign n10308 = ~n9003 & ~n9528 ;
  assign n10309 = ~n9539 & ~n10308 ;
  assign n10313 = ~n10307 & ~n10309 ;
  assign n10314 = ~n10312 & n10313 ;
  assign n10315 = ~n8988 & ~n10314 ;
  assign n10316 = ~n8963 & n9531 ;
  assign n10317 = ~n8972 & n9012 ;
  assign n10318 = ~n10316 & ~n10317 ;
  assign n10319 = ~n8944 & ~n10318 ;
  assign n10320 = n9532 & n9946 ;
  assign n10321 = n8963 & ~n10320 ;
  assign n10322 = n8974 & n10306 ;
  assign n10323 = ~n9538 & ~n10322 ;
  assign n10324 = ~n10321 & n10323 ;
  assign n10325 = n8988 & ~n10324 ;
  assign n10326 = ~n10319 & ~n10325 ;
  assign n10327 = ~n10315 & n10326 ;
  assign n10328 = ~\u2_L11_reg[9]/NET0131  & ~n10327 ;
  assign n10329 = \u2_L11_reg[9]/NET0131  & n10327 ;
  assign n10330 = ~n10328 & ~n10329 ;
  assign n10337 = n9665 & ~n9745 ;
  assign n10333 = n9629 & n9649 ;
  assign n10334 = n9642 & ~n9665 ;
  assign n10335 = ~n9744 & n10334 ;
  assign n10336 = ~n10333 & n10335 ;
  assign n10338 = n9683 & ~n9772 ;
  assign n10339 = ~n10336 & n10338 ;
  assign n10340 = ~n10337 & n10339 ;
  assign n10331 = n9635 & ~n9665 ;
  assign n10343 = n9642 & n9649 ;
  assign n10344 = ~n9749 & n10343 ;
  assign n10345 = ~n10331 & n10344 ;
  assign n10341 = ~n9642 & ~n9739 ;
  assign n10342 = n9758 & n10341 ;
  assign n10346 = ~n9765 & ~n10342 ;
  assign n10347 = ~n10345 & n10346 ;
  assign n10348 = n9689 & n10347 ;
  assign n10349 = ~n10340 & ~n10348 ;
  assign n10332 = n9656 & n10331 ;
  assign n10350 = n9642 & n10333 ;
  assign n10351 = ~n9891 & ~n10350 ;
  assign n10352 = n9665 & ~n10351 ;
  assign n10353 = ~n10332 & ~n10352 ;
  assign n10354 = ~n10349 & n10353 ;
  assign n10355 = ~\u2_L11_reg[18]/P0001  & ~n10354 ;
  assign n10356 = \u2_L11_reg[18]/P0001  & n10354 ;
  assign n10357 = ~n10355 & ~n10356 ;
  assign n10400 = decrypt_pad & ~\u2_uk_K_r10_reg[5]/NET0131  ;
  assign n10401 = ~decrypt_pad & ~\u2_uk_K_r10_reg[39]/NET0131  ;
  assign n10402 = ~n10400 & ~n10401 ;
  assign n10403 = \u2_R10_reg[4]/NET0131  & ~n10402 ;
  assign n10404 = ~\u2_R10_reg[4]/NET0131  & n10402 ;
  assign n10405 = ~n10403 & ~n10404 ;
  assign n10377 = decrypt_pad & ~\u2_uk_K_r10_reg[3]/NET0131  ;
  assign n10378 = ~decrypt_pad & ~\u2_uk_K_r10_reg[12]/NET0131  ;
  assign n10379 = ~n10377 & ~n10378 ;
  assign n10380 = \u2_R10_reg[1]/NET0131  & ~n10379 ;
  assign n10381 = ~\u2_R10_reg[1]/NET0131  & n10379 ;
  assign n10382 = ~n10380 & ~n10381 ;
  assign n10358 = decrypt_pad & ~\u2_uk_K_r10_reg[27]/NET0131  ;
  assign n10359 = ~decrypt_pad & ~\u2_uk_K_r10_reg[4]/NET0131  ;
  assign n10360 = ~n10358 & ~n10359 ;
  assign n10361 = \u2_R10_reg[3]/NET0131  & ~n10360 ;
  assign n10362 = ~\u2_R10_reg[3]/NET0131  & n10360 ;
  assign n10363 = ~n10361 & ~n10362 ;
  assign n10364 = decrypt_pad & ~\u2_uk_K_r10_reg[18]/NET0131  ;
  assign n10365 = ~decrypt_pad & ~\u2_uk_K_r10_reg[27]/NET0131  ;
  assign n10366 = ~n10364 & ~n10365 ;
  assign n10367 = \u2_R10_reg[2]/NET0131  & ~n10366 ;
  assign n10368 = ~\u2_R10_reg[2]/NET0131  & n10366 ;
  assign n10369 = ~n10367 & ~n10368 ;
  assign n10370 = decrypt_pad & ~\u2_uk_K_r10_reg[33]/NET0131  ;
  assign n10371 = ~decrypt_pad & ~\u2_uk_K_r10_reg[10]/NET0131  ;
  assign n10372 = ~n10370 & ~n10371 ;
  assign n10373 = \u2_R10_reg[5]/NET0131  & ~n10372 ;
  assign n10374 = ~\u2_R10_reg[5]/NET0131  & n10372 ;
  assign n10375 = ~n10373 & ~n10374 ;
  assign n10384 = decrypt_pad & ~\u2_uk_K_r10_reg[39]/NET0131  ;
  assign n10385 = ~decrypt_pad & ~\u2_uk_K_r10_reg[48]/NET0131  ;
  assign n10386 = ~n10384 & ~n10385 ;
  assign n10387 = \u2_R10_reg[32]/NET0131  & ~n10386 ;
  assign n10388 = ~\u2_R10_reg[32]/NET0131  & n10386 ;
  assign n10389 = ~n10387 & ~n10388 ;
  assign n10390 = n10375 & ~n10389 ;
  assign n10391 = n10369 & n10390 ;
  assign n10439 = n10363 & n10391 ;
  assign n10376 = ~n10369 & ~n10375 ;
  assign n10440 = n10376 & ~n10389 ;
  assign n10441 = ~n10439 & ~n10440 ;
  assign n10442 = n10382 & ~n10441 ;
  assign n10407 = n10369 & n10382 ;
  assign n10434 = ~n10375 & n10407 ;
  assign n10435 = n10389 & n10434 ;
  assign n10432 = ~n10369 & n10389 ;
  assign n10436 = n10375 & n10432 ;
  assign n10437 = ~n10435 & ~n10436 ;
  assign n10438 = n10363 & ~n10437 ;
  assign n10396 = n10375 & ~n10382 ;
  assign n10443 = n10396 & n10432 ;
  assign n10444 = ~n10438 & ~n10443 ;
  assign n10445 = ~n10442 & n10444 ;
  assign n10446 = ~n10405 & ~n10445 ;
  assign n10419 = ~n10375 & ~n10389 ;
  assign n10420 = n10369 & n10419 ;
  assign n10421 = ~n10396 & ~n10420 ;
  assign n10422 = n10363 & ~n10421 ;
  assign n10414 = ~n10363 & n10382 ;
  assign n10415 = ~n10369 & ~n10382 ;
  assign n10416 = ~n10375 & n10415 ;
  assign n10417 = ~n10414 & ~n10416 ;
  assign n10418 = n10389 & ~n10417 ;
  assign n10423 = n10363 & ~n10369 ;
  assign n10424 = n10382 & ~n10423 ;
  assign n10425 = ~n10376 & ~n10389 ;
  assign n10426 = ~n10424 & n10425 ;
  assign n10427 = ~n10418 & ~n10426 ;
  assign n10428 = ~n10422 & n10427 ;
  assign n10429 = n10405 & ~n10428 ;
  assign n10393 = ~n10375 & ~n10382 ;
  assign n10394 = n10389 & n10393 ;
  assign n10395 = n10369 & n10394 ;
  assign n10397 = ~n10369 & ~n10389 ;
  assign n10398 = ~n10396 & n10397 ;
  assign n10399 = ~n10395 & ~n10398 ;
  assign n10406 = ~n10399 & ~n10405 ;
  assign n10392 = ~n10382 & n10391 ;
  assign n10383 = n10376 & n10382 ;
  assign n10408 = n10375 & n10389 ;
  assign n10409 = n10407 & n10408 ;
  assign n10410 = ~n10383 & ~n10409 ;
  assign n10411 = ~n10392 & n10410 ;
  assign n10412 = ~n10406 & n10411 ;
  assign n10413 = ~n10363 & ~n10412 ;
  assign n10430 = n10363 & ~n10382 ;
  assign n10431 = n10420 & n10430 ;
  assign n10433 = n10430 & n10432 ;
  assign n10447 = ~n10431 & ~n10433 ;
  assign n10448 = ~n10413 & n10447 ;
  assign n10449 = ~n10429 & n10448 ;
  assign n10450 = ~n10446 & n10449 ;
  assign n10451 = ~\u2_L10_reg[31]/NET0131  & ~n10450 ;
  assign n10452 = \u2_L10_reg[31]/NET0131  & n10450 ;
  assign n10453 = ~n10451 & ~n10452 ;
  assign n10510 = decrypt_pad & ~\u2_uk_K_r10_reg[36]/NET0131  ;
  assign n10511 = ~decrypt_pad & ~\u2_uk_K_r10_reg[45]/P0001  ;
  assign n10512 = ~n10510 & ~n10511 ;
  assign n10513 = \u2_R10_reg[28]/NET0131  & ~n10512 ;
  assign n10514 = ~\u2_R10_reg[28]/NET0131  & n10512 ;
  assign n10515 = ~n10513 & ~n10514 ;
  assign n10467 = decrypt_pad & ~\u2_uk_K_r10_reg[49]/NET0131  ;
  assign n10468 = ~decrypt_pad & ~\u2_uk_K_r10_reg[30]/NET0131  ;
  assign n10469 = ~n10467 & ~n10468 ;
  assign n10470 = \u2_R10_reg[27]/NET0131  & ~n10469 ;
  assign n10471 = ~\u2_R10_reg[27]/NET0131  & n10469 ;
  assign n10472 = ~n10470 & ~n10471 ;
  assign n10483 = decrypt_pad & ~\u2_uk_K_r10_reg[16]/NET0131  ;
  assign n10484 = ~decrypt_pad & ~\u2_uk_K_r10_reg[21]/NET0131  ;
  assign n10485 = ~n10483 & ~n10484 ;
  assign n10486 = \u2_R10_reg[26]/NET0131  & ~n10485 ;
  assign n10487 = ~\u2_R10_reg[26]/NET0131  & n10485 ;
  assign n10488 = ~n10486 & ~n10487 ;
  assign n10460 = decrypt_pad & ~\u2_uk_K_r10_reg[51]/NET0131  ;
  assign n10461 = ~decrypt_pad & ~\u2_uk_K_r10_reg[1]/NET0131  ;
  assign n10462 = ~n10460 & ~n10461 ;
  assign n10463 = \u2_R10_reg[24]/NET0131  & ~n10462 ;
  assign n10464 = ~\u2_R10_reg[24]/NET0131  & n10462 ;
  assign n10465 = ~n10463 & ~n10464 ;
  assign n10454 = decrypt_pad & ~\u2_uk_K_r10_reg[28]/NET0131  ;
  assign n10455 = ~decrypt_pad & ~\u2_uk_K_r10_reg[9]/NET0131  ;
  assign n10456 = ~n10454 & ~n10455 ;
  assign n10457 = \u2_R10_reg[29]/NET0131  & ~n10456 ;
  assign n10458 = ~\u2_R10_reg[29]/NET0131  & n10456 ;
  assign n10459 = ~n10457 & ~n10458 ;
  assign n10474 = decrypt_pad & ~\u2_uk_K_r10_reg[0]/NET0131  ;
  assign n10475 = ~decrypt_pad & ~\u2_uk_K_r10_reg[36]/NET0131  ;
  assign n10476 = ~n10474 & ~n10475 ;
  assign n10477 = \u2_R10_reg[25]/NET0131  & ~n10476 ;
  assign n10478 = ~\u2_R10_reg[25]/NET0131  & n10476 ;
  assign n10479 = ~n10477 & ~n10478 ;
  assign n10528 = n10459 & ~n10479 ;
  assign n10529 = n10465 & n10528 ;
  assign n10530 = ~n10488 & n10529 ;
  assign n10505 = n10459 & n10479 ;
  assign n10531 = ~n10465 & n10505 ;
  assign n10532 = ~n10530 & ~n10531 ;
  assign n10533 = ~n10472 & ~n10532 ;
  assign n10499 = ~n10479 & ~n10488 ;
  assign n10534 = n10479 & n10488 ;
  assign n10535 = ~n10499 & ~n10534 ;
  assign n10490 = ~n10459 & n10479 ;
  assign n10500 = n10465 & n10472 ;
  assign n10536 = ~n10490 & n10500 ;
  assign n10537 = n10535 & n10536 ;
  assign n10466 = n10459 & ~n10465 ;
  assign n10495 = ~n10479 & n10488 ;
  assign n10524 = n10466 & n10495 ;
  assign n10480 = ~n10459 & ~n10479 ;
  assign n10502 = ~n10465 & ~n10488 ;
  assign n10538 = n10480 & n10502 ;
  assign n10539 = ~n10524 & ~n10538 ;
  assign n10540 = ~n10537 & n10539 ;
  assign n10541 = ~n10533 & n10540 ;
  assign n10542 = n10515 & ~n10541 ;
  assign n10491 = n10459 & n10488 ;
  assign n10492 = ~n10490 & ~n10491 ;
  assign n10493 = n10465 & ~n10492 ;
  assign n10494 = ~n10459 & ~n10465 ;
  assign n10496 = n10494 & n10495 ;
  assign n10497 = ~n10493 & ~n10496 ;
  assign n10498 = ~n10472 & ~n10497 ;
  assign n10473 = n10466 & ~n10472 ;
  assign n10481 = n10465 & n10480 ;
  assign n10482 = ~n10473 & ~n10481 ;
  assign n10489 = ~n10482 & ~n10488 ;
  assign n10501 = n10499 & n10500 ;
  assign n10503 = n10465 & n10488 ;
  assign n10504 = ~n10502 & ~n10503 ;
  assign n10506 = ~n10504 & n10505 ;
  assign n10507 = ~n10501 & ~n10506 ;
  assign n10508 = ~n10489 & n10507 ;
  assign n10509 = ~n10498 & n10508 ;
  assign n10516 = ~n10509 & ~n10515 ;
  assign n10522 = ~n10465 & n10490 ;
  assign n10523 = n10488 & n10522 ;
  assign n10525 = ~n10481 & ~n10524 ;
  assign n10526 = ~n10523 & n10525 ;
  assign n10527 = n10472 & ~n10526 ;
  assign n10517 = ~n10472 & n10479 ;
  assign n10518 = ~n10504 & n10517 ;
  assign n10519 = n10472 & ~n10479 ;
  assign n10520 = ~n10459 & ~n10488 ;
  assign n10521 = n10519 & n10520 ;
  assign n10543 = ~n10518 & ~n10521 ;
  assign n10544 = ~n10527 & n10543 ;
  assign n10545 = ~n10516 & n10544 ;
  assign n10546 = ~n10542 & n10545 ;
  assign n10547 = ~\u2_L10_reg[22]/NET0131  & ~n10546 ;
  assign n10548 = \u2_L10_reg[22]/NET0131  & n10546 ;
  assign n10549 = ~n10547 & ~n10548 ;
  assign n10591 = decrypt_pad & ~\u2_uk_K_r10_reg[29]/NET0131  ;
  assign n10592 = ~decrypt_pad & ~\u2_uk_K_r10_reg[38]/NET0131  ;
  assign n10593 = ~n10591 & ~n10592 ;
  assign n10594 = \u2_R10_reg[24]/NET0131  & ~n10593 ;
  assign n10595 = ~\u2_R10_reg[24]/NET0131  & n10593 ;
  assign n10596 = ~n10594 & ~n10595 ;
  assign n10550 = decrypt_pad & ~\u2_uk_K_r10_reg[31]/NET0131  ;
  assign n10551 = ~decrypt_pad & ~\u2_uk_K_r10_reg[8]/NET0131  ;
  assign n10552 = ~n10550 & ~n10551 ;
  assign n10553 = \u2_R10_reg[23]/NET0131  & ~n10552 ;
  assign n10554 = ~\u2_R10_reg[23]/NET0131  & n10552 ;
  assign n10555 = ~n10553 & ~n10554 ;
  assign n10563 = decrypt_pad & ~\u2_uk_K_r10_reg[8]/NET0131  ;
  assign n10564 = ~decrypt_pad & ~\u2_uk_K_r10_reg[44]/NET0131  ;
  assign n10565 = ~n10563 & ~n10564 ;
  assign n10566 = \u2_R10_reg[20]/NET0131  & ~n10565 ;
  assign n10567 = ~\u2_R10_reg[20]/NET0131  & n10565 ;
  assign n10568 = ~n10566 & ~n10567 ;
  assign n10576 = decrypt_pad & ~\u2_uk_K_r10_reg[52]/NET0131  ;
  assign n10577 = ~decrypt_pad & ~\u2_uk_K_r10_reg[29]/NET0131  ;
  assign n10578 = ~n10576 & ~n10577 ;
  assign n10579 = \u2_R10_reg[25]/NET0131  & ~n10578 ;
  assign n10580 = ~\u2_R10_reg[25]/NET0131  & n10578 ;
  assign n10581 = ~n10579 & ~n10580 ;
  assign n10613 = n10568 & n10581 ;
  assign n10556 = decrypt_pad & ~\u2_uk_K_r10_reg[14]/NET0131  ;
  assign n10557 = ~decrypt_pad & ~\u2_uk_K_r10_reg[50]/NET0131  ;
  assign n10558 = ~n10556 & ~n10557 ;
  assign n10559 = \u2_R10_reg[22]/NET0131  & ~n10558 ;
  assign n10560 = ~\u2_R10_reg[22]/NET0131  & n10558 ;
  assign n10561 = ~n10559 & ~n10560 ;
  assign n10569 = decrypt_pad & ~\u2_uk_K_r10_reg[23]/NET0131  ;
  assign n10570 = ~decrypt_pad & ~\u2_uk_K_r10_reg[28]/NET0131  ;
  assign n10571 = ~n10569 & ~n10570 ;
  assign n10572 = \u2_R10_reg[21]/NET0131  & ~n10571 ;
  assign n10573 = ~\u2_R10_reg[21]/NET0131  & n10571 ;
  assign n10574 = ~n10572 & ~n10573 ;
  assign n10604 = ~n10568 & n10574 ;
  assign n10629 = n10561 & ~n10604 ;
  assign n10630 = ~n10613 & n10629 ;
  assign n10631 = n10581 & n10604 ;
  assign n10632 = ~n10561 & n10631 ;
  assign n10633 = ~n10630 & ~n10632 ;
  assign n10634 = ~n10555 & ~n10633 ;
  assign n10586 = n10568 & ~n10581 ;
  assign n10623 = ~n10574 & n10586 ;
  assign n10624 = ~n10561 & n10623 ;
  assign n10615 = ~n10561 & ~n10568 ;
  assign n10625 = n10574 & ~n10586 ;
  assign n10626 = ~n10615 & n10625 ;
  assign n10627 = ~n10624 & ~n10626 ;
  assign n10628 = n10555 & ~n10627 ;
  assign n10562 = ~n10555 & ~n10561 ;
  assign n10635 = n10562 & n10613 ;
  assign n10636 = ~n10574 & n10635 ;
  assign n10637 = ~n10628 & ~n10636 ;
  assign n10638 = ~n10634 & n10637 ;
  assign n10639 = n10596 & ~n10638 ;
  assign n10605 = n10561 & n10604 ;
  assign n10597 = ~n10561 & n10574 ;
  assign n10606 = n10568 & n10597 ;
  assign n10607 = ~n10605 & ~n10606 ;
  assign n10608 = ~n10555 & ~n10607 ;
  assign n10599 = n10562 & n10586 ;
  assign n10600 = n10568 & ~n10574 ;
  assign n10601 = n10561 & n10600 ;
  assign n10602 = n10581 & n10601 ;
  assign n10603 = ~n10599 & ~n10602 ;
  assign n10575 = ~n10568 & ~n10574 ;
  assign n10584 = n10555 & n10581 ;
  assign n10585 = n10575 & n10584 ;
  assign n10598 = n10586 & n10597 ;
  assign n10609 = ~n10585 & ~n10598 ;
  assign n10610 = n10603 & n10609 ;
  assign n10611 = ~n10608 & n10610 ;
  assign n10612 = ~n10596 & ~n10611 ;
  assign n10616 = ~n10601 & ~n10615 ;
  assign n10617 = ~n10596 & ~n10616 ;
  assign n10614 = n10561 & n10613 ;
  assign n10618 = ~n10581 & n10604 ;
  assign n10619 = ~n10561 & n10618 ;
  assign n10620 = ~n10614 & ~n10619 ;
  assign n10621 = ~n10617 & n10620 ;
  assign n10622 = n10555 & ~n10621 ;
  assign n10582 = n10575 & ~n10581 ;
  assign n10583 = n10562 & n10582 ;
  assign n10587 = n10574 & n10586 ;
  assign n10588 = ~n10555 & n10587 ;
  assign n10589 = ~n10585 & ~n10588 ;
  assign n10590 = ~n10561 & ~n10589 ;
  assign n10640 = ~n10583 & ~n10590 ;
  assign n10641 = ~n10622 & n10640 ;
  assign n10642 = ~n10612 & n10641 ;
  assign n10643 = ~n10639 & n10642 ;
  assign n10644 = \u2_L10_reg[11]/NET0131  & ~n10643 ;
  assign n10645 = ~\u2_L10_reg[11]/NET0131  & n10643 ;
  assign n10646 = ~n10644 & ~n10645 ;
  assign n10647 = decrypt_pad & ~\u2_uk_K_r10_reg[32]/NET0131  ;
  assign n10648 = ~decrypt_pad & ~\u2_uk_K_r10_reg[41]/NET0131  ;
  assign n10649 = ~n10647 & ~n10648 ;
  assign n10650 = \u2_R10_reg[16]/NET0131  & ~n10649 ;
  assign n10651 = ~\u2_R10_reg[16]/NET0131  & n10649 ;
  assign n10652 = ~n10650 & ~n10651 ;
  assign n10673 = decrypt_pad & ~\u2_uk_K_r10_reg[24]/NET0131  ;
  assign n10674 = ~decrypt_pad & ~\u2_uk_K_r10_reg[33]/NET0131  ;
  assign n10675 = ~n10673 & ~n10674 ;
  assign n10676 = \u2_R10_reg[15]/NET0131  & ~n10675 ;
  assign n10677 = ~\u2_R10_reg[15]/NET0131  & n10675 ;
  assign n10678 = ~n10676 & ~n10677 ;
  assign n10682 = decrypt_pad & ~\u2_uk_K_r10_reg[48]/NET0131  ;
  assign n10683 = ~decrypt_pad & ~\u2_uk_K_r10_reg[25]/NET0131  ;
  assign n10684 = ~n10682 & ~n10683 ;
  assign n10685 = \u2_R10_reg[14]/NET0131  & ~n10684 ;
  assign n10686 = ~\u2_R10_reg[14]/NET0131  & n10684 ;
  assign n10687 = ~n10685 & ~n10686 ;
  assign n10712 = ~n10678 & ~n10687 ;
  assign n10653 = decrypt_pad & ~\u2_uk_K_r10_reg[53]/NET0131  ;
  assign n10654 = ~decrypt_pad & ~\u2_uk_K_r10_reg[5]/NET0131  ;
  assign n10655 = ~n10653 & ~n10654 ;
  assign n10656 = \u2_R10_reg[12]/NET0131  & ~n10655 ;
  assign n10657 = ~\u2_R10_reg[12]/NET0131  & n10655 ;
  assign n10658 = ~n10656 & ~n10657 ;
  assign n10666 = decrypt_pad & ~\u2_uk_K_r10_reg[47]/NET0131  ;
  assign n10667 = ~decrypt_pad & ~\u2_uk_K_r10_reg[24]/NET0131  ;
  assign n10668 = ~n10666 & ~n10667 ;
  assign n10669 = \u2_R10_reg[13]/NET0131  & ~n10668 ;
  assign n10670 = ~\u2_R10_reg[13]/NET0131  & n10668 ;
  assign n10671 = ~n10669 & ~n10670 ;
  assign n10680 = ~n10658 & n10671 ;
  assign n10703 = n10658 & ~n10671 ;
  assign n10724 = ~n10680 & ~n10703 ;
  assign n10725 = n10712 & ~n10724 ;
  assign n10659 = decrypt_pad & ~\u2_uk_K_r10_reg[12]/NET0131  ;
  assign n10660 = ~decrypt_pad & ~\u2_uk_K_r10_reg[46]/NET0131  ;
  assign n10661 = ~n10659 & ~n10660 ;
  assign n10662 = \u2_R10_reg[17]/NET0131  & ~n10661 ;
  assign n10663 = ~\u2_R10_reg[17]/NET0131  & n10661 ;
  assign n10664 = ~n10662 & ~n10663 ;
  assign n10721 = ~n10658 & n10664 ;
  assign n10722 = n10678 & n10721 ;
  assign n10723 = ~n10671 & n10722 ;
  assign n10693 = n10658 & ~n10664 ;
  assign n10698 = n10671 & n10678 ;
  assign n10732 = n10693 & n10698 ;
  assign n10733 = ~n10723 & ~n10732 ;
  assign n10734 = ~n10725 & n10733 ;
  assign n10665 = n10658 & n10664 ;
  assign n10672 = n10665 & n10671 ;
  assign n10726 = n10672 & n10687 ;
  assign n10727 = n10671 & n10721 ;
  assign n10728 = ~n10687 & n10727 ;
  assign n10729 = ~n10726 & ~n10728 ;
  assign n10689 = ~n10664 & ~n10671 ;
  assign n10701 = ~n10658 & n10689 ;
  assign n10730 = ~n10678 & n10701 ;
  assign n10731 = n10687 & n10730 ;
  assign n10735 = n10729 & ~n10731 ;
  assign n10736 = n10734 & n10735 ;
  assign n10737 = n10652 & ~n10736 ;
  assign n10679 = n10672 & n10678 ;
  assign n10699 = n10687 & n10698 ;
  assign n10700 = ~n10658 & n10699 ;
  assign n10706 = ~n10679 & ~n10700 ;
  assign n10702 = n10678 & n10701 ;
  assign n10704 = ~n10687 & n10703 ;
  assign n10705 = n10664 & n10704 ;
  assign n10707 = ~n10702 & ~n10705 ;
  assign n10708 = n10706 & n10707 ;
  assign n10681 = ~n10664 & n10680 ;
  assign n10688 = n10681 & n10687 ;
  assign n10690 = ~n10658 & ~n10687 ;
  assign n10691 = n10689 & n10690 ;
  assign n10692 = ~n10688 & ~n10691 ;
  assign n10694 = n10687 & n10693 ;
  assign n10695 = n10664 & ~n10671 ;
  assign n10696 = ~n10694 & ~n10695 ;
  assign n10697 = ~n10678 & ~n10696 ;
  assign n10709 = n10692 & ~n10697 ;
  assign n10710 = n10708 & n10709 ;
  assign n10711 = ~n10652 & ~n10710 ;
  assign n10715 = ~n10671 & n10687 ;
  assign n10716 = n10693 & n10715 ;
  assign n10717 = ~n10691 & ~n10716 ;
  assign n10718 = n10678 & ~n10717 ;
  assign n10713 = n10664 & n10712 ;
  assign n10714 = n10680 & n10713 ;
  assign n10719 = ~n10687 & n10693 ;
  assign n10720 = n10698 & n10719 ;
  assign n10738 = ~n10714 & ~n10720 ;
  assign n10739 = ~n10718 & n10738 ;
  assign n10740 = ~n10711 & n10739 ;
  assign n10741 = ~n10737 & n10740 ;
  assign n10742 = ~\u2_L10_reg[20]/NET0131  & ~n10741 ;
  assign n10743 = \u2_L10_reg[20]/NET0131  & n10741 ;
  assign n10744 = ~n10742 & ~n10743 ;
  assign n10745 = decrypt_pad & ~\u2_uk_K_r10_reg[6]/NET0131  ;
  assign n10746 = ~decrypt_pad & ~\u2_uk_K_r10_reg[40]/NET0131  ;
  assign n10747 = ~n10745 & ~n10746 ;
  assign n10748 = \u2_R10_reg[8]/NET0131  & ~n10747 ;
  assign n10749 = ~\u2_R10_reg[8]/NET0131  & n10747 ;
  assign n10750 = ~n10748 & ~n10749 ;
  assign n10751 = decrypt_pad & ~\u2_uk_K_r10_reg[40]/NET0131  ;
  assign n10752 = ~decrypt_pad & ~\u2_uk_K_r10_reg[17]/NET0131  ;
  assign n10753 = ~n10751 & ~n10752 ;
  assign n10754 = \u2_R10_reg[7]/NET0131  & ~n10753 ;
  assign n10755 = ~\u2_R10_reg[7]/NET0131  & n10753 ;
  assign n10756 = ~n10754 & ~n10755 ;
  assign n10770 = decrypt_pad & ~\u2_uk_K_r10_reg[55]/NET0131  ;
  assign n10771 = ~decrypt_pad & ~\u2_uk_K_r10_reg[32]/NET0131  ;
  assign n10772 = ~n10770 & ~n10771 ;
  assign n10773 = \u2_R10_reg[5]/NET0131  & ~n10772 ;
  assign n10774 = ~\u2_R10_reg[5]/NET0131  & n10772 ;
  assign n10775 = ~n10773 & ~n10774 ;
  assign n10757 = decrypt_pad & ~\u2_uk_K_r10_reg[19]/NET0131  ;
  assign n10758 = ~decrypt_pad & ~\u2_uk_K_r10_reg[53]/NET0131  ;
  assign n10759 = ~n10757 & ~n10758 ;
  assign n10760 = \u2_R10_reg[4]/NET0131  & ~n10759 ;
  assign n10761 = ~\u2_R10_reg[4]/NET0131  & n10759 ;
  assign n10762 = ~n10760 & ~n10761 ;
  assign n10763 = decrypt_pad & ~\u2_uk_K_r10_reg[11]/NET0131  ;
  assign n10764 = ~decrypt_pad & ~\u2_uk_K_r10_reg[20]/NET0131  ;
  assign n10765 = ~n10763 & ~n10764 ;
  assign n10766 = \u2_R10_reg[9]/NET0131  & ~n10765 ;
  assign n10767 = ~\u2_R10_reg[9]/NET0131  & n10765 ;
  assign n10768 = ~n10766 & ~n10767 ;
  assign n10785 = ~n10762 & n10768 ;
  assign n10786 = ~n10775 & n10785 ;
  assign n10777 = decrypt_pad & ~\u2_uk_K_r10_reg[46]/NET0131  ;
  assign n10778 = ~decrypt_pad & ~\u2_uk_K_r10_reg[55]/NET0131  ;
  assign n10779 = ~n10777 & ~n10778 ;
  assign n10780 = \u2_R10_reg[6]/NET0131  & ~n10779 ;
  assign n10781 = ~\u2_R10_reg[6]/NET0131  & n10779 ;
  assign n10782 = ~n10780 & ~n10781 ;
  assign n10787 = n10762 & ~n10768 ;
  assign n10788 = n10762 & n10775 ;
  assign n10789 = ~n10787 & ~n10788 ;
  assign n10790 = n10782 & ~n10789 ;
  assign n10791 = ~n10786 & ~n10790 ;
  assign n10792 = ~n10756 & ~n10791 ;
  assign n10796 = n10782 & n10785 ;
  assign n10797 = n10775 & n10796 ;
  assign n10798 = ~n10775 & ~n10782 ;
  assign n10799 = ~n10756 & n10768 ;
  assign n10800 = n10798 & n10799 ;
  assign n10801 = ~n10797 & ~n10800 ;
  assign n10769 = n10762 & n10768 ;
  assign n10776 = n10769 & ~n10775 ;
  assign n10783 = n10776 & n10782 ;
  assign n10784 = n10756 & n10783 ;
  assign n10793 = ~n10768 & n10775 ;
  assign n10794 = ~n10786 & ~n10793 ;
  assign n10795 = ~n10782 & ~n10794 ;
  assign n10802 = ~n10784 & ~n10795 ;
  assign n10803 = n10801 & n10802 ;
  assign n10804 = ~n10792 & n10803 ;
  assign n10805 = ~n10750 & ~n10804 ;
  assign n10823 = ~n10762 & ~n10768 ;
  assign n10824 = ~n10783 & ~n10823 ;
  assign n10825 = n10750 & ~n10824 ;
  assign n10806 = ~n10775 & n10782 ;
  assign n10826 = n10785 & ~n10806 ;
  assign n10827 = ~n10825 & ~n10826 ;
  assign n10809 = n10775 & ~n10782 ;
  assign n10828 = ~n10756 & ~n10809 ;
  assign n10829 = ~n10827 & n10828 ;
  assign n10807 = ~n10768 & n10806 ;
  assign n10808 = ~n10762 & n10807 ;
  assign n10810 = n10762 & n10809 ;
  assign n10811 = ~n10808 & ~n10810 ;
  assign n10812 = n10756 & ~n10811 ;
  assign n10818 = ~n10775 & n10787 ;
  assign n10819 = ~n10782 & n10818 ;
  assign n10813 = n10768 & n10788 ;
  assign n10814 = ~n10782 & n10813 ;
  assign n10815 = ~n10762 & n10782 ;
  assign n10816 = n10756 & n10775 ;
  assign n10817 = ~n10815 & n10816 ;
  assign n10820 = ~n10814 & ~n10817 ;
  assign n10821 = ~n10819 & n10820 ;
  assign n10822 = n10750 & ~n10821 ;
  assign n10830 = ~n10812 & ~n10822 ;
  assign n10831 = ~n10829 & n10830 ;
  assign n10832 = ~n10805 & n10831 ;
  assign n10833 = \u2_L10_reg[2]/NET0131  & n10832 ;
  assign n10834 = ~\u2_L10_reg[2]/NET0131  & ~n10832 ;
  assign n10835 = ~n10833 & ~n10834 ;
  assign n10844 = n10561 & n10587 ;
  assign n10860 = ~n10561 & ~n10575 ;
  assign n10861 = ~n10586 & n10860 ;
  assign n10862 = ~n10844 & ~n10861 ;
  assign n10863 = ~n10555 & ~n10862 ;
  assign n10853 = n10561 & n10581 ;
  assign n10854 = n10575 & n10853 ;
  assign n10855 = n10574 & n10613 ;
  assign n10856 = ~n10623 & ~n10855 ;
  assign n10840 = ~n10581 & ~n10597 ;
  assign n10857 = ~n10629 & n10840 ;
  assign n10858 = n10856 & ~n10857 ;
  assign n10859 = n10555 & ~n10858 ;
  assign n10864 = ~n10854 & ~n10859 ;
  assign n10865 = ~n10863 & n10864 ;
  assign n10866 = ~n10596 & ~n10865 ;
  assign n10836 = n10561 & ~n10581 ;
  assign n10845 = n10604 & ~n10836 ;
  assign n10846 = ~n10844 & ~n10845 ;
  assign n10847 = n10555 & ~n10846 ;
  assign n10841 = ~n10568 & n10840 ;
  assign n10842 = ~n10614 & ~n10841 ;
  assign n10843 = ~n10555 & ~n10842 ;
  assign n10837 = ~n10561 & n10581 ;
  assign n10838 = ~n10836 & ~n10837 ;
  assign n10839 = n10575 & ~n10838 ;
  assign n10848 = n10603 & ~n10839 ;
  assign n10849 = ~n10843 & n10848 ;
  assign n10850 = ~n10847 & n10849 ;
  assign n10851 = n10596 & ~n10850 ;
  assign n10852 = n10584 & n10597 ;
  assign n10867 = ~n10624 & ~n10852 ;
  assign n10868 = ~n10851 & n10867 ;
  assign n10869 = ~n10866 & n10868 ;
  assign n10870 = \u2_L10_reg[29]/NET0131  & ~n10869 ;
  assign n10871 = ~\u2_L10_reg[29]/NET0131  & n10869 ;
  assign n10872 = ~n10870 & ~n10871 ;
  assign n10925 = decrypt_pad & ~\u2_uk_K_r10_reg[1]/NET0131  ;
  assign n10926 = ~decrypt_pad & ~\u2_uk_K_r10_reg[37]/NET0131  ;
  assign n10927 = ~n10925 & ~n10926 ;
  assign n10928 = \u2_R10_reg[32]/NET0131  & ~n10927 ;
  assign n10929 = ~\u2_R10_reg[32]/NET0131  & n10927 ;
  assign n10930 = ~n10928 & ~n10929 ;
  assign n10899 = decrypt_pad & ~\u2_uk_K_r10_reg[50]/NET0131  ;
  assign n10900 = ~decrypt_pad & ~\u2_uk_K_r10_reg[0]/NET0131  ;
  assign n10901 = ~n10899 & ~n10900 ;
  assign n10902 = \u2_R10_reg[31]/P0001  & ~n10901 ;
  assign n10903 = ~\u2_R10_reg[31]/P0001  & n10901 ;
  assign n10904 = ~n10902 & ~n10903 ;
  assign n10879 = decrypt_pad & ~\u2_uk_K_r10_reg[7]/NET0131  ;
  assign n10880 = ~decrypt_pad & ~\u2_uk_K_r10_reg[43]/NET0131  ;
  assign n10881 = ~n10879 & ~n10880 ;
  assign n10882 = \u2_R10_reg[30]/NET0131  & ~n10881 ;
  assign n10883 = ~\u2_R10_reg[30]/NET0131  & n10881 ;
  assign n10884 = ~n10882 & ~n10883 ;
  assign n10873 = decrypt_pad & ~\u2_uk_K_r10_reg[38]/NET0131  ;
  assign n10874 = ~decrypt_pad & ~\u2_uk_K_r10_reg[15]/NET0131  ;
  assign n10875 = ~n10873 & ~n10874 ;
  assign n10876 = \u2_R10_reg[28]/NET0131  & ~n10875 ;
  assign n10877 = ~\u2_R10_reg[28]/NET0131  & n10875 ;
  assign n10878 = ~n10876 & ~n10877 ;
  assign n10885 = decrypt_pad & ~\u2_uk_K_r10_reg[37]/NET0131  ;
  assign n10886 = ~decrypt_pad & ~\u2_uk_K_r10_reg[42]/NET0131  ;
  assign n10887 = ~n10885 & ~n10886 ;
  assign n10888 = \u2_R10_reg[29]/NET0131  & ~n10887 ;
  assign n10889 = ~\u2_R10_reg[29]/NET0131  & n10887 ;
  assign n10890 = ~n10888 & ~n10889 ;
  assign n10933 = n10878 & ~n10890 ;
  assign n10892 = decrypt_pad & ~\u2_uk_K_r10_reg[22]/NET0131  ;
  assign n10893 = ~decrypt_pad & ~\u2_uk_K_r10_reg[31]/NET0131  ;
  assign n10894 = ~n10892 & ~n10893 ;
  assign n10895 = \u2_R10_reg[1]/NET0131  & ~n10894 ;
  assign n10896 = ~\u2_R10_reg[1]/NET0131  & n10894 ;
  assign n10897 = ~n10895 & ~n10896 ;
  assign n10951 = n10878 & n10897 ;
  assign n10952 = ~n10933 & ~n10951 ;
  assign n10953 = ~n10884 & ~n10952 ;
  assign n10906 = n10884 & n10890 ;
  assign n10950 = ~n10897 & n10906 ;
  assign n10918 = ~n10878 & ~n10897 ;
  assign n10954 = n10890 & n10918 ;
  assign n10955 = ~n10950 & ~n10954 ;
  assign n10956 = ~n10953 & n10955 ;
  assign n10957 = n10904 & ~n10956 ;
  assign n10938 = ~n10878 & n10906 ;
  assign n10949 = n10897 & n10938 ;
  assign n10940 = ~n10884 & ~n10890 ;
  assign n10958 = ~n10878 & n10940 ;
  assign n10959 = ~n10904 & n10958 ;
  assign n10960 = ~n10949 & ~n10959 ;
  assign n10961 = ~n10957 & n10960 ;
  assign n10962 = n10930 & ~n10961 ;
  assign n10907 = n10897 & n10906 ;
  assign n10891 = ~n10884 & n10890 ;
  assign n10898 = n10891 & ~n10897 ;
  assign n10905 = ~n10884 & ~n10904 ;
  assign n10908 = ~n10898 & ~n10905 ;
  assign n10909 = ~n10907 & n10908 ;
  assign n10910 = n10878 & ~n10909 ;
  assign n10913 = n10884 & ~n10890 ;
  assign n10914 = n10878 & ~n10897 ;
  assign n10915 = n10913 & n10914 ;
  assign n10911 = ~n10878 & n10897 ;
  assign n10912 = ~n10890 & n10911 ;
  assign n10916 = n10904 & ~n10912 ;
  assign n10917 = ~n10915 & n10916 ;
  assign n10919 = n10884 & n10918 ;
  assign n10920 = n10890 & n10897 ;
  assign n10921 = ~n10904 & ~n10920 ;
  assign n10922 = ~n10919 & n10921 ;
  assign n10923 = ~n10917 & ~n10922 ;
  assign n10924 = ~n10910 & ~n10923 ;
  assign n10931 = ~n10924 & ~n10930 ;
  assign n10939 = ~n10897 & n10938 ;
  assign n10941 = n10897 & n10940 ;
  assign n10942 = n10878 & n10941 ;
  assign n10943 = ~n10939 & ~n10942 ;
  assign n10944 = n10918 & n10940 ;
  assign n10945 = n10884 & n10912 ;
  assign n10946 = ~n10944 & ~n10945 ;
  assign n10947 = n10943 & n10946 ;
  assign n10948 = n10904 & ~n10947 ;
  assign n10932 = n10884 & ~n10904 ;
  assign n10934 = n10930 & n10932 ;
  assign n10935 = n10933 & n10934 ;
  assign n10936 = n10890 & n10914 ;
  assign n10937 = n10905 & n10936 ;
  assign n10963 = ~n10935 & ~n10937 ;
  assign n10964 = ~n10948 & n10963 ;
  assign n10965 = ~n10931 & n10964 ;
  assign n10966 = ~n10962 & n10965 ;
  assign n10967 = \u2_L10_reg[5]/NET0131  & ~n10966 ;
  assign n10968 = ~\u2_L10_reg[5]/NET0131  & n10966 ;
  assign n10969 = ~n10967 & ~n10968 ;
  assign n10979 = n10581 & ~n10616 ;
  assign n10980 = n10555 & ~n10587 ;
  assign n10981 = ~n10979 & n10980 ;
  assign n10982 = ~n10555 & ~n10618 ;
  assign n10983 = ~n10854 & n10982 ;
  assign n10984 = ~n10981 & ~n10983 ;
  assign n10985 = ~n10624 & ~n10635 ;
  assign n10986 = ~n10984 & n10985 ;
  assign n10987 = ~n10596 & ~n10986 ;
  assign n10992 = n10561 & ~n10856 ;
  assign n10993 = ~n10615 & ~n10992 ;
  assign n10994 = ~n10555 & ~n10837 ;
  assign n10995 = ~n10993 & n10994 ;
  assign n10971 = ~n10581 & n10597 ;
  assign n10972 = ~n10615 & ~n10971 ;
  assign n10973 = ~n10555 & ~n10972 ;
  assign n10970 = n10625 & n10838 ;
  assign n10974 = n10555 & ~n10561 ;
  assign n10975 = n10613 & n10974 ;
  assign n10976 = ~n10970 & ~n10975 ;
  assign n10977 = ~n10973 & n10976 ;
  assign n10978 = n10596 & ~n10977 ;
  assign n10988 = ~n10582 & ~n10631 ;
  assign n10989 = ~n10587 & n10988 ;
  assign n10990 = n10555 & n10561 ;
  assign n10991 = ~n10989 & n10990 ;
  assign n10996 = ~n10978 & ~n10991 ;
  assign n10997 = ~n10995 & n10996 ;
  assign n10998 = ~n10987 & n10997 ;
  assign n10999 = ~\u2_L10_reg[4]/NET0131  & ~n10998 ;
  assign n11000 = \u2_L10_reg[4]/NET0131  & n10998 ;
  assign n11001 = ~n10999 & ~n11000 ;
  assign n11006 = n10383 & n10389 ;
  assign n11007 = n10405 & ~n11006 ;
  assign n11002 = ~n10389 & ~n10415 ;
  assign n11003 = ~n10443 & ~n11002 ;
  assign n11004 = n10363 & ~n11003 ;
  assign n11005 = n10375 & n10407 ;
  assign n11008 = ~n10363 & ~n10432 ;
  assign n11009 = ~n11002 & n11008 ;
  assign n11010 = ~n11005 & ~n11009 ;
  assign n11011 = ~n11004 & n11010 ;
  assign n11012 = n11007 & n11011 ;
  assign n11017 = ~n10369 & n10390 ;
  assign n11018 = ~n10420 & ~n11017 ;
  assign n11019 = n10382 & ~n11018 ;
  assign n11020 = n10382 & n10408 ;
  assign n11021 = ~n10394 & ~n11020 ;
  assign n11022 = ~n11019 & n11021 ;
  assign n11023 = n10363 & ~n11022 ;
  assign n11013 = ~n10408 & ~n10419 ;
  assign n11014 = ~n10382 & ~n11013 ;
  assign n11015 = ~n10440 & ~n11014 ;
  assign n11016 = ~n10363 & ~n11015 ;
  assign n11024 = ~n10392 & ~n10405 ;
  assign n11025 = ~n10435 & n11024 ;
  assign n11026 = ~n11016 & n11025 ;
  assign n11027 = ~n11023 & n11026 ;
  assign n11028 = ~n11012 & ~n11027 ;
  assign n11029 = ~\u2_L10_reg[17]/NET0131  & n11028 ;
  assign n11030 = \u2_L10_reg[17]/NET0131  & ~n11028 ;
  assign n11031 = ~n11029 & ~n11030 ;
  assign n11036 = ~n10555 & ~n10988 ;
  assign n11032 = n10568 & ~n10597 ;
  assign n11033 = ~n10618 & ~n11032 ;
  assign n11034 = n10555 & ~n11033 ;
  assign n11035 = n10561 & n10855 ;
  assign n11037 = ~n10596 & ~n11035 ;
  assign n11038 = ~n11034 & n11037 ;
  assign n11039 = ~n11036 & n11038 ;
  assign n11043 = ~n10585 & n10596 ;
  assign n11041 = ~n10555 & n10600 ;
  assign n11044 = ~n10971 & ~n11041 ;
  assign n11045 = n11043 & n11044 ;
  assign n11042 = n10555 & n10606 ;
  assign n11040 = n10561 & n10631 ;
  assign n11046 = ~n10839 & ~n11040 ;
  assign n11047 = ~n11042 & n11046 ;
  assign n11048 = n11045 & n11047 ;
  assign n11049 = ~n11039 & ~n11048 ;
  assign n11050 = ~n10590 & ~n10636 ;
  assign n11051 = ~n11049 & n11050 ;
  assign n11052 = ~\u2_L10_reg[19]/NET0131  & ~n11051 ;
  assign n11053 = \u2_L10_reg[19]/NET0131  & n11051 ;
  assign n11054 = ~n11052 & ~n11053 ;
  assign n11072 = ~n10664 & n10690 ;
  assign n11073 = n10678 & ~n10716 ;
  assign n11074 = ~n11072 & n11073 ;
  assign n11075 = n10658 & n10695 ;
  assign n11076 = ~n10678 & ~n10719 ;
  assign n11077 = ~n11075 & n11076 ;
  assign n11078 = ~n11074 & ~n11077 ;
  assign n11079 = n10671 & n10719 ;
  assign n11080 = n10729 & ~n11079 ;
  assign n11081 = ~n11078 & n11080 ;
  assign n11082 = ~n10652 & ~n11081 ;
  assign n11065 = n10671 & ~n10687 ;
  assign n11066 = ~n10693 & n11065 ;
  assign n11067 = ~n10727 & ~n11066 ;
  assign n11068 = ~n10678 & ~n11067 ;
  assign n11055 = ~n10658 & n10715 ;
  assign n11063 = n10671 & n10694 ;
  assign n11069 = ~n11055 & ~n11063 ;
  assign n11070 = ~n11068 & n11069 ;
  assign n11071 = n10652 & ~n11070 ;
  assign n11056 = n10664 & n11055 ;
  assign n11057 = ~n10726 & ~n11056 ;
  assign n11058 = ~n10688 & n11057 ;
  assign n11059 = n10678 & ~n11058 ;
  assign n11064 = ~n10678 & n11063 ;
  assign n11060 = ~n10695 & ~n10704 ;
  assign n11061 = n10652 & n10678 ;
  assign n11062 = ~n11060 & n11061 ;
  assign n11083 = ~n10731 & ~n11062 ;
  assign n11084 = ~n11064 & n11083 ;
  assign n11085 = ~n11059 & n11084 ;
  assign n11086 = ~n11071 & n11085 ;
  assign n11087 = ~n11082 & n11086 ;
  assign n11088 = ~\u2_L10_reg[1]/NET0131  & ~n11087 ;
  assign n11089 = \u2_L10_reg[1]/NET0131  & n11087 ;
  assign n11090 = ~n11088 & ~n11089 ;
  assign n11096 = ~n10904 & n10954 ;
  assign n11091 = ~n10891 & ~n10905 ;
  assign n11092 = n10951 & ~n11091 ;
  assign n11098 = ~n10915 & ~n10930 ;
  assign n11101 = ~n11092 & n11098 ;
  assign n11102 = ~n11096 & n11101 ;
  assign n11093 = n10884 & n10933 ;
  assign n11094 = ~n10936 & ~n11093 ;
  assign n11095 = n10904 & ~n11094 ;
  assign n11097 = n10911 & n10932 ;
  assign n11099 = ~n10938 & ~n10944 ;
  assign n11100 = ~n11097 & n11099 ;
  assign n11103 = ~n11095 & n11100 ;
  assign n11104 = n11102 & n11103 ;
  assign n11111 = n10904 & ~n10941 ;
  assign n11109 = n10878 & n10906 ;
  assign n11110 = n10890 & n10911 ;
  assign n11112 = ~n11109 & ~n11110 ;
  assign n11113 = n11111 & n11112 ;
  assign n11115 = ~n10884 & n10914 ;
  assign n11114 = n10913 & n10951 ;
  assign n11116 = ~n10904 & ~n11114 ;
  assign n11117 = ~n11115 & n11116 ;
  assign n11118 = ~n11113 & ~n11117 ;
  assign n11106 = ~n10890 & n10918 ;
  assign n11107 = ~n10936 & ~n11106 ;
  assign n11108 = n10884 & ~n11107 ;
  assign n11105 = ~n10884 & n10912 ;
  assign n11119 = n10930 & ~n11105 ;
  assign n11120 = ~n11108 & n11119 ;
  assign n11121 = ~n11118 & n11120 ;
  assign n11122 = ~n11104 & ~n11121 ;
  assign n11123 = n10904 & n10958 ;
  assign n11124 = n10878 & n10905 ;
  assign n11125 = n10920 & n11124 ;
  assign n11126 = ~n11123 & ~n11125 ;
  assign n11127 = ~n11122 & n11126 ;
  assign n11128 = ~\u2_L10_reg[21]/NET0131  & ~n11127 ;
  assign n11129 = \u2_L10_reg[21]/NET0131  & n11127 ;
  assign n11130 = ~n11128 & ~n11129 ;
  assign n11132 = n10382 & n10419 ;
  assign n11151 = ~n10382 & n10390 ;
  assign n11152 = ~n11132 & ~n11151 ;
  assign n11153 = ~n10395 & n11152 ;
  assign n11154 = n10405 & ~n11153 ;
  assign n11155 = n10390 & n10415 ;
  assign n11156 = ~n11006 & ~n11155 ;
  assign n11157 = ~n11154 & n11156 ;
  assign n11158 = ~n10363 & ~n11157 ;
  assign n11145 = n10382 & n10390 ;
  assign n11146 = ~n10435 & ~n11145 ;
  assign n11147 = n10363 & ~n11146 ;
  assign n11148 = ~n10431 & ~n10443 ;
  assign n11149 = ~n11147 & n11148 ;
  assign n11150 = n10405 & ~n11149 ;
  assign n11133 = ~n10391 & ~n11132 ;
  assign n11134 = n10363 & ~n11133 ;
  assign n11137 = ~n10416 & ~n11005 ;
  assign n11131 = n10389 & n10414 ;
  assign n11135 = ~n10363 & n10369 ;
  assign n11136 = n10408 & n11135 ;
  assign n11138 = ~n11131 & ~n11136 ;
  assign n11139 = n11137 & n11138 ;
  assign n11140 = ~n11134 & n11139 ;
  assign n11141 = ~n10405 & ~n11140 ;
  assign n11142 = n10363 & n10440 ;
  assign n11143 = ~n11136 & ~n11142 ;
  assign n11144 = n10382 & ~n11143 ;
  assign n11159 = ~n10433 & ~n11144 ;
  assign n11160 = ~n11141 & n11159 ;
  assign n11161 = ~n11150 & n11160 ;
  assign n11162 = ~n11158 & n11161 ;
  assign n11163 = \u2_L10_reg[23]/NET0131  & ~n11162 ;
  assign n11164 = ~\u2_L10_reg[23]/NET0131  & n11162 ;
  assign n11165 = ~n11163 & ~n11164 ;
  assign n11198 = decrypt_pad & ~\u2_uk_K_r10_reg[2]/NET0131  ;
  assign n11199 = ~decrypt_pad & ~\u2_uk_K_r10_reg[7]/NET0131  ;
  assign n11200 = ~n11198 & ~n11199 ;
  assign n11201 = \u2_R10_reg[19]/NET0131  & ~n11200 ;
  assign n11202 = ~\u2_R10_reg[19]/NET0131  & n11200 ;
  assign n11203 = ~n11201 & ~n11202 ;
  assign n11166 = decrypt_pad & ~\u2_uk_K_r10_reg[15]/NET0131  ;
  assign n11167 = ~decrypt_pad & ~\u2_uk_K_r10_reg[51]/NET0131  ;
  assign n11168 = ~n11166 & ~n11167 ;
  assign n11169 = \u2_R10_reg[18]/NET0131  & ~n11168 ;
  assign n11170 = ~\u2_R10_reg[18]/NET0131  & n11168 ;
  assign n11171 = ~n11169 & ~n11170 ;
  assign n11179 = decrypt_pad & ~\u2_uk_K_r10_reg[21]/NET0131  ;
  assign n11180 = ~decrypt_pad & ~\u2_uk_K_r10_reg[2]/NET0131  ;
  assign n11181 = ~n11179 & ~n11180 ;
  assign n11182 = \u2_R10_reg[17]/NET0131  & ~n11181 ;
  assign n11183 = ~\u2_R10_reg[17]/NET0131  & n11181 ;
  assign n11184 = ~n11182 & ~n11183 ;
  assign n11193 = ~n11171 & n11184 ;
  assign n11172 = decrypt_pad & ~\u2_uk_K_r10_reg[42]/NET0131  ;
  assign n11173 = ~decrypt_pad & ~\u2_uk_K_r10_reg[23]/NET0131  ;
  assign n11174 = ~n11172 & ~n11173 ;
  assign n11175 = \u2_R10_reg[21]/NET0131  & ~n11174 ;
  assign n11176 = ~\u2_R10_reg[21]/NET0131  & n11174 ;
  assign n11177 = ~n11175 & ~n11176 ;
  assign n11205 = ~n11171 & ~n11177 ;
  assign n11185 = decrypt_pad & ~\u2_uk_K_r10_reg[30]/NET0131  ;
  assign n11186 = ~decrypt_pad & ~\u2_uk_K_r10_reg[35]/NET0131  ;
  assign n11187 = ~n11185 & ~n11186 ;
  assign n11188 = \u2_R10_reg[16]/NET0131  & ~n11187 ;
  assign n11189 = ~\u2_R10_reg[16]/NET0131  & n11187 ;
  assign n11190 = ~n11188 & ~n11189 ;
  assign n11206 = ~n11177 & ~n11190 ;
  assign n11207 = ~n11205 & ~n11206 ;
  assign n11208 = ~n11193 & ~n11207 ;
  assign n11209 = ~n11184 & ~n11190 ;
  assign n11191 = n11184 & n11190 ;
  assign n11210 = n11177 & n11191 ;
  assign n11211 = ~n11209 & ~n11210 ;
  assign n11212 = ~n11208 & n11211 ;
  assign n11213 = n11203 & ~n11212 ;
  assign n11194 = ~n11190 & n11193 ;
  assign n11195 = n11177 & n11190 ;
  assign n11196 = ~n11184 & n11195 ;
  assign n11197 = ~n11194 & ~n11196 ;
  assign n11204 = ~n11197 & ~n11203 ;
  assign n11178 = ~n11171 & n11177 ;
  assign n11214 = ~n11177 & n11190 ;
  assign n11215 = ~n11178 & ~n11214 ;
  assign n11216 = n11184 & ~n11205 ;
  assign n11217 = ~n11215 & n11216 ;
  assign n11218 = ~n11204 & ~n11217 ;
  assign n11219 = ~n11213 & n11218 ;
  assign n11220 = decrypt_pad & ~\u2_uk_K_r10_reg[45]/P0001  ;
  assign n11221 = ~decrypt_pad & ~\u2_uk_K_r10_reg[22]/NET0131  ;
  assign n11222 = ~n11220 & ~n11221 ;
  assign n11223 = \u2_R10_reg[20]/NET0131  & ~n11222 ;
  assign n11224 = ~\u2_R10_reg[20]/NET0131  & n11222 ;
  assign n11225 = ~n11223 & ~n11224 ;
  assign n11226 = ~n11219 & n11225 ;
  assign n11240 = ~n11184 & n11206 ;
  assign n11241 = ~n11177 & n11191 ;
  assign n11242 = ~n11240 & ~n11241 ;
  assign n11243 = n11171 & ~n11242 ;
  assign n11244 = n11177 & n11209 ;
  assign n11245 = ~n11171 & n11244 ;
  assign n11246 = ~n11243 & ~n11245 ;
  assign n11247 = n11203 & ~n11246 ;
  assign n11227 = n11184 & ~n11190 ;
  assign n11228 = n11171 & n11227 ;
  assign n11229 = ~n11184 & n11214 ;
  assign n11230 = ~n11228 & ~n11229 ;
  assign n11231 = ~n11177 & n11203 ;
  assign n11232 = ~n11230 & ~n11231 ;
  assign n11234 = ~n11177 & n11184 ;
  assign n11235 = n11203 & ~n11234 ;
  assign n11233 = ~n11203 & ~n11209 ;
  assign n11236 = ~n11171 & ~n11233 ;
  assign n11237 = ~n11235 & n11236 ;
  assign n11238 = ~n11232 & ~n11237 ;
  assign n11239 = ~n11225 & ~n11238 ;
  assign n11192 = n11178 & n11191 ;
  assign n11248 = ~n11184 & n11190 ;
  assign n11249 = n11171 & ~n11203 ;
  assign n11250 = n11248 & n11249 ;
  assign n11251 = ~n11192 & ~n11250 ;
  assign n11252 = ~n11239 & n11251 ;
  assign n11253 = ~n11247 & n11252 ;
  assign n11254 = ~n11226 & n11253 ;
  assign n11255 = ~\u2_L10_reg[25]/NET0131  & ~n11254 ;
  assign n11256 = \u2_L10_reg[25]/NET0131  & n11254 ;
  assign n11257 = ~n11255 & ~n11256 ;
  assign n11259 = ~n10652 & ~n10704 ;
  assign n11260 = ~n10732 & n11259 ;
  assign n11258 = n10699 & ~n10721 ;
  assign n11261 = ~n10728 & ~n11258 ;
  assign n11262 = n11260 & n11261 ;
  assign n11268 = n10671 & n10693 ;
  assign n11269 = ~n10722 & ~n10727 ;
  assign n11270 = ~n11268 & n11269 ;
  assign n11271 = n10687 & ~n11270 ;
  assign n11264 = n10665 & n10687 ;
  assign n11265 = n10690 & n10695 ;
  assign n11266 = ~n11264 & ~n11265 ;
  assign n11267 = ~n10678 & ~n11266 ;
  assign n11263 = n10681 & ~n10687 ;
  assign n11272 = n10652 & ~n10702 ;
  assign n11273 = ~n11263 & n11272 ;
  assign n11274 = ~n11267 & n11273 ;
  assign n11275 = ~n11271 & n11274 ;
  assign n11276 = ~n11262 & ~n11275 ;
  assign n11277 = ~n10664 & ~n10724 ;
  assign n11278 = ~n10672 & ~n11277 ;
  assign n11279 = ~n10687 & ~n11278 ;
  assign n11280 = ~n10689 & ~n11055 ;
  assign n11281 = ~n10652 & ~n11280 ;
  assign n11282 = ~n10678 & ~n11281 ;
  assign n11283 = ~n11279 & n11282 ;
  assign n11284 = n10678 & ~n10705 ;
  assign n11285 = ~n10728 & n11284 ;
  assign n11286 = ~n11283 & ~n11285 ;
  assign n11287 = ~n11276 & ~n11286 ;
  assign n11288 = ~\u2_L10_reg[26]/NET0131  & ~n11287 ;
  assign n11289 = \u2_L10_reg[26]/NET0131  & n11287 ;
  assign n11290 = ~n11288 & ~n11289 ;
  assign n11315 = n10793 & n10815 ;
  assign n11316 = ~n10813 & ~n10818 ;
  assign n11317 = ~n11315 & n11316 ;
  assign n11318 = n10756 & ~n11317 ;
  assign n11300 = n10775 & n10785 ;
  assign n11301 = ~n10782 & n10823 ;
  assign n11302 = ~n11300 & ~n11301 ;
  assign n11314 = ~n10756 & ~n11302 ;
  assign n11311 = n10756 & n10762 ;
  assign n11312 = ~n10776 & ~n11311 ;
  assign n11313 = ~n10782 & ~n11312 ;
  assign n11319 = n10785 & n10806 ;
  assign n11320 = ~n11313 & ~n11319 ;
  assign n11321 = ~n11314 & n11320 ;
  assign n11322 = ~n11318 & n11321 ;
  assign n11323 = n10750 & ~n11322 ;
  assign n11291 = ~n10768 & n10788 ;
  assign n11292 = n10782 & n11291 ;
  assign n11293 = ~n10775 & n10815 ;
  assign n11294 = ~n11292 & ~n11293 ;
  assign n11295 = ~n10756 & ~n11294 ;
  assign n11304 = ~n10775 & ~n10785 ;
  assign n11305 = ~n10787 & n11304 ;
  assign n11306 = ~n11291 & ~n11305 ;
  assign n11307 = n10782 & ~n11306 ;
  assign n11296 = ~n10782 & n10787 ;
  assign n11297 = ~n10786 & ~n10788 ;
  assign n11298 = ~n11296 & n11297 ;
  assign n11299 = ~n10756 & ~n11298 ;
  assign n11303 = n10756 & ~n11302 ;
  assign n11308 = ~n11299 & ~n11303 ;
  assign n11309 = ~n11307 & n11308 ;
  assign n11310 = ~n10750 & ~n11309 ;
  assign n11324 = ~n11295 & ~n11310 ;
  assign n11325 = ~n11323 & n11324 ;
  assign n11326 = ~\u2_L10_reg[28]/NET0131  & ~n11325 ;
  assign n11327 = \u2_L10_reg[28]/NET0131  & n11325 ;
  assign n11328 = ~n11326 & ~n11327 ;
  assign n11329 = n11171 & n11229 ;
  assign n11330 = ~n11203 & ~n11329 ;
  assign n11331 = n11171 & n11244 ;
  assign n11333 = n11178 & n11227 ;
  assign n11332 = n11171 & n11234 ;
  assign n11334 = n11203 & ~n11332 ;
  assign n11335 = ~n11333 & n11334 ;
  assign n11336 = ~n11331 & n11335 ;
  assign n11337 = ~n11330 & ~n11336 ;
  assign n11343 = ~n11177 & n11228 ;
  assign n11344 = ~n11331 & ~n11343 ;
  assign n11340 = n11205 & n11209 ;
  assign n11341 = ~n11196 & ~n11340 ;
  assign n11342 = n11203 & ~n11341 ;
  assign n11338 = ~n11171 & ~n11203 ;
  assign n11339 = n11190 & n11338 ;
  assign n11345 = n11225 & ~n11339 ;
  assign n11346 = ~n11342 & n11345 ;
  assign n11347 = n11344 & n11346 ;
  assign n11348 = n11205 & n11248 ;
  assign n11349 = n11203 & ~n11348 ;
  assign n11350 = ~n11196 & ~n11203 ;
  assign n11351 = n11177 & n11227 ;
  assign n11352 = n11178 & ~n11190 ;
  assign n11353 = ~n11351 & ~n11352 ;
  assign n11354 = n11350 & n11353 ;
  assign n11355 = ~n11349 & ~n11354 ;
  assign n11356 = n11203 & n11210 ;
  assign n11357 = ~n11194 & ~n11225 ;
  assign n11358 = ~n11356 & n11357 ;
  assign n11359 = ~n11243 & n11358 ;
  assign n11360 = ~n11355 & n11359 ;
  assign n11361 = ~n11347 & ~n11360 ;
  assign n11362 = ~n11337 & ~n11361 ;
  assign n11363 = ~\u2_L10_reg[8]/NET0131  & ~n11362 ;
  assign n11364 = \u2_L10_reg[8]/NET0131  & n11362 ;
  assign n11365 = ~n11363 & ~n11364 ;
  assign n11368 = n10693 & ~n11065 ;
  assign n11369 = ~n10728 & ~n11368 ;
  assign n11370 = ~n10678 & ~n11369 ;
  assign n11366 = ~n10681 & ~n10705 ;
  assign n11367 = n10678 & ~n11366 ;
  assign n11371 = n11057 & ~n11367 ;
  assign n11372 = ~n11370 & n11371 ;
  assign n11373 = n10652 & ~n11372 ;
  assign n11374 = ~n10689 & ~n10715 ;
  assign n11375 = n10678 & ~n11374 ;
  assign n11376 = ~n10713 & ~n11065 ;
  assign n11377 = ~n11375 & n11376 ;
  assign n11378 = n10658 & ~n11377 ;
  assign n11379 = ~n10687 & n10722 ;
  assign n11380 = ~n10730 & ~n11379 ;
  assign n11381 = n10692 & n11380 ;
  assign n11382 = ~n11378 & n11381 ;
  assign n11383 = ~n10652 & ~n11382 ;
  assign n11384 = ~n10691 & n11057 ;
  assign n11385 = ~n10678 & ~n11384 ;
  assign n11386 = ~n10700 & ~n10720 ;
  assign n11387 = ~n11385 & n11386 ;
  assign n11388 = ~n11383 & n11387 ;
  assign n11389 = ~n11373 & n11388 ;
  assign n11390 = ~\u2_L10_reg[10]/NET0131  & ~n11389 ;
  assign n11391 = \u2_L10_reg[10]/NET0131  & n11389 ;
  assign n11392 = ~n11390 & ~n11391 ;
  assign n11393 = ~n10488 & n10522 ;
  assign n11401 = ~n10515 & ~n11393 ;
  assign n11394 = n10480 & n10504 ;
  assign n11395 = n10472 & ~n10528 ;
  assign n11396 = n10503 & ~n11395 ;
  assign n11402 = ~n11394 & ~n11396 ;
  assign n11397 = ~n10519 & ~n10534 ;
  assign n11398 = n10466 & ~n11397 ;
  assign n11399 = ~n10472 & ~n10490 ;
  assign n11400 = ~n10528 & n11399 ;
  assign n11403 = ~n11398 & ~n11400 ;
  assign n11404 = n11402 & n11403 ;
  assign n11405 = n11401 & n11404 ;
  assign n11410 = n10502 & n10505 ;
  assign n11414 = n10515 & ~n11410 ;
  assign n11415 = ~n10523 & n11414 ;
  assign n11416 = ~n10530 & n11415 ;
  assign n11407 = ~n10479 & ~n10494 ;
  assign n11406 = ~n10465 & ~n10499 ;
  assign n11408 = n10472 & ~n11406 ;
  assign n11409 = ~n11407 & n11408 ;
  assign n11411 = ~n10459 & n10465 ;
  assign n11412 = ~n10473 & ~n11411 ;
  assign n11413 = n10495 & ~n11412 ;
  assign n11417 = ~n11409 & ~n11413 ;
  assign n11418 = n11416 & n11417 ;
  assign n11419 = ~n11405 & ~n11418 ;
  assign n11420 = \u2_L10_reg[12]/NET0131  & n11419 ;
  assign n11421 = ~\u2_L10_reg[12]/NET0131  & ~n11419 ;
  assign n11422 = ~n11420 & ~n11421 ;
  assign n11429 = ~n11192 & ~n11244 ;
  assign n11430 = ~n11332 & ~n11348 ;
  assign n11431 = n11429 & n11430 ;
  assign n11432 = ~n11203 & ~n11431 ;
  assign n11423 = n11171 & n11195 ;
  assign n11424 = ~n11194 & ~n11423 ;
  assign n11425 = ~n11240 & n11424 ;
  assign n11426 = n11203 & ~n11425 ;
  assign n11427 = ~n11193 & ~n11248 ;
  assign n11428 = n11215 & ~n11427 ;
  assign n11433 = ~n11426 & ~n11428 ;
  assign n11434 = ~n11432 & n11433 ;
  assign n11435 = ~n11225 & ~n11434 ;
  assign n11438 = n11191 & n11205 ;
  assign n11444 = ~n11329 & ~n11438 ;
  assign n11436 = ~n11171 & n11196 ;
  assign n11437 = n11210 & n11249 ;
  assign n11445 = ~n11436 & ~n11437 ;
  assign n11446 = n11444 & n11445 ;
  assign n11439 = ~n11240 & ~n11351 ;
  assign n11440 = n11338 & ~n11439 ;
  assign n11441 = ~n11177 & ~n11191 ;
  assign n11442 = n11203 & ~n11441 ;
  assign n11443 = n11424 & n11442 ;
  assign n11447 = ~n11440 & ~n11443 ;
  assign n11448 = n11446 & n11447 ;
  assign n11449 = n11225 & ~n11448 ;
  assign n11450 = n11171 & ~n11184 ;
  assign n11451 = n11206 & n11450 ;
  assign n11452 = ~n11438 & ~n11451 ;
  assign n11453 = n11203 & ~n11452 ;
  assign n11454 = ~n11203 & ~n11344 ;
  assign n11455 = ~n11453 & ~n11454 ;
  assign n11456 = ~n11449 & n11455 ;
  assign n11457 = ~n11435 & n11456 ;
  assign n11458 = ~\u2_L10_reg[14]/NET0131  & ~n11457 ;
  assign n11459 = \u2_L10_reg[14]/NET0131  & n11457 ;
  assign n11460 = ~n11458 & ~n11459 ;
  assign n11479 = ~n10768 & n10798 ;
  assign n11480 = n10756 & ~n10796 ;
  assign n11481 = ~n11479 & n11480 ;
  assign n11482 = ~n10756 & ~n10776 ;
  assign n11483 = ~n10807 & n11482 ;
  assign n11484 = ~n11481 & ~n11483 ;
  assign n11461 = ~n10814 & ~n11292 ;
  assign n11485 = n10775 & n11301 ;
  assign n11486 = n10801 & ~n11485 ;
  assign n11487 = n11461 & n11486 ;
  assign n11488 = ~n11484 & n11487 ;
  assign n11489 = n10750 & ~n11488 ;
  assign n11462 = ~n10762 & n10793 ;
  assign n11463 = ~n11319 & ~n11462 ;
  assign n11464 = ~n10819 & n11463 ;
  assign n11465 = ~n10750 & ~n11464 ;
  assign n11466 = n11461 & ~n11465 ;
  assign n11467 = ~n10756 & ~n11466 ;
  assign n11468 = n10787 & n10809 ;
  assign n11469 = ~n11305 & ~n11468 ;
  assign n11470 = n10756 & ~n11469 ;
  assign n11471 = n10782 & ~n10793 ;
  assign n11472 = n11311 & n11471 ;
  assign n11473 = ~n10756 & ~n10775 ;
  assign n11474 = ~n10782 & n10785 ;
  assign n11475 = ~n11473 & n11474 ;
  assign n11476 = ~n11472 & ~n11475 ;
  assign n11477 = ~n11470 & n11476 ;
  assign n11478 = ~n10750 & ~n11477 ;
  assign n11490 = ~n11467 & ~n11478 ;
  assign n11491 = ~n11489 & n11490 ;
  assign n11492 = ~\u2_L10_reg[13]/NET0131  & n11491 ;
  assign n11493 = \u2_L10_reg[13]/NET0131  & ~n11491 ;
  assign n11494 = ~n11492 & ~n11493 ;
  assign n11495 = n10878 & n10890 ;
  assign n11496 = ~n10898 & ~n11495 ;
  assign n11497 = ~n10912 & n11496 ;
  assign n11498 = n10904 & ~n11497 ;
  assign n11499 = n10914 & n10940 ;
  assign n11500 = ~n11498 & ~n11499 ;
  assign n11501 = ~n10930 & ~n11500 ;
  assign n11511 = ~n10891 & n10897 ;
  assign n11512 = ~n10898 & ~n11511 ;
  assign n11513 = ~n10878 & ~n10913 ;
  assign n11514 = n11512 & n11513 ;
  assign n11515 = ~n10904 & ~n11093 ;
  assign n11516 = ~n11514 & n11515 ;
  assign n11517 = n10904 & ~n10949 ;
  assign n11518 = ~n11105 & n11517 ;
  assign n11519 = ~n11516 & ~n11518 ;
  assign n11505 = ~n10884 & n11495 ;
  assign n11503 = n10897 & ~n10904 ;
  assign n11504 = n10913 & n11503 ;
  assign n11506 = ~n11114 & ~n11504 ;
  assign n11507 = ~n11505 & n11506 ;
  assign n11502 = n10904 & n11106 ;
  assign n11508 = ~n10939 & ~n11502 ;
  assign n11509 = n11507 & n11508 ;
  assign n11510 = n10930 & ~n11509 ;
  assign n11520 = ~n10904 & ~n10930 ;
  assign n11521 = n10933 & n11520 ;
  assign n11522 = ~n11510 & ~n11521 ;
  assign n11523 = ~n11519 & n11522 ;
  assign n11524 = ~n11501 & n11523 ;
  assign n11525 = ~\u2_L10_reg[15]/NET0131  & ~n11524 ;
  assign n11526 = \u2_L10_reg[15]/NET0131  & n11524 ;
  assign n11527 = ~n11525 & ~n11526 ;
  assign n11538 = n10904 & ~n10938 ;
  assign n11539 = n11512 & n11538 ;
  assign n11540 = n10932 & n10951 ;
  assign n11541 = ~n10945 & ~n11540 ;
  assign n11542 = ~n11096 & n11541 ;
  assign n11543 = ~n11539 & n11542 ;
  assign n11544 = ~n10930 & ~n11543 ;
  assign n11528 = ~n10936 & ~n10958 ;
  assign n11529 = ~n11110 & n11528 ;
  assign n11530 = ~n10904 & ~n11529 ;
  assign n11531 = n10904 & ~n10914 ;
  assign n11532 = ~n11496 & n11531 ;
  assign n11533 = ~n10915 & ~n10941 ;
  assign n11534 = ~n10949 & n11533 ;
  assign n11535 = ~n11532 & n11534 ;
  assign n11536 = ~n11530 & n11535 ;
  assign n11537 = n10930 & ~n11536 ;
  assign n11547 = ~n10904 & ~n10943 ;
  assign n11545 = ~n10897 & n10904 ;
  assign n11546 = n10913 & n11545 ;
  assign n11548 = ~n10937 & ~n11546 ;
  assign n11549 = ~n11547 & n11548 ;
  assign n11550 = ~n11537 & n11549 ;
  assign n11551 = ~n11544 & n11550 ;
  assign n11552 = ~\u2_L10_reg[27]/NET0131  & ~n11551 ;
  assign n11553 = \u2_L10_reg[27]/NET0131  & n11551 ;
  assign n11554 = ~n11552 & ~n11553 ;
  assign n11555 = ~n10466 & ~n11411 ;
  assign n11556 = n10499 & ~n11555 ;
  assign n11557 = n10503 & n10528 ;
  assign n11558 = ~n10472 & ~n10522 ;
  assign n11559 = ~n11557 & n11558 ;
  assign n11560 = ~n11556 & n11559 ;
  assign n11561 = n10492 & ~n11407 ;
  assign n11562 = n10488 & n11411 ;
  assign n11563 = n10472 & ~n11562 ;
  assign n11564 = ~n11561 & n11563 ;
  assign n11565 = ~n11560 & ~n11564 ;
  assign n11566 = n10479 & n11562 ;
  assign n11567 = ~n11565 & ~n11566 ;
  assign n11568 = n10515 & ~n11567 ;
  assign n11572 = n10465 & n10520 ;
  assign n11573 = n11400 & ~n11572 ;
  assign n11570 = ~n10534 & ~n11555 ;
  assign n11571 = ~n10492 & n11570 ;
  assign n11569 = n10534 & n11555 ;
  assign n11574 = ~n10520 & ~n10528 ;
  assign n11575 = n10500 & ~n11574 ;
  assign n11576 = ~n11569 & ~n11575 ;
  assign n11577 = ~n11571 & n11576 ;
  assign n11578 = ~n11573 & n11577 ;
  assign n11579 = ~n10515 & ~n11578 ;
  assign n11580 = n10472 & n10524 ;
  assign n11581 = n10517 & ~n11411 ;
  assign n11582 = n10504 & n11581 ;
  assign n11583 = ~n11580 & ~n11582 ;
  assign n11584 = ~n11579 & n11583 ;
  assign n11585 = ~n11568 & n11584 ;
  assign n11586 = \u2_L10_reg[32]/NET0131  & n11585 ;
  assign n11587 = ~\u2_L10_reg[32]/NET0131  & ~n11585 ;
  assign n11588 = ~n11586 & ~n11587 ;
  assign n11590 = ~n11215 & n11350 ;
  assign n11591 = n11203 & ~n11241 ;
  assign n11592 = ~n11352 & n11591 ;
  assign n11593 = ~n11590 & ~n11592 ;
  assign n11589 = ~n11214 & n11450 ;
  assign n11594 = ~n11225 & ~n11589 ;
  assign n11595 = ~n11593 & n11594 ;
  assign n11597 = n11178 & n11190 ;
  assign n11598 = n11184 & n11206 ;
  assign n11599 = ~n11597 & ~n11598 ;
  assign n11600 = n11203 & ~n11599 ;
  assign n11596 = ~n11203 & n11351 ;
  assign n11601 = ~n11192 & n11225 ;
  assign n11602 = ~n11329 & n11601 ;
  assign n11603 = ~n11596 & n11602 ;
  assign n11604 = ~n11600 & n11603 ;
  assign n11605 = ~n11595 & ~n11604 ;
  assign n11606 = ~n11331 & n11349 ;
  assign n11607 = n11171 & n11196 ;
  assign n11608 = ~n11203 & ~n11340 ;
  assign n11609 = ~n11438 & n11608 ;
  assign n11610 = ~n11607 & n11609 ;
  assign n11611 = ~n11606 & ~n11610 ;
  assign n11612 = ~n11605 & ~n11611 ;
  assign n11613 = ~\u2_L10_reg[3]/NET0131  & ~n11612 ;
  assign n11614 = \u2_L10_reg[3]/NET0131  & n11612 ;
  assign n11615 = ~n11613 & ~n11614 ;
  assign n11616 = decrypt_pad & ~\u2_uk_K_r10_reg[25]/NET0131  ;
  assign n11617 = ~decrypt_pad & ~\u2_uk_K_r10_reg[34]/NET0131  ;
  assign n11618 = ~n11616 & ~n11617 ;
  assign n11619 = \u2_R10_reg[10]/NET0131  & ~n11618 ;
  assign n11620 = ~\u2_R10_reg[10]/NET0131  & n11618 ;
  assign n11621 = ~n11619 & ~n11620 ;
  assign n11622 = decrypt_pad & ~\u2_uk_K_r10_reg[17]/NET0131  ;
  assign n11623 = ~decrypt_pad & ~\u2_uk_K_r10_reg[26]/NET0131  ;
  assign n11624 = ~n11622 & ~n11623 ;
  assign n11625 = \u2_R10_reg[9]/NET0131  & ~n11624 ;
  assign n11626 = ~\u2_R10_reg[9]/NET0131  & n11624 ;
  assign n11627 = ~n11625 & ~n11626 ;
  assign n11628 = n11621 & ~n11627 ;
  assign n11629 = decrypt_pad & ~\u2_uk_K_r10_reg[54]/NET0131  ;
  assign n11630 = ~decrypt_pad & ~\u2_uk_K_r10_reg[6]/NET0131  ;
  assign n11631 = ~n11629 & ~n11630 ;
  assign n11632 = \u2_R10_reg[13]/NET0131  & ~n11631 ;
  assign n11633 = ~\u2_R10_reg[13]/NET0131  & n11631 ;
  assign n11634 = ~n11632 & ~n11633 ;
  assign n11635 = n11628 & n11634 ;
  assign n11636 = decrypt_pad & ~\u2_uk_K_r10_reg[20]/NET0131  ;
  assign n11637 = ~decrypt_pad & ~\u2_uk_K_r10_reg[54]/NET0131  ;
  assign n11638 = ~n11636 & ~n11637 ;
  assign n11639 = \u2_R10_reg[8]/NET0131  & ~n11638 ;
  assign n11640 = ~\u2_R10_reg[8]/NET0131  & n11638 ;
  assign n11641 = ~n11639 & ~n11640 ;
  assign n11642 = ~n11634 & ~n11641 ;
  assign n11643 = ~n11621 & ~n11627 ;
  assign n11644 = n11642 & n11643 ;
  assign n11645 = ~n11635 & ~n11644 ;
  assign n11646 = decrypt_pad & ~\u2_uk_K_r10_reg[26]/NET0131  ;
  assign n11647 = ~decrypt_pad & ~\u2_uk_K_r10_reg[3]/NET0131  ;
  assign n11648 = ~n11646 & ~n11647 ;
  assign n11649 = \u2_R10_reg[11]/NET0131  & ~n11648 ;
  assign n11650 = ~\u2_R10_reg[11]/NET0131  & n11648 ;
  assign n11651 = ~n11649 & ~n11650 ;
  assign n11652 = ~n11645 & n11651 ;
  assign n11657 = ~n11621 & ~n11641 ;
  assign n11658 = n11634 & n11641 ;
  assign n11659 = ~n11642 & ~n11658 ;
  assign n11660 = ~n11657 & n11659 ;
  assign n11661 = n11627 & ~n11660 ;
  assign n11656 = ~n11627 & ~n11634 ;
  assign n11662 = n11651 & ~n11656 ;
  assign n11663 = ~n11661 & n11662 ;
  assign n11653 = n11621 & ~n11641 ;
  assign n11664 = n11627 & n11634 ;
  assign n11665 = ~n11653 & n11664 ;
  assign n11666 = ~n11627 & n11641 ;
  assign n11667 = ~n11634 & n11666 ;
  assign n11668 = ~n11665 & ~n11667 ;
  assign n11669 = ~n11651 & ~n11668 ;
  assign n11654 = n11627 & ~n11634 ;
  assign n11655 = n11653 & n11654 ;
  assign n11670 = decrypt_pad & ~\u2_uk_K_r10_reg[41]/NET0131  ;
  assign n11671 = ~decrypt_pad & ~\u2_uk_K_r10_reg[18]/NET0131  ;
  assign n11672 = ~n11670 & ~n11671 ;
  assign n11673 = \u2_R10_reg[12]/NET0131  & ~n11672 ;
  assign n11674 = ~\u2_R10_reg[12]/NET0131  & n11672 ;
  assign n11675 = ~n11673 & ~n11674 ;
  assign n11676 = ~n11655 & n11675 ;
  assign n11677 = ~n11669 & n11676 ;
  assign n11678 = ~n11663 & n11677 ;
  assign n11686 = n11628 & ~n11659 ;
  assign n11679 = ~n11651 & n11664 ;
  assign n11680 = n11653 & n11679 ;
  assign n11687 = n11621 & n11641 ;
  assign n11688 = n11654 & n11687 ;
  assign n11689 = ~n11675 & ~n11688 ;
  assign n11690 = ~n11680 & n11689 ;
  assign n11691 = ~n11686 & n11690 ;
  assign n11681 = ~n11641 & n11651 ;
  assign n11682 = n11659 & ~n11681 ;
  assign n11683 = n11643 & n11682 ;
  assign n11684 = ~n11621 & n11627 ;
  assign n11685 = ~n11682 & n11684 ;
  assign n11692 = ~n11683 & ~n11685 ;
  assign n11693 = n11691 & n11692 ;
  assign n11694 = ~n11678 & ~n11693 ;
  assign n11695 = ~n11652 & ~n11694 ;
  assign n11696 = ~\u2_L10_reg[6]/NET0131  & ~n11695 ;
  assign n11697 = \u2_L10_reg[6]/NET0131  & n11695 ;
  assign n11698 = ~n11696 & ~n11697 ;
  assign n11700 = ~n10465 & ~n10535 ;
  assign n11699 = n10479 & ~n11555 ;
  assign n11701 = ~n11562 & ~n11699 ;
  assign n11702 = ~n11700 & n11701 ;
  assign n11703 = ~n10472 & ~n11702 ;
  assign n11704 = ~n10529 & ~n11699 ;
  assign n11705 = n10488 & ~n11704 ;
  assign n11706 = ~n10480 & ~n10488 ;
  assign n11707 = n11555 & n11706 ;
  assign n11708 = n10472 & n11707 ;
  assign n11709 = ~n11705 & ~n11708 ;
  assign n11710 = ~n11703 & n11709 ;
  assign n11711 = n10515 & ~n11710 ;
  assign n11712 = n10488 & ~n10528 ;
  assign n11713 = n11555 & n11712 ;
  assign n11714 = ~n11570 & ~n11713 ;
  assign n11715 = n10472 & ~n11714 ;
  assign n11716 = ~n10472 & n11707 ;
  assign n11717 = ~n10496 & ~n11716 ;
  assign n11718 = ~n11715 & n11717 ;
  assign n11719 = ~n10515 & ~n11718 ;
  assign n11720 = n10472 & n10496 ;
  assign n11721 = ~n10472 & n11705 ;
  assign n11722 = ~n11720 & ~n11721 ;
  assign n11723 = ~n11719 & n11722 ;
  assign n11724 = ~n11711 & n11723 ;
  assign n11725 = ~\u2_L10_reg[7]/NET0131  & ~n11724 ;
  assign n11726 = \u2_L10_reg[7]/NET0131  & n11724 ;
  assign n11727 = ~n11725 & ~n11726 ;
  assign n11728 = ~n10391 & ~n10436 ;
  assign n11729 = n10414 & ~n11728 ;
  assign n11732 = n11021 & n11152 ;
  assign n11733 = n10369 & ~n11732 ;
  assign n11730 = ~n10393 & ~n11145 ;
  assign n11731 = n10423 & ~n11730 ;
  assign n11734 = n11007 & ~n11731 ;
  assign n11735 = ~n11733 & n11734 ;
  assign n11736 = ~n10396 & ~n10434 ;
  assign n11737 = ~n11132 & n11736 ;
  assign n11738 = n10363 & ~n11737 ;
  assign n11741 = ~n10363 & ~n11730 ;
  assign n11740 = n10369 & n11014 ;
  assign n11739 = ~n10369 & n11020 ;
  assign n11742 = ~n10405 & ~n11739 ;
  assign n11743 = ~n11740 & n11742 ;
  assign n11744 = ~n11741 & n11743 ;
  assign n11745 = ~n11738 & n11744 ;
  assign n11746 = ~n11735 & ~n11745 ;
  assign n11747 = ~n11729 & ~n11746 ;
  assign n11748 = ~\u2_L10_reg[9]/NET0131  & ~n11747 ;
  assign n11749 = \u2_L10_reg[9]/NET0131  & n11747 ;
  assign n11750 = ~n11748 & ~n11749 ;
  assign n11754 = n10756 & ~n10794 ;
  assign n11751 = n10769 & ~n10782 ;
  assign n11752 = ~n10818 & ~n11751 ;
  assign n11753 = ~n10756 & ~n11752 ;
  assign n11755 = ~n10808 & ~n11753 ;
  assign n11756 = ~n11754 & n11755 ;
  assign n11757 = n10750 & ~n11756 ;
  assign n11758 = n10769 & n10816 ;
  assign n11762 = ~n11479 & ~n11758 ;
  assign n11763 = ~n10783 & n11762 ;
  assign n11759 = ~n10762 & ~n10806 ;
  assign n11760 = ~n10809 & ~n10816 ;
  assign n11761 = n11759 & n11760 ;
  assign n11764 = ~n11292 & ~n11761 ;
  assign n11765 = n11763 & n11764 ;
  assign n11766 = ~n10750 & ~n11765 ;
  assign n11767 = ~n10756 & n11300 ;
  assign n11768 = n10769 & n10782 ;
  assign n11769 = ~n11485 & ~n11768 ;
  assign n11770 = n10756 & ~n11769 ;
  assign n11771 = ~n11767 & ~n11770 ;
  assign n11772 = ~n11766 & n11771 ;
  assign n11773 = ~n11757 & n11772 ;
  assign n11774 = ~\u2_L10_reg[18]/P0001  & ~n11773 ;
  assign n11775 = \u2_L10_reg[18]/P0001  & n11773 ;
  assign n11776 = ~n11774 & ~n11775 ;
  assign n11778 = n11643 & ~n11659 ;
  assign n11779 = n11660 & ~n11666 ;
  assign n11780 = ~n11778 & ~n11779 ;
  assign n11781 = ~n11651 & ~n11780 ;
  assign n11782 = ~n11675 & ~n11781 ;
  assign n11783 = ~n11621 & n11651 ;
  assign n11784 = ~n11656 & ~n11666 ;
  assign n11785 = n11783 & ~n11784 ;
  assign n11791 = n11675 & ~n11785 ;
  assign n11786 = ~n11642 & n11651 ;
  assign n11787 = n11621 & ~n11666 ;
  assign n11788 = n11786 & n11787 ;
  assign n11789 = ~n11643 & ~n11651 ;
  assign n11790 = ~n11659 & n11789 ;
  assign n11792 = ~n11788 & ~n11790 ;
  assign n11793 = n11791 & n11792 ;
  assign n11794 = ~n11683 & n11793 ;
  assign n11795 = ~n11782 & ~n11794 ;
  assign n11796 = n11634 & n11657 ;
  assign n11797 = ~n11634 & n11653 ;
  assign n11798 = ~n11796 & ~n11797 ;
  assign n11799 = n11627 & n11642 ;
  assign n11800 = ~n11627 & n11687 ;
  assign n11801 = ~n11799 & ~n11800 ;
  assign n11802 = n11798 & n11801 ;
  assign n11803 = n11651 & ~n11802 ;
  assign n11804 = ~n11634 & n11800 ;
  assign n11805 = ~n11803 & ~n11804 ;
  assign n11806 = ~n11675 & ~n11805 ;
  assign n11777 = n11679 & n11687 ;
  assign n11807 = ~n11664 & ~n11666 ;
  assign n11808 = ~n11658 & n11783 ;
  assign n11809 = ~n11807 & n11808 ;
  assign n11810 = ~n11777 & ~n11809 ;
  assign n11811 = ~n11806 & n11810 ;
  assign n11812 = ~n11795 & n11811 ;
  assign n11813 = ~\u2_L10_reg[24]/NET0131  & ~n11812 ;
  assign n11814 = \u2_L10_reg[24]/NET0131  & n11812 ;
  assign n11815 = ~n11813 & ~n11814 ;
  assign n11818 = ~n11621 & n11667 ;
  assign n11819 = n11798 & ~n11818 ;
  assign n11820 = n11675 & ~n11819 ;
  assign n11821 = ~n11654 & ~n11687 ;
  assign n11816 = n11621 & n11654 ;
  assign n11822 = ~n11675 & ~n11816 ;
  assign n11823 = ~n11821 & n11822 ;
  assign n11824 = ~n11820 & ~n11823 ;
  assign n11825 = n11651 & ~n11824 ;
  assign n11826 = n11627 & ~n11658 ;
  assign n11827 = n11621 & n11826 ;
  assign n11828 = ~n11687 & ~n11799 ;
  assign n11829 = ~n11651 & ~n11828 ;
  assign n11830 = ~n11827 & ~n11829 ;
  assign n11831 = n11675 & ~n11830 ;
  assign n11832 = ~n11651 & ~n11687 ;
  assign n11833 = ~n11807 & n11832 ;
  assign n11834 = ~n11778 & ~n11833 ;
  assign n11835 = ~n11675 & ~n11834 ;
  assign n11817 = ~n11651 & n11816 ;
  assign n11836 = ~n11641 & n11675 ;
  assign n11837 = n11641 & ~n11651 ;
  assign n11838 = ~n11836 & ~n11837 ;
  assign n11839 = n11635 & n11838 ;
  assign n11840 = ~n11817 & ~n11839 ;
  assign n11841 = ~n11835 & n11840 ;
  assign n11842 = ~n11831 & n11841 ;
  assign n11843 = ~n11825 & n11842 ;
  assign n11844 = \u2_L10_reg[30]/NET0131  & ~n11843 ;
  assign n11845 = ~\u2_L10_reg[30]/NET0131  & n11843 ;
  assign n11846 = ~n11844 & ~n11845 ;
  assign n11848 = ~n11627 & n11658 ;
  assign n11849 = ~n11826 & ~n11848 ;
  assign n11850 = ~n11642 & n11849 ;
  assign n11851 = n11654 & n11681 ;
  assign n11852 = ~n11850 & ~n11851 ;
  assign n11853 = ~n11621 & ~n11852 ;
  assign n11847 = n11653 & n11664 ;
  assign n11854 = ~n11634 & ~n11657 ;
  assign n11855 = n11832 & n11854 ;
  assign n11856 = ~n11847 & ~n11855 ;
  assign n11857 = ~n11853 & n11856 ;
  assign n11858 = n11675 & ~n11857 ;
  assign n11859 = n11784 & ~n11826 ;
  assign n11860 = ~n11634 & n11657 ;
  assign n11861 = ~n11859 & ~n11860 ;
  assign n11862 = ~n11675 & ~n11861 ;
  assign n11863 = ~n11800 & ~n11862 ;
  assign n11864 = ~n11651 & ~n11863 ;
  assign n11865 = n11628 & n11642 ;
  assign n11866 = ~n11688 & ~n11865 ;
  assign n11867 = n11651 & ~n11866 ;
  assign n11868 = n11786 & ~n11849 ;
  assign n11869 = ~n11644 & ~n11868 ;
  assign n11870 = ~n11675 & ~n11869 ;
  assign n11871 = ~n11867 & ~n11870 ;
  assign n11872 = ~n11864 & n11871 ;
  assign n11873 = ~n11858 & n11872 ;
  assign n11874 = ~\u2_L10_reg[16]/NET0131  & ~n11873 ;
  assign n11875 = \u2_L10_reg[16]/NET0131  & n11873 ;
  assign n11876 = ~n11874 & ~n11875 ;
  assign n11925 = decrypt_pad & ~\u2_uk_K_r9_reg[50]/NET0131  ;
  assign n11926 = ~decrypt_pad & ~\u2_uk_K_r9_reg[31]/P0001  ;
  assign n11927 = ~n11925 & ~n11926 ;
  assign n11928 = \u2_R9_reg[28]/NET0131  & ~n11927 ;
  assign n11929 = ~\u2_R9_reg[28]/NET0131  & n11927 ;
  assign n11930 = ~n11928 & ~n11929 ;
  assign n11890 = decrypt_pad & ~\u2_uk_K_r9_reg[8]/NET0131  ;
  assign n11891 = ~decrypt_pad & ~\u2_uk_K_r9_reg[16]/NET0131  ;
  assign n11892 = ~n11890 & ~n11891 ;
  assign n11893 = \u2_R9_reg[27]/NET0131  & ~n11892 ;
  assign n11894 = ~\u2_R9_reg[27]/NET0131  & n11892 ;
  assign n11895 = ~n11893 & ~n11894 ;
  assign n11877 = decrypt_pad & ~\u2_uk_K_r9_reg[30]/NET0131  ;
  assign n11878 = ~decrypt_pad & ~\u2_uk_K_r9_reg[7]/NET0131  ;
  assign n11879 = ~n11877 & ~n11878 ;
  assign n11880 = \u2_R9_reg[26]/NET0131  & ~n11879 ;
  assign n11881 = ~\u2_R9_reg[26]/NET0131  & n11879 ;
  assign n11882 = ~n11880 & ~n11881 ;
  assign n11896 = decrypt_pad & ~\u2_uk_K_r9_reg[38]/NET0131  ;
  assign n11897 = ~decrypt_pad & ~\u2_uk_K_r9_reg[42]/NET0131  ;
  assign n11898 = ~n11896 & ~n11897 ;
  assign n11899 = \u2_R9_reg[24]/NET0131  & ~n11898 ;
  assign n11900 = ~\u2_R9_reg[24]/NET0131  & n11898 ;
  assign n11901 = ~n11899 & ~n11900 ;
  assign n11883 = decrypt_pad & ~\u2_uk_K_r9_reg[14]/NET0131  ;
  assign n11884 = ~decrypt_pad & ~\u2_uk_K_r9_reg[22]/NET0131  ;
  assign n11885 = ~n11883 & ~n11884 ;
  assign n11886 = \u2_R9_reg[25]/NET0131  & ~n11885 ;
  assign n11887 = ~\u2_R9_reg[25]/NET0131  & n11885 ;
  assign n11888 = ~n11886 & ~n11887 ;
  assign n11907 = decrypt_pad & ~\u2_uk_K_r9_reg[42]/NET0131  ;
  assign n11908 = ~decrypt_pad & ~\u2_uk_K_r9_reg[50]/NET0131  ;
  assign n11909 = ~n11907 & ~n11908 ;
  assign n11910 = \u2_R9_reg[29]/NET0131  & ~n11909 ;
  assign n11911 = ~\u2_R9_reg[29]/NET0131  & n11909 ;
  assign n11912 = ~n11910 & ~n11911 ;
  assign n11947 = ~n11888 & n11912 ;
  assign n11948 = n11901 & n11947 ;
  assign n11949 = ~n11882 & n11948 ;
  assign n11935 = ~n11901 & n11912 ;
  assign n11950 = n11888 & n11935 ;
  assign n11951 = ~n11949 & ~n11950 ;
  assign n11952 = ~n11895 & ~n11951 ;
  assign n11889 = ~n11882 & ~n11888 ;
  assign n11953 = n11882 & n11888 ;
  assign n11954 = ~n11889 & ~n11953 ;
  assign n11902 = n11895 & n11901 ;
  assign n11932 = ~n11882 & ~n11912 ;
  assign n11955 = n11902 & ~n11932 ;
  assign n11956 = n11954 & n11955 ;
  assign n11915 = n11882 & ~n11888 ;
  assign n11936 = n11915 & n11935 ;
  assign n11918 = ~n11901 & ~n11912 ;
  assign n11946 = n11889 & n11918 ;
  assign n11957 = ~n11936 & ~n11946 ;
  assign n11958 = ~n11956 & n11957 ;
  assign n11959 = ~n11952 & n11958 ;
  assign n11960 = n11930 & ~n11959 ;
  assign n11904 = ~n11882 & ~n11901 ;
  assign n11905 = n11882 & n11901 ;
  assign n11906 = ~n11904 & ~n11905 ;
  assign n11913 = ~n11906 & n11912 ;
  assign n11916 = n11901 & ~n11912 ;
  assign n11917 = ~n11915 & n11916 ;
  assign n11919 = n11915 & n11918 ;
  assign n11920 = ~n11917 & ~n11919 ;
  assign n11921 = ~n11913 & n11920 ;
  assign n11922 = ~n11895 & ~n11921 ;
  assign n11903 = n11889 & n11902 ;
  assign n11914 = n11888 & n11913 ;
  assign n11923 = ~n11903 & ~n11914 ;
  assign n11924 = ~n11922 & n11923 ;
  assign n11931 = ~n11924 & ~n11930 ;
  assign n11937 = n11888 & n11918 ;
  assign n11938 = n11882 & n11937 ;
  assign n11939 = ~n11936 & ~n11938 ;
  assign n11940 = ~n11888 & ~n11912 ;
  assign n11941 = n11901 & n11940 ;
  assign n11942 = n11939 & ~n11941 ;
  assign n11943 = n11895 & ~n11942 ;
  assign n11933 = ~n11888 & n11895 ;
  assign n11934 = n11932 & n11933 ;
  assign n11944 = n11888 & ~n11895 ;
  assign n11945 = ~n11906 & n11944 ;
  assign n11961 = ~n11934 & ~n11945 ;
  assign n11962 = ~n11943 & n11961 ;
  assign n11963 = ~n11931 & n11962 ;
  assign n11964 = ~n11960 & n11963 ;
  assign n11965 = ~\u2_L9_reg[22]/NET0131  & ~n11964 ;
  assign n11966 = \u2_L9_reg[22]/NET0131  & n11964 ;
  assign n11967 = ~n11965 & ~n11966 ;
  assign n11968 = decrypt_pad & ~\u2_uk_K_r9_reg[41]/NET0131  ;
  assign n11969 = ~decrypt_pad & ~\u2_uk_K_r9_reg[47]/NET0131  ;
  assign n11970 = ~n11968 & ~n11969 ;
  assign n11971 = \u2_R9_reg[3]/NET0131  & ~n11970 ;
  assign n11972 = ~\u2_R9_reg[3]/NET0131  & n11970 ;
  assign n11973 = ~n11971 & ~n11972 ;
  assign n12012 = decrypt_pad & ~\u2_uk_K_r9_reg[19]/NET0131  ;
  assign n12013 = ~decrypt_pad & ~\u2_uk_K_r9_reg[25]/NET0131  ;
  assign n12014 = ~n12012 & ~n12013 ;
  assign n12015 = \u2_R9_reg[4]/NET0131  & ~n12014 ;
  assign n12016 = ~\u2_R9_reg[4]/NET0131  & n12014 ;
  assign n12017 = ~n12015 & ~n12016 ;
  assign n11987 = decrypt_pad & ~\u2_uk_K_r9_reg[32]/NET0131  ;
  assign n11988 = ~decrypt_pad & ~\u2_uk_K_r9_reg[13]/NET0131  ;
  assign n11989 = ~n11987 & ~n11988 ;
  assign n11990 = \u2_R9_reg[2]/NET0131  & ~n11989 ;
  assign n11991 = ~\u2_R9_reg[2]/NET0131  & n11989 ;
  assign n11992 = ~n11990 & ~n11991 ;
  assign n11981 = decrypt_pad & ~\u2_uk_K_r9_reg[47]/NET0131  ;
  assign n11982 = ~decrypt_pad & ~\u2_uk_K_r9_reg[53]/NET0131  ;
  assign n11983 = ~n11981 & ~n11982 ;
  assign n11984 = \u2_R9_reg[5]/NET0131  & ~n11983 ;
  assign n11985 = ~\u2_R9_reg[5]/NET0131  & n11983 ;
  assign n11986 = ~n11984 & ~n11985 ;
  assign n11974 = decrypt_pad & ~\u2_uk_K_r9_reg[17]/NET0131  ;
  assign n11975 = ~decrypt_pad & ~\u2_uk_K_r9_reg[55]/NET0131  ;
  assign n11976 = ~n11974 & ~n11975 ;
  assign n11977 = \u2_R9_reg[1]/NET0131  & ~n11976 ;
  assign n11978 = ~\u2_R9_reg[1]/NET0131  & n11976 ;
  assign n11979 = ~n11977 & ~n11978 ;
  assign n11996 = decrypt_pad & ~\u2_uk_K_r9_reg[53]/NET0131  ;
  assign n11997 = ~decrypt_pad & ~\u2_uk_K_r9_reg[34]/NET0131  ;
  assign n11998 = ~n11996 & ~n11997 ;
  assign n11999 = \u2_R9_reg[32]/NET0131  & ~n11998 ;
  assign n12000 = ~\u2_R9_reg[32]/NET0131  & n11998 ;
  assign n12001 = ~n11999 & ~n12000 ;
  assign n12043 = ~n11979 & n12001 ;
  assign n12044 = ~n11986 & n12043 ;
  assign n12045 = n11992 & n12044 ;
  assign n12007 = ~n11979 & n11986 ;
  assign n12024 = ~n11992 & ~n12001 ;
  assign n12046 = ~n12007 & n12024 ;
  assign n12047 = ~n12045 & ~n12046 ;
  assign n12048 = ~n12017 & ~n12047 ;
  assign n12022 = n11986 & ~n12001 ;
  assign n12049 = ~n11979 & n12022 ;
  assign n12050 = n11992 & n12049 ;
  assign n12028 = n11979 & n11992 ;
  assign n12041 = n11986 & n12028 ;
  assign n12042 = n12001 & n12041 ;
  assign n11993 = ~n11986 & ~n11992 ;
  assign n12051 = n11979 & n11993 ;
  assign n12052 = ~n12042 & ~n12051 ;
  assign n12053 = ~n12050 & n12052 ;
  assign n12054 = ~n12048 & n12053 ;
  assign n12055 = ~n11973 & ~n12054 ;
  assign n12008 = ~n11986 & ~n12001 ;
  assign n12009 = n11992 & n12008 ;
  assign n12010 = ~n12007 & ~n12009 ;
  assign n12011 = n11973 & ~n12010 ;
  assign n11980 = ~n11973 & n11979 ;
  assign n11994 = ~n11979 & n11993 ;
  assign n11995 = ~n11980 & ~n11994 ;
  assign n12002 = ~n11995 & n12001 ;
  assign n12003 = n11973 & ~n11992 ;
  assign n12004 = n11979 & ~n12003 ;
  assign n12005 = ~n11993 & ~n12001 ;
  assign n12006 = ~n12004 & n12005 ;
  assign n12018 = ~n12006 & n12017 ;
  assign n12019 = ~n12002 & n12018 ;
  assign n12020 = ~n12011 & n12019 ;
  assign n12029 = ~n11986 & n12028 ;
  assign n12030 = n12001 & n12029 ;
  assign n12031 = n11986 & n12001 ;
  assign n12032 = ~n11992 & n12031 ;
  assign n12033 = ~n12030 & ~n12032 ;
  assign n12034 = n11973 & ~n12033 ;
  assign n12021 = n11973 & n11992 ;
  assign n12023 = n12021 & n12022 ;
  assign n12025 = ~n11986 & n12024 ;
  assign n12026 = ~n12023 & ~n12025 ;
  assign n12027 = n11979 & ~n12026 ;
  assign n12035 = ~n11992 & n12001 ;
  assign n12036 = n12007 & n12035 ;
  assign n12037 = ~n12017 & ~n12036 ;
  assign n12038 = ~n12027 & n12037 ;
  assign n12039 = ~n12034 & n12038 ;
  assign n12040 = ~n12020 & ~n12039 ;
  assign n12056 = n12003 & n12043 ;
  assign n12057 = ~n11979 & n12008 ;
  assign n12058 = n12021 & n12057 ;
  assign n12059 = ~n12056 & ~n12058 ;
  assign n12060 = ~n12040 & n12059 ;
  assign n12061 = ~n12055 & n12060 ;
  assign n12062 = ~\u2_L9_reg[31]/NET0131  & ~n12061 ;
  assign n12063 = \u2_L9_reg[31]/NET0131  & n12061 ;
  assign n12064 = ~n12062 & ~n12063 ;
  assign n12116 = decrypt_pad & ~\u2_uk_K_r9_reg[43]/NET0131  ;
  assign n12117 = ~decrypt_pad & ~\u2_uk_K_r9_reg[51]/NET0131  ;
  assign n12118 = ~n12116 & ~n12117 ;
  assign n12119 = \u2_R9_reg[24]/NET0131  & ~n12118 ;
  assign n12120 = ~\u2_R9_reg[24]/NET0131  & n12118 ;
  assign n12121 = ~n12119 & ~n12120 ;
  assign n12071 = decrypt_pad & ~\u2_uk_K_r9_reg[22]/NET0131  ;
  assign n12072 = ~decrypt_pad & ~\u2_uk_K_r9_reg[30]/NET0131  ;
  assign n12073 = ~n12071 & ~n12072 ;
  assign n12074 = \u2_R9_reg[20]/NET0131  & ~n12073 ;
  assign n12075 = ~\u2_R9_reg[20]/NET0131  & n12073 ;
  assign n12076 = ~n12074 & ~n12075 ;
  assign n12084 = decrypt_pad & ~\u2_uk_K_r9_reg[28]/NET0131  ;
  assign n12085 = ~decrypt_pad & ~\u2_uk_K_r9_reg[36]/NET0131  ;
  assign n12086 = ~n12084 & ~n12085 ;
  assign n12087 = \u2_R9_reg[22]/NET0131  & ~n12086 ;
  assign n12088 = ~\u2_R9_reg[22]/NET0131  & n12086 ;
  assign n12089 = ~n12087 & ~n12088 ;
  assign n12090 = decrypt_pad & ~\u2_uk_K_r9_reg[37]/NET0131  ;
  assign n12091 = ~decrypt_pad & ~\u2_uk_K_r9_reg[14]/NET0131  ;
  assign n12092 = ~n12090 & ~n12091 ;
  assign n12093 = \u2_R9_reg[21]/NET0131  & ~n12092 ;
  assign n12094 = ~\u2_R9_reg[21]/NET0131  & n12092 ;
  assign n12095 = ~n12093 & ~n12094 ;
  assign n12125 = ~n12089 & n12095 ;
  assign n12141 = n12076 & n12125 ;
  assign n12065 = decrypt_pad & ~\u2_uk_K_r9_reg[45]/NET0131  ;
  assign n12066 = ~decrypt_pad & ~\u2_uk_K_r9_reg[49]/NET0131  ;
  assign n12067 = ~n12065 & ~n12066 ;
  assign n12068 = \u2_R9_reg[23]/NET0131  & ~n12067 ;
  assign n12069 = ~\u2_R9_reg[23]/NET0131  & n12067 ;
  assign n12070 = ~n12068 & ~n12069 ;
  assign n12098 = ~n12076 & n12095 ;
  assign n12099 = n12089 & n12098 ;
  assign n12142 = ~n12070 & ~n12099 ;
  assign n12143 = ~n12141 & n12142 ;
  assign n12077 = decrypt_pad & ~\u2_uk_K_r9_reg[7]/NET0131  ;
  assign n12078 = ~decrypt_pad & ~\u2_uk_K_r9_reg[15]/NET0131  ;
  assign n12079 = ~n12077 & ~n12078 ;
  assign n12080 = \u2_R9_reg[25]/NET0131  & ~n12079 ;
  assign n12081 = ~\u2_R9_reg[25]/NET0131  & n12079 ;
  assign n12082 = ~n12080 & ~n12081 ;
  assign n12133 = n12082 & ~n12095 ;
  assign n12134 = ~n12076 & n12133 ;
  assign n12135 = n12070 & ~n12134 ;
  assign n12144 = n12089 & ~n12095 ;
  assign n12145 = n12076 & n12144 ;
  assign n12146 = ~n12076 & ~n12089 ;
  assign n12147 = ~n12145 & ~n12146 ;
  assign n12148 = n12135 & n12147 ;
  assign n12149 = ~n12143 & ~n12148 ;
  assign n12100 = n12076 & n12082 ;
  assign n12111 = ~n12095 & n12100 ;
  assign n12138 = n12089 & n12111 ;
  assign n12083 = n12076 & ~n12082 ;
  assign n12105 = ~n12070 & ~n12089 ;
  assign n12139 = ~n12105 & ~n12125 ;
  assign n12140 = n12083 & ~n12139 ;
  assign n12150 = ~n12138 & ~n12140 ;
  assign n12151 = ~n12149 & n12150 ;
  assign n12152 = ~n12121 & ~n12151 ;
  assign n12101 = n12095 & n12100 ;
  assign n12096 = ~n12089 & ~n12095 ;
  assign n12097 = n12083 & n12096 ;
  assign n12102 = ~n12097 & ~n12099 ;
  assign n12103 = ~n12101 & n12102 ;
  assign n12104 = n12070 & ~n12103 ;
  assign n12106 = ~n12098 & ~n12100 ;
  assign n12107 = ~n12070 & n12106 ;
  assign n12108 = ~n12105 & ~n12107 ;
  assign n12109 = n12082 & n12095 ;
  assign n12110 = ~n12076 & n12109 ;
  assign n12112 = ~n12089 & ~n12110 ;
  assign n12113 = ~n12111 & n12112 ;
  assign n12114 = ~n12108 & ~n12113 ;
  assign n12115 = ~n12104 & ~n12114 ;
  assign n12122 = ~n12115 & n12121 ;
  assign n12131 = n12083 & n12095 ;
  assign n12132 = ~n12070 & ~n12131 ;
  assign n12136 = ~n12089 & ~n12132 ;
  assign n12137 = ~n12135 & n12136 ;
  assign n12126 = ~n12100 & ~n12125 ;
  assign n12123 = ~n12076 & ~n12082 ;
  assign n12124 = ~n12089 & ~n12123 ;
  assign n12127 = n12070 & ~n12124 ;
  assign n12128 = ~n12126 & n12127 ;
  assign n12129 = ~n12095 & n12123 ;
  assign n12130 = n12105 & n12129 ;
  assign n12153 = ~n12128 & ~n12130 ;
  assign n12154 = ~n12137 & n12153 ;
  assign n12155 = ~n12122 & n12154 ;
  assign n12156 = ~n12152 & n12155 ;
  assign n12157 = \u2_L9_reg[11]/NET0131  & ~n12156 ;
  assign n12158 = ~\u2_L9_reg[11]/NET0131  & n12156 ;
  assign n12159 = ~n12157 & ~n12158 ;
  assign n12160 = decrypt_pad & ~\u2_uk_K_r9_reg[4]/NET0131  ;
  assign n12161 = ~decrypt_pad & ~\u2_uk_K_r9_reg[10]/NET0131  ;
  assign n12162 = ~n12160 & ~n12161 ;
  assign n12163 = \u2_R9_reg[13]/NET0131  & ~n12162 ;
  assign n12164 = ~\u2_R9_reg[13]/NET0131  & n12162 ;
  assign n12165 = ~n12163 & ~n12164 ;
  assign n12178 = decrypt_pad & ~\u2_uk_K_r9_reg[10]/NET0131  ;
  assign n12179 = ~decrypt_pad & ~\u2_uk_K_r9_reg[48]/NET0131  ;
  assign n12180 = ~n12178 & ~n12179 ;
  assign n12181 = \u2_R9_reg[12]/NET0131  & ~n12180 ;
  assign n12182 = ~\u2_R9_reg[12]/NET0131  & n12180 ;
  assign n12183 = ~n12181 & ~n12182 ;
  assign n12187 = n12165 & ~n12183 ;
  assign n12191 = ~n12165 & n12183 ;
  assign n12192 = ~n12187 & ~n12191 ;
  assign n12172 = decrypt_pad & ~\u2_uk_K_r9_reg[5]/NET0131  ;
  assign n12173 = ~decrypt_pad & ~\u2_uk_K_r9_reg[11]/NET0131  ;
  assign n12174 = ~n12172 & ~n12173 ;
  assign n12175 = \u2_R9_reg[14]/NET0131  & ~n12174 ;
  assign n12176 = ~\u2_R9_reg[14]/NET0131  & n12174 ;
  assign n12177 = ~n12175 & ~n12176 ;
  assign n12193 = decrypt_pad & ~\u2_uk_K_r9_reg[13]/NET0131  ;
  assign n12194 = ~decrypt_pad & ~\u2_uk_K_r9_reg[19]/NET0131  ;
  assign n12195 = ~n12193 & ~n12194 ;
  assign n12196 = \u2_R9_reg[15]/NET0131  & ~n12195 ;
  assign n12197 = ~\u2_R9_reg[15]/NET0131  & n12195 ;
  assign n12198 = ~n12196 & ~n12197 ;
  assign n12199 = ~n12177 & ~n12198 ;
  assign n12200 = ~n12192 & n12199 ;
  assign n12166 = decrypt_pad & ~\u2_uk_K_r9_reg[26]/NET0131  ;
  assign n12167 = ~decrypt_pad & ~\u2_uk_K_r9_reg[32]/NET0131  ;
  assign n12168 = ~n12166 & ~n12167 ;
  assign n12169 = \u2_R9_reg[17]/NET0131  & ~n12168 ;
  assign n12170 = ~\u2_R9_reg[17]/NET0131  & n12168 ;
  assign n12171 = ~n12169 & ~n12170 ;
  assign n12208 = ~n12171 & n12183 ;
  assign n12209 = n12165 & n12198 ;
  assign n12210 = n12208 & n12209 ;
  assign n12205 = ~n12165 & n12198 ;
  assign n12206 = n12171 & ~n12183 ;
  assign n12207 = n12205 & n12206 ;
  assign n12211 = decrypt_pad & ~\u2_uk_K_r9_reg[46]/NET0131  ;
  assign n12212 = ~decrypt_pad & ~\u2_uk_K_r9_reg[27]/NET0131  ;
  assign n12213 = ~n12211 & ~n12212 ;
  assign n12214 = \u2_R9_reg[16]/NET0131  & ~n12213 ;
  assign n12215 = ~\u2_R9_reg[16]/NET0131  & n12213 ;
  assign n12216 = ~n12214 & ~n12215 ;
  assign n12217 = ~n12207 & n12216 ;
  assign n12218 = ~n12210 & n12217 ;
  assign n12219 = ~n12200 & n12218 ;
  assign n12184 = n12177 & n12183 ;
  assign n12185 = n12171 & n12184 ;
  assign n12186 = n12165 & n12185 ;
  assign n12188 = n12171 & ~n12177 ;
  assign n12189 = n12187 & n12188 ;
  assign n12190 = ~n12186 & ~n12189 ;
  assign n12201 = ~n12165 & ~n12171 ;
  assign n12202 = ~n12183 & n12201 ;
  assign n12203 = ~n12198 & n12202 ;
  assign n12204 = n12177 & n12203 ;
  assign n12220 = n12190 & ~n12204 ;
  assign n12221 = n12219 & n12220 ;
  assign n12223 = ~n12177 & ~n12183 ;
  assign n12224 = ~n12208 & n12209 ;
  assign n12225 = ~n12223 & n12224 ;
  assign n12222 = n12198 & n12202 ;
  assign n12234 = n12188 & n12191 ;
  assign n12235 = ~n12216 & ~n12234 ;
  assign n12236 = ~n12222 & n12235 ;
  assign n12237 = ~n12225 & n12236 ;
  assign n12226 = ~n12171 & n12187 ;
  assign n12227 = n12177 & n12226 ;
  assign n12228 = n12201 & n12223 ;
  assign n12229 = ~n12227 & ~n12228 ;
  assign n12230 = n12177 & n12208 ;
  assign n12231 = ~n12165 & n12171 ;
  assign n12232 = ~n12230 & ~n12231 ;
  assign n12233 = ~n12198 & ~n12232 ;
  assign n12238 = n12229 & ~n12233 ;
  assign n12239 = n12237 & n12238 ;
  assign n12240 = ~n12221 & ~n12239 ;
  assign n12242 = ~n12171 & n12223 ;
  assign n12243 = ~n12230 & ~n12242 ;
  assign n12244 = n12205 & ~n12243 ;
  assign n12241 = ~n12177 & n12210 ;
  assign n12245 = n12188 & ~n12198 ;
  assign n12246 = n12187 & n12245 ;
  assign n12247 = ~n12241 & ~n12246 ;
  assign n12248 = ~n12244 & n12247 ;
  assign n12249 = ~n12240 & n12248 ;
  assign n12250 = ~\u2_L9_reg[20]/NET0131  & ~n12249 ;
  assign n12251 = \u2_L9_reg[20]/NET0131  & n12249 ;
  assign n12252 = ~n12250 & ~n12251 ;
  assign n12281 = decrypt_pad & ~\u2_uk_K_r9_reg[9]/NET0131  ;
  assign n12282 = ~decrypt_pad & ~\u2_uk_K_r9_reg[45]/NET0131  ;
  assign n12283 = ~n12281 & ~n12282 ;
  assign n12284 = \u2_R9_reg[31]/P0001  & ~n12283 ;
  assign n12285 = ~\u2_R9_reg[31]/P0001  & n12283 ;
  assign n12286 = ~n12284 & ~n12285 ;
  assign n12272 = decrypt_pad & ~\u2_uk_K_r9_reg[36]/NET0131  ;
  assign n12273 = ~decrypt_pad & ~\u2_uk_K_r9_reg[44]/NET0131  ;
  assign n12274 = ~n12272 & ~n12273 ;
  assign n12275 = \u2_R9_reg[1]/NET0131  & ~n12274 ;
  assign n12276 = ~\u2_R9_reg[1]/NET0131  & n12274 ;
  assign n12277 = ~n12275 & ~n12276 ;
  assign n12265 = decrypt_pad & ~\u2_uk_K_r9_reg[21]/NET0131  ;
  assign n12266 = ~decrypt_pad & ~\u2_uk_K_r9_reg[29]/NET0131  ;
  assign n12267 = ~n12265 & ~n12266 ;
  assign n12268 = \u2_R9_reg[30]/NET0131  & ~n12267 ;
  assign n12269 = ~\u2_R9_reg[30]/NET0131  & n12267 ;
  assign n12270 = ~n12268 & ~n12269 ;
  assign n12253 = decrypt_pad & ~\u2_uk_K_r9_reg[52]/NET0131  ;
  assign n12254 = ~decrypt_pad & ~\u2_uk_K_r9_reg[1]/NET0131  ;
  assign n12255 = ~n12253 & ~n12254 ;
  assign n12256 = \u2_R9_reg[28]/NET0131  & ~n12255 ;
  assign n12257 = ~\u2_R9_reg[28]/NET0131  & n12255 ;
  assign n12258 = ~n12256 & ~n12257 ;
  assign n12259 = decrypt_pad & ~\u2_uk_K_r9_reg[51]/NET0131  ;
  assign n12260 = ~decrypt_pad & ~\u2_uk_K_r9_reg[28]/NET0131  ;
  assign n12261 = ~n12259 & ~n12260 ;
  assign n12262 = \u2_R9_reg[29]/NET0131  & ~n12261 ;
  assign n12263 = ~\u2_R9_reg[29]/NET0131  & n12261 ;
  assign n12264 = ~n12262 & ~n12263 ;
  assign n12291 = n12258 & ~n12264 ;
  assign n12292 = n12270 & n12291 ;
  assign n12293 = ~n12277 & n12292 ;
  assign n12294 = ~n12258 & n12277 ;
  assign n12295 = ~n12264 & n12294 ;
  assign n12296 = ~n12293 & ~n12295 ;
  assign n12297 = n12286 & ~n12296 ;
  assign n12279 = n12264 & n12270 ;
  assign n12280 = n12277 & n12279 ;
  assign n12271 = n12264 & ~n12270 ;
  assign n12278 = n12271 & ~n12277 ;
  assign n12287 = ~n12270 & ~n12286 ;
  assign n12288 = ~n12278 & ~n12287 ;
  assign n12289 = ~n12280 & n12288 ;
  assign n12290 = n12258 & ~n12289 ;
  assign n12298 = ~n12264 & n12277 ;
  assign n12301 = ~n12286 & ~n12298 ;
  assign n12299 = ~n12270 & ~n12277 ;
  assign n12300 = n12258 & ~n12277 ;
  assign n12302 = ~n12299 & ~n12300 ;
  assign n12303 = n12301 & n12302 ;
  assign n12304 = ~n12290 & ~n12303 ;
  assign n12305 = ~n12297 & n12304 ;
  assign n12306 = decrypt_pad & ~\u2_uk_K_r9_reg[15]/NET0131  ;
  assign n12307 = ~decrypt_pad & ~\u2_uk_K_r9_reg[23]/NET0131  ;
  assign n12308 = ~n12306 & ~n12307 ;
  assign n12309 = \u2_R9_reg[32]/NET0131  & ~n12308 ;
  assign n12310 = ~\u2_R9_reg[32]/NET0131  & n12308 ;
  assign n12311 = ~n12309 & ~n12310 ;
  assign n12312 = ~n12305 & ~n12311 ;
  assign n12322 = ~n12258 & ~n12277 ;
  assign n12331 = n12270 & ~n12277 ;
  assign n12332 = ~n12322 & ~n12331 ;
  assign n12333 = n12264 & ~n12332 ;
  assign n12318 = n12258 & n12277 ;
  assign n12319 = ~n12270 & n12318 ;
  assign n12334 = ~n12270 & n12291 ;
  assign n12335 = ~n12319 & ~n12334 ;
  assign n12336 = ~n12333 & n12335 ;
  assign n12337 = n12286 & ~n12336 ;
  assign n12330 = ~n12258 & n12280 ;
  assign n12324 = ~n12264 & ~n12270 ;
  assign n12338 = ~n12258 & n12324 ;
  assign n12339 = ~n12286 & n12338 ;
  assign n12340 = ~n12330 & ~n12339 ;
  assign n12341 = ~n12337 & n12340 ;
  assign n12342 = n12311 & ~n12341 ;
  assign n12323 = n12279 & n12322 ;
  assign n12325 = n12322 & n12324 ;
  assign n12326 = ~n12323 & ~n12325 ;
  assign n12320 = ~n12264 & n12319 ;
  assign n12321 = n12270 & n12295 ;
  assign n12327 = ~n12320 & ~n12321 ;
  assign n12328 = n12326 & n12327 ;
  assign n12329 = n12286 & ~n12328 ;
  assign n12313 = n12270 & ~n12286 ;
  assign n12314 = n12291 & n12311 ;
  assign n12315 = n12313 & n12314 ;
  assign n12316 = n12264 & n12300 ;
  assign n12317 = n12287 & n12316 ;
  assign n12343 = ~n12315 & ~n12317 ;
  assign n12344 = ~n12329 & n12343 ;
  assign n12345 = ~n12342 & n12344 ;
  assign n12346 = ~n12312 & n12345 ;
  assign n12347 = \u2_L9_reg[5]/NET0131  & ~n12346 ;
  assign n12348 = ~\u2_L9_reg[5]/NET0131  & n12346 ;
  assign n12349 = ~n12347 & ~n12348 ;
  assign n12369 = ~n12188 & n12205 ;
  assign n12360 = n12165 & ~n12177 ;
  assign n12370 = ~n12245 & ~n12360 ;
  assign n12371 = ~n12369 & n12370 ;
  assign n12372 = n12183 & ~n12371 ;
  assign n12367 = n12188 & n12198 ;
  assign n12368 = ~n12183 & n12367 ;
  assign n12373 = ~n12203 & ~n12368 ;
  assign n12374 = n12229 & n12373 ;
  assign n12375 = ~n12372 & n12374 ;
  assign n12376 = ~n12216 & ~n12375 ;
  assign n12361 = n12208 & ~n12360 ;
  assign n12362 = ~n12189 & ~n12361 ;
  assign n12363 = ~n12198 & ~n12362 ;
  assign n12350 = n12177 & ~n12183 ;
  assign n12351 = n12231 & n12350 ;
  assign n12352 = ~n12186 & ~n12351 ;
  assign n12358 = ~n12226 & ~n12234 ;
  assign n12359 = n12198 & ~n12358 ;
  assign n12364 = n12352 & ~n12359 ;
  assign n12365 = ~n12363 & n12364 ;
  assign n12366 = n12216 & ~n12365 ;
  assign n12353 = ~n12228 & n12352 ;
  assign n12354 = ~n12198 & ~n12353 ;
  assign n12355 = ~n12177 & n12208 ;
  assign n12356 = ~n12350 & ~n12355 ;
  assign n12357 = n12209 & ~n12356 ;
  assign n12377 = ~n12354 & ~n12357 ;
  assign n12378 = ~n12366 & n12377 ;
  assign n12379 = ~n12376 & n12378 ;
  assign n12380 = ~\u2_L9_reg[10]/NET0131  & ~n12379 ;
  assign n12381 = \u2_L9_reg[10]/NET0131  & n12379 ;
  assign n12382 = ~n12380 & ~n12381 ;
  assign n12391 = n11930 & ~n11938 ;
  assign n12390 = ~n11895 & n11936 ;
  assign n12392 = ~n11949 & ~n12390 ;
  assign n12393 = n12391 & n12392 ;
  assign n12383 = n11888 & n11901 ;
  assign n12384 = ~n11946 & ~n12383 ;
  assign n12385 = n11895 & ~n12384 ;
  assign n12386 = n11882 & n11912 ;
  assign n12387 = ~n11932 & ~n12386 ;
  assign n12388 = ~n11906 & n11954 ;
  assign n12389 = n12387 & n12388 ;
  assign n12394 = ~n12385 & ~n12389 ;
  assign n12395 = n12393 & n12394 ;
  assign n12396 = ~n11937 & ~n11941 ;
  assign n12397 = ~n11882 & ~n12396 ;
  assign n12405 = ~n11919 & ~n11930 ;
  assign n12400 = n11905 & n11947 ;
  assign n12401 = ~n11895 & n11905 ;
  assign n12406 = ~n12400 & ~n12401 ;
  assign n12407 = n12405 & n12406 ;
  assign n12398 = ~n11933 & ~n11953 ;
  assign n12399 = n11935 & ~n12398 ;
  assign n12402 = n11888 & ~n11912 ;
  assign n12403 = ~n11895 & ~n11947 ;
  assign n12404 = ~n12402 & n12403 ;
  assign n12408 = ~n12399 & ~n12404 ;
  assign n12409 = n12407 & n12408 ;
  assign n12410 = ~n12397 & n12409 ;
  assign n12411 = ~n12395 & ~n12410 ;
  assign n12412 = \u2_L9_reg[12]/NET0131  & n12411 ;
  assign n12413 = ~\u2_L9_reg[12]/NET0131  & ~n12411 ;
  assign n12414 = ~n12412 & ~n12413 ;
  assign n12472 = decrypt_pad & ~\u2_uk_K_r9_reg[0]/P0001  ;
  assign n12473 = ~decrypt_pad & ~\u2_uk_K_r9_reg[8]/NET0131  ;
  assign n12474 = ~n12472 & ~n12473 ;
  assign n12475 = \u2_R9_reg[20]/NET0131  & ~n12474 ;
  assign n12476 = ~\u2_R9_reg[20]/NET0131  & n12474 ;
  assign n12477 = ~n12475 & ~n12476 ;
  assign n12421 = decrypt_pad & ~\u2_uk_K_r9_reg[29]/NET0131  ;
  assign n12422 = ~decrypt_pad & ~\u2_uk_K_r9_reg[37]/NET0131  ;
  assign n12423 = ~n12421 & ~n12422 ;
  assign n12424 = \u2_R9_reg[18]/NET0131  & ~n12423 ;
  assign n12425 = ~\u2_R9_reg[18]/NET0131  & n12423 ;
  assign n12426 = ~n12424 & ~n12425 ;
  assign n12415 = decrypt_pad & ~\u2_uk_K_r9_reg[35]/NET0131  ;
  assign n12416 = ~decrypt_pad & ~\u2_uk_K_r9_reg[43]/NET0131  ;
  assign n12417 = ~n12415 & ~n12416 ;
  assign n12418 = \u2_R9_reg[17]/NET0131  & ~n12417 ;
  assign n12419 = ~\u2_R9_reg[17]/NET0131  & n12417 ;
  assign n12420 = ~n12418 & ~n12419 ;
  assign n12428 = decrypt_pad & ~\u2_uk_K_r9_reg[44]/NET0131  ;
  assign n12429 = ~decrypt_pad & ~\u2_uk_K_r9_reg[21]/NET0131  ;
  assign n12430 = ~n12428 & ~n12429 ;
  assign n12431 = \u2_R9_reg[16]/NET0131  & ~n12430 ;
  assign n12432 = ~\u2_R9_reg[16]/NET0131  & n12430 ;
  assign n12433 = ~n12431 & ~n12432 ;
  assign n12436 = decrypt_pad & ~\u2_uk_K_r9_reg[1]/NET0131  ;
  assign n12437 = ~decrypt_pad & ~\u2_uk_K_r9_reg[9]/NET0131  ;
  assign n12438 = ~n12436 & ~n12437 ;
  assign n12439 = \u2_R9_reg[21]/NET0131  & ~n12438 ;
  assign n12440 = ~\u2_R9_reg[21]/NET0131  & n12438 ;
  assign n12441 = ~n12439 & ~n12440 ;
  assign n12454 = n12433 & n12441 ;
  assign n12465 = n12420 & n12454 ;
  assign n12444 = n12433 & ~n12441 ;
  assign n12467 = ~n12420 & n12444 ;
  assign n12482 = ~n12465 & ~n12467 ;
  assign n12483 = ~n12426 & ~n12482 ;
  assign n12456 = ~n12420 & ~n12433 ;
  assign n12481 = n12441 & n12456 ;
  assign n12447 = decrypt_pad & ~\u2_uk_K_r9_reg[16]/NET0131  ;
  assign n12448 = ~decrypt_pad & ~\u2_uk_K_r9_reg[52]/NET0131  ;
  assign n12449 = ~n12447 & ~n12448 ;
  assign n12450 = \u2_R9_reg[19]/NET0131  & ~n12449 ;
  assign n12451 = ~\u2_R9_reg[19]/NET0131  & n12449 ;
  assign n12452 = ~n12450 & ~n12451 ;
  assign n12479 = n12420 & ~n12441 ;
  assign n12480 = n12426 & n12479 ;
  assign n12484 = ~n12452 & ~n12480 ;
  assign n12485 = ~n12481 & n12484 ;
  assign n12486 = ~n12483 & n12485 ;
  assign n12435 = n12426 & n12433 ;
  assign n12442 = ~n12435 & n12441 ;
  assign n12487 = ~n12444 & ~n12479 ;
  assign n12488 = ~n12442 & n12487 ;
  assign n12427 = n12420 & ~n12426 ;
  assign n12434 = n12427 & ~n12433 ;
  assign n12489 = ~n12434 & n12452 ;
  assign n12490 = ~n12488 & n12489 ;
  assign n12491 = ~n12486 & ~n12490 ;
  assign n12455 = ~n12420 & n12454 ;
  assign n12492 = n12426 & n12455 ;
  assign n12493 = n12434 & ~n12441 ;
  assign n12494 = ~n12492 & ~n12493 ;
  assign n12495 = ~n12491 & n12494 ;
  assign n12496 = ~n12477 & ~n12495 ;
  assign n12443 = ~n12434 & n12442 ;
  assign n12445 = n12420 & n12444 ;
  assign n12446 = ~n12443 & ~n12445 ;
  assign n12453 = ~n12446 & n12452 ;
  assign n12457 = ~n12441 & n12456 ;
  assign n12458 = ~n12433 & n12441 ;
  assign n12459 = n12420 & n12458 ;
  assign n12460 = ~n12457 & ~n12459 ;
  assign n12461 = ~n12452 & ~n12460 ;
  assign n12462 = ~n12426 & ~n12445 ;
  assign n12463 = ~n12455 & n12462 ;
  assign n12464 = ~n12461 & n12463 ;
  assign n12466 = ~n12452 & n12465 ;
  assign n12468 = n12426 & ~n12467 ;
  assign n12469 = ~n12466 & n12468 ;
  assign n12470 = ~n12464 & ~n12469 ;
  assign n12471 = ~n12453 & ~n12470 ;
  assign n12478 = ~n12471 & n12477 ;
  assign n12497 = ~n12420 & n12426 ;
  assign n12498 = n12458 & n12497 ;
  assign n12499 = ~n12480 & ~n12498 ;
  assign n12500 = ~n12433 & ~n12499 ;
  assign n12501 = ~n12452 & n12500 ;
  assign n12502 = n12426 & n12457 ;
  assign n12503 = ~n12426 & n12445 ;
  assign n12504 = ~n12502 & ~n12503 ;
  assign n12505 = n12452 & ~n12504 ;
  assign n12506 = ~n12501 & ~n12505 ;
  assign n12507 = ~n12478 & n12506 ;
  assign n12508 = ~n12496 & n12507 ;
  assign n12509 = ~\u2_L9_reg[14]/NET0131  & ~n12508 ;
  assign n12510 = \u2_L9_reg[14]/NET0131  & n12508 ;
  assign n12511 = ~n12509 & ~n12510 ;
  assign n12513 = n12258 & n12264 ;
  assign n12514 = ~n12278 & ~n12513 ;
  assign n12515 = ~n12295 & n12514 ;
  assign n12516 = n12286 & ~n12515 ;
  assign n12512 = n12291 & n12299 ;
  assign n12517 = ~n12311 & ~n12512 ;
  assign n12518 = ~n12516 & n12517 ;
  assign n12524 = n12311 & ~n12323 ;
  assign n12522 = n12298 & n12313 ;
  assign n12523 = n12258 & n12271 ;
  assign n12525 = ~n12522 & ~n12523 ;
  assign n12526 = n12524 & n12525 ;
  assign n12519 = ~n12264 & n12322 ;
  assign n12520 = n12286 & n12519 ;
  assign n12521 = n12277 & n12292 ;
  assign n12527 = ~n12520 & ~n12521 ;
  assign n12528 = n12526 & n12527 ;
  assign n12529 = ~n12518 & ~n12528 ;
  assign n12532 = ~n12286 & ~n12292 ;
  assign n12530 = n12271 & n12294 ;
  assign n12531 = n12291 & ~n12311 ;
  assign n12533 = ~n12530 & ~n12531 ;
  assign n12534 = n12532 & n12533 ;
  assign n12535 = n12326 & n12534 ;
  assign n12536 = ~n12270 & n12295 ;
  assign n12537 = n12286 & ~n12330 ;
  assign n12538 = ~n12536 & n12537 ;
  assign n12539 = ~n12535 & ~n12538 ;
  assign n12540 = ~n12529 & ~n12539 ;
  assign n12541 = ~\u2_L9_reg[15]/NET0131  & ~n12540 ;
  assign n12542 = \u2_L9_reg[15]/NET0131  & n12540 ;
  assign n12543 = ~n12541 & ~n12542 ;
  assign n12560 = ~n11979 & ~n11992 ;
  assign n12561 = ~n12001 & ~n12560 ;
  assign n12562 = ~n12036 & ~n12561 ;
  assign n12563 = n11973 & ~n12562 ;
  assign n12564 = ~n11973 & ~n12035 ;
  assign n12565 = ~n12561 & n12564 ;
  assign n12559 = n12001 & n12051 ;
  assign n12566 = ~n12041 & ~n12559 ;
  assign n12567 = ~n12565 & n12566 ;
  assign n12568 = ~n12563 & n12567 ;
  assign n12569 = n12017 & ~n12568 ;
  assign n12544 = n11986 & n12024 ;
  assign n12545 = ~n12009 & ~n12544 ;
  assign n12546 = n11973 & n11979 ;
  assign n12547 = ~n12545 & n12546 ;
  assign n12548 = ~n12008 & ~n12031 ;
  assign n12549 = ~n11979 & ~n12548 ;
  assign n12550 = ~n12025 & ~n12549 ;
  assign n12551 = ~n11973 & ~n12550 ;
  assign n12552 = n11979 & n12031 ;
  assign n12553 = ~n12044 & ~n12552 ;
  assign n12554 = n11973 & ~n12553 ;
  assign n12555 = ~n12030 & ~n12050 ;
  assign n12556 = ~n12554 & n12555 ;
  assign n12557 = ~n12551 & n12556 ;
  assign n12558 = ~n12017 & ~n12557 ;
  assign n12570 = ~n12547 & ~n12558 ;
  assign n12571 = ~n12569 & n12570 ;
  assign n12572 = ~\u2_L9_reg[17]/NET0131  & ~n12571 ;
  assign n12573 = \u2_L9_reg[17]/NET0131  & n12571 ;
  assign n12574 = ~n12572 & ~n12573 ;
  assign n12591 = n12183 & n12231 ;
  assign n12592 = ~n12198 & ~n12355 ;
  assign n12593 = ~n12591 & n12592 ;
  assign n12594 = n12184 & n12201 ;
  assign n12595 = n12198 & ~n12242 ;
  assign n12596 = ~n12594 & n12595 ;
  assign n12597 = ~n12593 & ~n12596 ;
  assign n12598 = n12165 & n12355 ;
  assign n12599 = n12190 & ~n12598 ;
  assign n12600 = ~n12597 & n12599 ;
  assign n12601 = ~n12216 & ~n12600 ;
  assign n12585 = n12177 & ~n12206 ;
  assign n12581 = n12165 & ~n12198 ;
  assign n12586 = ~n12208 & n12581 ;
  assign n12587 = ~n12585 & n12586 ;
  assign n12583 = n12165 & n12230 ;
  assign n12584 = ~n12165 & n12350 ;
  assign n12588 = ~n12583 & ~n12584 ;
  assign n12589 = ~n12587 & n12588 ;
  assign n12590 = n12216 & ~n12589 ;
  assign n12575 = ~n12227 & n12352 ;
  assign n12576 = n12198 & ~n12575 ;
  assign n12577 = ~n12177 & n12191 ;
  assign n12578 = ~n12231 & ~n12577 ;
  assign n12579 = n12198 & n12216 ;
  assign n12580 = ~n12578 & n12579 ;
  assign n12582 = n12230 & n12581 ;
  assign n12602 = ~n12204 & ~n12582 ;
  assign n12603 = ~n12580 & n12602 ;
  assign n12604 = ~n12576 & n12603 ;
  assign n12605 = ~n12590 & n12604 ;
  assign n12606 = ~n12601 & n12605 ;
  assign n12607 = ~\u2_L9_reg[1]/NET0131  & ~n12606 ;
  assign n12608 = \u2_L9_reg[1]/NET0131  & n12606 ;
  assign n12609 = ~n12607 & ~n12608 ;
  assign n12635 = n12258 & n12299 ;
  assign n12636 = ~n12521 & ~n12635 ;
  assign n12637 = ~n12286 & ~n12636 ;
  assign n12631 = n12270 & n12513 ;
  assign n12629 = n12277 & n12324 ;
  assign n12630 = n12264 & n12294 ;
  assign n12632 = ~n12629 & ~n12630 ;
  assign n12633 = ~n12631 & n12632 ;
  assign n12634 = n12286 & ~n12633 ;
  assign n12627 = ~n12316 & ~n12519 ;
  assign n12628 = n12270 & ~n12627 ;
  assign n12638 = ~n12536 & ~n12628 ;
  assign n12639 = ~n12634 & n12638 ;
  assign n12640 = ~n12637 & n12639 ;
  assign n12641 = n12311 & ~n12640 ;
  assign n12610 = ~n12292 & ~n12316 ;
  assign n12611 = n12286 & ~n12610 ;
  assign n12612 = ~n12258 & n12279 ;
  assign n12618 = ~n12325 & ~n12612 ;
  assign n12613 = n12294 & n12313 ;
  assign n12614 = n12264 & ~n12286 ;
  assign n12615 = n12322 & n12614 ;
  assign n12619 = ~n12613 & ~n12615 ;
  assign n12620 = n12618 & n12619 ;
  assign n12616 = ~n12264 & n12286 ;
  assign n12617 = n12319 & ~n12616 ;
  assign n12621 = ~n12293 & ~n12617 ;
  assign n12622 = n12620 & n12621 ;
  assign n12623 = ~n12611 & n12622 ;
  assign n12624 = ~n12311 & ~n12623 ;
  assign n12625 = n12286 & n12338 ;
  assign n12626 = n12319 & n12614 ;
  assign n12642 = ~n12625 & ~n12626 ;
  assign n12643 = ~n12624 & n12642 ;
  assign n12644 = ~n12641 & n12643 ;
  assign n12645 = ~\u2_L9_reg[21]/NET0131  & ~n12644 ;
  assign n12646 = \u2_L9_reg[21]/NET0131  & n12644 ;
  assign n12647 = ~n12645 & ~n12646 ;
  assign n12669 = ~n12427 & ~n12441 ;
  assign n12670 = ~n12435 & n12669 ;
  assign n12671 = ~n12456 & ~n12465 ;
  assign n12672 = ~n12670 & n12671 ;
  assign n12673 = n12452 & ~n12672 ;
  assign n12674 = ~n12434 & ~n12455 ;
  assign n12675 = ~n12452 & ~n12674 ;
  assign n12648 = n12433 & n12480 ;
  assign n12666 = n12427 & n12441 ;
  assign n12676 = ~n12648 & ~n12666 ;
  assign n12677 = ~n12675 & n12676 ;
  assign n12678 = ~n12673 & n12677 ;
  assign n12679 = n12477 & ~n12678 ;
  assign n12653 = ~n12427 & ~n12433 ;
  assign n12654 = ~n12497 & n12653 ;
  assign n12655 = ~n12467 & ~n12654 ;
  assign n12656 = ~n12452 & ~n12655 ;
  assign n12659 = n12426 & ~n12458 ;
  assign n12658 = ~n12426 & n12441 ;
  assign n12657 = ~n12426 & ~n12452 ;
  assign n12660 = n12420 & ~n12657 ;
  assign n12661 = ~n12658 & n12660 ;
  assign n12662 = ~n12659 & n12661 ;
  assign n12663 = ~n12656 & ~n12662 ;
  assign n12664 = ~n12477 & ~n12663 ;
  assign n12649 = ~n12502 & ~n12648 ;
  assign n12650 = ~n12426 & n12481 ;
  assign n12651 = n12649 & ~n12650 ;
  assign n12652 = n12452 & ~n12651 ;
  assign n12665 = ~n12452 & n12497 ;
  assign n12667 = ~n12665 & ~n12666 ;
  assign n12668 = n12433 & ~n12667 ;
  assign n12680 = ~n12652 & ~n12668 ;
  assign n12681 = ~n12664 & n12680 ;
  assign n12682 = ~n12679 & n12681 ;
  assign n12683 = ~\u2_L9_reg[25]/NET0131  & ~n12682 ;
  assign n12684 = \u2_L9_reg[25]/NET0131  & n12682 ;
  assign n12685 = ~n12683 & ~n12684 ;
  assign n12692 = decrypt_pad & ~\u2_uk_K_r9_reg[12]/NET0131  ;
  assign n12693 = ~decrypt_pad & ~\u2_uk_K_r9_reg[18]/NET0131  ;
  assign n12694 = ~n12692 & ~n12693 ;
  assign n12695 = \u2_R9_reg[5]/NET0131  & ~n12694 ;
  assign n12696 = ~\u2_R9_reg[5]/NET0131  & n12694 ;
  assign n12697 = ~n12695 & ~n12696 ;
  assign n12699 = decrypt_pad & ~\u2_uk_K_r9_reg[33]/NET0131  ;
  assign n12700 = ~decrypt_pad & ~\u2_uk_K_r9_reg[39]/NET0131  ;
  assign n12701 = ~n12699 & ~n12700 ;
  assign n12702 = \u2_R9_reg[4]/NET0131  & ~n12701 ;
  assign n12703 = ~\u2_R9_reg[4]/NET0131  & n12701 ;
  assign n12704 = ~n12702 & ~n12703 ;
  assign n12706 = decrypt_pad & ~\u2_uk_K_r9_reg[25]/NET0131  ;
  assign n12707 = ~decrypt_pad & ~\u2_uk_K_r9_reg[6]/NET0131  ;
  assign n12708 = ~n12706 & ~n12707 ;
  assign n12709 = \u2_R9_reg[9]/NET0131  & ~n12708 ;
  assign n12710 = ~\u2_R9_reg[9]/NET0131  & n12708 ;
  assign n12711 = ~n12709 & ~n12710 ;
  assign n12713 = n12704 & ~n12711 ;
  assign n12714 = ~n12697 & ~n12713 ;
  assign n12715 = n12697 & n12704 ;
  assign n12716 = ~n12711 & n12715 ;
  assign n12717 = ~n12714 & ~n12716 ;
  assign n12718 = ~n12704 & n12711 ;
  assign n12686 = decrypt_pad & ~\u2_uk_K_r9_reg[3]/NET0131  ;
  assign n12687 = ~decrypt_pad & ~\u2_uk_K_r9_reg[41]/NET0131  ;
  assign n12688 = ~n12686 & ~n12687 ;
  assign n12689 = \u2_R9_reg[6]/NET0131  & ~n12688 ;
  assign n12690 = ~\u2_R9_reg[6]/NET0131  & n12688 ;
  assign n12691 = ~n12689 & ~n12690 ;
  assign n12719 = ~n12691 & ~n12704 ;
  assign n12720 = ~n12718 & ~n12719 ;
  assign n12721 = n12717 & n12720 ;
  assign n12722 = decrypt_pad & ~\u2_uk_K_r9_reg[54]/NET0131  ;
  assign n12723 = ~decrypt_pad & ~\u2_uk_K_r9_reg[3]/NET0131  ;
  assign n12724 = ~n12722 & ~n12723 ;
  assign n12725 = \u2_R9_reg[7]/NET0131  & ~n12724 ;
  assign n12726 = ~\u2_R9_reg[7]/NET0131  & n12724 ;
  assign n12727 = ~n12725 & ~n12726 ;
  assign n12728 = ~n12721 & n12727 ;
  assign n12729 = ~n12697 & n12711 ;
  assign n12730 = ~n12720 & ~n12729 ;
  assign n12731 = n12691 & n12716 ;
  assign n12698 = n12691 & ~n12697 ;
  assign n12705 = n12698 & ~n12704 ;
  assign n12732 = ~n12705 & ~n12727 ;
  assign n12733 = ~n12731 & n12732 ;
  assign n12734 = ~n12730 & n12733 ;
  assign n12735 = ~n12728 & ~n12734 ;
  assign n12736 = n12704 & n12729 ;
  assign n12737 = ~n12727 & ~n12736 ;
  assign n12738 = ~n12691 & n12704 ;
  assign n12739 = ~n12737 & n12738 ;
  assign n12712 = n12705 & n12711 ;
  assign n12740 = decrypt_pad & ~\u2_uk_K_r9_reg[20]/NET0131  ;
  assign n12741 = ~decrypt_pad & ~\u2_uk_K_r9_reg[26]/NET0131  ;
  assign n12742 = ~n12740 & ~n12741 ;
  assign n12743 = \u2_R9_reg[8]/NET0131  & ~n12742 ;
  assign n12744 = ~\u2_R9_reg[8]/NET0131  & n12742 ;
  assign n12745 = ~n12743 & ~n12744 ;
  assign n12746 = ~n12712 & n12745 ;
  assign n12747 = ~n12739 & n12746 ;
  assign n12748 = ~n12735 & n12747 ;
  assign n12752 = n12727 & ~n12730 ;
  assign n12753 = n12704 & ~n12729 ;
  assign n12754 = ~n12698 & n12753 ;
  assign n12755 = ~n12704 & n12729 ;
  assign n12756 = ~n12754 & ~n12755 ;
  assign n12757 = n12733 & n12756 ;
  assign n12758 = ~n12752 & ~n12757 ;
  assign n12749 = n12691 & ~n12718 ;
  assign n12750 = n12714 & n12749 ;
  assign n12751 = ~n12731 & ~n12745 ;
  assign n12759 = ~n12750 & n12751 ;
  assign n12760 = ~n12758 & n12759 ;
  assign n12761 = ~n12748 & ~n12760 ;
  assign n12762 = ~\u2_L9_reg[28]/NET0131  & n12761 ;
  assign n12763 = \u2_L9_reg[28]/NET0131  & ~n12761 ;
  assign n12764 = ~n12762 & ~n12763 ;
  assign n12781 = n12083 & ~n12095 ;
  assign n12782 = ~n12101 & ~n12781 ;
  assign n12783 = ~n12096 & ~n12099 ;
  assign n12784 = ~n12082 & ~n12783 ;
  assign n12785 = n12782 & ~n12784 ;
  assign n12786 = n12070 & ~n12785 ;
  assign n12765 = n12089 & n12131 ;
  assign n12772 = ~n12089 & ~n12106 ;
  assign n12787 = ~n12765 & ~n12772 ;
  assign n12788 = ~n12070 & ~n12787 ;
  assign n12789 = n12089 & n12134 ;
  assign n12790 = ~n12788 & ~n12789 ;
  assign n12791 = ~n12786 & n12790 ;
  assign n12792 = ~n12121 & ~n12791 ;
  assign n12766 = n12095 & n12146 ;
  assign n12767 = ~n12110 & ~n12766 ;
  assign n12768 = ~n12765 & n12767 ;
  assign n12769 = n12070 & ~n12768 ;
  assign n12773 = n12070 & ~n12133 ;
  assign n12774 = ~n12144 & n12773 ;
  assign n12770 = n12089 & ~n12100 ;
  assign n12771 = ~n12123 & n12770 ;
  assign n12775 = ~n12771 & ~n12772 ;
  assign n12776 = ~n12774 & n12775 ;
  assign n12777 = ~n12769 & ~n12776 ;
  assign n12778 = n12121 & ~n12777 ;
  assign n12779 = n12070 & n12082 ;
  assign n12780 = n12125 & n12779 ;
  assign n12793 = ~n12097 & ~n12780 ;
  assign n12794 = ~n12778 & n12793 ;
  assign n12795 = ~n12792 & n12794 ;
  assign n12796 = \u2_L9_reg[29]/NET0131  & ~n12795 ;
  assign n12797 = ~\u2_L9_reg[29]/NET0131  & n12795 ;
  assign n12798 = ~n12796 & ~n12797 ;
  assign n12804 = n12165 & n12208 ;
  assign n12805 = ~n12165 & ~n12198 ;
  assign n12806 = n12206 & ~n12805 ;
  assign n12807 = ~n12804 & ~n12806 ;
  assign n12808 = n12177 & ~n12807 ;
  assign n12801 = n12223 & n12231 ;
  assign n12802 = ~n12185 & ~n12801 ;
  assign n12803 = ~n12198 & ~n12802 ;
  assign n12800 = ~n12177 & n12226 ;
  assign n12809 = ~n12222 & ~n12800 ;
  assign n12810 = ~n12803 & n12809 ;
  assign n12811 = ~n12808 & n12810 ;
  assign n12812 = n12216 & ~n12811 ;
  assign n12821 = n12209 & n12585 ;
  assign n12822 = ~n12189 & ~n12210 ;
  assign n12823 = ~n12577 & n12822 ;
  assign n12824 = ~n12821 & n12823 ;
  assign n12825 = ~n12216 & ~n12824 ;
  assign n12799 = ~n12192 & n12367 ;
  assign n12813 = ~n12201 & ~n12584 ;
  assign n12814 = ~n12216 & ~n12813 ;
  assign n12815 = ~n12165 & ~n12208 ;
  assign n12816 = ~n12177 & ~n12206 ;
  assign n12817 = ~n12804 & n12816 ;
  assign n12818 = ~n12815 & n12817 ;
  assign n12819 = ~n12814 & ~n12818 ;
  assign n12820 = ~n12198 & ~n12819 ;
  assign n12826 = ~n12799 & ~n12820 ;
  assign n12827 = ~n12825 & n12826 ;
  assign n12828 = ~n12812 & n12827 ;
  assign n12829 = ~\u2_L9_reg[26]/NET0131  & ~n12828 ;
  assign n12830 = \u2_L9_reg[26]/NET0131  & n12828 ;
  assign n12831 = ~n12829 & ~n12830 ;
  assign n12832 = n12691 & n12727 ;
  assign n12833 = n12736 & n12832 ;
  assign n12834 = n12691 & n12704 ;
  assign n12835 = ~n12729 & ~n12834 ;
  assign n12836 = n12737 & ~n12835 ;
  assign n12846 = ~n12833 & ~n12836 ;
  assign n12837 = n12697 & ~n12711 ;
  assign n12838 = ~n12755 & ~n12837 ;
  assign n12839 = ~n12691 & ~n12838 ;
  assign n12840 = n12691 & n12718 ;
  assign n12841 = n12697 & n12840 ;
  assign n12842 = ~n12691 & ~n12697 ;
  assign n12843 = n12711 & ~n12727 ;
  assign n12844 = n12842 & n12843 ;
  assign n12845 = ~n12841 & ~n12844 ;
  assign n12847 = ~n12839 & n12845 ;
  assign n12848 = n12846 & n12847 ;
  assign n12849 = ~n12745 & ~n12848 ;
  assign n12855 = ~n12697 & ~n12711 ;
  assign n12856 = ~n12749 & ~n12855 ;
  assign n12857 = ~n12753 & ~n12856 ;
  assign n12850 = ~n12691 & n12697 ;
  assign n12853 = n12704 & n12850 ;
  assign n12854 = n12711 & n12853 ;
  assign n12858 = ~n12711 & n12842 ;
  assign n12859 = n12704 & n12858 ;
  assign n12860 = ~n12854 & ~n12859 ;
  assign n12861 = ~n12857 & n12860 ;
  assign n12862 = n12745 & ~n12861 ;
  assign n12851 = ~n12698 & ~n12850 ;
  assign n12852 = n12718 & n12851 ;
  assign n12863 = ~n12727 & ~n12852 ;
  assign n12864 = ~n12862 & n12863 ;
  assign n12866 = n12691 & ~n12715 ;
  assign n12867 = ~n12714 & n12745 ;
  assign n12868 = ~n12866 & n12867 ;
  assign n12865 = n12705 & ~n12711 ;
  assign n12869 = n12727 & ~n12853 ;
  assign n12870 = ~n12865 & n12869 ;
  assign n12871 = ~n12868 & n12870 ;
  assign n12872 = ~n12864 & ~n12871 ;
  assign n12873 = ~n12849 & ~n12872 ;
  assign n12874 = \u2_L9_reg[2]/NET0131  & n12873 ;
  assign n12875 = ~\u2_L9_reg[2]/NET0131  & ~n12873 ;
  assign n12876 = ~n12874 & ~n12875 ;
  assign n12880 = n12082 & n12146 ;
  assign n12881 = ~n12131 & ~n12880 ;
  assign n12882 = ~n12138 & n12881 ;
  assign n12883 = n12070 & ~n12882 ;
  assign n12877 = n12095 & n12123 ;
  assign n12878 = ~n12789 & ~n12877 ;
  assign n12879 = ~n12070 & ~n12878 ;
  assign n12884 = n12100 & n12105 ;
  assign n12885 = ~n12097 & ~n12884 ;
  assign n12886 = ~n12879 & n12885 ;
  assign n12887 = ~n12883 & n12886 ;
  assign n12888 = ~n12121 & ~n12887 ;
  assign n12892 = n12070 & n12100 ;
  assign n12893 = ~n12877 & ~n12892 ;
  assign n12894 = ~n12089 & ~n12893 ;
  assign n12889 = ~n12082 & n12125 ;
  assign n12890 = ~n12146 & ~n12889 ;
  assign n12891 = ~n12070 & ~n12890 ;
  assign n12895 = n12089 & n12109 ;
  assign n12896 = ~n12891 & ~n12895 ;
  assign n12897 = ~n12894 & n12896 ;
  assign n12898 = n12121 & ~n12897 ;
  assign n12899 = n12089 & n12782 ;
  assign n12900 = ~n12070 & ~n12124 ;
  assign n12901 = ~n12899 & n12900 ;
  assign n12902 = ~n12110 & ~n12129 ;
  assign n12903 = ~n12131 & n12902 ;
  assign n12904 = n12070 & n12089 ;
  assign n12905 = ~n12903 & n12904 ;
  assign n12906 = ~n12901 & ~n12905 ;
  assign n12907 = ~n12898 & n12906 ;
  assign n12908 = ~n12888 & n12907 ;
  assign n12909 = ~\u2_L9_reg[4]/NET0131  & ~n12908 ;
  assign n12910 = \u2_L9_reg[4]/NET0131  & n12908 ;
  assign n12911 = ~n12909 & ~n12910 ;
  assign n12913 = n12698 & ~n12711 ;
  assign n12914 = n12737 & ~n12913 ;
  assign n12915 = n12727 & ~n12840 ;
  assign n12916 = ~n12858 & n12915 ;
  assign n12917 = ~n12914 & ~n12916 ;
  assign n12912 = n12719 & n12837 ;
  assign n12918 = n12745 & ~n12912 ;
  assign n12919 = n12845 & n12918 ;
  assign n12920 = ~n12917 & n12919 ;
  assign n12922 = n12718 & ~n12851 ;
  assign n12921 = ~n12704 & n12837 ;
  assign n12923 = ~n12727 & ~n12745 ;
  assign n12924 = ~n12921 & n12923 ;
  assign n12925 = ~n12859 & n12924 ;
  assign n12926 = ~n12922 & n12925 ;
  assign n12927 = ~n12920 & ~n12926 ;
  assign n12928 = ~n12731 & ~n12854 ;
  assign n12929 = ~n12927 & n12928 ;
  assign n12932 = ~n12691 & ~n12717 ;
  assign n12930 = n12749 & ~n12837 ;
  assign n12931 = n12718 & n12850 ;
  assign n12933 = n12727 & ~n12745 ;
  assign n12934 = ~n12931 & n12933 ;
  assign n12935 = ~n12930 & n12934 ;
  assign n12936 = ~n12932 & n12935 ;
  assign n12937 = ~n12929 & ~n12936 ;
  assign n12938 = ~\u2_L9_reg[13]/NET0131  & ~n12937 ;
  assign n12939 = \u2_L9_reg[13]/NET0131  & n12937 ;
  assign n12940 = ~n12938 & ~n12939 ;
  assign n12941 = ~n12070 & n12076 ;
  assign n12942 = ~n12880 & ~n12941 ;
  assign n12943 = ~n12095 & ~n12942 ;
  assign n12947 = n12121 & ~n12889 ;
  assign n12948 = ~n12943 & n12947 ;
  assign n12944 = n12089 & ~n12902 ;
  assign n12945 = ~n12134 & ~n12141 ;
  assign n12946 = n12070 & ~n12945 ;
  assign n12949 = ~n12944 & ~n12946 ;
  assign n12950 = n12948 & n12949 ;
  assign n12953 = n12076 & ~n12125 ;
  assign n12954 = ~n12877 & ~n12953 ;
  assign n12955 = n12070 & ~n12954 ;
  assign n12952 = ~n12070 & ~n12902 ;
  assign n12951 = n12089 & n12101 ;
  assign n12956 = ~n12121 & ~n12951 ;
  assign n12957 = ~n12952 & n12956 ;
  assign n12958 = ~n12955 & n12957 ;
  assign n12959 = ~n12950 & ~n12958 ;
  assign n12960 = ~n12095 & n12884 ;
  assign n12961 = ~n12137 & ~n12960 ;
  assign n12962 = ~n12959 & n12961 ;
  assign n12963 = ~\u2_L9_reg[19]/NET0131  & ~n12962 ;
  assign n12964 = \u2_L9_reg[19]/NET0131  & n12962 ;
  assign n12965 = ~n12963 & ~n12964 ;
  assign n12974 = ~n12035 & n12546 ;
  assign n12975 = n12548 & n12974 ;
  assign n12976 = n12017 & ~n12036 ;
  assign n12977 = ~n12058 & n12976 ;
  assign n12978 = ~n12975 & n12977 ;
  assign n12980 = ~n11973 & n11992 ;
  assign n12981 = n11986 & n12980 ;
  assign n12982 = ~n11980 & ~n12981 ;
  assign n12983 = n12001 & ~n12982 ;
  assign n12984 = ~n11994 & ~n12017 ;
  assign n12979 = n12008 & n12546 ;
  assign n12985 = ~n12023 & ~n12041 ;
  assign n12986 = ~n12979 & n12985 ;
  assign n12987 = n12984 & n12986 ;
  assign n12988 = ~n12983 & n12987 ;
  assign n12989 = ~n12978 & ~n12988 ;
  assign n12966 = n11979 & n12008 ;
  assign n12967 = ~n12049 & ~n12966 ;
  assign n12968 = ~n12045 & n12967 ;
  assign n12969 = n12017 & ~n12968 ;
  assign n12970 = ~n11979 & n12544 ;
  assign n12971 = ~n12559 & ~n12970 ;
  assign n12972 = ~n12969 & n12971 ;
  assign n12973 = ~n11973 & ~n12972 ;
  assign n12990 = n12552 & n12980 ;
  assign n12991 = ~n12043 & ~n12966 ;
  assign n12992 = n12003 & ~n12991 ;
  assign n12993 = ~n12990 & ~n12992 ;
  assign n12994 = ~n12973 & n12993 ;
  assign n12995 = ~n12989 & n12994 ;
  assign n12996 = \u2_L9_reg[23]/NET0131  & ~n12995 ;
  assign n12997 = ~\u2_L9_reg[23]/NET0131  & n12995 ;
  assign n12998 = ~n12996 & ~n12997 ;
  assign n13001 = ~n12316 & ~n12338 ;
  assign n13002 = ~n12630 & n13001 ;
  assign n13003 = ~n12286 & ~n13002 ;
  assign n12999 = n12286 & ~n12300 ;
  assign n13000 = ~n12514 & n12999 ;
  assign n13004 = ~n12293 & ~n12629 ;
  assign n13005 = ~n12330 & n13004 ;
  assign n13006 = ~n13000 & n13005 ;
  assign n13007 = ~n13003 & n13006 ;
  assign n13008 = n12311 & ~n13007 ;
  assign n13012 = ~n12278 & n12286 ;
  assign n13011 = ~n12271 & n12277 ;
  assign n13013 = ~n12612 & ~n13011 ;
  assign n13014 = n13012 & n13013 ;
  assign n13010 = n12313 & n12318 ;
  assign n13015 = ~n12615 & ~n13010 ;
  assign n13016 = ~n12321 & n13015 ;
  assign n13017 = ~n13014 & n13016 ;
  assign n13018 = ~n12311 & ~n13017 ;
  assign n13019 = ~n12320 & ~n12323 ;
  assign n13020 = ~n12286 & ~n13019 ;
  assign n13009 = n12331 & n12616 ;
  assign n13021 = ~n12317 & ~n13009 ;
  assign n13022 = ~n13020 & n13021 ;
  assign n13023 = ~n13018 & n13022 ;
  assign n13024 = ~n13008 & n13023 ;
  assign n13025 = ~\u2_L9_reg[27]/NET0131  & ~n13024 ;
  assign n13026 = \u2_L9_reg[27]/NET0131  & n13024 ;
  assign n13027 = ~n13025 & ~n13026 ;
  assign n13035 = ~n11932 & ~n11947 ;
  assign n13036 = ~n12386 & n13035 ;
  assign n13037 = ~n11918 & ~n13036 ;
  assign n13038 = n11895 & ~n11937 ;
  assign n13039 = ~n13037 & n13038 ;
  assign n13028 = n11905 & ~n11912 ;
  assign n13029 = n11888 & n13028 ;
  assign n13030 = ~n11916 & ~n11935 ;
  assign n13031 = n11889 & ~n13030 ;
  assign n13032 = ~n11937 & ~n12400 ;
  assign n13033 = ~n13031 & n13032 ;
  assign n13034 = ~n11895 & ~n13033 ;
  assign n13040 = ~n13029 & ~n13034 ;
  assign n13041 = ~n13039 & n13040 ;
  assign n13042 = n11930 & ~n13041 ;
  assign n13044 = ~n11882 & n11916 ;
  assign n13045 = n12404 & ~n13044 ;
  assign n13043 = n11902 & ~n13035 ;
  assign n13046 = n12383 & ~n12387 ;
  assign n13047 = ~n13043 & ~n13046 ;
  assign n13048 = n11939 & n13047 ;
  assign n13049 = ~n13045 & n13048 ;
  assign n13050 = ~n11930 & ~n13049 ;
  assign n13051 = n11895 & n11936 ;
  assign n13052 = ~n11932 & n11944 ;
  assign n13053 = n11906 & n13052 ;
  assign n13054 = ~n13051 & ~n13053 ;
  assign n13055 = ~n13050 & n13054 ;
  assign n13056 = ~n13042 & n13055 ;
  assign n13057 = \u2_L9_reg[32]/NET0131  & n13056 ;
  assign n13058 = ~\u2_L9_reg[32]/NET0131  & ~n13056 ;
  assign n13059 = ~n13057 & ~n13058 ;
  assign n13093 = decrypt_pad & ~\u2_uk_K_r9_reg[55]/NET0131  ;
  assign n13094 = ~decrypt_pad & ~\u2_uk_K_r9_reg[4]/NET0131  ;
  assign n13095 = ~n13093 & ~n13094 ;
  assign n13096 = \u2_R9_reg[12]/NET0131  & ~n13095 ;
  assign n13097 = ~\u2_R9_reg[12]/NET0131  & n13095 ;
  assign n13098 = ~n13096 & ~n13097 ;
  assign n13060 = decrypt_pad & ~\u2_uk_K_r9_reg[11]/NET0131  ;
  assign n13061 = ~decrypt_pad & ~\u2_uk_K_r9_reg[17]/NET0131  ;
  assign n13062 = ~n13060 & ~n13061 ;
  assign n13063 = \u2_R9_reg[13]/NET0131  & ~n13062 ;
  assign n13064 = ~\u2_R9_reg[13]/NET0131  & n13062 ;
  assign n13065 = ~n13063 & ~n13064 ;
  assign n13073 = decrypt_pad & ~\u2_uk_K_r9_reg[34]/NET0131  ;
  assign n13074 = ~decrypt_pad & ~\u2_uk_K_r9_reg[40]/NET0131  ;
  assign n13075 = ~n13073 & ~n13074 ;
  assign n13076 = \u2_R9_reg[8]/NET0131  & ~n13075 ;
  assign n13077 = ~\u2_R9_reg[8]/NET0131  & n13075 ;
  assign n13078 = ~n13076 & ~n13077 ;
  assign n13080 = ~n13065 & ~n13078 ;
  assign n13081 = n13065 & n13078 ;
  assign n13082 = ~n13080 & ~n13081 ;
  assign n13066 = decrypt_pad & ~\u2_uk_K_r9_reg[6]/NET0131  ;
  assign n13067 = ~decrypt_pad & ~\u2_uk_K_r9_reg[12]/NET0131  ;
  assign n13068 = ~n13066 & ~n13067 ;
  assign n13069 = \u2_R9_reg[9]/NET0131  & ~n13068 ;
  assign n13070 = ~\u2_R9_reg[9]/NET0131  & n13068 ;
  assign n13071 = ~n13069 & ~n13070 ;
  assign n13083 = decrypt_pad & ~\u2_uk_K_r9_reg[39]/NET0131  ;
  assign n13084 = ~decrypt_pad & ~\u2_uk_K_r9_reg[20]/NET0131  ;
  assign n13085 = ~n13083 & ~n13084 ;
  assign n13086 = \u2_R9_reg[10]/NET0131  & ~n13085 ;
  assign n13087 = ~\u2_R9_reg[10]/NET0131  & n13085 ;
  assign n13088 = ~n13086 & ~n13087 ;
  assign n13134 = ~n13071 & n13088 ;
  assign n13135 = ~n13082 & n13134 ;
  assign n13123 = n13065 & ~n13078 ;
  assign n13124 = n13071 & n13123 ;
  assign n13105 = decrypt_pad & ~\u2_uk_K_r9_reg[40]/NET0131  ;
  assign n13106 = ~decrypt_pad & ~\u2_uk_K_r9_reg[46]/NET0131  ;
  assign n13107 = ~n13105 & ~n13106 ;
  assign n13108 = \u2_R9_reg[11]/NET0131  & ~n13107 ;
  assign n13109 = ~\u2_R9_reg[11]/NET0131  & n13107 ;
  assign n13110 = ~n13108 & ~n13109 ;
  assign n13125 = n13088 & ~n13110 ;
  assign n13126 = n13124 & n13125 ;
  assign n13131 = ~n13065 & n13071 ;
  assign n13132 = n13088 & n13131 ;
  assign n13133 = n13078 & n13132 ;
  assign n13136 = ~n13126 & ~n13133 ;
  assign n13137 = ~n13135 & n13136 ;
  assign n13116 = n13071 & ~n13088 ;
  assign n13127 = n13065 & n13110 ;
  assign n13128 = n13082 & ~n13127 ;
  assign n13129 = n13116 & ~n13128 ;
  assign n13100 = ~n13071 & ~n13088 ;
  assign n13130 = n13100 & n13128 ;
  assign n13138 = ~n13129 & ~n13130 ;
  assign n13139 = n13137 & n13138 ;
  assign n13140 = ~n13098 & ~n13139 ;
  assign n13072 = n13065 & ~n13071 ;
  assign n13079 = ~n13071 & n13078 ;
  assign n13089 = ~n13078 & ~n13088 ;
  assign n13090 = ~n13079 & ~n13089 ;
  assign n13091 = n13082 & n13090 ;
  assign n13092 = ~n13072 & ~n13091 ;
  assign n13099 = ~n13092 & n13098 ;
  assign n13101 = n13080 & n13100 ;
  assign n13102 = n13072 & n13088 ;
  assign n13103 = ~n13101 & ~n13102 ;
  assign n13104 = ~n13099 & n13103 ;
  assign n13111 = ~n13104 & n13110 ;
  assign n13112 = n13088 & n13098 ;
  assign n13113 = n13071 & n13080 ;
  assign n13114 = n13112 & n13113 ;
  assign n13115 = n13098 & ~n13110 ;
  assign n13117 = n13065 & n13116 ;
  assign n13118 = ~n13065 & n13079 ;
  assign n13119 = n13071 & n13081 ;
  assign n13120 = ~n13118 & ~n13119 ;
  assign n13121 = ~n13117 & n13120 ;
  assign n13122 = n13115 & ~n13121 ;
  assign n13141 = ~n13114 & ~n13122 ;
  assign n13142 = ~n13111 & n13141 ;
  assign n13143 = ~n13140 & n13142 ;
  assign n13144 = ~\u2_L9_reg[6]/NET0131  & ~n13143 ;
  assign n13145 = \u2_L9_reg[6]/NET0131  & n13143 ;
  assign n13146 = ~n13144 & ~n13145 ;
  assign n13151 = ~n11901 & ~n11954 ;
  assign n13147 = n11888 & ~n13030 ;
  assign n13152 = ~n13028 & ~n13147 ;
  assign n13153 = ~n13151 & n13152 ;
  assign n13154 = ~n11895 & ~n13153 ;
  assign n13148 = ~n11948 & ~n13147 ;
  assign n13149 = n11882 & ~n13148 ;
  assign n13155 = ~n11882 & ~n11940 ;
  assign n13156 = n13030 & n13155 ;
  assign n13157 = n11895 & n13156 ;
  assign n13158 = ~n13149 & ~n13157 ;
  assign n13159 = ~n13154 & n13158 ;
  assign n13160 = n11930 & ~n13159 ;
  assign n13161 = ~n11895 & n13156 ;
  assign n13162 = ~n11919 & ~n13161 ;
  assign n13163 = ~n11930 & ~n13162 ;
  assign n13150 = ~n11895 & n13149 ;
  assign n13164 = n11953 & ~n13030 ;
  assign n13168 = n11895 & ~n13164 ;
  assign n13165 = n11882 & ~n11947 ;
  assign n13166 = n13030 & ~n13165 ;
  assign n13167 = ~n11919 & n11930 ;
  assign n13169 = ~n13166 & ~n13167 ;
  assign n13170 = n13168 & n13169 ;
  assign n13171 = ~n13150 & ~n13170 ;
  assign n13172 = ~n13163 & n13171 ;
  assign n13173 = ~n13160 & n13172 ;
  assign n13174 = ~\u2_L9_reg[7]/NET0131  & ~n13173 ;
  assign n13175 = \u2_L9_reg[7]/NET0131  & n13173 ;
  assign n13176 = ~n13174 & ~n13175 ;
  assign n13178 = ~n12426 & n12467 ;
  assign n13179 = ~n12465 & ~n13178 ;
  assign n13180 = n12452 & ~n13179 ;
  assign n13181 = n12458 & ~n12497 ;
  assign n13182 = ~n12455 & ~n13181 ;
  assign n13183 = ~n12452 & ~n13182 ;
  assign n13184 = ~n12434 & n12649 ;
  assign n13185 = ~n13183 & n13184 ;
  assign n13186 = ~n13180 & n13185 ;
  assign n13187 = ~n12477 & ~n13186 ;
  assign n13191 = ~n12426 & n12457 ;
  assign n13192 = ~n12455 & ~n13191 ;
  assign n13193 = n12452 & ~n13192 ;
  assign n13194 = n12433 & n12657 ;
  assign n13195 = ~n12500 & ~n13194 ;
  assign n13196 = ~n13193 & n13195 ;
  assign n13197 = n12477 & ~n13196 ;
  assign n13177 = n12444 & n12665 ;
  assign n13188 = n12434 & n12441 ;
  assign n13189 = n12499 & ~n13188 ;
  assign n13190 = n12452 & ~n13189 ;
  assign n13198 = ~n13177 & ~n13190 ;
  assign n13199 = ~n13197 & n13198 ;
  assign n13200 = ~n13187 & n13199 ;
  assign n13201 = ~\u2_L9_reg[8]/NET0131  & ~n13200 ;
  assign n13202 = \u2_L9_reg[8]/NET0131  & n13200 ;
  assign n13203 = ~n13201 & ~n13202 ;
  assign n13204 = n13088 & ~n13124 ;
  assign n13206 = n13110 & n13113 ;
  assign n13205 = n13072 & ~n13078 ;
  assign n13207 = ~n13088 & ~n13205 ;
  assign n13208 = n13120 & n13207 ;
  assign n13209 = ~n13206 & n13208 ;
  assign n13210 = ~n13204 & ~n13209 ;
  assign n13211 = n13080 & n13088 ;
  assign n13212 = ~n13071 & n13211 ;
  assign n13213 = n13110 & ~n13133 ;
  assign n13214 = ~n13212 & n13213 ;
  assign n13215 = n13078 & n13088 ;
  assign n13216 = ~n13065 & ~n13089 ;
  assign n13217 = ~n13215 & n13216 ;
  assign n13218 = ~n13214 & n13217 ;
  assign n13219 = ~n13210 & ~n13218 ;
  assign n13220 = n13098 & ~n13219 ;
  assign n13221 = ~n13071 & n13215 ;
  assign n13222 = ~n13110 & ~n13221 ;
  assign n13223 = ~n13214 & ~n13222 ;
  assign n13228 = n13080 & ~n13088 ;
  assign n13229 = ~n13119 & ~n13205 ;
  assign n13230 = ~n13228 & n13229 ;
  assign n13231 = ~n13110 & ~n13230 ;
  assign n13225 = ~n13080 & n13110 ;
  assign n13224 = ~n13071 & ~n13081 ;
  assign n13226 = ~n13119 & ~n13224 ;
  assign n13227 = n13225 & n13226 ;
  assign n13232 = ~n13101 & ~n13227 ;
  assign n13233 = ~n13231 & n13232 ;
  assign n13234 = ~n13098 & ~n13233 ;
  assign n13235 = ~n13223 & ~n13234 ;
  assign n13236 = ~n13220 & n13235 ;
  assign n13237 = ~\u2_L9_reg[16]/NET0131  & ~n13236 ;
  assign n13238 = \u2_L9_reg[16]/NET0131  & n13236 ;
  assign n13239 = ~n13237 & ~n13238 ;
  assign n13249 = ~n13088 & n13110 ;
  assign n13260 = ~n13071 & ~n13123 ;
  assign n13261 = n13249 & n13260 ;
  assign n13256 = ~n13100 & ~n13110 ;
  assign n13257 = ~n13082 & n13256 ;
  assign n13258 = ~n13079 & n13088 ;
  assign n13259 = n13225 & n13258 ;
  assign n13262 = ~n13257 & ~n13259 ;
  assign n13263 = ~n13261 & n13262 ;
  assign n13264 = ~n13130 & n13263 ;
  assign n13265 = n13098 & ~n13264 ;
  assign n13240 = n13065 & n13089 ;
  assign n13241 = ~n13211 & ~n13240 ;
  assign n13242 = ~n13113 & ~n13221 ;
  assign n13243 = n13241 & n13242 ;
  assign n13244 = n13110 & ~n13243 ;
  assign n13245 = ~n13065 & n13221 ;
  assign n13246 = ~n13244 & ~n13245 ;
  assign n13247 = ~n13098 & ~n13246 ;
  assign n13252 = ~n13082 & n13100 ;
  assign n13253 = ~n13091 & ~n13252 ;
  assign n13254 = ~n13098 & ~n13110 ;
  assign n13255 = ~n13253 & n13254 ;
  assign n13248 = n13119 & n13125 ;
  assign n13250 = ~n13118 & ~n13124 ;
  assign n13251 = n13249 & ~n13250 ;
  assign n13266 = ~n13248 & ~n13251 ;
  assign n13267 = ~n13255 & n13266 ;
  assign n13268 = ~n13247 & n13267 ;
  assign n13269 = ~n13265 & n13268 ;
  assign n13270 = ~\u2_L9_reg[24]/NET0131  & ~n13269 ;
  assign n13271 = \u2_L9_reg[24]/NET0131  & n13269 ;
  assign n13272 = ~n13270 & ~n13271 ;
  assign n13274 = ~n13088 & n13118 ;
  assign n13275 = n13241 & ~n13274 ;
  assign n13276 = n13098 & ~n13275 ;
  assign n13277 = ~n13131 & ~n13215 ;
  assign n13278 = ~n13098 & ~n13132 ;
  assign n13279 = ~n13277 & n13278 ;
  assign n13280 = ~n13276 & ~n13279 ;
  assign n13281 = n13110 & ~n13280 ;
  assign n13285 = n13088 & n13205 ;
  assign n13282 = ~n13071 & ~n13078 ;
  assign n13283 = ~n13110 & ~n13282 ;
  assign n13284 = n13277 & n13283 ;
  assign n13286 = ~n13252 & ~n13284 ;
  assign n13287 = ~n13285 & n13286 ;
  assign n13288 = ~n13098 & ~n13287 ;
  assign n13289 = ~n13113 & ~n13215 ;
  assign n13290 = n13115 & ~n13289 ;
  assign n13292 = n13071 & ~n13081 ;
  assign n13293 = n13112 & n13292 ;
  assign n13273 = n13125 & n13131 ;
  assign n13291 = n13127 & n13221 ;
  assign n13294 = ~n13273 & ~n13291 ;
  assign n13295 = ~n13293 & n13294 ;
  assign n13296 = ~n13290 & n13295 ;
  assign n13297 = ~n13288 & n13296 ;
  assign n13298 = ~n13281 & n13297 ;
  assign n13299 = \u2_L9_reg[30]/NET0131  & ~n13298 ;
  assign n13300 = ~\u2_L9_reg[30]/NET0131  & n13298 ;
  assign n13301 = ~n13299 & ~n13300 ;
  assign n13302 = n12420 & n12442 ;
  assign n13303 = n12444 & n12497 ;
  assign n13304 = n12477 & ~n13303 ;
  assign n13305 = ~n13302 & n13304 ;
  assign n13306 = ~n12444 & n12497 ;
  assign n13307 = ~n12477 & ~n13306 ;
  assign n13308 = ~n12444 & ~n12658 ;
  assign n13309 = ~n12455 & ~n13308 ;
  assign n13310 = n13307 & n13309 ;
  assign n13311 = ~n13305 & ~n13310 ;
  assign n13312 = ~n12452 & ~n12492 ;
  assign n13313 = ~n12503 & ~n13191 ;
  assign n13314 = n13312 & n13313 ;
  assign n13315 = ~n13311 & n13314 ;
  assign n13316 = n12433 & n12658 ;
  assign n13317 = ~n12433 & n12479 ;
  assign n13318 = ~n13316 & ~n13317 ;
  assign n13319 = n13304 & n13318 ;
  assign n13320 = ~n12433 & n12658 ;
  assign n13321 = ~n12445 & ~n13320 ;
  assign n13322 = n13307 & n13321 ;
  assign n13323 = ~n13319 & ~n13322 ;
  assign n13324 = n12452 & ~n12498 ;
  assign n13325 = ~n13178 & n13324 ;
  assign n13326 = ~n13323 & n13325 ;
  assign n13327 = ~n13315 & ~n13326 ;
  assign n13328 = ~\u2_L9_reg[3]/NET0131  & n13327 ;
  assign n13329 = \u2_L9_reg[3]/NET0131  & ~n13327 ;
  assign n13330 = ~n13328 & ~n13329 ;
  assign n13336 = ~n12007 & ~n12029 ;
  assign n13337 = ~n12966 & n13336 ;
  assign n13338 = n11973 & ~n13337 ;
  assign n13331 = n11979 & ~n12022 ;
  assign n13332 = ~n12007 & ~n13331 ;
  assign n13333 = ~n11973 & n13332 ;
  assign n13334 = ~n12032 & ~n12549 ;
  assign n13335 = ~n12560 & ~n13334 ;
  assign n13339 = ~n13333 & ~n13335 ;
  assign n13340 = ~n13338 & n13339 ;
  assign n13341 = ~n12017 & ~n13340 ;
  assign n13342 = ~n11992 & n12552 ;
  assign n13343 = ~n12001 & n12041 ;
  assign n13344 = ~n13342 & ~n13343 ;
  assign n13345 = ~n11973 & ~n13344 ;
  assign n13346 = n12553 & n12967 ;
  assign n13347 = n11992 & ~n13346 ;
  assign n13348 = n12003 & n13332 ;
  assign n13349 = ~n12559 & ~n13348 ;
  assign n13350 = ~n13347 & n13349 ;
  assign n13351 = n12017 & ~n13350 ;
  assign n13352 = ~n13345 & ~n13351 ;
  assign n13353 = ~n13341 & n13352 ;
  assign n13354 = ~\u2_L9_reg[9]/NET0131  & ~n13353 ;
  assign n13355 = \u2_L9_reg[9]/NET0131  & n13353 ;
  assign n13356 = ~n13354 & ~n13355 ;
  assign n13363 = n12727 & ~n12838 ;
  assign n13359 = n12691 & n12711 ;
  assign n13360 = n12704 & ~n12727 ;
  assign n13361 = ~n12837 & n13360 ;
  assign n13362 = ~n13359 & n13361 ;
  assign n13364 = n12745 & ~n12865 ;
  assign n13365 = ~n13362 & n13364 ;
  assign n13366 = ~n13363 & n13365 ;
  assign n13357 = n12697 & ~n12727 ;
  assign n13369 = n12704 & n12711 ;
  assign n13370 = ~n12842 & n13369 ;
  assign n13371 = ~n13357 & n13370 ;
  assign n13367 = ~n12704 & ~n12832 ;
  assign n13368 = n12851 & n13367 ;
  assign n13372 = ~n12858 & ~n13368 ;
  assign n13373 = ~n13371 & n13372 ;
  assign n13374 = n12751 & n13373 ;
  assign n13375 = ~n13366 & ~n13374 ;
  assign n13358 = n12718 & n13357 ;
  assign n13376 = n12704 & n13359 ;
  assign n13377 = ~n12912 & ~n13376 ;
  assign n13378 = n12727 & ~n13377 ;
  assign n13379 = ~n13358 & ~n13378 ;
  assign n13380 = ~n13375 & n13379 ;
  assign n13381 = ~\u2_L9_reg[18]/P0001  & ~n13380 ;
  assign n13382 = \u2_L9_reg[18]/P0001  & n13380 ;
  assign n13383 = ~n13381 & ~n13382 ;
  assign n13411 = decrypt_pad & ~\u2_uk_K_r8_reg[33]/NET0131  ;
  assign n13412 = ~decrypt_pad & ~\u2_uk_K_r8_reg[11]/NET0131  ;
  assign n13413 = ~n13411 & ~n13412 ;
  assign n13414 = \u2_R8_reg[4]/NET0131  & ~n13413 ;
  assign n13415 = ~\u2_R8_reg[4]/NET0131  & n13413 ;
  assign n13416 = ~n13414 & ~n13415 ;
  assign n13397 = decrypt_pad & ~\u2_uk_K_r8_reg[46]/NET0131  ;
  assign n13398 = ~decrypt_pad & ~\u2_uk_K_r8_reg[24]/NET0131  ;
  assign n13399 = ~n13397 & ~n13398 ;
  assign n13400 = \u2_R8_reg[2]/NET0131  & ~n13399 ;
  assign n13401 = ~\u2_R8_reg[2]/NET0131  & n13399 ;
  assign n13402 = ~n13400 & ~n13401 ;
  assign n13417 = decrypt_pad & ~\u2_uk_K_r8_reg[4]/NET0131  ;
  assign n13418 = ~decrypt_pad & ~\u2_uk_K_r8_reg[39]/NET0131  ;
  assign n13419 = ~n13417 & ~n13418 ;
  assign n13420 = \u2_R8_reg[5]/NET0131  & ~n13419 ;
  assign n13421 = ~\u2_R8_reg[5]/NET0131  & n13419 ;
  assign n13422 = ~n13420 & ~n13421 ;
  assign n13431 = ~n13402 & ~n13422 ;
  assign n13432 = n13402 & n13422 ;
  assign n13433 = ~n13431 & ~n13432 ;
  assign n13403 = decrypt_pad & ~\u2_uk_K_r8_reg[55]/NET0131  ;
  assign n13404 = ~decrypt_pad & ~\u2_uk_K_r8_reg[33]/NET0131  ;
  assign n13405 = ~n13403 & ~n13404 ;
  assign n13406 = \u2_R8_reg[3]/NET0131  & ~n13405 ;
  assign n13407 = ~\u2_R8_reg[3]/NET0131  & n13405 ;
  assign n13408 = ~n13406 & ~n13407 ;
  assign n13434 = ~n13408 & n13422 ;
  assign n13384 = decrypt_pad & ~\u2_uk_K_r8_reg[10]/NET0131  ;
  assign n13385 = ~decrypt_pad & ~\u2_uk_K_r8_reg[20]/NET0131  ;
  assign n13386 = ~n13384 & ~n13385 ;
  assign n13387 = \u2_R8_reg[32]/NET0131  & ~n13386 ;
  assign n13388 = ~\u2_R8_reg[32]/NET0131  & n13386 ;
  assign n13389 = ~n13387 & ~n13388 ;
  assign n13390 = decrypt_pad & ~\u2_uk_K_r8_reg[6]/NET0131  ;
  assign n13391 = ~decrypt_pad & ~\u2_uk_K_r8_reg[41]/NET0131  ;
  assign n13392 = ~n13390 & ~n13391 ;
  assign n13393 = \u2_R8_reg[1]/NET0131  & ~n13392 ;
  assign n13394 = ~\u2_R8_reg[1]/NET0131  & n13392 ;
  assign n13395 = ~n13393 & ~n13394 ;
  assign n13435 = ~n13389 & n13395 ;
  assign n13436 = ~n13434 & n13435 ;
  assign n13437 = ~n13433 & n13436 ;
  assign n13423 = n13402 & ~n13422 ;
  assign n13424 = n13389 & n13395 ;
  assign n13425 = n13423 & n13424 ;
  assign n13426 = n13408 & n13425 ;
  assign n13427 = n13395 & ~n13408 ;
  assign n13428 = n13389 & ~n13402 ;
  assign n13429 = n13422 & n13428 ;
  assign n13430 = ~n13427 & n13429 ;
  assign n13438 = ~n13426 & ~n13430 ;
  assign n13439 = ~n13437 & n13438 ;
  assign n13440 = ~n13416 & ~n13439 ;
  assign n13396 = n13389 & ~n13395 ;
  assign n13409 = ~n13402 & n13408 ;
  assign n13410 = n13396 & n13409 ;
  assign n13465 = ~n13395 & ~n13422 ;
  assign n13464 = ~n13389 & n13408 ;
  assign n13466 = n13402 & n13464 ;
  assign n13467 = n13465 & n13466 ;
  assign n13468 = ~n13410 & ~n13467 ;
  assign n13469 = ~n13440 & n13468 ;
  assign n13441 = ~n13395 & n13422 ;
  assign n13444 = ~n13389 & ~n13402 ;
  assign n13445 = ~n13441 & n13444 ;
  assign n13446 = n13396 & n13423 ;
  assign n13447 = ~n13445 & ~n13446 ;
  assign n13448 = ~n13416 & ~n13447 ;
  assign n13442 = ~n13389 & n13402 ;
  assign n13443 = n13441 & n13442 ;
  assign n13449 = n13395 & ~n13442 ;
  assign n13450 = ~n13433 & n13449 ;
  assign n13451 = ~n13443 & ~n13450 ;
  assign n13452 = ~n13448 & n13451 ;
  assign n13453 = ~n13408 & ~n13452 ;
  assign n13458 = n13408 & ~n13432 ;
  assign n13459 = n13395 & ~n13458 ;
  assign n13460 = ~n13431 & ~n13459 ;
  assign n13461 = ~n13389 & ~n13460 ;
  assign n13454 = ~n13395 & ~n13423 ;
  assign n13455 = ~n13434 & n13454 ;
  assign n13456 = n13389 & ~n13427 ;
  assign n13457 = ~n13455 & n13456 ;
  assign n13462 = n13416 & ~n13457 ;
  assign n13463 = ~n13461 & n13462 ;
  assign n13470 = ~n13453 & ~n13463 ;
  assign n13471 = n13469 & n13470 ;
  assign n13472 = ~\u2_L8_reg[31]/NET0131  & ~n13471 ;
  assign n13473 = \u2_L8_reg[31]/NET0131  & n13471 ;
  assign n13474 = ~n13472 & ~n13473 ;
  assign n13526 = decrypt_pad & ~\u2_uk_K_r8_reg[2]/NET0131  ;
  assign n13527 = ~decrypt_pad & ~\u2_uk_K_r8_reg[37]/P0001  ;
  assign n13528 = ~n13526 & ~n13527 ;
  assign n13529 = \u2_R8_reg[24]/NET0131  & ~n13528 ;
  assign n13530 = ~\u2_R8_reg[24]/NET0131  & n13528 ;
  assign n13531 = ~n13529 & ~n13530 ;
  assign n13481 = decrypt_pad & ~\u2_uk_K_r8_reg[36]/NET0131  ;
  assign n13482 = ~decrypt_pad & ~\u2_uk_K_r8_reg[16]/NET0131  ;
  assign n13483 = ~n13481 & ~n13482 ;
  assign n13484 = \u2_R8_reg[20]/NET0131  & ~n13483 ;
  assign n13485 = ~\u2_R8_reg[20]/NET0131  & n13483 ;
  assign n13486 = ~n13484 & ~n13485 ;
  assign n13494 = decrypt_pad & ~\u2_uk_K_r8_reg[42]/NET0131  ;
  assign n13495 = ~decrypt_pad & ~\u2_uk_K_r8_reg[22]/NET0131  ;
  assign n13496 = ~n13494 & ~n13495 ;
  assign n13497 = \u2_R8_reg[22]/NET0131  & ~n13496 ;
  assign n13498 = ~\u2_R8_reg[22]/NET0131  & n13496 ;
  assign n13499 = ~n13497 & ~n13498 ;
  assign n13500 = decrypt_pad & ~\u2_uk_K_r8_reg[51]/NET0131  ;
  assign n13501 = ~decrypt_pad & ~\u2_uk_K_r8_reg[0]/NET0131  ;
  assign n13502 = ~n13500 & ~n13501 ;
  assign n13503 = \u2_R8_reg[21]/NET0131  & ~n13502 ;
  assign n13504 = ~\u2_R8_reg[21]/NET0131  & n13502 ;
  assign n13505 = ~n13503 & ~n13504 ;
  assign n13535 = ~n13499 & n13505 ;
  assign n13551 = n13486 & n13535 ;
  assign n13475 = decrypt_pad & ~\u2_uk_K_r8_reg[0]/NET0131  ;
  assign n13476 = ~decrypt_pad & ~\u2_uk_K_r8_reg[35]/NET0131  ;
  assign n13477 = ~n13475 & ~n13476 ;
  assign n13478 = \u2_R8_reg[23]/NET0131  & ~n13477 ;
  assign n13479 = ~\u2_R8_reg[23]/NET0131  & n13477 ;
  assign n13480 = ~n13478 & ~n13479 ;
  assign n13508 = ~n13486 & n13505 ;
  assign n13509 = n13499 & n13508 ;
  assign n13552 = ~n13480 & ~n13509 ;
  assign n13553 = ~n13551 & n13552 ;
  assign n13487 = decrypt_pad & ~\u2_uk_K_r8_reg[21]/NET0131  ;
  assign n13488 = ~decrypt_pad & ~\u2_uk_K_r8_reg[1]/NET0131  ;
  assign n13489 = ~n13487 & ~n13488 ;
  assign n13490 = \u2_R8_reg[25]/NET0131  & ~n13489 ;
  assign n13491 = ~\u2_R8_reg[25]/NET0131  & n13489 ;
  assign n13492 = ~n13490 & ~n13491 ;
  assign n13543 = n13492 & ~n13505 ;
  assign n13544 = ~n13486 & n13543 ;
  assign n13545 = n13480 & ~n13544 ;
  assign n13554 = n13499 & ~n13505 ;
  assign n13555 = n13486 & n13554 ;
  assign n13556 = ~n13486 & ~n13499 ;
  assign n13557 = ~n13555 & ~n13556 ;
  assign n13558 = n13545 & n13557 ;
  assign n13559 = ~n13553 & ~n13558 ;
  assign n13510 = n13486 & n13492 ;
  assign n13521 = ~n13505 & n13510 ;
  assign n13548 = n13499 & n13521 ;
  assign n13493 = n13486 & ~n13492 ;
  assign n13515 = ~n13480 & ~n13499 ;
  assign n13549 = ~n13515 & ~n13535 ;
  assign n13550 = n13493 & ~n13549 ;
  assign n13560 = ~n13548 & ~n13550 ;
  assign n13561 = ~n13559 & n13560 ;
  assign n13562 = ~n13531 & ~n13561 ;
  assign n13511 = n13505 & n13510 ;
  assign n13506 = ~n13499 & ~n13505 ;
  assign n13507 = n13493 & n13506 ;
  assign n13512 = ~n13507 & ~n13509 ;
  assign n13513 = ~n13511 & n13512 ;
  assign n13514 = n13480 & ~n13513 ;
  assign n13516 = ~n13508 & ~n13510 ;
  assign n13517 = ~n13480 & n13516 ;
  assign n13518 = ~n13515 & ~n13517 ;
  assign n13519 = n13492 & n13505 ;
  assign n13520 = ~n13486 & n13519 ;
  assign n13522 = ~n13499 & ~n13520 ;
  assign n13523 = ~n13521 & n13522 ;
  assign n13524 = ~n13518 & ~n13523 ;
  assign n13525 = ~n13514 & ~n13524 ;
  assign n13532 = ~n13525 & n13531 ;
  assign n13541 = n13493 & n13505 ;
  assign n13542 = ~n13480 & ~n13541 ;
  assign n13546 = ~n13499 & ~n13542 ;
  assign n13547 = ~n13545 & n13546 ;
  assign n13536 = ~n13510 & ~n13535 ;
  assign n13533 = ~n13486 & ~n13492 ;
  assign n13534 = ~n13499 & ~n13533 ;
  assign n13537 = n13480 & ~n13534 ;
  assign n13538 = ~n13536 & n13537 ;
  assign n13539 = ~n13505 & n13533 ;
  assign n13540 = n13515 & n13539 ;
  assign n13563 = ~n13538 & ~n13540 ;
  assign n13564 = ~n13547 & n13563 ;
  assign n13565 = ~n13532 & n13564 ;
  assign n13566 = ~n13562 & n13565 ;
  assign n13567 = \u2_L8_reg[11]/NET0131  & ~n13566 ;
  assign n13568 = ~\u2_L8_reg[11]/NET0131  & n13566 ;
  assign n13569 = ~n13567 & ~n13568 ;
  assign n13570 = decrypt_pad & ~\u2_uk_K_r8_reg[22]/NET0131  ;
  assign n13571 = ~decrypt_pad & ~\u2_uk_K_r8_reg[2]/NET0131  ;
  assign n13572 = ~n13570 & ~n13571 ;
  assign n13573 = \u2_R8_reg[27]/NET0131  & ~n13572 ;
  assign n13574 = ~\u2_R8_reg[27]/NET0131  & n13572 ;
  assign n13575 = ~n13573 & ~n13574 ;
  assign n13589 = decrypt_pad & ~\u2_uk_K_r8_reg[52]/NET0131  ;
  assign n13590 = ~decrypt_pad & ~\u2_uk_K_r8_reg[28]/NET0131  ;
  assign n13591 = ~n13589 & ~n13590 ;
  assign n13592 = \u2_R8_reg[24]/NET0131  & ~n13591 ;
  assign n13593 = ~\u2_R8_reg[24]/NET0131  & n13591 ;
  assign n13594 = ~n13592 & ~n13593 ;
  assign n13576 = decrypt_pad & ~\u2_uk_K_r8_reg[28]/NET0131  ;
  assign n13577 = ~decrypt_pad & ~\u2_uk_K_r8_reg[8]/NET0131  ;
  assign n13578 = ~n13576 & ~n13577 ;
  assign n13579 = \u2_R8_reg[25]/NET0131  & ~n13578 ;
  assign n13580 = ~\u2_R8_reg[25]/NET0131  & n13578 ;
  assign n13581 = ~n13579 & ~n13580 ;
  assign n13595 = decrypt_pad & ~\u2_uk_K_r8_reg[1]/NET0131  ;
  assign n13596 = ~decrypt_pad & ~\u2_uk_K_r8_reg[36]/NET0131  ;
  assign n13597 = ~n13595 & ~n13596 ;
  assign n13598 = \u2_R8_reg[29]/NET0131  & ~n13597 ;
  assign n13599 = ~\u2_R8_reg[29]/NET0131  & n13597 ;
  assign n13600 = ~n13598 & ~n13599 ;
  assign n13643 = ~n13581 & ~n13600 ;
  assign n13619 = decrypt_pad & ~\u2_uk_K_r8_reg[9]/NET0131  ;
  assign n13620 = ~decrypt_pad & ~\u2_uk_K_r8_reg[44]/NET0131  ;
  assign n13621 = ~n13619 & ~n13620 ;
  assign n13622 = \u2_R8_reg[28]/NET0131  & ~n13621 ;
  assign n13623 = ~\u2_R8_reg[28]/NET0131  & n13621 ;
  assign n13624 = ~n13622 & ~n13623 ;
  assign n13582 = decrypt_pad & ~\u2_uk_K_r8_reg[44]/NET0131  ;
  assign n13583 = ~decrypt_pad & ~\u2_uk_K_r8_reg[52]/NET0131  ;
  assign n13584 = ~n13582 & ~n13583 ;
  assign n13585 = \u2_R8_reg[26]/NET0131  & ~n13584 ;
  assign n13586 = ~\u2_R8_reg[26]/NET0131  & n13584 ;
  assign n13587 = ~n13585 & ~n13586 ;
  assign n13588 = ~n13581 & n13587 ;
  assign n13644 = n13581 & ~n13587 ;
  assign n13645 = n13600 & n13644 ;
  assign n13646 = ~n13588 & ~n13645 ;
  assign n13647 = n13624 & ~n13646 ;
  assign n13648 = ~n13643 & ~n13647 ;
  assign n13649 = n13594 & ~n13648 ;
  assign n13634 = ~n13594 & n13600 ;
  assign n13635 = n13588 & n13634 ;
  assign n13601 = ~n13594 & ~n13600 ;
  assign n13640 = n13587 & n13601 ;
  assign n13641 = n13581 & n13640 ;
  assign n13642 = ~n13635 & ~n13641 ;
  assign n13613 = ~n13581 & ~n13587 ;
  assign n13650 = ~n13600 & n13613 ;
  assign n13651 = n13642 & ~n13650 ;
  assign n13652 = ~n13649 & n13651 ;
  assign n13653 = n13575 & ~n13652 ;
  assign n13603 = n13587 & n13594 ;
  assign n13604 = ~n13587 & ~n13594 ;
  assign n13605 = ~n13603 & ~n13604 ;
  assign n13606 = n13600 & ~n13605 ;
  assign n13602 = n13588 & n13601 ;
  assign n13607 = n13594 & ~n13600 ;
  assign n13608 = n13581 & n13607 ;
  assign n13609 = ~n13602 & ~n13608 ;
  assign n13610 = ~n13606 & n13609 ;
  assign n13611 = ~n13575 & ~n13610 ;
  assign n13612 = n13581 & n13606 ;
  assign n13614 = ~n13575 & n13600 ;
  assign n13615 = n13594 & n13613 ;
  assign n13616 = ~n13614 & n13615 ;
  assign n13617 = ~n13612 & ~n13616 ;
  assign n13618 = ~n13611 & n13617 ;
  assign n13625 = ~n13618 & ~n13624 ;
  assign n13626 = ~n13575 & n13581 ;
  assign n13627 = ~n13605 & n13626 ;
  assign n13628 = n13594 & n13600 ;
  assign n13629 = n13613 & n13628 ;
  assign n13630 = n13581 & n13600 ;
  assign n13631 = ~n13594 & n13630 ;
  assign n13632 = ~n13629 & ~n13631 ;
  assign n13633 = ~n13575 & ~n13632 ;
  assign n13636 = n13601 & n13613 ;
  assign n13637 = ~n13635 & ~n13636 ;
  assign n13638 = ~n13633 & n13637 ;
  assign n13639 = n13624 & ~n13638 ;
  assign n13654 = ~n13627 & ~n13639 ;
  assign n13655 = ~n13625 & n13654 ;
  assign n13656 = ~n13653 & n13655 ;
  assign n13657 = ~\u2_L8_reg[22]/NET0131  & ~n13656 ;
  assign n13658 = \u2_L8_reg[22]/NET0131  & n13656 ;
  assign n13659 = ~n13657 & ~n13658 ;
  assign n13664 = ~n13435 & ~n13442 ;
  assign n13665 = n13428 & n13441 ;
  assign n13666 = n13664 & ~n13665 ;
  assign n13667 = n13408 & ~n13666 ;
  assign n13668 = ~n13408 & ~n13428 ;
  assign n13669 = n13664 & n13668 ;
  assign n13660 = n13424 & n13431 ;
  assign n13661 = n13416 & ~n13660 ;
  assign n13662 = n13395 & n13422 ;
  assign n13663 = n13402 & n13662 ;
  assign n13670 = n13661 & ~n13663 ;
  assign n13671 = ~n13669 & n13670 ;
  assign n13672 = ~n13667 & n13671 ;
  assign n13675 = n13433 & n13435 ;
  assign n13673 = ~n13465 & ~n13662 ;
  assign n13674 = n13389 & ~n13673 ;
  assign n13676 = n13408 & ~n13674 ;
  assign n13677 = ~n13675 & n13676 ;
  assign n13678 = n13389 & n13422 ;
  assign n13679 = ~n13389 & ~n13422 ;
  assign n13680 = ~n13678 & ~n13679 ;
  assign n13681 = ~n13395 & ~n13680 ;
  assign n13682 = ~n13402 & n13679 ;
  assign n13683 = ~n13408 & ~n13682 ;
  assign n13684 = ~n13681 & n13683 ;
  assign n13685 = ~n13677 & ~n13684 ;
  assign n13686 = ~n13416 & ~n13425 ;
  assign n13687 = ~n13443 & n13686 ;
  assign n13688 = ~n13685 & n13687 ;
  assign n13689 = ~n13672 & ~n13688 ;
  assign n13690 = ~\u2_L8_reg[17]/NET0131  & n13689 ;
  assign n13691 = \u2_L8_reg[17]/NET0131  & ~n13689 ;
  assign n13692 = ~n13690 & ~n13691 ;
  assign n13699 = decrypt_pad & ~\u2_uk_K_r8_reg[27]/NET0131  ;
  assign n13700 = ~decrypt_pad & ~\u2_uk_K_r8_reg[5]/NET0131  ;
  assign n13701 = ~n13699 & ~n13700 ;
  assign n13702 = \u2_R8_reg[15]/NET0131  & ~n13701 ;
  assign n13703 = ~\u2_R8_reg[15]/NET0131  & n13701 ;
  assign n13704 = ~n13702 & ~n13703 ;
  assign n13693 = decrypt_pad & ~\u2_uk_K_r8_reg[18]/NET0131  ;
  assign n13694 = ~decrypt_pad & ~\u2_uk_K_r8_reg[53]/NET0131  ;
  assign n13695 = ~n13693 & ~n13694 ;
  assign n13696 = \u2_R8_reg[13]/NET0131  & ~n13695 ;
  assign n13697 = ~\u2_R8_reg[13]/NET0131  & n13695 ;
  assign n13698 = ~n13696 & ~n13697 ;
  assign n13706 = decrypt_pad & ~\u2_uk_K_r8_reg[24]/NET0131  ;
  assign n13707 = ~decrypt_pad & ~\u2_uk_K_r8_reg[34]/NET0131  ;
  assign n13708 = ~n13706 & ~n13707 ;
  assign n13709 = \u2_R8_reg[12]/NET0131  & ~n13708 ;
  assign n13710 = ~\u2_R8_reg[12]/NET0131  & n13708 ;
  assign n13711 = ~n13709 & ~n13710 ;
  assign n13745 = ~n13698 & ~n13711 ;
  assign n13748 = n13698 & n13711 ;
  assign n13749 = ~n13745 & ~n13748 ;
  assign n13712 = decrypt_pad & ~\u2_uk_K_r8_reg[40]/NET0131  ;
  assign n13713 = ~decrypt_pad & ~\u2_uk_K_r8_reg[18]/NET0131  ;
  assign n13714 = ~n13712 & ~n13713 ;
  assign n13715 = \u2_R8_reg[17]/NET0131  & ~n13714 ;
  assign n13716 = ~\u2_R8_reg[17]/NET0131  & n13714 ;
  assign n13717 = ~n13715 & ~n13716 ;
  assign n13726 = ~n13711 & ~n13717 ;
  assign n13750 = n13711 & n13717 ;
  assign n13751 = ~n13726 & ~n13750 ;
  assign n13752 = ~n13749 & ~n13751 ;
  assign n13753 = n13704 & ~n13752 ;
  assign n13718 = n13711 & ~n13717 ;
  assign n13719 = decrypt_pad & ~\u2_uk_K_r8_reg[19]/NET0131  ;
  assign n13720 = ~decrypt_pad & ~\u2_uk_K_r8_reg[54]/NET0131  ;
  assign n13721 = ~n13719 & ~n13720 ;
  assign n13722 = \u2_R8_reg[14]/NET0131  & ~n13721 ;
  assign n13723 = ~\u2_R8_reg[14]/NET0131  & n13721 ;
  assign n13724 = ~n13722 & ~n13723 ;
  assign n13725 = n13718 & n13724 ;
  assign n13754 = ~n13698 & n13717 ;
  assign n13755 = ~n13704 & ~n13754 ;
  assign n13756 = ~n13725 & n13755 ;
  assign n13757 = ~n13753 & ~n13756 ;
  assign n13742 = n13698 & n13726 ;
  assign n13743 = n13724 & n13742 ;
  assign n13744 = ~n13717 & ~n13724 ;
  assign n13746 = n13744 & n13745 ;
  assign n13747 = ~n13743 & ~n13746 ;
  assign n13739 = n13711 & ~n13724 ;
  assign n13740 = ~n13698 & n13739 ;
  assign n13741 = n13717 & n13740 ;
  assign n13730 = decrypt_pad & ~\u2_uk_K_r8_reg[3]/NET0131  ;
  assign n13731 = ~decrypt_pad & ~\u2_uk_K_r8_reg[13]/P0001  ;
  assign n13732 = ~n13730 & ~n13731 ;
  assign n13733 = \u2_R8_reg[16]/NET0131  & ~n13732 ;
  assign n13734 = ~\u2_R8_reg[16]/NET0131  & n13732 ;
  assign n13735 = ~n13733 & ~n13734 ;
  assign n13736 = n13698 & n13704 ;
  assign n13737 = n13724 & n13736 ;
  assign n13738 = ~n13711 & n13737 ;
  assign n13758 = ~n13735 & ~n13738 ;
  assign n13759 = ~n13741 & n13758 ;
  assign n13760 = n13747 & n13759 ;
  assign n13761 = ~n13757 & n13760 ;
  assign n13762 = n13718 & n13736 ;
  assign n13763 = ~n13711 & n13717 ;
  assign n13764 = n13698 & n13763 ;
  assign n13765 = ~n13724 & n13764 ;
  assign n13766 = ~n13762 & ~n13765 ;
  assign n13767 = ~n13704 & ~n13717 ;
  assign n13768 = n13745 & n13767 ;
  assign n13769 = n13724 & n13768 ;
  assign n13770 = n13717 & n13724 ;
  assign n13771 = n13748 & n13770 ;
  assign n13776 = n13735 & ~n13771 ;
  assign n13777 = ~n13769 & n13776 ;
  assign n13772 = n13704 & n13763 ;
  assign n13773 = ~n13698 & n13772 ;
  assign n13774 = ~n13704 & ~n13724 ;
  assign n13775 = n13749 & n13774 ;
  assign n13778 = ~n13773 & ~n13775 ;
  assign n13779 = n13777 & n13778 ;
  assign n13780 = n13766 & n13779 ;
  assign n13781 = ~n13761 & ~n13780 ;
  assign n13783 = ~n13704 & n13765 ;
  assign n13705 = ~n13698 & n13704 ;
  assign n13727 = ~n13724 & n13726 ;
  assign n13728 = ~n13725 & ~n13727 ;
  assign n13729 = n13705 & ~n13728 ;
  assign n13782 = ~n13724 & n13762 ;
  assign n13784 = ~n13729 & ~n13782 ;
  assign n13785 = ~n13783 & n13784 ;
  assign n13786 = ~n13781 & n13785 ;
  assign n13787 = ~\u2_L8_reg[20]/NET0131  & ~n13786 ;
  assign n13788 = \u2_L8_reg[20]/NET0131  & n13786 ;
  assign n13789 = ~n13787 & ~n13788 ;
  assign n13796 = decrypt_pad & ~\u2_uk_K_r8_reg[39]/NET0131  ;
  assign n13797 = ~decrypt_pad & ~\u2_uk_K_r8_reg[17]/NET0131  ;
  assign n13798 = ~n13796 & ~n13797 ;
  assign n13799 = \u2_R8_reg[9]/NET0131  & ~n13798 ;
  assign n13800 = ~\u2_R8_reg[9]/NET0131  & n13798 ;
  assign n13801 = ~n13799 & ~n13800 ;
  assign n13802 = decrypt_pad & ~\u2_uk_K_r8_reg[47]/NET0131  ;
  assign n13803 = ~decrypt_pad & ~\u2_uk_K_r8_reg[25]/NET0131  ;
  assign n13804 = ~n13802 & ~n13803 ;
  assign n13805 = \u2_R8_reg[4]/NET0131  & ~n13804 ;
  assign n13806 = ~\u2_R8_reg[4]/NET0131  & n13804 ;
  assign n13807 = ~n13805 & ~n13806 ;
  assign n13808 = ~n13801 & n13807 ;
  assign n13835 = n13801 & ~n13807 ;
  assign n13836 = ~n13808 & ~n13835 ;
  assign n13790 = decrypt_pad & ~\u2_uk_K_r8_reg[26]/NET0131  ;
  assign n13791 = ~decrypt_pad & ~\u2_uk_K_r8_reg[4]/NET0131  ;
  assign n13792 = ~n13790 & ~n13791 ;
  assign n13793 = \u2_R8_reg[5]/NET0131  & ~n13792 ;
  assign n13794 = ~\u2_R8_reg[5]/NET0131  & n13792 ;
  assign n13795 = ~n13793 & ~n13794 ;
  assign n13809 = decrypt_pad & ~\u2_uk_K_r8_reg[17]/NET0131  ;
  assign n13810 = ~decrypt_pad & ~\u2_uk_K_r8_reg[27]/NET0131  ;
  assign n13811 = ~n13809 & ~n13810 ;
  assign n13812 = \u2_R8_reg[6]/NET0131  & ~n13811 ;
  assign n13813 = ~\u2_R8_reg[6]/NET0131  & n13811 ;
  assign n13814 = ~n13812 & ~n13813 ;
  assign n13826 = ~n13807 & n13814 ;
  assign n13827 = n13795 & ~n13826 ;
  assign n13828 = decrypt_pad & ~\u2_uk_K_r8_reg[11]/NET0131  ;
  assign n13829 = ~decrypt_pad & ~\u2_uk_K_r8_reg[46]/NET0131  ;
  assign n13830 = ~n13828 & ~n13829 ;
  assign n13831 = \u2_R8_reg[7]/NET0131  & ~n13830 ;
  assign n13832 = ~\u2_R8_reg[7]/NET0131  & n13830 ;
  assign n13833 = ~n13831 & ~n13832 ;
  assign n13837 = n13807 & ~n13814 ;
  assign n13838 = ~n13833 & ~n13837 ;
  assign n13839 = ~n13827 & n13838 ;
  assign n13840 = n13836 & n13839 ;
  assign n13815 = n13808 & ~n13814 ;
  assign n13816 = ~n13795 & n13815 ;
  assign n13820 = decrypt_pad & ~\u2_uk_K_r8_reg[34]/NET0131  ;
  assign n13821 = ~decrypt_pad & ~\u2_uk_K_r8_reg[12]/NET0131  ;
  assign n13822 = ~n13820 & ~n13821 ;
  assign n13823 = \u2_R8_reg[8]/NET0131  & ~n13822 ;
  assign n13824 = ~\u2_R8_reg[8]/NET0131  & n13822 ;
  assign n13825 = ~n13823 & ~n13824 ;
  assign n13841 = ~n13816 & n13825 ;
  assign n13817 = n13795 & n13807 ;
  assign n13818 = ~n13814 & n13817 ;
  assign n13819 = n13801 & n13818 ;
  assign n13834 = n13827 & n13833 ;
  assign n13842 = ~n13819 & ~n13834 ;
  assign n13843 = n13841 & n13842 ;
  assign n13844 = ~n13840 & n13843 ;
  assign n13845 = n13795 & ~n13801 ;
  assign n13846 = ~n13795 & n13801 ;
  assign n13847 = ~n13807 & n13846 ;
  assign n13848 = ~n13845 & ~n13847 ;
  assign n13849 = ~n13814 & ~n13848 ;
  assign n13857 = n13807 & n13814 ;
  assign n13861 = n13833 & n13857 ;
  assign n13862 = n13846 & n13861 ;
  assign n13863 = ~n13825 & ~n13862 ;
  assign n13864 = ~n13849 & n13863 ;
  assign n13851 = n13795 & n13835 ;
  assign n13852 = n13814 & ~n13851 ;
  assign n13850 = ~n13801 & ~n13814 ;
  assign n13853 = ~n13795 & ~n13833 ;
  assign n13854 = ~n13814 & ~n13853 ;
  assign n13855 = ~n13850 & ~n13854 ;
  assign n13856 = ~n13852 & n13855 ;
  assign n13858 = ~n13846 & n13857 ;
  assign n13859 = ~n13847 & ~n13858 ;
  assign n13860 = ~n13833 & ~n13859 ;
  assign n13865 = ~n13856 & ~n13860 ;
  assign n13866 = n13864 & n13865 ;
  assign n13867 = ~n13844 & ~n13866 ;
  assign n13868 = ~n13795 & n13814 ;
  assign n13869 = ~n13807 & n13868 ;
  assign n13870 = ~n13801 & n13869 ;
  assign n13871 = ~n13818 & ~n13870 ;
  assign n13872 = n13833 & ~n13871 ;
  assign n13873 = n13814 & ~n13833 ;
  assign n13874 = ~n13853 & ~n13873 ;
  assign n13875 = n13835 & ~n13868 ;
  assign n13876 = ~n13874 & n13875 ;
  assign n13877 = ~n13872 & ~n13876 ;
  assign n13878 = ~n13867 & n13877 ;
  assign n13879 = \u2_L8_reg[2]/NET0131  & n13878 ;
  assign n13880 = ~\u2_L8_reg[2]/NET0131  & ~n13878 ;
  assign n13881 = ~n13879 & ~n13880 ;
  assign n13898 = n13493 & ~n13505 ;
  assign n13899 = ~n13511 & ~n13898 ;
  assign n13900 = ~n13506 & ~n13509 ;
  assign n13901 = ~n13492 & ~n13900 ;
  assign n13902 = n13899 & ~n13901 ;
  assign n13903 = n13480 & ~n13902 ;
  assign n13882 = n13499 & n13541 ;
  assign n13889 = ~n13499 & ~n13516 ;
  assign n13904 = ~n13882 & ~n13889 ;
  assign n13905 = ~n13480 & ~n13904 ;
  assign n13906 = n13499 & n13544 ;
  assign n13907 = ~n13905 & ~n13906 ;
  assign n13908 = ~n13903 & n13907 ;
  assign n13909 = ~n13531 & ~n13908 ;
  assign n13883 = n13505 & n13556 ;
  assign n13884 = ~n13520 & ~n13883 ;
  assign n13885 = ~n13882 & n13884 ;
  assign n13886 = n13480 & ~n13885 ;
  assign n13890 = n13480 & ~n13543 ;
  assign n13891 = ~n13554 & n13890 ;
  assign n13887 = n13499 & ~n13510 ;
  assign n13888 = ~n13533 & n13887 ;
  assign n13892 = ~n13888 & ~n13889 ;
  assign n13893 = ~n13891 & n13892 ;
  assign n13894 = ~n13886 & ~n13893 ;
  assign n13895 = n13531 & ~n13894 ;
  assign n13896 = n13480 & n13492 ;
  assign n13897 = n13535 & n13896 ;
  assign n13910 = ~n13507 & ~n13897 ;
  assign n13911 = ~n13895 & n13910 ;
  assign n13912 = ~n13909 & n13911 ;
  assign n13913 = \u2_L8_reg[29]/NET0131  & ~n13912 ;
  assign n13914 = ~\u2_L8_reg[29]/NET0131  & n13912 ;
  assign n13915 = ~n13913 & ~n13914 ;
  assign n13919 = n13492 & n13556 ;
  assign n13920 = ~n13541 & ~n13919 ;
  assign n13921 = ~n13548 & n13920 ;
  assign n13922 = n13480 & ~n13921 ;
  assign n13916 = n13505 & n13533 ;
  assign n13917 = ~n13906 & ~n13916 ;
  assign n13918 = ~n13480 & ~n13917 ;
  assign n13923 = n13510 & n13515 ;
  assign n13924 = ~n13507 & ~n13923 ;
  assign n13925 = ~n13918 & n13924 ;
  assign n13926 = ~n13922 & n13925 ;
  assign n13927 = ~n13531 & ~n13926 ;
  assign n13931 = n13480 & n13510 ;
  assign n13932 = ~n13916 & ~n13931 ;
  assign n13933 = ~n13499 & ~n13932 ;
  assign n13928 = ~n13492 & n13535 ;
  assign n13929 = ~n13556 & ~n13928 ;
  assign n13930 = ~n13480 & ~n13929 ;
  assign n13934 = n13499 & n13519 ;
  assign n13935 = ~n13930 & ~n13934 ;
  assign n13936 = ~n13933 & n13935 ;
  assign n13937 = n13531 & ~n13936 ;
  assign n13938 = n13499 & n13899 ;
  assign n13939 = ~n13480 & ~n13534 ;
  assign n13940 = ~n13938 & n13939 ;
  assign n13941 = ~n13520 & ~n13539 ;
  assign n13942 = ~n13541 & n13941 ;
  assign n13943 = n13480 & n13499 ;
  assign n13944 = ~n13942 & n13943 ;
  assign n13945 = ~n13940 & ~n13944 ;
  assign n13946 = ~n13937 & n13945 ;
  assign n13947 = ~n13927 & n13946 ;
  assign n13948 = ~\u2_L8_reg[4]/NET0131  & ~n13947 ;
  assign n13949 = \u2_L8_reg[4]/NET0131  & n13947 ;
  assign n13950 = ~n13948 & ~n13949 ;
  assign n13995 = decrypt_pad & ~\u2_uk_K_r8_reg[29]/NET0131  ;
  assign n13996 = ~decrypt_pad & ~\u2_uk_K_r8_reg[9]/NET0131  ;
  assign n13997 = ~n13995 & ~n13996 ;
  assign n13998 = \u2_R8_reg[32]/NET0131  & ~n13997 ;
  assign n13999 = ~\u2_R8_reg[32]/NET0131  & n13997 ;
  assign n14000 = ~n13998 & ~n13999 ;
  assign n13971 = decrypt_pad & ~\u2_uk_K_r8_reg[23]/NET0131  ;
  assign n13972 = ~decrypt_pad & ~\u2_uk_K_r8_reg[31]/NET0131  ;
  assign n13973 = ~n13971 & ~n13972 ;
  assign n13974 = \u2_R8_reg[31]/P0001  & ~n13973 ;
  assign n13975 = ~\u2_R8_reg[31]/P0001  & n13973 ;
  assign n13976 = ~n13974 & ~n13975 ;
  assign n13979 = decrypt_pad & ~\u2_uk_K_r8_reg[50]/NET0131  ;
  assign n13980 = ~decrypt_pad & ~\u2_uk_K_r8_reg[30]/NET0131  ;
  assign n13981 = ~n13979 & ~n13980 ;
  assign n13982 = \u2_R8_reg[1]/NET0131  & ~n13981 ;
  assign n13983 = ~\u2_R8_reg[1]/NET0131  & n13981 ;
  assign n13984 = ~n13982 & ~n13983 ;
  assign n13951 = decrypt_pad & ~\u2_uk_K_r8_reg[35]/NET0131  ;
  assign n13952 = ~decrypt_pad & ~\u2_uk_K_r8_reg[15]/NET0131  ;
  assign n13953 = ~n13951 & ~n13952 ;
  assign n13954 = \u2_R8_reg[30]/NET0131  & ~n13953 ;
  assign n13955 = ~\u2_R8_reg[30]/NET0131  & n13953 ;
  assign n13956 = ~n13954 & ~n13955 ;
  assign n13957 = decrypt_pad & ~\u2_uk_K_r8_reg[7]/NET0131  ;
  assign n13958 = ~decrypt_pad & ~\u2_uk_K_r8_reg[42]/NET0131  ;
  assign n13959 = ~n13957 & ~n13958 ;
  assign n13960 = \u2_R8_reg[28]/NET0131  & ~n13959 ;
  assign n13961 = ~\u2_R8_reg[28]/NET0131  & n13959 ;
  assign n13962 = ~n13960 & ~n13961 ;
  assign n13964 = decrypt_pad & ~\u2_uk_K_r8_reg[38]/NET0131  ;
  assign n13965 = ~decrypt_pad & ~\u2_uk_K_r8_reg[14]/NET0131  ;
  assign n13966 = ~n13964 & ~n13965 ;
  assign n13967 = \u2_R8_reg[29]/NET0131  & ~n13966 ;
  assign n13968 = ~\u2_R8_reg[29]/NET0131  & n13966 ;
  assign n13969 = ~n13967 & ~n13968 ;
  assign n14002 = n13962 & ~n13969 ;
  assign n14003 = n13956 & n14002 ;
  assign n14004 = ~n13984 & n14003 ;
  assign n14005 = ~n13969 & n13984 ;
  assign n14006 = ~n13962 & n14005 ;
  assign n14007 = ~n14004 & ~n14006 ;
  assign n14008 = n13976 & ~n14007 ;
  assign n14013 = ~n13956 & ~n13984 ;
  assign n14014 = ~n13976 & ~n14013 ;
  assign n14012 = n13962 & ~n13984 ;
  assign n14015 = ~n14005 & ~n14012 ;
  assign n14016 = n14014 & n14015 ;
  assign n13991 = n13956 & n13969 ;
  assign n14010 = n13962 & n13984 ;
  assign n14011 = n13991 & n14010 ;
  assign n13978 = ~n13956 & n13962 ;
  assign n13985 = n13969 & ~n13984 ;
  assign n13987 = n13978 & n13985 ;
  assign n14009 = ~n13976 & n13978 ;
  assign n14017 = ~n13987 & ~n14009 ;
  assign n14018 = ~n14011 & n14017 ;
  assign n14019 = ~n14016 & n14018 ;
  assign n14020 = ~n14008 & n14019 ;
  assign n14021 = ~n14000 & ~n14020 ;
  assign n13963 = ~n13956 & ~n13962 ;
  assign n13970 = n13963 & ~n13969 ;
  assign n13977 = ~n13970 & ~n13976 ;
  assign n13986 = ~n13978 & ~n13985 ;
  assign n13988 = ~n13986 & ~n13987 ;
  assign n13989 = n13976 & ~n13988 ;
  assign n13990 = ~n13977 & ~n13989 ;
  assign n13992 = ~n13962 & n13991 ;
  assign n13993 = n13984 & n13992 ;
  assign n13994 = ~n13990 & ~n13993 ;
  assign n14001 = ~n13994 & n14000 ;
  assign n14025 = ~n13956 & n13969 ;
  assign n14026 = ~n14012 & ~n14025 ;
  assign n14027 = ~n13986 & n14026 ;
  assign n14022 = ~n13969 & ~n13984 ;
  assign n14023 = n13963 & n14022 ;
  assign n14024 = n13956 & n14006 ;
  assign n14028 = ~n14023 & ~n14024 ;
  assign n14029 = ~n14027 & n14028 ;
  assign n14030 = n13976 & ~n14029 ;
  assign n14031 = ~n13976 & n13987 ;
  assign n14032 = n13956 & ~n13976 ;
  assign n14033 = n14000 & n14002 ;
  assign n14034 = n14032 & n14033 ;
  assign n14035 = ~n14031 & ~n14034 ;
  assign n14036 = ~n14030 & n14035 ;
  assign n14037 = ~n14001 & n14036 ;
  assign n14038 = ~n14021 & n14037 ;
  assign n14039 = \u2_L8_reg[5]/NET0131  & ~n14038 ;
  assign n14040 = ~\u2_L8_reg[5]/NET0131  & n14038 ;
  assign n14041 = ~n14039 & ~n14040 ;
  assign n14058 = ~n13741 & ~n13742 ;
  assign n14059 = n13704 & ~n14058 ;
  assign n14043 = n13698 & ~n13724 ;
  assign n14055 = n13718 & ~n14043 ;
  assign n14056 = ~n13765 & ~n14055 ;
  assign n14057 = ~n13704 & ~n14056 ;
  assign n14060 = ~n13749 & n13770 ;
  assign n14061 = ~n14057 & ~n14060 ;
  assign n14062 = ~n14059 & n14061 ;
  assign n14063 = n13735 & ~n14062 ;
  assign n14044 = n13711 & n14043 ;
  assign n14042 = n13750 & n13774 ;
  assign n14049 = ~n13768 & ~n14042 ;
  assign n14050 = ~n14044 & n14049 ;
  assign n14045 = n13717 & ~n13724 ;
  assign n14046 = n13705 & n13711 ;
  assign n14047 = ~n14045 & n14046 ;
  assign n14048 = ~n13724 & n13772 ;
  assign n14051 = ~n14047 & ~n14048 ;
  assign n14052 = n14050 & n14051 ;
  assign n14053 = n13747 & n14052 ;
  assign n14054 = ~n13735 & ~n14053 ;
  assign n14064 = ~n13746 & ~n14060 ;
  assign n14065 = ~n13704 & ~n14064 ;
  assign n14066 = ~n13738 & ~n13782 ;
  assign n14067 = ~n14065 & n14066 ;
  assign n14068 = ~n14054 & n14067 ;
  assign n14069 = ~n14063 & n14068 ;
  assign n14070 = ~\u2_L8_reg[10]/NET0131  & ~n14069 ;
  assign n14071 = \u2_L8_reg[10]/NET0131  & n14069 ;
  assign n14072 = ~n14070 & ~n14071 ;
  assign n14074 = ~n13588 & ~n13644 ;
  assign n14075 = n13601 & ~n14074 ;
  assign n14073 = n13607 & n13613 ;
  assign n14076 = n13588 & n13628 ;
  assign n14085 = ~n14073 & ~n14076 ;
  assign n14086 = ~n14075 & n14085 ;
  assign n14082 = n13575 & ~n13624 ;
  assign n14083 = ~n13603 & ~n13624 ;
  assign n14084 = ~n14082 & ~n14083 ;
  assign n14077 = ~n13575 & ~n13581 ;
  assign n14078 = n13634 & ~n13644 ;
  assign n14079 = ~n14077 & n14078 ;
  assign n14080 = ~n13630 & ~n13643 ;
  assign n14081 = ~n13575 & ~n14080 ;
  assign n14087 = ~n14079 & ~n14081 ;
  assign n14088 = ~n14084 & n14087 ;
  assign n14089 = n14086 & n14088 ;
  assign n14094 = n13581 & n13594 ;
  assign n14095 = ~n13636 & ~n14094 ;
  assign n14096 = n13575 & ~n14095 ;
  assign n14098 = n13624 & ~n13629 ;
  assign n14099 = ~n13641 & n14098 ;
  assign n14091 = ~n13607 & ~n13634 ;
  assign n14090 = n13575 & ~n13594 ;
  assign n14092 = n13588 & ~n14090 ;
  assign n14093 = ~n14091 & n14092 ;
  assign n14097 = ~n13587 & n13631 ;
  assign n14100 = ~n14093 & ~n14097 ;
  assign n14101 = n14099 & n14100 ;
  assign n14102 = ~n14096 & n14101 ;
  assign n14103 = ~n14089 & ~n14102 ;
  assign n14104 = \u2_L8_reg[12]/NET0131  & n14103 ;
  assign n14105 = ~\u2_L8_reg[12]/NET0131  & ~n14103 ;
  assign n14106 = ~n14104 & ~n14105 ;
  assign n14107 = n13845 & n13857 ;
  assign n14108 = ~n13819 & ~n14107 ;
  assign n14109 = ~n13807 & n13845 ;
  assign n14110 = ~n13826 & ~n13837 ;
  assign n14111 = ~n13795 & ~n13836 ;
  assign n14112 = ~n14110 & n14111 ;
  assign n14113 = ~n14109 & ~n14112 ;
  assign n14114 = ~n13825 & ~n14113 ;
  assign n14115 = n14108 & ~n14114 ;
  assign n14116 = ~n13833 & ~n14115 ;
  assign n14118 = ~n13795 & ~n13835 ;
  assign n14119 = ~n13815 & ~n14118 ;
  assign n14117 = ~n13795 & n13808 ;
  assign n14120 = n13833 & ~n14117 ;
  assign n14121 = ~n14119 & n14120 ;
  assign n14123 = n13835 & n13854 ;
  assign n14122 = ~n13845 & n13861 ;
  assign n14124 = ~n13825 & ~n14122 ;
  assign n14125 = ~n14123 & n14124 ;
  assign n14126 = ~n14121 & n14125 ;
  assign n14127 = ~n13850 & n14118 ;
  assign n14128 = ~n13833 & ~n14127 ;
  assign n14130 = n13801 & n13826 ;
  assign n14129 = ~n13795 & n13850 ;
  assign n14131 = n13833 & ~n14129 ;
  assign n14132 = ~n14130 & n14131 ;
  assign n14133 = ~n14128 & ~n14132 ;
  assign n14134 = ~n13807 & n13850 ;
  assign n14135 = n13795 & n14134 ;
  assign n14136 = n13825 & ~n14135 ;
  assign n14137 = ~n13856 & n14136 ;
  assign n14138 = n14108 & n14137 ;
  assign n14139 = ~n14133 & n14138 ;
  assign n14140 = ~n14126 & ~n14139 ;
  assign n14141 = ~n14116 & ~n14140 ;
  assign n14142 = ~\u2_L8_reg[13]/NET0131  & n14141 ;
  assign n14143 = \u2_L8_reg[13]/NET0131  & ~n14141 ;
  assign n14144 = ~n14142 & ~n14143 ;
  assign n14205 = decrypt_pad & ~\u2_uk_K_r8_reg[14]/NET0131  ;
  assign n14206 = ~decrypt_pad & ~\u2_uk_K_r8_reg[49]/NET0131  ;
  assign n14207 = ~n14205 & ~n14206 ;
  assign n14208 = \u2_R8_reg[20]/NET0131  & ~n14207 ;
  assign n14209 = ~\u2_R8_reg[20]/NET0131  & n14207 ;
  assign n14210 = ~n14208 & ~n14209 ;
  assign n14170 = decrypt_pad & ~\u2_uk_K_r8_reg[30]/NET0131  ;
  assign n14171 = ~decrypt_pad & ~\u2_uk_K_r8_reg[38]/NET0131  ;
  assign n14172 = ~n14170 & ~n14171 ;
  assign n14173 = \u2_R8_reg[19]/NET0131  & ~n14172 ;
  assign n14174 = ~\u2_R8_reg[19]/NET0131  & n14172 ;
  assign n14175 = ~n14173 & ~n14174 ;
  assign n14145 = decrypt_pad & ~\u2_uk_K_r8_reg[31]/NET0131  ;
  assign n14146 = ~decrypt_pad & ~\u2_uk_K_r8_reg[7]/NET0131  ;
  assign n14147 = ~n14145 & ~n14146 ;
  assign n14148 = \u2_R8_reg[16]/NET0131  & ~n14147 ;
  assign n14149 = ~\u2_R8_reg[16]/NET0131  & n14147 ;
  assign n14150 = ~n14148 & ~n14149 ;
  assign n14158 = decrypt_pad & ~\u2_uk_K_r8_reg[49]/NET0131  ;
  assign n14159 = ~decrypt_pad & ~\u2_uk_K_r8_reg[29]/NET0131  ;
  assign n14160 = ~n14158 & ~n14159 ;
  assign n14161 = \u2_R8_reg[17]/NET0131  & ~n14160 ;
  assign n14162 = ~\u2_R8_reg[17]/NET0131  & n14160 ;
  assign n14163 = ~n14161 & ~n14162 ;
  assign n14151 = decrypt_pad & ~\u2_uk_K_r8_reg[15]/NET0131  ;
  assign n14152 = ~decrypt_pad & ~\u2_uk_K_r8_reg[50]/NET0131  ;
  assign n14153 = ~n14151 & ~n14152 ;
  assign n14154 = \u2_R8_reg[21]/NET0131  & ~n14153 ;
  assign n14155 = ~\u2_R8_reg[21]/NET0131  & n14153 ;
  assign n14156 = ~n14154 & ~n14155 ;
  assign n14178 = decrypt_pad & ~\u2_uk_K_r8_reg[43]/NET0131  ;
  assign n14179 = ~decrypt_pad & ~\u2_uk_K_r8_reg[23]/NET0131  ;
  assign n14180 = ~n14178 & ~n14179 ;
  assign n14181 = \u2_R8_reg[18]/NET0131  & ~n14180 ;
  assign n14182 = ~\u2_R8_reg[18]/NET0131  & n14180 ;
  assign n14183 = ~n14181 & ~n14182 ;
  assign n14212 = n14156 & ~n14183 ;
  assign n14213 = n14163 & n14212 ;
  assign n14214 = n14150 & n14213 ;
  assign n14157 = n14150 & ~n14156 ;
  assign n14186 = ~n14163 & ~n14183 ;
  assign n14216 = n14157 & n14186 ;
  assign n14193 = ~n14150 & n14156 ;
  assign n14194 = ~n14163 & n14193 ;
  assign n14187 = n14163 & n14183 ;
  assign n14215 = ~n14156 & n14187 ;
  assign n14217 = ~n14194 & ~n14215 ;
  assign n14218 = ~n14216 & n14217 ;
  assign n14219 = ~n14214 & n14218 ;
  assign n14220 = ~n14175 & ~n14219 ;
  assign n14167 = ~n14150 & n14163 ;
  assign n14221 = n14167 & ~n14183 ;
  assign n14222 = ~n14167 & ~n14212 ;
  assign n14223 = ~n14157 & ~n14193 ;
  assign n14224 = n14222 & n14223 ;
  assign n14225 = ~n14221 & ~n14224 ;
  assign n14226 = n14175 & ~n14225 ;
  assign n14227 = ~n14157 & ~n14212 ;
  assign n14165 = ~n14150 & ~n14163 ;
  assign n14228 = ~n14165 & ~n14187 ;
  assign n14229 = n14227 & n14228 ;
  assign n14230 = ~n14226 & ~n14229 ;
  assign n14231 = ~n14220 & n14230 ;
  assign n14232 = ~n14210 & ~n14231 ;
  assign n14164 = n14157 & n14163 ;
  assign n14166 = ~n14156 & n14165 ;
  assign n14168 = n14156 & n14167 ;
  assign n14169 = ~n14166 & ~n14168 ;
  assign n14176 = ~n14169 & ~n14175 ;
  assign n14177 = ~n14164 & ~n14176 ;
  assign n14184 = ~n14177 & ~n14183 ;
  assign n14198 = ~n14164 & ~n14194 ;
  assign n14185 = n14150 & n14156 ;
  assign n14195 = ~n14183 & n14185 ;
  assign n14196 = ~n14150 & n14183 ;
  assign n14197 = n14156 & n14196 ;
  assign n14199 = ~n14195 & ~n14197 ;
  assign n14200 = n14198 & n14199 ;
  assign n14201 = n14175 & ~n14200 ;
  assign n14188 = ~n14175 & n14187 ;
  assign n14189 = ~n14186 & ~n14188 ;
  assign n14190 = n14185 & ~n14189 ;
  assign n14191 = ~n14163 & n14183 ;
  assign n14192 = n14157 & n14191 ;
  assign n14202 = ~n14190 & ~n14192 ;
  assign n14203 = ~n14201 & n14202 ;
  assign n14204 = ~n14184 & n14203 ;
  assign n14211 = ~n14204 & n14210 ;
  assign n14233 = ~n14163 & n14197 ;
  assign n14234 = ~n14215 & ~n14233 ;
  assign n14235 = ~n14150 & ~n14234 ;
  assign n14236 = ~n14175 & n14235 ;
  assign n14237 = n14164 & ~n14183 ;
  assign n14238 = n14166 & n14183 ;
  assign n14239 = ~n14237 & ~n14238 ;
  assign n14240 = n14175 & ~n14239 ;
  assign n14241 = ~n14236 & ~n14240 ;
  assign n14242 = ~n14211 & n14241 ;
  assign n14243 = ~n14232 & n14242 ;
  assign n14244 = ~\u2_L8_reg[14]/NET0131  & ~n14243 ;
  assign n14245 = \u2_L8_reg[14]/NET0131  & n14243 ;
  assign n14246 = ~n14244 & ~n14245 ;
  assign n14247 = ~n13962 & ~n14013 ;
  assign n14248 = n13969 & ~n14247 ;
  assign n14249 = ~n14006 & ~n14248 ;
  assign n14250 = n13976 & ~n14249 ;
  assign n14251 = n14002 & n14013 ;
  assign n14252 = ~n14250 & ~n14251 ;
  assign n14253 = ~n14000 & ~n14252 ;
  assign n14256 = ~n13962 & n14022 ;
  assign n14257 = n13976 & n14256 ;
  assign n14254 = n13969 & n13978 ;
  assign n14255 = n14005 & n14032 ;
  assign n14260 = ~n14254 & ~n14255 ;
  assign n14261 = ~n14257 & n14260 ;
  assign n14258 = ~n13984 & n13992 ;
  assign n14259 = n13984 & n14003 ;
  assign n14262 = ~n14258 & ~n14259 ;
  assign n14263 = n14261 & n14262 ;
  assign n14264 = n14000 & ~n14263 ;
  assign n14268 = ~n13956 & n14000 ;
  assign n14269 = n14002 & ~n14268 ;
  assign n14270 = ~n13976 & ~n14023 ;
  assign n14271 = ~n14269 & n14270 ;
  assign n14265 = n13969 & n13984 ;
  assign n14266 = ~n13962 & n14265 ;
  assign n14267 = ~n13956 & n14266 ;
  assign n14272 = ~n14258 & ~n14267 ;
  assign n14273 = n14271 & n14272 ;
  assign n14274 = n13970 & n13984 ;
  assign n14275 = n13976 & ~n13993 ;
  assign n14276 = ~n14274 & n14275 ;
  assign n14277 = ~n14273 & ~n14276 ;
  assign n14278 = ~n14264 & ~n14277 ;
  assign n14279 = ~n14253 & n14278 ;
  assign n14280 = ~\u2_L8_reg[15]/NET0131  & ~n14279 ;
  assign n14281 = \u2_L8_reg[15]/NET0131  & n14279 ;
  assign n14282 = ~n14280 & ~n14281 ;
  assign n14283 = ~n13744 & ~n13754 ;
  assign n14284 = n13711 & ~n14283 ;
  assign n14285 = ~n13704 & ~n14284 ;
  assign n14286 = ~n13698 & n13725 ;
  assign n14287 = n13704 & ~n13727 ;
  assign n14288 = ~n14286 & n14287 ;
  assign n14289 = ~n14285 & ~n14288 ;
  assign n14290 = n13751 & n14043 ;
  assign n14291 = ~n13771 & ~n14290 ;
  assign n14292 = ~n14289 & n14291 ;
  assign n14293 = ~n13735 & ~n14292 ;
  assign n14303 = ~n13740 & ~n13754 ;
  assign n14304 = n13735 & ~n14303 ;
  assign n14305 = ~n13743 & ~n14060 ;
  assign n14306 = ~n14304 & n14305 ;
  assign n14307 = n13704 & ~n14306 ;
  assign n14294 = ~n13718 & n14043 ;
  assign n14295 = ~n13764 & ~n14294 ;
  assign n14296 = ~n13704 & ~n14295 ;
  assign n14297 = n13724 & n13745 ;
  assign n14298 = n13698 & n13725 ;
  assign n14299 = ~n14297 & ~n14298 ;
  assign n14300 = ~n14296 & n14299 ;
  assign n14301 = n13735 & ~n14300 ;
  assign n14302 = ~n13704 & n14298 ;
  assign n14308 = ~n13769 & ~n14302 ;
  assign n14309 = ~n14301 & n14308 ;
  assign n14310 = ~n14307 & n14309 ;
  assign n14311 = ~n14293 & n14310 ;
  assign n14312 = ~\u2_L8_reg[1]/NET0131  & ~n14311 ;
  assign n14313 = \u2_L8_reg[1]/NET0131  & n14311 ;
  assign n14314 = ~n14312 & ~n14313 ;
  assign n14315 = ~n13480 & n13486 ;
  assign n14316 = ~n13919 & ~n14315 ;
  assign n14317 = ~n13505 & ~n14316 ;
  assign n14321 = n13531 & ~n13928 ;
  assign n14322 = ~n14317 & n14321 ;
  assign n14318 = n13499 & ~n13941 ;
  assign n14319 = ~n13544 & ~n13551 ;
  assign n14320 = n13480 & ~n14319 ;
  assign n14323 = ~n14318 & ~n14320 ;
  assign n14324 = n14322 & n14323 ;
  assign n14327 = n13486 & ~n13535 ;
  assign n14328 = ~n13916 & ~n14327 ;
  assign n14329 = n13480 & ~n14328 ;
  assign n14326 = ~n13480 & ~n13941 ;
  assign n14325 = n13499 & n13511 ;
  assign n14330 = ~n13531 & ~n14325 ;
  assign n14331 = ~n14326 & n14330 ;
  assign n14332 = ~n14329 & n14331 ;
  assign n14333 = ~n14324 & ~n14332 ;
  assign n14334 = ~n13505 & n13923 ;
  assign n14335 = ~n13547 & ~n14334 ;
  assign n14336 = ~n14333 & n14335 ;
  assign n14337 = ~\u2_L8_reg[19]/NET0131  & ~n14336 ;
  assign n14338 = \u2_L8_reg[19]/NET0131  & n14336 ;
  assign n14339 = ~n14337 & ~n14338 ;
  assign n14345 = ~n13962 & ~n13976 ;
  assign n14346 = ~n14014 & ~n14345 ;
  assign n14347 = ~n14259 & ~n14346 ;
  assign n14350 = n13976 & ~n14266 ;
  assign n14348 = n13962 & n13991 ;
  assign n14349 = ~n13956 & n14005 ;
  assign n14351 = ~n14348 & ~n14349 ;
  assign n14352 = n14350 & n14351 ;
  assign n14353 = ~n14347 & ~n14352 ;
  assign n14342 = n13969 & n14012 ;
  assign n14343 = ~n14256 & ~n14342 ;
  assign n14344 = n13956 & ~n14343 ;
  assign n14354 = n14000 & ~n14274 ;
  assign n14355 = ~n14344 & n14354 ;
  assign n14356 = ~n14353 & n14355 ;
  assign n14365 = ~n14004 & ~n14023 ;
  assign n14361 = n13956 & n13984 ;
  assign n14362 = ~n13985 & ~n14361 ;
  assign n14363 = n14345 & ~n14362 ;
  assign n14364 = ~n13992 & ~n14000 ;
  assign n14366 = ~n14363 & n14364 ;
  assign n14367 = n14365 & n14366 ;
  assign n14357 = ~n14003 & ~n14342 ;
  assign n14358 = n13976 & ~n14357 ;
  assign n14359 = ~n14009 & ~n14254 ;
  assign n14360 = n13984 & ~n14359 ;
  assign n14368 = ~n14358 & ~n14360 ;
  assign n14369 = n14367 & n14368 ;
  assign n14370 = ~n14356 & ~n14369 ;
  assign n14340 = n13970 & n13976 ;
  assign n14341 = n14009 & n14265 ;
  assign n14371 = ~n14340 & ~n14341 ;
  assign n14372 = ~n14370 & n14371 ;
  assign n14373 = ~\u2_L8_reg[21]/NET0131  & ~n14372 ;
  assign n14374 = \u2_L8_reg[21]/NET0131  & n14372 ;
  assign n14375 = ~n14373 & ~n14374 ;
  assign n14387 = ~n13395 & ~n13402 ;
  assign n14388 = n13389 & ~n13465 ;
  assign n14389 = ~n14387 & n14388 ;
  assign n14390 = ~n13408 & ~n14389 ;
  assign n14391 = n13422 & n13442 ;
  assign n14376 = ~n13422 & n13435 ;
  assign n14392 = n13408 & ~n14376 ;
  assign n14393 = ~n14391 & n14392 ;
  assign n14394 = ~n14390 & ~n14393 ;
  assign n14395 = ~n13422 & n14387 ;
  assign n14396 = ~n13416 & ~n13663 ;
  assign n14397 = ~n14395 & n14396 ;
  assign n14398 = ~n14394 & n14397 ;
  assign n14399 = n13464 & n13662 ;
  assign n14400 = n13416 & ~n13665 ;
  assign n14401 = ~n14399 & n14400 ;
  assign n14402 = ~n13426 & ~n13467 ;
  assign n14403 = n14401 & n14402 ;
  assign n14404 = ~n14398 & ~n14403 ;
  assign n14377 = ~n13396 & ~n14376 ;
  assign n14378 = n13409 & ~n14377 ;
  assign n14380 = ~n13389 & n13673 ;
  assign n14381 = ~n13446 & ~n14380 ;
  assign n14382 = n13416 & ~n14381 ;
  assign n14379 = n13424 & ~n13433 ;
  assign n14383 = n13441 & n13444 ;
  assign n14384 = ~n14379 & ~n14383 ;
  assign n14385 = ~n14382 & n14384 ;
  assign n14386 = ~n13408 & ~n14385 ;
  assign n14405 = ~n14378 & ~n14386 ;
  assign n14406 = ~n14404 & n14405 ;
  assign n14407 = \u2_L8_reg[23]/NET0131  & ~n14406 ;
  assign n14408 = ~\u2_L8_reg[23]/NET0131  & n14406 ;
  assign n14409 = ~n14407 & ~n14408 ;
  assign n14430 = ~n14186 & ~n14196 ;
  assign n14431 = ~n14156 & ~n14430 ;
  assign n14429 = n14163 & n14185 ;
  assign n14432 = ~n14165 & ~n14429 ;
  assign n14433 = ~n14431 & n14432 ;
  assign n14434 = n14175 & ~n14433 ;
  assign n14410 = ~n14163 & n14185 ;
  assign n14435 = ~n14221 & ~n14410 ;
  assign n14436 = ~n14175 & ~n14435 ;
  assign n14422 = n14164 & n14183 ;
  assign n14437 = ~n14213 & ~n14422 ;
  assign n14438 = ~n14436 & n14437 ;
  assign n14439 = ~n14434 & n14438 ;
  assign n14440 = n14210 & ~n14439 ;
  assign n14411 = ~n14175 & ~n14410 ;
  assign n14416 = n14196 & n14411 ;
  assign n14414 = ~n14156 & ~n14183 ;
  assign n14415 = n14175 & n14414 ;
  assign n14417 = n14163 & ~n14197 ;
  assign n14418 = ~n14415 & n14417 ;
  assign n14419 = ~n14416 & n14418 ;
  assign n14412 = ~n14196 & n14411 ;
  assign n14413 = ~n14163 & ~n14412 ;
  assign n14420 = ~n14210 & ~n14413 ;
  assign n14421 = ~n14419 & n14420 ;
  assign n14423 = ~n14238 & ~n14422 ;
  assign n14424 = n14186 & n14193 ;
  assign n14425 = n14423 & ~n14424 ;
  assign n14426 = n14175 & ~n14425 ;
  assign n14427 = n14150 & ~n14175 ;
  assign n14428 = n14191 & n14427 ;
  assign n14441 = ~n14214 & ~n14428 ;
  assign n14442 = ~n14426 & n14441 ;
  assign n14443 = ~n14421 & n14442 ;
  assign n14444 = ~n14440 & n14443 ;
  assign n14445 = ~\u2_L8_reg[25]/NET0131  & ~n14444 ;
  assign n14446 = \u2_L8_reg[25]/NET0131  & n14444 ;
  assign n14447 = ~n14445 & ~n14446 ;
  assign n14459 = ~n13705 & ~n14043 ;
  assign n14460 = n13726 & ~n14459 ;
  assign n14467 = n13735 & ~n14298 ;
  assign n14468 = ~n14460 & n14467 ;
  assign n14461 = ~n13764 & ~n13772 ;
  assign n14462 = n13724 & ~n14461 ;
  assign n14463 = ~n13698 & n14045 ;
  assign n14464 = ~n13750 & ~n14463 ;
  assign n14465 = ~n13704 & ~n13739 ;
  assign n14466 = ~n14464 & n14465 ;
  assign n14469 = ~n14462 & ~n14466 ;
  assign n14470 = n14468 & n14469 ;
  assign n14471 = n13737 & ~n13763 ;
  assign n14472 = ~n13735 & ~n14471 ;
  assign n14473 = n13766 & n14472 ;
  assign n14474 = ~n14470 & ~n14473 ;
  assign n14448 = n13735 & ~n13767 ;
  assign n14449 = n13740 & ~n14448 ;
  assign n14450 = ~n13698 & ~n13717 ;
  assign n14451 = ~n14297 & ~n14450 ;
  assign n14452 = ~n13735 & ~n14451 ;
  assign n14453 = ~n13751 & n14043 ;
  assign n14454 = ~n13704 & ~n14453 ;
  assign n14455 = ~n14452 & n14454 ;
  assign n14456 = n13704 & ~n13741 ;
  assign n14457 = ~n13765 & n14456 ;
  assign n14458 = ~n14455 & ~n14457 ;
  assign n14475 = ~n14449 & ~n14458 ;
  assign n14476 = ~n14474 & n14475 ;
  assign n14477 = ~\u2_L8_reg[26]/NET0131  & ~n14476 ;
  assign n14478 = \u2_L8_reg[26]/NET0131  & n14476 ;
  assign n14479 = ~n14477 & ~n14478 ;
  assign n14481 = ~n13845 & ~n13846 ;
  assign n14482 = n14110 & ~n14481 ;
  assign n14483 = ~n13807 & ~n13845 ;
  assign n14484 = ~n14482 & ~n14483 ;
  assign n14485 = n13833 & ~n14484 ;
  assign n14487 = ~n13851 & ~n14134 ;
  assign n14486 = ~n13833 & ~n13869 ;
  assign n14488 = ~n14107 & n14486 ;
  assign n14489 = n14487 & n14488 ;
  assign n14490 = ~n14485 & ~n14489 ;
  assign n14480 = n13846 & ~n14110 ;
  assign n14491 = n13825 & ~n14480 ;
  assign n14492 = ~n14490 & n14491 ;
  assign n14493 = n13833 & n14487 ;
  assign n14494 = ~n13815 & ~n13817 ;
  assign n14495 = ~n13847 & n14494 ;
  assign n14496 = n14486 & n14495 ;
  assign n14497 = ~n14493 & ~n14496 ;
  assign n14498 = n13836 & n13868 ;
  assign n14499 = ~n13825 & ~n14107 ;
  assign n14500 = ~n14498 & n14499 ;
  assign n14501 = ~n14497 & n14500 ;
  assign n14502 = ~n14492 & ~n14501 ;
  assign n14503 = ~\u2_L8_reg[28]/NET0131  & n14502 ;
  assign n14504 = \u2_L8_reg[28]/NET0131  & ~n14502 ;
  assign n14505 = ~n14503 & ~n14504 ;
  assign n14517 = n14175 & ~n14216 ;
  assign n14518 = ~n14429 & n14517 ;
  assign n14519 = ~n14191 & n14193 ;
  assign n14520 = n14411 & ~n14519 ;
  assign n14521 = ~n14518 & ~n14520 ;
  assign n14522 = ~n14221 & n14423 ;
  assign n14523 = ~n14521 & n14522 ;
  assign n14524 = ~n14210 & ~n14523 ;
  assign n14507 = n14165 & n14414 ;
  assign n14508 = ~n14410 & ~n14507 ;
  assign n14509 = n14175 & ~n14508 ;
  assign n14510 = ~n14183 & n14427 ;
  assign n14511 = ~n14509 & ~n14510 ;
  assign n14512 = ~n14235 & n14511 ;
  assign n14513 = n14210 & ~n14512 ;
  assign n14506 = ~n14156 & n14428 ;
  assign n14514 = n14167 & n14212 ;
  assign n14515 = n14234 & ~n14514 ;
  assign n14516 = n14175 & ~n14515 ;
  assign n14525 = ~n14506 & ~n14516 ;
  assign n14526 = ~n14513 & n14525 ;
  assign n14527 = ~n14524 & n14526 ;
  assign n14528 = ~\u2_L8_reg[8]/NET0131  & ~n14527 ;
  assign n14529 = \u2_L8_reg[8]/NET0131  & n14527 ;
  assign n14530 = ~n14528 & ~n14529 ;
  assign n14544 = ~n14012 & n14248 ;
  assign n14545 = n13976 & ~n14544 ;
  assign n14546 = ~n14266 & ~n14342 ;
  assign n14547 = n13977 & n14546 ;
  assign n14548 = ~n14545 & ~n14547 ;
  assign n14549 = ~n13993 & ~n14349 ;
  assign n14550 = ~n14004 & n14549 ;
  assign n14551 = ~n14548 & n14550 ;
  assign n14552 = n14000 & ~n14551 ;
  assign n14531 = n14022 & ~n14268 ;
  assign n14532 = ~n14005 & ~n14013 ;
  assign n14533 = ~n14361 & n14532 ;
  assign n14534 = n14364 & n14533 ;
  assign n14535 = ~n14531 & ~n14534 ;
  assign n14536 = n13976 & ~n14535 ;
  assign n14537 = n13985 & n14345 ;
  assign n14538 = n14010 & n14032 ;
  assign n14539 = ~n14537 & ~n14538 ;
  assign n14540 = ~n14024 & n14539 ;
  assign n14541 = ~n14000 & ~n14540 ;
  assign n14542 = ~n13987 & ~n14027 ;
  assign n14543 = ~n13976 & ~n14542 ;
  assign n14553 = ~n14541 & ~n14543 ;
  assign n14554 = ~n14536 & n14553 ;
  assign n14555 = ~n14552 & n14554 ;
  assign n14556 = ~\u2_L8_reg[27]/NET0131  & ~n14555 ;
  assign n14557 = \u2_L8_reg[27]/NET0131  & n14555 ;
  assign n14558 = ~n14556 & ~n14557 ;
  assign n14576 = ~n13613 & n14080 ;
  assign n14577 = n14091 & ~n14576 ;
  assign n14578 = ~n13613 & ~n14091 ;
  assign n14579 = ~n13575 & ~n14578 ;
  assign n14580 = ~n14577 & n14579 ;
  assign n14571 = n13587 & n13607 ;
  assign n14572 = ~n14077 & n14571 ;
  assign n14573 = ~n13594 & n13643 ;
  assign n14574 = ~n13645 & ~n14573 ;
  assign n14575 = n13575 & ~n14574 ;
  assign n14581 = ~n14572 & ~n14575 ;
  assign n14582 = ~n14580 & n14581 ;
  assign n14583 = n13624 & ~n14582 ;
  assign n14559 = ~n13587 & n13607 ;
  assign n14560 = n13581 & n14559 ;
  assign n14561 = n13603 & n13630 ;
  assign n14566 = ~n14560 & ~n14561 ;
  assign n14567 = n13642 & n14566 ;
  assign n14562 = ~n13581 & n13628 ;
  assign n14563 = ~n14559 & ~n14562 ;
  assign n14564 = n13575 & ~n14563 ;
  assign n14565 = n14081 & ~n14559 ;
  assign n14568 = ~n14564 & ~n14565 ;
  assign n14569 = n14567 & n14568 ;
  assign n14570 = ~n13624 & ~n14569 ;
  assign n14584 = n13575 & n13635 ;
  assign n14585 = ~n13607 & n13626 ;
  assign n14586 = n13605 & n14585 ;
  assign n14587 = ~n14584 & ~n14586 ;
  assign n14588 = ~n14570 & n14587 ;
  assign n14589 = ~n14583 & n14588 ;
  assign n14590 = \u2_L8_reg[32]/NET0131  & n14589 ;
  assign n14591 = ~\u2_L8_reg[32]/NET0131  & ~n14589 ;
  assign n14592 = ~n14590 & ~n14591 ;
  assign n14593 = ~n14157 & n14191 ;
  assign n14594 = ~n14210 & ~n14593 ;
  assign n14595 = ~n14227 & ~n14410 ;
  assign n14596 = n14594 & n14595 ;
  assign n14597 = ~n14192 & n14210 ;
  assign n14598 = ~n14168 & ~n14214 ;
  assign n14599 = n14597 & n14598 ;
  assign n14600 = ~n14596 & ~n14599 ;
  assign n14601 = n14183 & n14410 ;
  assign n14602 = ~n14175 & ~n14507 ;
  assign n14603 = ~n14237 & n14602 ;
  assign n14604 = ~n14601 & n14603 ;
  assign n14605 = ~n14600 & n14604 ;
  assign n14606 = ~n14193 & ~n14222 ;
  assign n14607 = n14597 & ~n14606 ;
  assign n14608 = ~n14183 & n14193 ;
  assign n14609 = ~n14164 & ~n14608 ;
  assign n14610 = n14594 & n14609 ;
  assign n14611 = ~n14607 & ~n14610 ;
  assign n14612 = ~n14233 & n14517 ;
  assign n14613 = ~n14611 & n14612 ;
  assign n14614 = ~n14605 & ~n14613 ;
  assign n14615 = ~\u2_L8_reg[3]/NET0131  & n14614 ;
  assign n14616 = \u2_L8_reg[3]/NET0131  & ~n14614 ;
  assign n14617 = ~n14615 & ~n14616 ;
  assign n14618 = decrypt_pad & ~\u2_uk_K_r8_reg[25]/NET0131  ;
  assign n14619 = ~decrypt_pad & ~\u2_uk_K_r8_reg[3]/NET0131  ;
  assign n14620 = ~n14618 & ~n14619 ;
  assign n14621 = \u2_R8_reg[13]/NET0131  & ~n14620 ;
  assign n14622 = ~\u2_R8_reg[13]/NET0131  & n14620 ;
  assign n14623 = ~n14621 & ~n14622 ;
  assign n14631 = decrypt_pad & ~\u2_uk_K_r8_reg[20]/NET0131  ;
  assign n14632 = ~decrypt_pad & ~\u2_uk_K_r8_reg[55]/NET0131  ;
  assign n14633 = ~n14631 & ~n14632 ;
  assign n14634 = \u2_R8_reg[9]/NET0131  & ~n14633 ;
  assign n14635 = ~\u2_R8_reg[9]/NET0131  & n14633 ;
  assign n14636 = ~n14634 & ~n14635 ;
  assign n14645 = ~n14623 & n14636 ;
  assign n14646 = decrypt_pad & ~\u2_uk_K_r8_reg[54]/NET0131  ;
  assign n14647 = ~decrypt_pad & ~\u2_uk_K_r8_reg[32]/NET0131  ;
  assign n14648 = ~n14646 & ~n14647 ;
  assign n14649 = \u2_R8_reg[11]/NET0131  & ~n14648 ;
  assign n14650 = ~\u2_R8_reg[11]/NET0131  & n14648 ;
  assign n14651 = ~n14649 & ~n14650 ;
  assign n14652 = ~n14645 & ~n14651 ;
  assign n14637 = decrypt_pad & ~\u2_uk_K_r8_reg[53]/NET0131  ;
  assign n14638 = ~decrypt_pad & ~\u2_uk_K_r8_reg[6]/NET0131  ;
  assign n14639 = ~n14637 & ~n14638 ;
  assign n14640 = \u2_R8_reg[10]/NET0131  & ~n14639 ;
  assign n14641 = ~\u2_R8_reg[10]/NET0131  & n14639 ;
  assign n14642 = ~n14640 & ~n14641 ;
  assign n14653 = n14636 & ~n14642 ;
  assign n14624 = decrypt_pad & ~\u2_uk_K_r8_reg[48]/NET0131  ;
  assign n14625 = ~decrypt_pad & ~\u2_uk_K_r8_reg[26]/NET0131  ;
  assign n14626 = ~n14624 & ~n14625 ;
  assign n14627 = \u2_R8_reg[8]/NET0131  & ~n14626 ;
  assign n14628 = ~\u2_R8_reg[8]/NET0131  & n14626 ;
  assign n14629 = ~n14627 & ~n14628 ;
  assign n14654 = n14623 & ~n14636 ;
  assign n14655 = n14629 & ~n14654 ;
  assign n14656 = ~n14653 & ~n14655 ;
  assign n14657 = n14652 & ~n14656 ;
  assign n14630 = ~n14623 & ~n14629 ;
  assign n14643 = n14636 & n14642 ;
  assign n14644 = n14630 & n14643 ;
  assign n14658 = decrypt_pad & ~\u2_uk_K_r8_reg[12]/NET0131  ;
  assign n14659 = ~decrypt_pad & ~\u2_uk_K_r8_reg[47]/NET0131  ;
  assign n14660 = ~n14658 & ~n14659 ;
  assign n14661 = \u2_R8_reg[12]/NET0131  & ~n14660 ;
  assign n14662 = ~\u2_R8_reg[12]/NET0131  & n14660 ;
  assign n14663 = ~n14661 & ~n14662 ;
  assign n14664 = ~n14644 & n14663 ;
  assign n14665 = ~n14657 & n14664 ;
  assign n14670 = n14623 & n14629 ;
  assign n14671 = ~n14630 & ~n14670 ;
  assign n14672 = ~n14636 & ~n14642 ;
  assign n14675 = ~n14671 & ~n14672 ;
  assign n14676 = ~n14643 & n14675 ;
  assign n14678 = n14629 & n14642 ;
  assign n14679 = n14645 & n14678 ;
  assign n14669 = ~n14629 & n14651 ;
  assign n14677 = n14653 & n14669 ;
  assign n14680 = ~n14663 & ~n14677 ;
  assign n14681 = ~n14679 & n14680 ;
  assign n14666 = n14623 & ~n14629 ;
  assign n14667 = n14643 & n14666 ;
  assign n14668 = ~n14651 & n14667 ;
  assign n14673 = ~n14669 & n14672 ;
  assign n14674 = n14671 & n14673 ;
  assign n14682 = ~n14668 & ~n14674 ;
  assign n14683 = n14681 & n14682 ;
  assign n14684 = ~n14676 & n14683 ;
  assign n14685 = ~n14665 & ~n14684 ;
  assign n14687 = ~n14629 & ~n14642 ;
  assign n14688 = n14629 & ~n14636 ;
  assign n14689 = ~n14687 & ~n14688 ;
  assign n14690 = n14671 & n14689 ;
  assign n14691 = ~n14654 & ~n14690 ;
  assign n14692 = n14663 & ~n14691 ;
  assign n14686 = n14642 & n14654 ;
  assign n14693 = n14630 & ~n14642 ;
  assign n14694 = ~n14636 & n14693 ;
  assign n14695 = ~n14686 & ~n14694 ;
  assign n14696 = ~n14692 & n14695 ;
  assign n14697 = n14651 & ~n14696 ;
  assign n14698 = ~n14685 & ~n14697 ;
  assign n14699 = ~\u2_L8_reg[6]/NET0131  & ~n14698 ;
  assign n14700 = \u2_L8_reg[6]/NET0131  & n14698 ;
  assign n14701 = ~n14699 & ~n14700 ;
  assign n14704 = n13587 & n14091 ;
  assign n14702 = n13581 & n13587 ;
  assign n14703 = ~n14091 & ~n14702 ;
  assign n14705 = ~n13650 & ~n14703 ;
  assign n14706 = ~n14704 & n14705 ;
  assign n14707 = ~n13575 & n13624 ;
  assign n14708 = ~n14082 & ~n14707 ;
  assign n14709 = ~n13602 & n14708 ;
  assign n14710 = ~n14706 & n14709 ;
  assign n14712 = ~n13594 & n14074 ;
  assign n14711 = n13581 & ~n14091 ;
  assign n14713 = ~n14571 & n14707 ;
  assign n14714 = ~n14711 & n14713 ;
  assign n14715 = ~n14712 & n14714 ;
  assign n14716 = ~n14710 & ~n14715 ;
  assign n14717 = ~n14076 & ~n14716 ;
  assign n14718 = ~n13640 & n14082 ;
  assign n14719 = ~n14561 & n14718 ;
  assign n14720 = ~n14703 & n14719 ;
  assign n14721 = ~n14717 & ~n14720 ;
  assign n14722 = ~\u2_L8_reg[7]/NET0131  & n14721 ;
  assign n14723 = \u2_L8_reg[7]/NET0131  & ~n14721 ;
  assign n14724 = ~n14722 & ~n14723 ;
  assign n14725 = ~n13429 & ~n14391 ;
  assign n14726 = n13427 & ~n14725 ;
  assign n14729 = ~n13424 & ~n13673 ;
  assign n14730 = n13389 & n13431 ;
  assign n14731 = n13408 & ~n14730 ;
  assign n14732 = ~n14729 & ~n14731 ;
  assign n14733 = n13408 & ~n13673 ;
  assign n14734 = ~n14732 & ~n14733 ;
  assign n14727 = ~n13429 & ~n13681 ;
  assign n14728 = ~n14387 & ~n14727 ;
  assign n14735 = ~n13416 & ~n14728 ;
  assign n14736 = ~n14734 & n14735 ;
  assign n14738 = ~n13674 & ~n14380 ;
  assign n14739 = n13402 & ~n14738 ;
  assign n14737 = n13409 & n14729 ;
  assign n14740 = n13661 & ~n14737 ;
  assign n14741 = ~n14739 & n14740 ;
  assign n14742 = ~n14736 & ~n14741 ;
  assign n14743 = ~n14726 & ~n14742 ;
  assign n14744 = ~\u2_L8_reg[9]/NET0131  & ~n14743 ;
  assign n14745 = \u2_L8_reg[9]/NET0131  & n14743 ;
  assign n14746 = ~n14744 & ~n14745 ;
  assign n14749 = n14636 & ~n14670 ;
  assign n14750 = ~n14636 & n14670 ;
  assign n14751 = ~n14749 & ~n14750 ;
  assign n14752 = ~n14630 & n14751 ;
  assign n14753 = n14645 & n14669 ;
  assign n14754 = ~n14752 & ~n14753 ;
  assign n14755 = ~n14642 & ~n14754 ;
  assign n14756 = ~n14651 & ~n14678 ;
  assign n14757 = ~n14623 & ~n14687 ;
  assign n14758 = n14756 & n14757 ;
  assign n14759 = ~n14667 & ~n14758 ;
  assign n14760 = ~n14755 & n14759 ;
  assign n14761 = n14663 & ~n14760 ;
  assign n14762 = ~n14630 & n14651 ;
  assign n14763 = ~n14751 & n14762 ;
  assign n14764 = n14651 & ~n14694 ;
  assign n14765 = ~n14636 & ~n14666 ;
  assign n14766 = ~n14749 & ~n14765 ;
  assign n14767 = ~n14693 & ~n14766 ;
  assign n14768 = ~n14764 & ~n14767 ;
  assign n14769 = ~n14763 & ~n14768 ;
  assign n14770 = ~n14663 & ~n14769 ;
  assign n14747 = ~n14651 & n14678 ;
  assign n14748 = ~n14636 & n14747 ;
  assign n14771 = n14630 & n14642 ;
  assign n14772 = ~n14636 & n14771 ;
  assign n14773 = ~n14679 & ~n14772 ;
  assign n14774 = n14651 & ~n14773 ;
  assign n14775 = ~n14748 & ~n14774 ;
  assign n14776 = ~n14770 & n14775 ;
  assign n14777 = ~n14761 & n14776 ;
  assign n14778 = ~\u2_L8_reg[16]/NET0131  & ~n14777 ;
  assign n14779 = \u2_L8_reg[16]/NET0131  & n14777 ;
  assign n14780 = ~n14778 & ~n14779 ;
  assign n14798 = n13833 & ~n13848 ;
  assign n14795 = n13801 & n13837 ;
  assign n14796 = ~n14117 & ~n14795 ;
  assign n14797 = ~n13833 & ~n14796 ;
  assign n14799 = ~n13870 & ~n14797 ;
  assign n14800 = ~n14798 & n14799 ;
  assign n14801 = n13825 & ~n14800 ;
  assign n14784 = n13795 & ~n13873 ;
  assign n14785 = ~n13807 & ~n13868 ;
  assign n14786 = ~n14784 & n14785 ;
  assign n14783 = n13857 & ~n14481 ;
  assign n14781 = n13801 & n13833 ;
  assign n14782 = n13817 & n14781 ;
  assign n14787 = ~n14129 & ~n14782 ;
  assign n14788 = ~n14783 & n14787 ;
  assign n14789 = ~n14786 & n14788 ;
  assign n14790 = ~n13825 & ~n14789 ;
  assign n14791 = ~n13833 & n13851 ;
  assign n14792 = ~n13808 & n13833 ;
  assign n14793 = n14110 & n14792 ;
  assign n14794 = ~n14483 & n14793 ;
  assign n14802 = ~n14791 & ~n14794 ;
  assign n14803 = ~n14790 & n14802 ;
  assign n14804 = ~n14801 & n14803 ;
  assign n14805 = ~\u2_L8_reg[18]/P0001  & ~n14804 ;
  assign n14806 = \u2_L8_reg[18]/P0001  & n14804 ;
  assign n14807 = ~n14805 & ~n14806 ;
  assign n14815 = ~n14642 & n14666 ;
  assign n14816 = ~n14771 & ~n14815 ;
  assign n14817 = n14642 & n14688 ;
  assign n14814 = n14630 & n14636 ;
  assign n14818 = n14651 & ~n14814 ;
  assign n14819 = ~n14817 & n14818 ;
  assign n14820 = n14816 & n14819 ;
  assign n14823 = ~n14671 & n14672 ;
  assign n14821 = ~n14642 & ~n14645 ;
  assign n14822 = n14671 & ~n14821 ;
  assign n14824 = ~n14651 & ~n14822 ;
  assign n14825 = ~n14823 & n14824 ;
  assign n14826 = ~n14820 & ~n14825 ;
  assign n14827 = ~n14663 & ~n14826 ;
  assign n14828 = ~n14651 & n14675 ;
  assign n14832 = n14663 & ~n14674 ;
  assign n14829 = n14642 & ~n14688 ;
  assign n14830 = n14762 & n14829 ;
  assign n14810 = ~n14642 & n14651 ;
  assign n14831 = n14765 & n14810 ;
  assign n14833 = ~n14830 & ~n14831 ;
  assign n14834 = n14832 & n14833 ;
  assign n14835 = ~n14828 & n14834 ;
  assign n14836 = ~n14827 & ~n14835 ;
  assign n14808 = n14623 & n14636 ;
  assign n14809 = ~n14688 & ~n14808 ;
  assign n14811 = ~n14670 & n14810 ;
  assign n14812 = ~n14809 & n14811 ;
  assign n14813 = n14747 & n14808 ;
  assign n14837 = ~n14812 & ~n14813 ;
  assign n14838 = ~n14836 & n14837 ;
  assign n14839 = ~\u2_L8_reg[24]/NET0131  & ~n14838 ;
  assign n14840 = \u2_L8_reg[24]/NET0131  & n14838 ;
  assign n14841 = ~n14839 & ~n14840 ;
  assign n14858 = ~n14645 & n14678 ;
  assign n14853 = ~n14623 & ~n14642 ;
  assign n14857 = n14636 & n14853 ;
  assign n14859 = ~n14663 & ~n14857 ;
  assign n14860 = ~n14858 & n14859 ;
  assign n14854 = n14688 & n14853 ;
  assign n14855 = n14663 & ~n14854 ;
  assign n14856 = n14816 & n14855 ;
  assign n14861 = n14651 & ~n14856 ;
  assign n14862 = ~n14860 & n14861 ;
  assign n14843 = ~n14678 & ~n14814 ;
  assign n14844 = ~n14651 & ~n14843 ;
  assign n14842 = n14642 & n14749 ;
  assign n14845 = n14663 & ~n14842 ;
  assign n14846 = ~n14844 & n14845 ;
  assign n14849 = ~n14663 & ~n14823 ;
  assign n14847 = ~n14629 & n14686 ;
  assign n14848 = n14756 & ~n14809 ;
  assign n14850 = ~n14847 & ~n14848 ;
  assign n14851 = n14849 & n14850 ;
  assign n14852 = ~n14846 & ~n14851 ;
  assign n14863 = n14651 & ~n14750 ;
  assign n14864 = n14642 & ~n14652 ;
  assign n14865 = ~n14863 & n14864 ;
  assign n14866 = ~n14852 & ~n14865 ;
  assign n14867 = ~n14862 & n14866 ;
  assign n14868 = \u2_L8_reg[30]/NET0131  & ~n14867 ;
  assign n14869 = ~\u2_L8_reg[30]/NET0131  & n14867 ;
  assign n14870 = ~n14868 & ~n14869 ;
  assign n14871 = decrypt_pad & ~\u2_uk_K_r7_reg[31]/NET0131  ;
  assign n14872 = ~decrypt_pad & ~\u2_uk_K_r7_reg[38]/NET0131  ;
  assign n14873 = ~n14871 & ~n14872 ;
  assign n14874 = \u2_R7_reg[26]/NET0131  & ~n14873 ;
  assign n14875 = ~\u2_R7_reg[26]/NET0131  & n14873 ;
  assign n14876 = ~n14874 & ~n14875 ;
  assign n14877 = decrypt_pad & ~\u2_uk_K_r7_reg[42]/NET0131  ;
  assign n14878 = ~decrypt_pad & ~\u2_uk_K_r7_reg[49]/NET0131  ;
  assign n14879 = ~n14877 & ~n14878 ;
  assign n14880 = \u2_R7_reg[25]/NET0131  & ~n14879 ;
  assign n14881 = ~\u2_R7_reg[25]/NET0131  & n14879 ;
  assign n14882 = ~n14880 & ~n14881 ;
  assign n14883 = n14876 & ~n14882 ;
  assign n14884 = decrypt_pad & ~\u2_uk_K_r7_reg[7]/NET0131  ;
  assign n14885 = ~decrypt_pad & ~\u2_uk_K_r7_reg[14]/NET0131  ;
  assign n14886 = ~n14884 & ~n14885 ;
  assign n14887 = \u2_R7_reg[24]/NET0131  & ~n14886 ;
  assign n14888 = ~\u2_R7_reg[24]/NET0131  & n14886 ;
  assign n14889 = ~n14887 & ~n14888 ;
  assign n14890 = decrypt_pad & ~\u2_uk_K_r7_reg[15]/NET0131  ;
  assign n14891 = ~decrypt_pad & ~\u2_uk_K_r7_reg[22]/NET0131  ;
  assign n14892 = ~n14890 & ~n14891 ;
  assign n14893 = \u2_R7_reg[29]/NET0131  & ~n14892 ;
  assign n14894 = ~\u2_R7_reg[29]/NET0131  & n14892 ;
  assign n14895 = ~n14893 & ~n14894 ;
  assign n14896 = ~n14889 & n14895 ;
  assign n14897 = n14883 & n14896 ;
  assign n14898 = ~n14889 & ~n14895 ;
  assign n14899 = n14876 & n14898 ;
  assign n14900 = n14882 & n14899 ;
  assign n14901 = ~n14897 & ~n14900 ;
  assign n14902 = ~n14882 & ~n14895 ;
  assign n14903 = n14882 & n14895 ;
  assign n14904 = ~n14876 & n14903 ;
  assign n14905 = ~n14883 & ~n14904 ;
  assign n14906 = decrypt_pad & ~\u2_uk_K_r7_reg[23]/P0001  ;
  assign n14907 = ~decrypt_pad & ~\u2_uk_K_r7_reg[30]/P0001  ;
  assign n14908 = ~n14906 & ~n14907 ;
  assign n14909 = \u2_R7_reg[28]/NET0131  & ~n14908 ;
  assign n14910 = ~\u2_R7_reg[28]/NET0131  & n14908 ;
  assign n14911 = ~n14909 & ~n14910 ;
  assign n14912 = ~n14905 & n14911 ;
  assign n14913 = ~n14902 & ~n14912 ;
  assign n14914 = n14889 & ~n14913 ;
  assign n14915 = n14901 & ~n14914 ;
  assign n14916 = decrypt_pad & ~\u2_uk_K_r7_reg[36]/NET0131  ;
  assign n14917 = ~decrypt_pad & ~\u2_uk_K_r7_reg[43]/NET0131  ;
  assign n14918 = ~n14916 & ~n14917 ;
  assign n14919 = \u2_R7_reg[27]/NET0131  & ~n14918 ;
  assign n14920 = ~\u2_R7_reg[27]/NET0131  & n14918 ;
  assign n14921 = ~n14919 & ~n14920 ;
  assign n14922 = ~n14915 & n14921 ;
  assign n14923 = ~n14882 & n14921 ;
  assign n14924 = ~n14876 & n14923 ;
  assign n14925 = ~n14895 & ~n14921 ;
  assign n14926 = ~n14883 & n14925 ;
  assign n14927 = ~n14924 & ~n14926 ;
  assign n14928 = n14889 & ~n14927 ;
  assign n14929 = ~n14876 & ~n14889 ;
  assign n14930 = n14876 & n14889 ;
  assign n14931 = ~n14929 & ~n14930 ;
  assign n14932 = n14895 & ~n14931 ;
  assign n14933 = ~n14882 & n14899 ;
  assign n14934 = ~n14932 & ~n14933 ;
  assign n14935 = ~n14923 & ~n14934 ;
  assign n14936 = ~n14928 & ~n14935 ;
  assign n14937 = ~n14911 & ~n14936 ;
  assign n14941 = n14889 & n14895 ;
  assign n14942 = ~n14876 & ~n14882 ;
  assign n14943 = n14941 & n14942 ;
  assign n14944 = ~n14889 & n14903 ;
  assign n14945 = ~n14943 & ~n14944 ;
  assign n14946 = ~n14921 & ~n14945 ;
  assign n14947 = n14898 & n14942 ;
  assign n14948 = ~n14897 & ~n14947 ;
  assign n14949 = ~n14946 & n14948 ;
  assign n14950 = n14911 & ~n14949 ;
  assign n14938 = ~n14895 & n14924 ;
  assign n14939 = n14882 & ~n14921 ;
  assign n14940 = ~n14931 & n14939 ;
  assign n14951 = ~n14938 & ~n14940 ;
  assign n14952 = ~n14950 & n14951 ;
  assign n14953 = ~n14937 & n14952 ;
  assign n14954 = ~n14922 & n14953 ;
  assign n14955 = ~\u2_L7_reg[22]/NET0131  & ~n14954 ;
  assign n14956 = \u2_L7_reg[22]/NET0131  & n14954 ;
  assign n14957 = ~n14955 & ~n14956 ;
  assign n14985 = decrypt_pad & ~\u2_uk_K_r7_reg[47]/NET0131  ;
  assign n14986 = ~decrypt_pad & ~\u2_uk_K_r7_reg[54]/NET0131  ;
  assign n14987 = ~n14985 & ~n14986 ;
  assign n14988 = \u2_R7_reg[4]/NET0131  & ~n14987 ;
  assign n14989 = ~\u2_R7_reg[4]/NET0131  & n14987 ;
  assign n14990 = ~n14988 & ~n14989 ;
  assign n14971 = decrypt_pad & ~\u2_uk_K_r7_reg[12]/NET0131  ;
  assign n14972 = ~decrypt_pad & ~\u2_uk_K_r7_reg[19]/NET0131  ;
  assign n14973 = ~n14971 & ~n14972 ;
  assign n14974 = \u2_R7_reg[3]/NET0131  & ~n14973 ;
  assign n14975 = ~\u2_R7_reg[3]/NET0131  & n14973 ;
  assign n14976 = ~n14974 & ~n14975 ;
  assign n14964 = decrypt_pad & ~\u2_uk_K_r7_reg[20]/NET0131  ;
  assign n14965 = ~decrypt_pad & ~\u2_uk_K_r7_reg[27]/NET0131  ;
  assign n14966 = ~n14964 & ~n14965 ;
  assign n14967 = \u2_R7_reg[1]/NET0131  & ~n14966 ;
  assign n14968 = ~\u2_R7_reg[1]/NET0131  & n14966 ;
  assign n14969 = ~n14967 & ~n14968 ;
  assign n14992 = decrypt_pad & ~\u2_uk_K_r7_reg[18]/NET0131  ;
  assign n14993 = ~decrypt_pad & ~\u2_uk_K_r7_reg[25]/NET0131  ;
  assign n14994 = ~n14992 & ~n14993 ;
  assign n14995 = \u2_R7_reg[5]/NET0131  & ~n14994 ;
  assign n14996 = ~\u2_R7_reg[5]/NET0131  & n14994 ;
  assign n14997 = ~n14995 & ~n14996 ;
  assign n15006 = ~n14969 & n14997 ;
  assign n14977 = decrypt_pad & ~\u2_uk_K_r7_reg[3]/NET0131  ;
  assign n14978 = ~decrypt_pad & ~\u2_uk_K_r7_reg[10]/NET0131  ;
  assign n14979 = ~n14977 & ~n14978 ;
  assign n14980 = \u2_R7_reg[2]/NET0131  & ~n14979 ;
  assign n14981 = ~\u2_R7_reg[2]/NET0131  & n14979 ;
  assign n14982 = ~n14980 & ~n14981 ;
  assign n14958 = decrypt_pad & ~\u2_uk_K_r7_reg[24]/NET0131  ;
  assign n14959 = ~decrypt_pad & ~\u2_uk_K_r7_reg[6]/NET0131  ;
  assign n14960 = ~n14958 & ~n14959 ;
  assign n14961 = \u2_R7_reg[32]/NET0131  & ~n14960 ;
  assign n14962 = ~\u2_R7_reg[32]/NET0131  & n14960 ;
  assign n14963 = ~n14961 & ~n14962 ;
  assign n14999 = ~n14963 & ~n14997 ;
  assign n15019 = n14982 & n14999 ;
  assign n15020 = ~n14963 & n14997 ;
  assign n15021 = ~n14982 & n15020 ;
  assign n15022 = ~n15019 & ~n15021 ;
  assign n15023 = ~n15006 & n15022 ;
  assign n15024 = n14976 & ~n15023 ;
  assign n14970 = n14963 & ~n14969 ;
  assign n15025 = ~n14969 & n14982 ;
  assign n15026 = n14963 & ~n14976 ;
  assign n15027 = ~n15025 & ~n15026 ;
  assign n15028 = ~n14970 & ~n15027 ;
  assign n14998 = n14963 & n14997 ;
  assign n15000 = ~n14998 & ~n14999 ;
  assign n15003 = n14963 & n14982 ;
  assign n15029 = ~n14969 & ~n15003 ;
  assign n15030 = n15000 & n15029 ;
  assign n15031 = ~n15028 & ~n15030 ;
  assign n15032 = ~n15024 & n15031 ;
  assign n15033 = n14990 & ~n15032 ;
  assign n15011 = n14969 & ~n14976 ;
  assign n15012 = n14998 & ~n15011 ;
  assign n15013 = n14969 & n14999 ;
  assign n15014 = ~n15012 & ~n15013 ;
  assign n15015 = ~n14982 & ~n15014 ;
  assign n14991 = n14976 & n14982 ;
  assign n15001 = n14969 & n15000 ;
  assign n15002 = n14991 & n15001 ;
  assign n15004 = ~n14969 & ~n14997 ;
  assign n15005 = n15003 & n15004 ;
  assign n15007 = ~n14963 & ~n14982 ;
  assign n15008 = ~n15006 & n15007 ;
  assign n15009 = ~n15005 & ~n15008 ;
  assign n15010 = ~n14976 & ~n15009 ;
  assign n15016 = ~n15002 & ~n15010 ;
  assign n15017 = ~n15015 & n15016 ;
  assign n15018 = ~n14990 & ~n15017 ;
  assign n15040 = n15020 & n15025 ;
  assign n15036 = n14969 & n14997 ;
  assign n15037 = n15003 & n15036 ;
  assign n15038 = n14969 & ~n14997 ;
  assign n15039 = ~n14982 & n15038 ;
  assign n15041 = ~n15037 & ~n15039 ;
  assign n15042 = ~n15040 & n15041 ;
  assign n15043 = ~n14976 & ~n15042 ;
  assign n14983 = n14976 & ~n14982 ;
  assign n14984 = n14970 & n14983 ;
  assign n15034 = n14976 & n14999 ;
  assign n15035 = n15025 & n15034 ;
  assign n15044 = ~n14984 & ~n15035 ;
  assign n15045 = ~n15043 & n15044 ;
  assign n15046 = ~n15018 & n15045 ;
  assign n15047 = ~n15033 & n15046 ;
  assign n15048 = ~\u2_L7_reg[31]/NET0131  & ~n15047 ;
  assign n15049 = \u2_L7_reg[31]/NET0131  & n15047 ;
  assign n15050 = ~n15048 & ~n15049 ;
  assign n15051 = decrypt_pad & ~\u2_uk_K_r7_reg[16]/NET0131  ;
  assign n15052 = ~decrypt_pad & ~\u2_uk_K_r7_reg[23]/P0001  ;
  assign n15053 = ~n15051 & ~n15052 ;
  assign n15054 = \u2_R7_reg[24]/NET0131  & ~n15053 ;
  assign n15055 = ~\u2_R7_reg[24]/NET0131  & n15053 ;
  assign n15056 = ~n15054 & ~n15055 ;
  assign n15057 = decrypt_pad & ~\u2_uk_K_r7_reg[14]/NET0131  ;
  assign n15058 = ~decrypt_pad & ~\u2_uk_K_r7_reg[21]/NET0131  ;
  assign n15059 = ~n15057 & ~n15058 ;
  assign n15060 = \u2_R7_reg[23]/NET0131  & ~n15059 ;
  assign n15061 = ~\u2_R7_reg[23]/NET0131  & n15059 ;
  assign n15062 = ~n15060 & ~n15061 ;
  assign n15063 = decrypt_pad & ~\u2_uk_K_r7_reg[50]/NET0131  ;
  assign n15064 = ~decrypt_pad & ~\u2_uk_K_r7_reg[2]/NET0131  ;
  assign n15065 = ~n15063 & ~n15064 ;
  assign n15066 = \u2_R7_reg[20]/NET0131  & ~n15065 ;
  assign n15067 = ~\u2_R7_reg[20]/NET0131  & n15065 ;
  assign n15068 = ~n15066 & ~n15067 ;
  assign n15076 = decrypt_pad & ~\u2_uk_K_r7_reg[38]/NET0131  ;
  assign n15077 = ~decrypt_pad & ~\u2_uk_K_r7_reg[45]/NET0131  ;
  assign n15078 = ~n15076 & ~n15077 ;
  assign n15079 = \u2_R7_reg[21]/NET0131  & ~n15078 ;
  assign n15080 = ~\u2_R7_reg[21]/NET0131  & n15078 ;
  assign n15081 = ~n15079 & ~n15080 ;
  assign n15088 = ~n15068 & n15081 ;
  assign n15069 = decrypt_pad & ~\u2_uk_K_r7_reg[1]/NET0131  ;
  assign n15070 = ~decrypt_pad & ~\u2_uk_K_r7_reg[8]/NET0131  ;
  assign n15071 = ~n15069 & ~n15070 ;
  assign n15072 = \u2_R7_reg[22]/NET0131  & ~n15071 ;
  assign n15073 = ~\u2_R7_reg[22]/NET0131  & n15071 ;
  assign n15074 = ~n15072 & ~n15073 ;
  assign n15093 = decrypt_pad & ~\u2_uk_K_r7_reg[35]/NET0131  ;
  assign n15094 = ~decrypt_pad & ~\u2_uk_K_r7_reg[42]/NET0131  ;
  assign n15095 = ~n15093 & ~n15094 ;
  assign n15096 = \u2_R7_reg[25]/NET0131  & ~n15095 ;
  assign n15097 = ~\u2_R7_reg[25]/NET0131  & n15095 ;
  assign n15098 = ~n15096 & ~n15097 ;
  assign n15111 = n15068 & n15098 ;
  assign n15112 = n15074 & ~n15111 ;
  assign n15131 = ~n15088 & n15112 ;
  assign n15075 = ~n15068 & ~n15074 ;
  assign n15132 = n15075 & n15098 ;
  assign n15133 = n15081 & n15132 ;
  assign n15134 = ~n15131 & ~n15133 ;
  assign n15135 = ~n15062 & ~n15134 ;
  assign n15103 = n15068 & ~n15098 ;
  assign n15124 = ~n15081 & n15103 ;
  assign n15125 = ~n15074 & n15124 ;
  assign n15089 = n15074 & n15088 ;
  assign n15126 = n15081 & n15098 ;
  assign n15127 = n15068 & n15126 ;
  assign n15128 = ~n15089 & ~n15127 ;
  assign n15129 = ~n15125 & n15128 ;
  assign n15130 = n15062 & ~n15129 ;
  assign n15104 = ~n15062 & ~n15074 ;
  assign n15136 = n15104 & n15111 ;
  assign n15137 = ~n15081 & n15136 ;
  assign n15138 = ~n15130 & ~n15137 ;
  assign n15139 = ~n15135 & n15138 ;
  assign n15140 = n15056 & ~n15139 ;
  assign n15082 = n15068 & n15074 ;
  assign n15083 = ~n15081 & n15082 ;
  assign n15084 = n15062 & ~n15075 ;
  assign n15085 = ~n15083 & n15084 ;
  assign n15086 = ~n15074 & n15081 ;
  assign n15087 = n15068 & n15086 ;
  assign n15090 = ~n15062 & ~n15087 ;
  assign n15091 = ~n15089 & n15090 ;
  assign n15092 = ~n15085 & ~n15091 ;
  assign n15105 = ~n15086 & ~n15104 ;
  assign n15106 = n15103 & ~n15105 ;
  assign n15099 = n15083 & n15098 ;
  assign n15100 = ~n15068 & ~n15081 ;
  assign n15101 = n15098 & n15100 ;
  assign n15102 = n15062 & n15101 ;
  assign n15107 = ~n15099 & ~n15102 ;
  assign n15108 = ~n15106 & n15107 ;
  assign n15109 = ~n15092 & n15108 ;
  assign n15110 = ~n15056 & ~n15109 ;
  assign n15118 = n15081 & n15103 ;
  assign n15119 = ~n15062 & n15118 ;
  assign n15120 = ~n15102 & ~n15119 ;
  assign n15121 = ~n15074 & ~n15120 ;
  assign n15113 = ~n15068 & ~n15098 ;
  assign n15114 = n15081 & n15113 ;
  assign n15115 = ~n15074 & ~n15114 ;
  assign n15116 = n15062 & ~n15112 ;
  assign n15117 = ~n15115 & n15116 ;
  assign n15122 = ~n15081 & n15113 ;
  assign n15123 = n15104 & n15122 ;
  assign n15141 = ~n15117 & ~n15123 ;
  assign n15142 = ~n15121 & n15141 ;
  assign n15143 = ~n15110 & n15142 ;
  assign n15144 = ~n15140 & n15143 ;
  assign n15145 = \u2_L7_reg[11]/NET0131  & ~n15144 ;
  assign n15146 = ~\u2_L7_reg[11]/NET0131  & n15144 ;
  assign n15147 = ~n15145 & ~n15146 ;
  assign n15148 = decrypt_pad & ~\u2_uk_K_r7_reg[54]/NET0131  ;
  assign n15149 = ~decrypt_pad & ~\u2_uk_K_r7_reg[4]/NET0131  ;
  assign n15150 = ~n15148 & ~n15149 ;
  assign n15151 = \u2_R7_reg[17]/NET0131  & ~n15150 ;
  assign n15152 = ~\u2_R7_reg[17]/NET0131  & n15150 ;
  assign n15153 = ~n15151 & ~n15152 ;
  assign n15154 = decrypt_pad & ~\u2_uk_K_r7_reg[13]/NET0131  ;
  assign n15155 = ~decrypt_pad & ~\u2_uk_K_r7_reg[20]/NET0131  ;
  assign n15156 = ~n15154 & ~n15155 ;
  assign n15157 = \u2_R7_reg[12]/NET0131  & ~n15156 ;
  assign n15158 = ~\u2_R7_reg[12]/NET0131  & n15156 ;
  assign n15159 = ~n15157 & ~n15158 ;
  assign n15160 = ~n15153 & n15159 ;
  assign n15179 = decrypt_pad & ~\u2_uk_K_r7_reg[33]/NET0131  ;
  assign n15180 = ~decrypt_pad & ~\u2_uk_K_r7_reg[40]/NET0131  ;
  assign n15181 = ~n15179 & ~n15180 ;
  assign n15182 = \u2_R7_reg[14]/NET0131  & ~n15181 ;
  assign n15183 = ~\u2_R7_reg[14]/NET0131  & n15181 ;
  assign n15184 = ~n15182 & ~n15183 ;
  assign n15187 = ~n15159 & ~n15184 ;
  assign n15161 = decrypt_pad & ~\u2_uk_K_r7_reg[32]/NET0131  ;
  assign n15162 = ~decrypt_pad & ~\u2_uk_K_r7_reg[39]/NET0131  ;
  assign n15163 = ~n15161 & ~n15162 ;
  assign n15164 = \u2_R7_reg[13]/NET0131  & ~n15163 ;
  assign n15165 = ~\u2_R7_reg[13]/NET0131  & n15163 ;
  assign n15166 = ~n15164 & ~n15165 ;
  assign n15168 = decrypt_pad & ~\u2_uk_K_r7_reg[41]/NET0131  ;
  assign n15169 = ~decrypt_pad & ~\u2_uk_K_r7_reg[48]/NET0131  ;
  assign n15170 = ~n15168 & ~n15169 ;
  assign n15171 = \u2_R7_reg[15]/NET0131  & ~n15170 ;
  assign n15172 = ~\u2_R7_reg[15]/NET0131  & n15170 ;
  assign n15173 = ~n15171 & ~n15172 ;
  assign n15192 = n15166 & n15173 ;
  assign n15193 = ~n15187 & n15192 ;
  assign n15194 = ~n15160 & n15193 ;
  assign n15204 = ~n15159 & ~n15166 ;
  assign n15205 = ~n15153 & ~n15184 ;
  assign n15206 = n15204 & n15205 ;
  assign n15209 = decrypt_pad & ~\u2_uk_K_r7_reg[17]/NET0131  ;
  assign n15210 = ~decrypt_pad & ~\u2_uk_K_r7_reg[24]/NET0131  ;
  assign n15211 = ~n15209 & ~n15210 ;
  assign n15212 = \u2_R7_reg[16]/NET0131  & ~n15211 ;
  assign n15213 = ~\u2_R7_reg[16]/NET0131  & n15211 ;
  assign n15214 = ~n15212 & ~n15213 ;
  assign n15215 = ~n15206 & ~n15214 ;
  assign n15216 = ~n15194 & n15215 ;
  assign n15188 = n15159 & n15184 ;
  assign n15195 = ~n15153 & ~n15188 ;
  assign n15175 = n15153 & n15166 ;
  assign n15196 = ~n15173 & ~n15175 ;
  assign n15197 = ~n15195 & n15196 ;
  assign n15198 = ~n15159 & n15166 ;
  assign n15199 = ~n15153 & n15198 ;
  assign n15200 = n15184 & n15199 ;
  assign n15217 = ~n15197 & ~n15200 ;
  assign n15201 = n15159 & ~n15166 ;
  assign n15202 = ~n15184 & n15201 ;
  assign n15203 = n15153 & n15202 ;
  assign n15186 = ~n15153 & ~n15166 ;
  assign n15207 = ~n15159 & n15186 ;
  assign n15208 = n15173 & n15207 ;
  assign n15218 = ~n15203 & ~n15208 ;
  assign n15219 = n15217 & n15218 ;
  assign n15220 = n15216 & n15219 ;
  assign n15225 = ~n15198 & ~n15201 ;
  assign n15226 = ~n15184 & ~n15225 ;
  assign n15227 = n15184 & n15204 ;
  assign n15228 = ~n15153 & n15227 ;
  assign n15229 = ~n15226 & ~n15228 ;
  assign n15230 = ~n15173 & ~n15229 ;
  assign n15167 = n15160 & n15166 ;
  assign n15174 = n15167 & n15173 ;
  assign n15231 = ~n15174 & n15214 ;
  assign n15189 = ~n15187 & ~n15188 ;
  assign n15221 = n15175 & ~n15189 ;
  assign n15222 = n15153 & ~n15159 ;
  assign n15223 = n15173 & n15222 ;
  assign n15224 = ~n15166 & n15223 ;
  assign n15232 = ~n15221 & ~n15224 ;
  assign n15233 = n15231 & n15232 ;
  assign n15234 = ~n15230 & n15233 ;
  assign n15235 = ~n15220 & ~n15234 ;
  assign n15176 = ~n15159 & n15175 ;
  assign n15177 = ~n15173 & n15176 ;
  assign n15178 = ~n15174 & ~n15177 ;
  assign n15185 = ~n15178 & ~n15184 ;
  assign n15190 = n15173 & ~n15189 ;
  assign n15191 = n15186 & n15190 ;
  assign n15236 = ~n15185 & ~n15191 ;
  assign n15237 = ~n15235 & n15236 ;
  assign n15238 = ~\u2_L7_reg[20]/NET0131  & ~n15237 ;
  assign n15239 = \u2_L7_reg[20]/NET0131  & n15237 ;
  assign n15240 = ~n15238 & ~n15239 ;
  assign n15241 = decrypt_pad & ~\u2_uk_K_r7_reg[21]/NET0131  ;
  assign n15242 = ~decrypt_pad & ~\u2_uk_K_r7_reg[28]/NET0131  ;
  assign n15243 = ~n15241 & ~n15242 ;
  assign n15244 = \u2_R7_reg[28]/NET0131  & ~n15243 ;
  assign n15245 = ~\u2_R7_reg[28]/NET0131  & n15243 ;
  assign n15246 = ~n15244 & ~n15245 ;
  assign n15247 = decrypt_pad & ~\u2_uk_K_r7_reg[9]/NET0131  ;
  assign n15248 = ~decrypt_pad & ~\u2_uk_K_r7_reg[16]/NET0131  ;
  assign n15249 = ~n15247 & ~n15248 ;
  assign n15250 = \u2_R7_reg[1]/NET0131  & ~n15249 ;
  assign n15251 = ~\u2_R7_reg[1]/NET0131  & n15249 ;
  assign n15252 = ~n15250 & ~n15251 ;
  assign n15253 = n15246 & ~n15252 ;
  assign n15254 = decrypt_pad & ~\u2_uk_K_r7_reg[52]/NET0131  ;
  assign n15255 = ~decrypt_pad & ~\u2_uk_K_r7_reg[0]/NET0131  ;
  assign n15256 = ~n15254 & ~n15255 ;
  assign n15257 = \u2_R7_reg[29]/NET0131  & ~n15256 ;
  assign n15258 = ~\u2_R7_reg[29]/NET0131  & n15256 ;
  assign n15259 = ~n15257 & ~n15258 ;
  assign n15260 = decrypt_pad & ~\u2_uk_K_r7_reg[49]/NET0131  ;
  assign n15261 = ~decrypt_pad & ~\u2_uk_K_r7_reg[1]/NET0131  ;
  assign n15262 = ~n15260 & ~n15261 ;
  assign n15263 = \u2_R7_reg[30]/NET0131  & ~n15262 ;
  assign n15264 = ~\u2_R7_reg[30]/NET0131  & n15262 ;
  assign n15265 = ~n15263 & ~n15264 ;
  assign n15266 = ~n15259 & n15265 ;
  assign n15267 = n15253 & n15266 ;
  assign n15268 = ~n15246 & n15252 ;
  assign n15269 = ~n15259 & n15268 ;
  assign n15270 = ~n15267 & ~n15269 ;
  assign n15271 = decrypt_pad & ~\u2_uk_K_r7_reg[37]/NET0131  ;
  assign n15272 = ~decrypt_pad & ~\u2_uk_K_r7_reg[44]/NET0131  ;
  assign n15273 = ~n15271 & ~n15272 ;
  assign n15274 = \u2_R7_reg[31]/P0001  & ~n15273 ;
  assign n15275 = ~\u2_R7_reg[31]/P0001  & n15273 ;
  assign n15276 = ~n15274 & ~n15275 ;
  assign n15277 = ~n15270 & n15276 ;
  assign n15285 = ~n15253 & ~n15276 ;
  assign n15283 = ~n15252 & ~n15265 ;
  assign n15284 = n15252 & ~n15259 ;
  assign n15286 = ~n15283 & ~n15284 ;
  assign n15287 = n15285 & n15286 ;
  assign n15281 = n15246 & ~n15265 ;
  assign n15288 = ~n15252 & n15259 ;
  assign n15289 = n15281 & n15288 ;
  assign n15278 = n15259 & n15265 ;
  assign n15279 = n15246 & n15252 ;
  assign n15280 = n15278 & n15279 ;
  assign n15282 = ~n15276 & n15281 ;
  assign n15290 = ~n15280 & ~n15282 ;
  assign n15291 = ~n15289 & n15290 ;
  assign n15292 = ~n15287 & n15291 ;
  assign n15293 = ~n15277 & n15292 ;
  assign n15294 = decrypt_pad & ~\u2_uk_K_r7_reg[43]/NET0131  ;
  assign n15295 = ~decrypt_pad & ~\u2_uk_K_r7_reg[50]/NET0131  ;
  assign n15296 = ~n15294 & ~n15295 ;
  assign n15297 = \u2_R7_reg[32]/NET0131  & ~n15296 ;
  assign n15298 = ~\u2_R7_reg[32]/NET0131  & n15296 ;
  assign n15299 = ~n15297 & ~n15298 ;
  assign n15300 = ~n15293 & ~n15299 ;
  assign n15305 = ~n15281 & ~n15288 ;
  assign n15322 = n15276 & ~n15289 ;
  assign n15323 = ~n15305 & n15322 ;
  assign n15318 = ~n15246 & ~n15276 ;
  assign n15319 = ~n15259 & ~n15265 ;
  assign n15320 = n15318 & n15319 ;
  assign n15321 = n15268 & n15278 ;
  assign n15324 = ~n15320 & ~n15321 ;
  assign n15325 = ~n15323 & n15324 ;
  assign n15326 = n15299 & ~n15325 ;
  assign n15308 = n15265 & n15284 ;
  assign n15309 = ~n15246 & n15308 ;
  assign n15301 = ~n15246 & ~n15252 ;
  assign n15302 = ~n15259 & n15301 ;
  assign n15303 = ~n15265 & n15302 ;
  assign n15304 = n15259 & ~n15265 ;
  assign n15306 = ~n15253 & ~n15304 ;
  assign n15307 = ~n15305 & n15306 ;
  assign n15310 = ~n15303 & ~n15307 ;
  assign n15311 = ~n15309 & n15310 ;
  assign n15312 = n15276 & ~n15311 ;
  assign n15313 = ~n15276 & n15289 ;
  assign n15315 = n15246 & ~n15259 ;
  assign n15314 = n15265 & ~n15276 ;
  assign n15316 = n15299 & n15314 ;
  assign n15317 = n15315 & n15316 ;
  assign n15327 = ~n15313 & ~n15317 ;
  assign n15328 = ~n15312 & n15327 ;
  assign n15329 = ~n15326 & n15328 ;
  assign n15330 = ~n15300 & n15329 ;
  assign n15331 = \u2_L7_reg[5]/NET0131  & ~n15330 ;
  assign n15332 = ~\u2_L7_reg[5]/NET0131  & n15330 ;
  assign n15333 = ~n15331 & ~n15332 ;
  assign n15355 = n15166 & ~n15184 ;
  assign n15356 = n15160 & ~n15355 ;
  assign n15357 = n15176 & ~n15184 ;
  assign n15358 = ~n15356 & ~n15357 ;
  assign n15359 = ~n15173 & ~n15358 ;
  assign n15347 = n15153 & n15184 ;
  assign n15348 = n15225 & n15347 ;
  assign n15353 = ~n15199 & ~n15203 ;
  assign n15354 = n15173 & ~n15353 ;
  assign n15360 = ~n15348 & ~n15354 ;
  assign n15361 = ~n15359 & n15360 ;
  assign n15362 = n15214 & ~n15361 ;
  assign n15334 = n15173 & n15184 ;
  assign n15335 = ~n15207 & ~n15223 ;
  assign n15336 = ~n15334 & ~n15335 ;
  assign n15337 = ~n15166 & n15173 ;
  assign n15340 = n15159 & ~n15337 ;
  assign n15341 = ~n15184 & ~n15186 ;
  assign n15342 = n15340 & n15341 ;
  assign n15338 = ~n15160 & ~n15188 ;
  assign n15339 = n15337 & ~n15338 ;
  assign n15343 = ~n15200 & ~n15339 ;
  assign n15344 = ~n15342 & n15343 ;
  assign n15345 = ~n15336 & n15344 ;
  assign n15346 = ~n15214 & ~n15345 ;
  assign n15349 = ~n15206 & ~n15348 ;
  assign n15350 = ~n15173 & ~n15349 ;
  assign n15351 = n15159 & ~n15205 ;
  assign n15352 = n15193 & ~n15351 ;
  assign n15363 = ~n15350 & ~n15352 ;
  assign n15364 = ~n15346 & n15363 ;
  assign n15365 = ~n15362 & n15364 ;
  assign n15366 = ~\u2_L7_reg[10]/NET0131  & ~n15365 ;
  assign n15367 = \u2_L7_reg[10]/NET0131  & n15365 ;
  assign n15368 = ~n15366 & ~n15367 ;
  assign n15371 = n14876 & n14882 ;
  assign n15379 = ~n14942 & ~n15371 ;
  assign n15369 = n14889 & ~n14895 ;
  assign n15377 = ~n14896 & ~n15369 ;
  assign n15378 = n14882 & n14889 ;
  assign n15380 = n15377 & ~n15378 ;
  assign n15381 = n15379 & n15380 ;
  assign n15374 = ~n14903 & ~n14930 ;
  assign n15375 = ~n14902 & n15374 ;
  assign n15376 = ~n14921 & ~n15375 ;
  assign n15372 = ~n14923 & ~n15371 ;
  assign n15373 = n14896 & ~n15372 ;
  assign n15370 = n14942 & n15369 ;
  assign n15382 = ~n14911 & ~n15370 ;
  assign n15383 = ~n15373 & n15382 ;
  assign n15384 = ~n15376 & n15383 ;
  assign n15385 = ~n15381 & n15384 ;
  assign n15389 = ~n14947 & ~n15378 ;
  assign n15390 = n14921 & ~n15389 ;
  assign n15391 = n14911 & ~n14943 ;
  assign n15392 = ~n14900 & n15391 ;
  assign n15386 = n14897 & ~n14921 ;
  assign n15387 = ~n14941 & ~n15371 ;
  assign n15388 = ~n15374 & n15387 ;
  assign n15393 = ~n15386 & ~n15388 ;
  assign n15394 = n15392 & n15393 ;
  assign n15395 = ~n15390 & n15394 ;
  assign n15396 = ~n15385 & ~n15395 ;
  assign n15397 = \u2_L7_reg[12]/NET0131  & n15396 ;
  assign n15398 = ~\u2_L7_reg[12]/NET0131  & ~n15396 ;
  assign n15399 = ~n15397 & ~n15398 ;
  assign n15400 = ~n15246 & ~n15283 ;
  assign n15401 = n15259 & ~n15400 ;
  assign n15402 = ~n15269 & ~n15401 ;
  assign n15403 = n15276 & ~n15402 ;
  assign n15404 = n15283 & n15315 ;
  assign n15405 = ~n15403 & ~n15404 ;
  assign n15406 = ~n15299 & ~n15405 ;
  assign n15409 = n15246 & n15265 ;
  assign n15410 = ~n15314 & ~n15409 ;
  assign n15411 = n15284 & ~n15410 ;
  assign n15408 = n15276 & n15302 ;
  assign n15407 = n15259 & n15281 ;
  assign n15412 = n15278 & n15301 ;
  assign n15413 = ~n15407 & ~n15412 ;
  assign n15414 = ~n15408 & n15413 ;
  assign n15415 = ~n15411 & n15414 ;
  assign n15416 = n15299 & ~n15415 ;
  assign n15420 = ~n15276 & ~n15412 ;
  assign n15417 = n15268 & n15304 ;
  assign n15418 = ~n15265 & n15299 ;
  assign n15419 = n15315 & ~n15418 ;
  assign n15421 = ~n15417 & ~n15419 ;
  assign n15422 = n15420 & n15421 ;
  assign n15423 = ~n15303 & n15422 ;
  assign n15424 = n15268 & n15319 ;
  assign n15425 = n15276 & ~n15321 ;
  assign n15426 = ~n15424 & n15425 ;
  assign n15427 = ~n15423 & ~n15426 ;
  assign n15428 = ~n15416 & ~n15427 ;
  assign n15429 = ~n15406 & n15428 ;
  assign n15430 = ~\u2_L7_reg[15]/NET0131  & ~n15429 ;
  assign n15431 = \u2_L7_reg[15]/NET0131  & n15429 ;
  assign n15432 = ~n15430 & ~n15431 ;
  assign n15436 = ~n14969 & ~n14982 ;
  assign n15437 = ~n14963 & ~n15436 ;
  assign n15441 = n14998 & n15436 ;
  assign n15442 = ~n15437 & ~n15441 ;
  assign n15443 = n14976 & ~n15442 ;
  assign n15433 = n14963 & n15039 ;
  assign n15434 = n14990 & ~n15433 ;
  assign n15435 = n14963 & ~n14982 ;
  assign n15438 = ~n14976 & ~n15435 ;
  assign n15439 = ~n15437 & n15438 ;
  assign n15440 = n14982 & n15036 ;
  assign n15444 = ~n15439 & ~n15440 ;
  assign n15445 = n15434 & n15444 ;
  assign n15446 = ~n15443 & n15445 ;
  assign n15451 = ~n14969 & ~n15000 ;
  assign n15452 = ~n14982 & n14999 ;
  assign n15453 = ~n15451 & ~n15452 ;
  assign n15454 = ~n14976 & ~n15453 ;
  assign n15447 = ~n14976 & ~n15038 ;
  assign n15448 = n14963 & ~n15006 ;
  assign n15449 = ~n15039 & n15448 ;
  assign n15450 = ~n15447 & n15449 ;
  assign n15455 = ~n14990 & ~n15040 ;
  assign n15456 = ~n15450 & n15455 ;
  assign n15457 = ~n15454 & n15456 ;
  assign n15458 = ~n15446 & ~n15457 ;
  assign n15459 = n14969 & n14976 ;
  assign n15460 = ~n15022 & n15459 ;
  assign n15461 = ~n15458 & ~n15460 ;
  assign n15462 = ~\u2_L7_reg[17]/NET0131  & ~n15461 ;
  assign n15463 = \u2_L7_reg[17]/NET0131  & n15461 ;
  assign n15464 = ~n15462 & ~n15463 ;
  assign n15465 = decrypt_pad & ~\u2_uk_K_r7_reg[44]/NET0131  ;
  assign n15466 = ~decrypt_pad & ~\u2_uk_K_r7_reg[51]/NET0131  ;
  assign n15467 = ~n15465 & ~n15466 ;
  assign n15468 = \u2_R7_reg[19]/NET0131  & ~n15467 ;
  assign n15469 = ~\u2_R7_reg[19]/NET0131  & n15467 ;
  assign n15470 = ~n15468 & ~n15469 ;
  assign n15471 = decrypt_pad & ~\u2_uk_K_r7_reg[2]/NET0131  ;
  assign n15472 = ~decrypt_pad & ~\u2_uk_K_r7_reg[9]/NET0131  ;
  assign n15473 = ~n15471 & ~n15472 ;
  assign n15474 = \u2_R7_reg[18]/NET0131  & ~n15473 ;
  assign n15475 = ~\u2_R7_reg[18]/NET0131  & n15473 ;
  assign n15476 = ~n15474 & ~n15475 ;
  assign n15477 = decrypt_pad & ~\u2_uk_K_r7_reg[8]/NET0131  ;
  assign n15478 = ~decrypt_pad & ~\u2_uk_K_r7_reg[15]/NET0131  ;
  assign n15479 = ~n15477 & ~n15478 ;
  assign n15480 = \u2_R7_reg[17]/NET0131  & ~n15479 ;
  assign n15481 = ~\u2_R7_reg[17]/NET0131  & n15479 ;
  assign n15482 = ~n15480 & ~n15481 ;
  assign n15484 = decrypt_pad & ~\u2_uk_K_r7_reg[45]/NET0131  ;
  assign n15485 = ~decrypt_pad & ~\u2_uk_K_r7_reg[52]/NET0131  ;
  assign n15486 = ~n15484 & ~n15485 ;
  assign n15487 = \u2_R7_reg[16]/NET0131  & ~n15486 ;
  assign n15488 = ~\u2_R7_reg[16]/NET0131  & n15486 ;
  assign n15489 = ~n15487 & ~n15488 ;
  assign n15491 = decrypt_pad & ~\u2_uk_K_r7_reg[29]/NET0131  ;
  assign n15492 = ~decrypt_pad & ~\u2_uk_K_r7_reg[36]/NET0131  ;
  assign n15493 = ~n15491 & ~n15492 ;
  assign n15494 = \u2_R7_reg[21]/NET0131  & ~n15493 ;
  assign n15495 = ~\u2_R7_reg[21]/NET0131  & n15493 ;
  assign n15496 = ~n15494 & ~n15495 ;
  assign n15497 = n15489 & ~n15496 ;
  assign n15508 = ~n15482 & n15497 ;
  assign n15509 = ~n15476 & n15508 ;
  assign n15483 = ~n15476 & n15482 ;
  assign n15510 = n15489 & n15496 ;
  assign n15511 = n15483 & n15510 ;
  assign n15500 = n15482 & ~n15496 ;
  assign n15505 = n15476 & n15500 ;
  assign n15506 = ~n15489 & n15496 ;
  assign n15507 = ~n15482 & n15506 ;
  assign n15512 = ~n15505 & ~n15507 ;
  assign n15513 = ~n15511 & n15512 ;
  assign n15514 = ~n15509 & n15513 ;
  assign n15515 = ~n15470 & ~n15514 ;
  assign n15490 = n15483 & ~n15489 ;
  assign n15498 = n15476 & n15489 ;
  assign n15499 = n15496 & ~n15498 ;
  assign n15501 = ~n15497 & ~n15500 ;
  assign n15502 = ~n15499 & n15501 ;
  assign n15503 = ~n15490 & ~n15502 ;
  assign n15504 = n15470 & ~n15503 ;
  assign n15516 = ~n15476 & n15496 ;
  assign n15517 = ~n15497 & ~n15516 ;
  assign n15518 = ~n15482 & ~n15489 ;
  assign n15519 = n15476 & n15482 ;
  assign n15520 = ~n15518 & ~n15519 ;
  assign n15521 = n15517 & n15520 ;
  assign n15522 = ~n15504 & ~n15521 ;
  assign n15523 = ~n15515 & n15522 ;
  assign n15524 = decrypt_pad & ~\u2_uk_K_r7_reg[28]/NET0131  ;
  assign n15525 = ~decrypt_pad & ~\u2_uk_K_r7_reg[35]/NET0131  ;
  assign n15526 = ~n15524 & ~n15525 ;
  assign n15527 = \u2_R7_reg[20]/NET0131  & ~n15526 ;
  assign n15528 = ~\u2_R7_reg[20]/NET0131  & n15526 ;
  assign n15529 = ~n15527 & ~n15528 ;
  assign n15530 = ~n15523 & ~n15529 ;
  assign n15534 = ~n15490 & n15499 ;
  assign n15535 = n15489 & n15500 ;
  assign n15536 = ~n15534 & ~n15535 ;
  assign n15537 = n15470 & ~n15536 ;
  assign n15538 = n15482 & n15506 ;
  assign n15539 = ~n15496 & n15518 ;
  assign n15540 = ~n15538 & ~n15539 ;
  assign n15541 = ~n15470 & ~n15476 ;
  assign n15542 = ~n15540 & n15541 ;
  assign n15531 = n15476 & ~n15482 ;
  assign n15532 = ~n15483 & ~n15531 ;
  assign n15533 = n15497 & ~n15532 ;
  assign n15543 = n15470 & n15476 ;
  assign n15544 = n15510 & ~n15543 ;
  assign n15545 = n15532 & n15544 ;
  assign n15546 = ~n15533 & ~n15545 ;
  assign n15547 = ~n15542 & n15546 ;
  assign n15548 = ~n15537 & n15547 ;
  assign n15549 = n15529 & ~n15548 ;
  assign n15550 = n15476 & n15539 ;
  assign n15551 = ~n15476 & n15535 ;
  assign n15552 = ~n15550 & ~n15551 ;
  assign n15553 = n15470 & ~n15552 ;
  assign n15554 = n15476 & n15507 ;
  assign n15555 = ~n15489 & n15505 ;
  assign n15556 = ~n15554 & ~n15555 ;
  assign n15557 = ~n15470 & ~n15556 ;
  assign n15558 = ~n15553 & ~n15557 ;
  assign n15559 = ~n15549 & n15558 ;
  assign n15560 = ~n15530 & n15559 ;
  assign n15561 = ~\u2_L7_reg[14]/NET0131  & ~n15560 ;
  assign n15562 = \u2_L7_reg[14]/NET0131  & n15560 ;
  assign n15563 = ~n15561 & ~n15562 ;
  assign n15564 = ~n15186 & ~n15205 ;
  assign n15565 = n15190 & ~n15564 ;
  assign n15566 = n15153 & ~n15166 ;
  assign n15567 = ~n15205 & ~n15566 ;
  assign n15568 = n15340 & ~n15567 ;
  assign n15569 = ~n15214 & ~n15221 ;
  assign n15570 = ~n15568 & n15569 ;
  assign n15571 = ~n15565 & n15570 ;
  assign n15574 = ~n15176 & ~n15355 ;
  assign n15575 = ~n15160 & ~n15173 ;
  assign n15576 = ~n15574 & n15575 ;
  assign n15572 = n15167 & n15184 ;
  assign n15573 = n15214 & ~n15572 ;
  assign n15577 = ~n15227 & n15573 ;
  assign n15578 = ~n15576 & n15577 ;
  assign n15579 = ~n15571 & ~n15578 ;
  assign n15580 = ~n15173 & ~n15228 ;
  assign n15581 = ~n15572 & n15580 ;
  assign n15582 = ~n15202 & ~n15566 ;
  assign n15583 = n15214 & ~n15582 ;
  assign n15584 = n15173 & ~n15200 ;
  assign n15585 = ~n15348 & n15584 ;
  assign n15586 = ~n15583 & n15585 ;
  assign n15587 = ~n15581 & ~n15586 ;
  assign n15588 = ~n15579 & ~n15587 ;
  assign n15589 = ~\u2_L7_reg[1]/NET0131  & ~n15588 ;
  assign n15590 = \u2_L7_reg[1]/NET0131  & n15588 ;
  assign n15591 = ~n15589 & ~n15590 ;
  assign n15597 = n15288 & n15318 ;
  assign n15601 = ~n15267 & ~n15299 ;
  assign n15602 = ~n15597 & n15601 ;
  assign n15598 = ~n15266 & ~n15288 ;
  assign n15599 = n15246 & n15276 ;
  assign n15600 = ~n15598 & n15599 ;
  assign n15603 = ~n15303 & ~n15600 ;
  assign n15604 = n15602 & n15603 ;
  assign n15592 = ~n15282 & ~n15407 ;
  assign n15593 = n15252 & ~n15592 ;
  assign n15594 = n15252 & n15314 ;
  assign n15595 = ~n15278 & ~n15594 ;
  assign n15596 = ~n15246 & ~n15595 ;
  assign n15605 = ~n15593 & ~n15596 ;
  assign n15606 = n15604 & n15605 ;
  assign n15607 = n15253 & n15259 ;
  assign n15608 = ~n15302 & ~n15607 ;
  assign n15609 = n15265 & ~n15608 ;
  assign n15617 = n15299 & ~n15424 ;
  assign n15618 = ~n15609 & n15617 ;
  assign n15610 = ~n15266 & n15276 ;
  assign n15611 = ~n15283 & ~n15301 ;
  assign n15612 = n15610 & n15611 ;
  assign n15613 = ~n15407 & n15612 ;
  assign n15614 = ~n15283 & ~n15308 ;
  assign n15615 = n15246 & ~n15276 ;
  assign n15616 = ~n15614 & n15615 ;
  assign n15619 = ~n15613 & ~n15616 ;
  assign n15620 = n15618 & n15619 ;
  assign n15621 = ~n15606 & ~n15620 ;
  assign n15622 = ~n15276 & ~n15279 ;
  assign n15623 = n15259 & n15276 ;
  assign n15624 = ~n15265 & ~n15315 ;
  assign n15625 = ~n15623 & n15624 ;
  assign n15626 = ~n15622 & n15625 ;
  assign n15627 = ~n15621 & ~n15626 ;
  assign n15628 = ~\u2_L7_reg[21]/NET0131  & ~n15627 ;
  assign n15629 = \u2_L7_reg[21]/NET0131  & n15627 ;
  assign n15630 = ~n15628 & ~n15629 ;
  assign n15633 = ~n15483 & ~n15496 ;
  assign n15634 = ~n15498 & n15633 ;
  assign n15632 = n15482 & n15510 ;
  assign n15635 = ~n15518 & ~n15632 ;
  assign n15636 = ~n15634 & n15635 ;
  assign n15637 = n15470 & ~n15636 ;
  assign n15638 = ~n15482 & n15510 ;
  assign n15639 = ~n15490 & ~n15638 ;
  assign n15640 = ~n15470 & ~n15639 ;
  assign n15631 = n15482 & n15516 ;
  assign n15641 = n15498 & n15500 ;
  assign n15642 = ~n15631 & ~n15641 ;
  assign n15643 = ~n15640 & n15642 ;
  assign n15644 = ~n15637 & n15643 ;
  assign n15645 = n15529 & ~n15644 ;
  assign n15657 = ~n15550 & ~n15641 ;
  assign n15658 = ~n15476 & n15507 ;
  assign n15659 = n15657 & ~n15658 ;
  assign n15660 = n15470 & ~n15659 ;
  assign n15651 = n15470 & ~n15500 ;
  assign n15650 = ~n15470 & ~n15518 ;
  assign n15652 = ~n15476 & ~n15650 ;
  assign n15653 = ~n15651 & n15652 ;
  assign n15646 = ~n15470 & n15508 ;
  assign n15647 = n15470 & ~n15496 ;
  assign n15648 = ~n15489 & n15519 ;
  assign n15649 = ~n15647 & n15648 ;
  assign n15654 = ~n15646 & ~n15649 ;
  assign n15655 = ~n15653 & n15654 ;
  assign n15656 = ~n15529 & ~n15655 ;
  assign n15661 = ~n15470 & n15489 ;
  assign n15662 = n15531 & n15661 ;
  assign n15663 = ~n15511 & ~n15662 ;
  assign n15664 = ~n15656 & n15663 ;
  assign n15665 = ~n15660 & n15664 ;
  assign n15666 = ~n15645 & n15665 ;
  assign n15667 = ~\u2_L7_reg[25]/NET0131  & ~n15666 ;
  assign n15668 = \u2_L7_reg[25]/NET0131  & n15666 ;
  assign n15669 = ~n15667 & ~n15668 ;
  assign n15673 = n15153 & ~n15173 ;
  assign n15674 = ~n15198 & n15673 ;
  assign n15675 = ~n15189 & n15674 ;
  assign n15672 = n15198 & n15205 ;
  assign n15676 = ~n15208 & ~n15672 ;
  assign n15677 = ~n15675 & n15676 ;
  assign n15670 = ~n15176 & ~n15223 ;
  assign n15671 = n15184 & ~n15670 ;
  assign n15678 = n15573 & ~n15671 ;
  assign n15679 = n15677 & n15678 ;
  assign n15680 = ~n15186 & ~n15227 ;
  assign n15681 = ~n15173 & ~n15680 ;
  assign n15684 = ~n15202 & ~n15214 ;
  assign n15685 = ~n15174 & n15684 ;
  assign n15682 = n15166 & ~n15222 ;
  assign n15683 = n15334 & n15682 ;
  assign n15686 = ~n15357 & ~n15683 ;
  assign n15687 = n15685 & n15686 ;
  assign n15688 = ~n15681 & n15687 ;
  assign n15689 = ~n15679 & ~n15688 ;
  assign n15690 = ~n15160 & ~n15682 ;
  assign n15691 = ~n15173 & ~n15184 ;
  assign n15692 = ~n15167 & n15691 ;
  assign n15693 = ~n15690 & n15692 ;
  assign n15694 = n15153 & n15173 ;
  assign n15695 = n15226 & n15694 ;
  assign n15696 = ~n15693 & ~n15695 ;
  assign n15697 = ~n15689 & n15696 ;
  assign n15698 = ~\u2_L7_reg[26]/NET0131  & ~n15697 ;
  assign n15699 = \u2_L7_reg[26]/NET0131  & n15697 ;
  assign n15700 = ~n15698 & ~n15699 ;
  assign n15738 = decrypt_pad & ~\u2_uk_K_r7_reg[48]/NET0131  ;
  assign n15739 = ~decrypt_pad & ~\u2_uk_K_r7_reg[55]/P0001  ;
  assign n15740 = ~n15738 & ~n15739 ;
  assign n15741 = \u2_R7_reg[8]/NET0131  & ~n15740 ;
  assign n15742 = ~\u2_R7_reg[8]/NET0131  & n15740 ;
  assign n15743 = ~n15741 & ~n15742 ;
  assign n15731 = decrypt_pad & ~\u2_uk_K_r7_reg[25]/NET0131  ;
  assign n15732 = ~decrypt_pad & ~\u2_uk_K_r7_reg[32]/NET0131  ;
  assign n15733 = ~n15731 & ~n15732 ;
  assign n15734 = \u2_R7_reg[7]/NET0131  & ~n15733 ;
  assign n15735 = ~\u2_R7_reg[7]/NET0131  & n15733 ;
  assign n15736 = ~n15734 & ~n15735 ;
  assign n15707 = decrypt_pad & ~\u2_uk_K_r7_reg[6]/NET0131  ;
  assign n15708 = ~decrypt_pad & ~\u2_uk_K_r7_reg[13]/NET0131  ;
  assign n15709 = ~n15707 & ~n15708 ;
  assign n15710 = \u2_R7_reg[6]/NET0131  & ~n15709 ;
  assign n15711 = ~\u2_R7_reg[6]/NET0131  & n15709 ;
  assign n15712 = ~n15710 & ~n15711 ;
  assign n15714 = decrypt_pad & ~\u2_uk_K_r7_reg[4]/NET0131  ;
  assign n15715 = ~decrypt_pad & ~\u2_uk_K_r7_reg[11]/NET0131  ;
  assign n15716 = ~n15714 & ~n15715 ;
  assign n15717 = \u2_R7_reg[4]/NET0131  & ~n15716 ;
  assign n15718 = ~\u2_R7_reg[4]/NET0131  & n15716 ;
  assign n15719 = ~n15717 & ~n15718 ;
  assign n15721 = decrypt_pad & ~\u2_uk_K_r7_reg[53]/NET0131  ;
  assign n15722 = ~decrypt_pad & ~\u2_uk_K_r7_reg[3]/NET0131  ;
  assign n15723 = ~n15721 & ~n15722 ;
  assign n15724 = \u2_R7_reg[9]/NET0131  & ~n15723 ;
  assign n15725 = ~\u2_R7_reg[9]/NET0131  & n15723 ;
  assign n15726 = ~n15724 & ~n15725 ;
  assign n15748 = n15719 & ~n15726 ;
  assign n15773 = ~n15712 & n15748 ;
  assign n15701 = decrypt_pad & ~\u2_uk_K_r7_reg[40]/NET0131  ;
  assign n15702 = ~decrypt_pad & ~\u2_uk_K_r7_reg[47]/NET0131  ;
  assign n15703 = ~n15701 & ~n15702 ;
  assign n15704 = \u2_R7_reg[5]/NET0131  & ~n15703 ;
  assign n15705 = ~\u2_R7_reg[5]/NET0131  & n15703 ;
  assign n15706 = ~n15704 & ~n15705 ;
  assign n15771 = n15706 & n15719 ;
  assign n15744 = ~n15719 & n15726 ;
  assign n15772 = ~n15706 & n15744 ;
  assign n15774 = ~n15771 & ~n15772 ;
  assign n15775 = ~n15773 & n15774 ;
  assign n15776 = ~n15736 & ~n15775 ;
  assign n15755 = ~n15719 & ~n15726 ;
  assign n15756 = ~n15712 & n15755 ;
  assign n15757 = n15706 & n15744 ;
  assign n15758 = ~n15756 & ~n15757 ;
  assign n15777 = n15736 & ~n15758 ;
  assign n15727 = n15706 & ~n15726 ;
  assign n15728 = n15719 & n15727 ;
  assign n15729 = n15712 & n15728 ;
  assign n15768 = ~n15706 & ~n15748 ;
  assign n15769 = n15712 & ~n15744 ;
  assign n15770 = n15768 & n15769 ;
  assign n15778 = ~n15729 & ~n15770 ;
  assign n15779 = ~n15777 & n15778 ;
  assign n15780 = ~n15776 & n15779 ;
  assign n15781 = ~n15743 & ~n15780 ;
  assign n15713 = ~n15706 & n15712 ;
  assign n15720 = n15713 & ~n15719 ;
  assign n15730 = ~n15720 & ~n15729 ;
  assign n15737 = ~n15730 & ~n15736 ;
  assign n15746 = ~n15719 & n15727 ;
  assign n15747 = n15712 & n15746 ;
  assign n15749 = ~n15706 & n15748 ;
  assign n15750 = n15719 & n15726 ;
  assign n15751 = n15706 & n15750 ;
  assign n15752 = ~n15749 & ~n15751 ;
  assign n15753 = ~n15747 & n15752 ;
  assign n15754 = n15736 & ~n15753 ;
  assign n15759 = ~n15736 & ~n15758 ;
  assign n15745 = n15713 & n15744 ;
  assign n15760 = ~n15706 & n15726 ;
  assign n15761 = ~n15736 & ~n15760 ;
  assign n15762 = ~n15712 & n15719 ;
  assign n15763 = ~n15761 & n15762 ;
  assign n15764 = ~n15745 & ~n15763 ;
  assign n15765 = ~n15759 & n15764 ;
  assign n15766 = ~n15754 & n15765 ;
  assign n15767 = n15743 & ~n15766 ;
  assign n15782 = ~n15737 & ~n15767 ;
  assign n15783 = ~n15781 & n15782 ;
  assign n15784 = ~\u2_L7_reg[28]/NET0131  & ~n15783 ;
  assign n15785 = \u2_L7_reg[28]/NET0131  & n15783 ;
  assign n15786 = ~n15784 & ~n15785 ;
  assign n15796 = n15074 & n15118 ;
  assign n15797 = ~n15074 & ~n15100 ;
  assign n15798 = ~n15103 & n15797 ;
  assign n15799 = ~n15796 & ~n15798 ;
  assign n15800 = ~n15062 & ~n15799 ;
  assign n15789 = ~n15124 & ~n15127 ;
  assign n15790 = n15074 & ~n15088 ;
  assign n15791 = ~n15086 & ~n15098 ;
  assign n15792 = ~n15790 & n15791 ;
  assign n15793 = n15789 & ~n15792 ;
  assign n15794 = n15062 & ~n15793 ;
  assign n15795 = n15074 & n15101 ;
  assign n15801 = ~n15056 & ~n15795 ;
  assign n15802 = ~n15794 & n15801 ;
  assign n15803 = ~n15800 & n15802 ;
  assign n15809 = ~n15074 & ~n15098 ;
  assign n15810 = ~n15081 & ~n15809 ;
  assign n15811 = n15062 & ~n15810 ;
  assign n15808 = n15112 & ~n15113 ;
  assign n15812 = ~n15798 & ~n15808 ;
  assign n15813 = ~n15811 & n15812 ;
  assign n15804 = n15074 & ~n15098 ;
  assign n15805 = n15088 & ~n15804 ;
  assign n15806 = ~n15796 & ~n15805 ;
  assign n15807 = n15062 & ~n15806 ;
  assign n15814 = n15056 & ~n15807 ;
  assign n15815 = ~n15813 & n15814 ;
  assign n15816 = ~n15803 & ~n15815 ;
  assign n15787 = n15062 & ~n15074 ;
  assign n15788 = n15126 & n15787 ;
  assign n15817 = ~n15125 & ~n15788 ;
  assign n15818 = ~n15816 & n15817 ;
  assign n15819 = \u2_L7_reg[29]/NET0131  & ~n15818 ;
  assign n15820 = ~\u2_L7_reg[29]/NET0131  & n15818 ;
  assign n15821 = ~n15819 & ~n15820 ;
  assign n15854 = ~n15727 & ~n15772 ;
  assign n15855 = ~n15712 & ~n15854 ;
  assign n15845 = n15712 & n15757 ;
  assign n15846 = ~n15706 & ~n15712 ;
  assign n15847 = n15726 & ~n15736 ;
  assign n15848 = n15846 & n15847 ;
  assign n15849 = ~n15845 & ~n15848 ;
  assign n15829 = n15712 & n15719 ;
  assign n15850 = ~n15760 & ~n15829 ;
  assign n15851 = ~n15706 & n15750 ;
  assign n15852 = ~n15736 & ~n15851 ;
  assign n15853 = ~n15850 & n15852 ;
  assign n15856 = n15849 & ~n15853 ;
  assign n15857 = ~n15855 & n15856 ;
  assign n15858 = ~n15743 & ~n15857 ;
  assign n15822 = ~n15712 & ~n15752 ;
  assign n15823 = n15706 & ~n15712 ;
  assign n15824 = ~n15771 & ~n15823 ;
  assign n15825 = n15736 & ~n15824 ;
  assign n15826 = ~n15822 & ~n15825 ;
  assign n15827 = n15743 & ~n15826 ;
  assign n15832 = n15713 & ~n15726 ;
  assign n15833 = ~n15719 & n15832 ;
  assign n15830 = n15760 & n15829 ;
  assign n15831 = ~n15743 & n15830 ;
  assign n15828 = ~n15712 & n15771 ;
  assign n15834 = n15736 & ~n15828 ;
  assign n15835 = ~n15831 & n15834 ;
  assign n15836 = ~n15833 & n15835 ;
  assign n15837 = n15755 & ~n15823 ;
  assign n15838 = ~n15830 & ~n15837 ;
  assign n15839 = n15743 & ~n15838 ;
  assign n15840 = ~n15713 & ~n15823 ;
  assign n15841 = n15744 & n15840 ;
  assign n15842 = ~n15736 & ~n15841 ;
  assign n15843 = ~n15839 & n15842 ;
  assign n15844 = ~n15836 & ~n15843 ;
  assign n15859 = ~n15827 & ~n15844 ;
  assign n15860 = ~n15858 & n15859 ;
  assign n15861 = \u2_L7_reg[2]/NET0131  & n15860 ;
  assign n15862 = ~\u2_L7_reg[2]/NET0131  & ~n15860 ;
  assign n15863 = ~n15861 & ~n15862 ;
  assign n15880 = n15074 & ~n15126 ;
  assign n15881 = ~n15115 & ~n15880 ;
  assign n15882 = n15111 & n15787 ;
  assign n15883 = n15056 & ~n15882 ;
  assign n15884 = ~n15881 & n15883 ;
  assign n15885 = ~n15118 & ~n15132 ;
  assign n15886 = ~n15099 & n15885 ;
  assign n15887 = n15062 & ~n15886 ;
  assign n15888 = ~n15056 & ~n15136 ;
  assign n15889 = ~n15125 & n15888 ;
  assign n15890 = ~n15887 & n15889 ;
  assign n15891 = ~n15884 & ~n15890 ;
  assign n15865 = ~n15114 & ~n15795 ;
  assign n15866 = ~n15056 & ~n15865 ;
  assign n15864 = ~n15068 & n15809 ;
  assign n15867 = n15081 & n15809 ;
  assign n15868 = ~n15075 & ~n15867 ;
  assign n15869 = n15056 & ~n15868 ;
  assign n15870 = ~n15864 & ~n15869 ;
  assign n15871 = ~n15866 & n15870 ;
  assign n15872 = ~n15062 & ~n15871 ;
  assign n15877 = ~n15062 & n15789 ;
  assign n15873 = n15088 & n15098 ;
  assign n15874 = ~n15122 & ~n15873 ;
  assign n15875 = n15062 & ~n15118 ;
  assign n15876 = n15874 & n15875 ;
  assign n15878 = n15074 & ~n15876 ;
  assign n15879 = ~n15877 & n15878 ;
  assign n15892 = ~n15872 & ~n15879 ;
  assign n15893 = ~n15891 & n15892 ;
  assign n15894 = ~\u2_L7_reg[4]/NET0131  & ~n15893 ;
  assign n15895 = \u2_L7_reg[4]/NET0131  & n15893 ;
  assign n15896 = ~n15894 & ~n15895 ;
  assign n15898 = ~n15832 & n15852 ;
  assign n15900 = ~n15726 & n15846 ;
  assign n15899 = n15712 & n15744 ;
  assign n15901 = n15736 & ~n15899 ;
  assign n15902 = ~n15900 & n15901 ;
  assign n15903 = ~n15898 & ~n15902 ;
  assign n15897 = n15706 & n15756 ;
  assign n15904 = n15743 & ~n15897 ;
  assign n15905 = n15849 & n15904 ;
  assign n15906 = ~n15903 & n15905 ;
  assign n15908 = n15744 & ~n15840 ;
  assign n15907 = n15748 & n15846 ;
  assign n15909 = ~n15736 & ~n15743 ;
  assign n15910 = ~n15746 & n15909 ;
  assign n15911 = ~n15907 & n15910 ;
  assign n15912 = ~n15908 & n15911 ;
  assign n15913 = ~n15906 & ~n15912 ;
  assign n15914 = ~n15712 & n15750 ;
  assign n15915 = n15706 & n15914 ;
  assign n15916 = ~n15729 & ~n15915 ;
  assign n15917 = ~n15913 & n15916 ;
  assign n15918 = ~n15728 & ~n15744 ;
  assign n15919 = ~n15768 & n15918 ;
  assign n15920 = ~n15712 & ~n15919 ;
  assign n15921 = ~n15727 & n15769 ;
  assign n15922 = n15736 & ~n15743 ;
  assign n15923 = ~n15921 & n15922 ;
  assign n15924 = ~n15920 & n15923 ;
  assign n15925 = ~n15917 & ~n15924 ;
  assign n15926 = ~\u2_L7_reg[13]/NET0131  & ~n15925 ;
  assign n15927 = \u2_L7_reg[13]/NET0131  & n15925 ;
  assign n15928 = ~n15926 & ~n15927 ;
  assign n15941 = n15068 & ~n15086 ;
  assign n15942 = ~n15114 & ~n15941 ;
  assign n15943 = n15062 & ~n15942 ;
  assign n15939 = n15074 & n15127 ;
  assign n15940 = ~n15062 & ~n15874 ;
  assign n15944 = ~n15939 & ~n15940 ;
  assign n15945 = ~n15943 & n15944 ;
  assign n15946 = ~n15056 & ~n15945 ;
  assign n15929 = ~n15087 & ~n15101 ;
  assign n15930 = n15062 & ~n15929 ;
  assign n15935 = ~n15867 & ~n15930 ;
  assign n15931 = ~n15062 & n15068 ;
  assign n15932 = ~n15132 & ~n15931 ;
  assign n15933 = ~n15081 & ~n15932 ;
  assign n15934 = n15074 & ~n15874 ;
  assign n15936 = ~n15933 & ~n15934 ;
  assign n15937 = n15935 & n15936 ;
  assign n15938 = n15056 & ~n15937 ;
  assign n15947 = ~n15121 & ~n15137 ;
  assign n15948 = ~n15938 & n15947 ;
  assign n15949 = ~n15946 & n15948 ;
  assign n15950 = ~\u2_L7_reg[19]/NET0131  & ~n15949 ;
  assign n15951 = \u2_L7_reg[19]/NET0131  & n15949 ;
  assign n15952 = ~n15950 & ~n15951 ;
  assign n15969 = ~n15004 & ~n15036 ;
  assign n15970 = ~n14963 & n15969 ;
  assign n15971 = ~n15005 & ~n15970 ;
  assign n15972 = n14990 & ~n15971 ;
  assign n15973 = n15020 & n15436 ;
  assign n15974 = ~n15037 & ~n15973 ;
  assign n15975 = ~n15433 & n15974 ;
  assign n15976 = ~n15972 & n15975 ;
  assign n15977 = ~n14976 & ~n15976 ;
  assign n15964 = n14976 & ~n15435 ;
  assign n15965 = n15001 & n15964 ;
  assign n15966 = ~n15035 & ~n15441 ;
  assign n15967 = ~n15965 & n15966 ;
  assign n15968 = n14990 & ~n15967 ;
  assign n15954 = n15026 & ~n15436 ;
  assign n15955 = ~n15034 & ~n15954 ;
  assign n15956 = ~n15004 & ~n15955 ;
  assign n15957 = n14991 & n15020 ;
  assign n15953 = ~n14982 & n15004 ;
  assign n15958 = ~n15440 & ~n15953 ;
  assign n15959 = ~n15957 & n15958 ;
  assign n15960 = ~n15956 & n15959 ;
  assign n15961 = ~n14990 & ~n15960 ;
  assign n15962 = ~n14970 & ~n15013 ;
  assign n15963 = n14983 & ~n15962 ;
  assign n15978 = ~n15961 & ~n15963 ;
  assign n15979 = ~n15968 & n15978 ;
  assign n15980 = ~n15977 & n15979 ;
  assign n15981 = \u2_L7_reg[23]/NET0131  & ~n15980 ;
  assign n15982 = ~\u2_L7_reg[23]/NET0131  & n15980 ;
  assign n15983 = ~n15981 & ~n15982 ;
  assign n15984 = ~n15246 & n15598 ;
  assign n15985 = ~n15607 & ~n15984 ;
  assign n15986 = ~n15276 & ~n15985 ;
  assign n15988 = ~n15253 & n15276 ;
  assign n15989 = n15401 & n15988 ;
  assign n15987 = n15252 & n15319 ;
  assign n15990 = ~n15267 & ~n15321 ;
  assign n15991 = ~n15987 & n15990 ;
  assign n15992 = ~n15989 & n15991 ;
  assign n15993 = ~n15986 & n15992 ;
  assign n15994 = n15299 & ~n15993 ;
  assign n15997 = n15252 & ~n15304 ;
  assign n15996 = n15288 & ~n15409 ;
  assign n15998 = n15276 & ~n15996 ;
  assign n15999 = ~n15997 & n15998 ;
  assign n15995 = n15279 & n15314 ;
  assign n16000 = ~n15597 & ~n15995 ;
  assign n16001 = ~n15309 & n16000 ;
  assign n16002 = ~n15999 & n16001 ;
  assign n16003 = ~n15299 & ~n16002 ;
  assign n16006 = ~n15276 & n15307 ;
  assign n16004 = ~n15252 & n15276 ;
  assign n16005 = n15266 & n16004 ;
  assign n16007 = ~n15313 & ~n16005 ;
  assign n16008 = ~n16006 & n16007 ;
  assign n16009 = ~n16003 & n16008 ;
  assign n16010 = ~n15994 & n16009 ;
  assign n16011 = ~\u2_L7_reg[27]/NET0131  & ~n16010 ;
  assign n16012 = \u2_L7_reg[27]/NET0131  & n16010 ;
  assign n16013 = ~n16011 & ~n16012 ;
  assign n16031 = ~n14898 & ~n14942 ;
  assign n16032 = ~n14882 & n15377 ;
  assign n16033 = ~n16031 & ~n16032 ;
  assign n16018 = ~n14882 & n14941 ;
  assign n16034 = n14876 & n16018 ;
  assign n16035 = ~n16033 & ~n16034 ;
  assign n16036 = ~n14921 & ~n16035 ;
  assign n16037 = n14876 & n15369 ;
  assign n16038 = ~n14882 & ~n14921 ;
  assign n16039 = n16037 & ~n16038 ;
  assign n16040 = ~n14882 & n14898 ;
  assign n16041 = ~n14904 & ~n16040 ;
  assign n16042 = n14921 & ~n16041 ;
  assign n16043 = ~n16039 & ~n16042 ;
  assign n16044 = ~n16036 & n16043 ;
  assign n16045 = n14911 & ~n16044 ;
  assign n16014 = ~n14876 & n15369 ;
  assign n16015 = ~n14902 & ~n14903 ;
  assign n16016 = ~n16014 & ~n16015 ;
  assign n16017 = ~n14921 & ~n16016 ;
  assign n16019 = n14921 & ~n16014 ;
  assign n16020 = ~n16018 & n16019 ;
  assign n16021 = ~n16017 & ~n16020 ;
  assign n16022 = n14882 & n16014 ;
  assign n16023 = n14903 & n14930 ;
  assign n16024 = ~n16022 & ~n16023 ;
  assign n16025 = n14901 & n16024 ;
  assign n16026 = ~n16021 & n16025 ;
  assign n16027 = ~n14911 & ~n16026 ;
  assign n16028 = n14897 & n14921 ;
  assign n16029 = n14939 & ~n15369 ;
  assign n16030 = n14931 & n16029 ;
  assign n16046 = ~n16028 & ~n16030 ;
  assign n16047 = ~n16027 & n16046 ;
  assign n16048 = ~n16045 & n16047 ;
  assign n16049 = \u2_L7_reg[32]/NET0131  & n16048 ;
  assign n16050 = ~\u2_L7_reg[32]/NET0131  & ~n16048 ;
  assign n16051 = ~n16049 & ~n16050 ;
  assign n16052 = decrypt_pad & ~\u2_uk_K_r7_reg[26]/NET0131  ;
  assign n16053 = ~decrypt_pad & ~\u2_uk_K_r7_reg[33]/NET0131  ;
  assign n16054 = ~n16052 & ~n16053 ;
  assign n16055 = \u2_R7_reg[12]/NET0131  & ~n16054 ;
  assign n16056 = ~\u2_R7_reg[12]/NET0131  & n16054 ;
  assign n16057 = ~n16055 & ~n16056 ;
  assign n16064 = decrypt_pad & ~\u2_uk_K_r7_reg[11]/NET0131  ;
  assign n16065 = ~decrypt_pad & ~\u2_uk_K_r7_reg[18]/NET0131  ;
  assign n16066 = ~n16064 & ~n16065 ;
  assign n16067 = \u2_R7_reg[11]/NET0131  & ~n16066 ;
  assign n16068 = ~\u2_R7_reg[11]/NET0131  & n16066 ;
  assign n16069 = ~n16067 & ~n16068 ;
  assign n16080 = decrypt_pad & ~\u2_uk_K_r7_reg[34]/NET0131  ;
  assign n16081 = ~decrypt_pad & ~\u2_uk_K_r7_reg[41]/NET0131  ;
  assign n16082 = ~n16080 & ~n16081 ;
  assign n16083 = \u2_R7_reg[9]/NET0131  & ~n16082 ;
  assign n16084 = ~\u2_R7_reg[9]/NET0131  & n16082 ;
  assign n16085 = ~n16083 & ~n16084 ;
  assign n16086 = decrypt_pad & ~\u2_uk_K_r7_reg[10]/NET0131  ;
  assign n16087 = ~decrypt_pad & ~\u2_uk_K_r7_reg[17]/NET0131  ;
  assign n16088 = ~n16086 & ~n16087 ;
  assign n16089 = \u2_R7_reg[10]/NET0131  & ~n16088 ;
  assign n16090 = ~\u2_R7_reg[10]/NET0131  & n16088 ;
  assign n16091 = ~n16089 & ~n16090 ;
  assign n16058 = decrypt_pad & ~\u2_uk_K_r7_reg[5]/NET0131  ;
  assign n16059 = ~decrypt_pad & ~\u2_uk_K_r7_reg[12]/NET0131  ;
  assign n16060 = ~n16058 & ~n16059 ;
  assign n16061 = \u2_R7_reg[8]/NET0131  & ~n16060 ;
  assign n16062 = ~\u2_R7_reg[8]/NET0131  & n16060 ;
  assign n16063 = ~n16061 & ~n16062 ;
  assign n16071 = decrypt_pad & ~\u2_uk_K_r7_reg[39]/NET0131  ;
  assign n16072 = ~decrypt_pad & ~\u2_uk_K_r7_reg[46]/NET0131  ;
  assign n16073 = ~n16071 & ~n16072 ;
  assign n16074 = \u2_R7_reg[13]/NET0131  & ~n16073 ;
  assign n16075 = ~\u2_R7_reg[13]/NET0131  & n16073 ;
  assign n16076 = ~n16074 & ~n16075 ;
  assign n16098 = ~n16063 & n16076 ;
  assign n16099 = n16091 & n16098 ;
  assign n16100 = n16085 & n16099 ;
  assign n16101 = ~n16069 & n16100 ;
  assign n16095 = n16085 & n16091 ;
  assign n16077 = ~n16063 & ~n16076 ;
  assign n16078 = n16063 & n16076 ;
  assign n16079 = ~n16077 & ~n16078 ;
  assign n16092 = ~n16085 & ~n16091 ;
  assign n16096 = ~n16079 & ~n16092 ;
  assign n16097 = ~n16095 & n16096 ;
  assign n16070 = ~n16063 & n16069 ;
  assign n16093 = ~n16070 & n16092 ;
  assign n16094 = n16079 & n16093 ;
  assign n16102 = ~n16063 & n16085 ;
  assign n16103 = n16069 & ~n16091 ;
  assign n16104 = n16102 & n16103 ;
  assign n16105 = ~n16076 & n16085 ;
  assign n16106 = n16063 & n16091 ;
  assign n16107 = n16105 & n16106 ;
  assign n16108 = ~n16104 & ~n16107 ;
  assign n16109 = ~n16094 & n16108 ;
  assign n16110 = ~n16097 & n16109 ;
  assign n16111 = ~n16101 & n16110 ;
  assign n16112 = ~n16057 & ~n16111 ;
  assign n16113 = n16057 & n16091 ;
  assign n16114 = ~n16063 & n16105 ;
  assign n16115 = n16113 & n16114 ;
  assign n16116 = n16076 & ~n16085 ;
  assign n16117 = n16063 & n16105 ;
  assign n16118 = ~n16099 & ~n16117 ;
  assign n16119 = ~n16116 & n16118 ;
  assign n16120 = n16057 & n16069 ;
  assign n16121 = ~n16119 & n16120 ;
  assign n16136 = ~n16115 & ~n16121 ;
  assign n16122 = n16091 & n16116 ;
  assign n16123 = n16077 & ~n16091 ;
  assign n16124 = ~n16085 & n16123 ;
  assign n16125 = ~n16122 & ~n16124 ;
  assign n16126 = n16069 & ~n16125 ;
  assign n16127 = n16057 & ~n16069 ;
  assign n16132 = n16078 & n16085 ;
  assign n16128 = n16085 & ~n16091 ;
  assign n16129 = n16076 & n16128 ;
  assign n16130 = n16063 & ~n16085 ;
  assign n16131 = ~n16076 & n16130 ;
  assign n16133 = ~n16129 & ~n16131 ;
  assign n16134 = ~n16132 & n16133 ;
  assign n16135 = n16127 & ~n16134 ;
  assign n16137 = ~n16126 & ~n16135 ;
  assign n16138 = n16136 & n16137 ;
  assign n16139 = ~n16112 & n16138 ;
  assign n16140 = ~\u2_L7_reg[6]/NET0131  & ~n16139 ;
  assign n16141 = \u2_L7_reg[6]/NET0131  & n16139 ;
  assign n16142 = ~n16140 & ~n16141 ;
  assign n16143 = n14882 & ~n15377 ;
  assign n16144 = ~n16018 & ~n16143 ;
  assign n16145 = n14876 & ~n16144 ;
  assign n16146 = ~n14876 & ~n14902 ;
  assign n16147 = n15377 & n16146 ;
  assign n16148 = n14921 & ~n16147 ;
  assign n16149 = ~n14889 & ~n15379 ;
  assign n16150 = ~n14921 & ~n16037 ;
  assign n16151 = ~n16143 & n16150 ;
  assign n16152 = ~n16149 & n16151 ;
  assign n16153 = ~n16148 & ~n16152 ;
  assign n16154 = ~n16145 & ~n16153 ;
  assign n16155 = n14911 & ~n16154 ;
  assign n16163 = ~n14921 & n16147 ;
  assign n16164 = ~n14933 & ~n16163 ;
  assign n16165 = ~n14911 & ~n16164 ;
  assign n16157 = ~n15371 & ~n15377 ;
  assign n16158 = ~n14899 & ~n16023 ;
  assign n16159 = ~n16157 & n16158 ;
  assign n16156 = n14911 & ~n14933 ;
  assign n16160 = n14921 & ~n16156 ;
  assign n16161 = ~n16159 & n16160 ;
  assign n16162 = ~n14921 & n16145 ;
  assign n16166 = ~n16161 & ~n16162 ;
  assign n16167 = ~n16165 & n16166 ;
  assign n16168 = ~n16155 & n16167 ;
  assign n16169 = ~\u2_L7_reg[7]/NET0131  & ~n16168 ;
  assign n16170 = \u2_L7_reg[7]/NET0131  & n16168 ;
  assign n16171 = ~n16169 & ~n16170 ;
  assign n16183 = ~n15509 & ~n15632 ;
  assign n16184 = n15470 & ~n16183 ;
  assign n16185 = n15506 & ~n15531 ;
  assign n16186 = ~n15638 & ~n16185 ;
  assign n16187 = ~n15470 & ~n16186 ;
  assign n16188 = ~n15490 & n15657 ;
  assign n16189 = ~n16187 & n16188 ;
  assign n16190 = ~n16184 & n16189 ;
  assign n16191 = ~n15529 & ~n16190 ;
  assign n16176 = ~n15476 & n15539 ;
  assign n16177 = ~n15638 & ~n16176 ;
  assign n16178 = n15470 & ~n16177 ;
  assign n16179 = ~n15476 & n15661 ;
  assign n16180 = n15556 & ~n16179 ;
  assign n16181 = ~n16178 & n16180 ;
  assign n16182 = n15529 & ~n16181 ;
  assign n16172 = n15506 & ~n15532 ;
  assign n16173 = ~n15505 & ~n16172 ;
  assign n16174 = n15470 & ~n16173 ;
  assign n16175 = n15476 & n15646 ;
  assign n16192 = ~n16174 & ~n16175 ;
  assign n16193 = ~n16182 & n16192 ;
  assign n16194 = ~n16191 & n16193 ;
  assign n16195 = ~\u2_L7_reg[8]/NET0131  & ~n16194 ;
  assign n16196 = \u2_L7_reg[8]/NET0131  & n16194 ;
  assign n16197 = ~n16195 & ~n16196 ;
  assign n16206 = n16069 & n16114 ;
  assign n16204 = n16076 & ~n16102 ;
  assign n16205 = ~n16130 & n16204 ;
  assign n16207 = ~n16131 & ~n16205 ;
  assign n16208 = ~n16206 & n16207 ;
  assign n16209 = ~n16091 & ~n16208 ;
  assign n16198 = n16077 & n16091 ;
  assign n16210 = n16063 & ~n16091 ;
  assign n16211 = ~n16076 & n16210 ;
  assign n16212 = ~n16198 & ~n16211 ;
  assign n16213 = ~n16069 & ~n16212 ;
  assign n16214 = n16057 & ~n16100 ;
  assign n16215 = ~n16213 & n16214 ;
  assign n16216 = ~n16209 & n16215 ;
  assign n16217 = n16076 & n16130 ;
  assign n16218 = n16069 & ~n16217 ;
  assign n16219 = ~n16078 & n16085 ;
  assign n16220 = ~n16077 & n16219 ;
  assign n16221 = n16218 & ~n16220 ;
  assign n16222 = ~n16069 & ~n16123 ;
  assign n16223 = ~n16205 & n16222 ;
  assign n16224 = ~n16221 & ~n16223 ;
  assign n16225 = ~n16057 & ~n16124 ;
  assign n16226 = ~n16224 & n16225 ;
  assign n16227 = ~n16216 & ~n16226 ;
  assign n16199 = ~n16085 & n16198 ;
  assign n16200 = ~n16107 & ~n16199 ;
  assign n16201 = n16069 & ~n16200 ;
  assign n16202 = ~n16069 & n16091 ;
  assign n16203 = n16130 & n16202 ;
  assign n16228 = ~n16201 & ~n16203 ;
  assign n16229 = ~n16227 & n16228 ;
  assign n16230 = ~\u2_L7_reg[16]/NET0131  & ~n16229 ;
  assign n16231 = \u2_L7_reg[16]/NET0131  & n16229 ;
  assign n16232 = ~n16230 & ~n16231 ;
  assign n16243 = ~n16079 & n16092 ;
  assign n16244 = n16118 & ~n16243 ;
  assign n16245 = ~n16069 & ~n16244 ;
  assign n16246 = ~n16057 & ~n16245 ;
  assign n16249 = ~n16069 & n16096 ;
  assign n16253 = n16057 & ~n16094 ;
  assign n16247 = ~n16085 & ~n16098 ;
  assign n16248 = n16103 & n16247 ;
  assign n16250 = n16069 & n16091 ;
  assign n16251 = ~n16077 & n16250 ;
  assign n16252 = ~n16130 & n16251 ;
  assign n16254 = ~n16248 & ~n16252 ;
  assign n16255 = n16253 & n16254 ;
  assign n16256 = ~n16249 & n16255 ;
  assign n16257 = ~n16246 & ~n16256 ;
  assign n16234 = ~n16091 & n16098 ;
  assign n16235 = ~n16198 & ~n16234 ;
  assign n16236 = n16091 & n16130 ;
  assign n16237 = ~n16114 & ~n16236 ;
  assign n16238 = n16235 & n16237 ;
  assign n16239 = n16069 & ~n16238 ;
  assign n16240 = n16091 & n16131 ;
  assign n16241 = ~n16239 & ~n16240 ;
  assign n16242 = ~n16057 & ~n16241 ;
  assign n16259 = n16070 & n16129 ;
  assign n16233 = n16103 & n16131 ;
  assign n16258 = n16132 & n16202 ;
  assign n16260 = ~n16233 & ~n16258 ;
  assign n16261 = ~n16259 & n16260 ;
  assign n16262 = ~n16242 & n16261 ;
  assign n16263 = ~n16257 & n16262 ;
  assign n16264 = ~\u2_L7_reg[24]/NET0131  & ~n16263 ;
  assign n16265 = \u2_L7_reg[24]/NET0131  & n16263 ;
  assign n16266 = ~n16264 & ~n16265 ;
  assign n16267 = ~n16105 & n16106 ;
  assign n16268 = ~n16076 & n16128 ;
  assign n16269 = ~n16267 & ~n16268 ;
  assign n16270 = n16069 & ~n16269 ;
  assign n16274 = ~n16063 & n16122 ;
  assign n16271 = ~n16102 & ~n16210 ;
  assign n16272 = ~n16069 & ~n16105 ;
  assign n16273 = ~n16271 & n16272 ;
  assign n16275 = ~n16243 & ~n16273 ;
  assign n16276 = ~n16274 & n16275 ;
  assign n16277 = ~n16270 & n16276 ;
  assign n16278 = ~n16057 & ~n16277 ;
  assign n16279 = n16069 & ~n16235 ;
  assign n16280 = ~n16233 & ~n16279 ;
  assign n16281 = n16057 & ~n16280 ;
  assign n16285 = n16091 & ~n16272 ;
  assign n16286 = ~n16218 & n16285 ;
  assign n16282 = ~n16106 & ~n16114 ;
  assign n16283 = n16127 & ~n16282 ;
  assign n16284 = n16113 & n16219 ;
  assign n16287 = ~n16283 & ~n16284 ;
  assign n16288 = ~n16286 & n16287 ;
  assign n16289 = ~n16281 & n16288 ;
  assign n16290 = ~n16278 & n16289 ;
  assign n16291 = \u2_L7_reg[30]/NET0131  & ~n16290 ;
  assign n16292 = ~\u2_L7_reg[30]/NET0131  & n16290 ;
  assign n16293 = ~n16291 & ~n16292 ;
  assign n16297 = ~n15476 & n15506 ;
  assign n16298 = ~n15535 & ~n16297 ;
  assign n16299 = n15470 & ~n16298 ;
  assign n16294 = n15470 & ~n15531 ;
  assign n16295 = ~n15517 & ~n15638 ;
  assign n16296 = ~n16294 & ~n16295 ;
  assign n16300 = ~n15529 & ~n16296 ;
  assign n16301 = ~n16299 & n16300 ;
  assign n16304 = n15489 & ~n15516 ;
  assign n16303 = ~n15489 & ~n15500 ;
  assign n16305 = n15470 & ~n16303 ;
  assign n16306 = ~n16304 & n16305 ;
  assign n16307 = ~n15470 & n15538 ;
  assign n16302 = n15476 & n15508 ;
  assign n16308 = ~n15511 & n15529 ;
  assign n16309 = ~n16302 & n16308 ;
  assign n16310 = ~n16307 & n16309 ;
  assign n16311 = ~n16306 & n16310 ;
  assign n16312 = ~n16301 & ~n16311 ;
  assign n16313 = n15510 & n15531 ;
  assign n16314 = ~n15470 & ~n16313 ;
  assign n16315 = ~n15551 & n16314 ;
  assign n16316 = ~n16176 & n16315 ;
  assign n16317 = n15470 & ~n15509 ;
  assign n16318 = ~n15554 & n16317 ;
  assign n16319 = ~n16316 & ~n16318 ;
  assign n16320 = ~n16312 & ~n16319 ;
  assign n16321 = ~\u2_L7_reg[3]/NET0131  & ~n16320 ;
  assign n16322 = \u2_L7_reg[3]/NET0131  & n16320 ;
  assign n16323 = ~n16321 & ~n16322 ;
  assign n16327 = n14969 & n15435 ;
  assign n16330 = n14997 & n16327 ;
  assign n16324 = ~n15000 & n15025 ;
  assign n16331 = ~n14990 & ~n16324 ;
  assign n16332 = ~n16330 & n16331 ;
  assign n16325 = ~n14998 & ~n15969 ;
  assign n16326 = ~n14976 & n16325 ;
  assign n16328 = n14976 & n15969 ;
  assign n16329 = ~n16327 & n16328 ;
  assign n16333 = ~n16326 & ~n16329 ;
  assign n16334 = n16332 & n16333 ;
  assign n16336 = n14982 & ~n15001 ;
  assign n16337 = ~n15451 & n16336 ;
  assign n16335 = n14983 & n16325 ;
  assign n16338 = n15434 & ~n16335 ;
  assign n16339 = ~n16337 & n16338 ;
  assign n16340 = ~n16334 & ~n16339 ;
  assign n16341 = ~n14976 & ~n15003 ;
  assign n16342 = ~n15007 & n15036 ;
  assign n16343 = n16341 & n16342 ;
  assign n16344 = ~n16340 & ~n16343 ;
  assign n16345 = ~\u2_L7_reg[9]/NET0131  & ~n16344 ;
  assign n16346 = \u2_L7_reg[9]/NET0131  & n16344 ;
  assign n16347 = ~n16345 & ~n16346 ;
  assign n16350 = n15736 & ~n15854 ;
  assign n16348 = ~n15749 & ~n15914 ;
  assign n16349 = ~n15736 & ~n16348 ;
  assign n16351 = ~n15833 & ~n16349 ;
  assign n16352 = ~n16350 & n16351 ;
  assign n16353 = n15743 & ~n16352 ;
  assign n16358 = ~n15830 & ~n15900 ;
  assign n16359 = ~n15729 & n16358 ;
  assign n16354 = n15736 & n15751 ;
  assign n16355 = n15712 & n15736 ;
  assign n16356 = ~n15719 & ~n16355 ;
  assign n16357 = n15840 & n16356 ;
  assign n16360 = ~n16354 & ~n16357 ;
  assign n16361 = n16359 & n16360 ;
  assign n16362 = ~n15743 & ~n16361 ;
  assign n16363 = ~n15736 & n15757 ;
  assign n16364 = n15712 & n15750 ;
  assign n16365 = ~n15897 & ~n16364 ;
  assign n16366 = n15736 & ~n16365 ;
  assign n16367 = ~n16363 & ~n16366 ;
  assign n16368 = ~n16362 & n16367 ;
  assign n16369 = ~n16353 & n16368 ;
  assign n16370 = ~\u2_L7_reg[18]/P0001  & ~n16369 ;
  assign n16371 = \u2_L7_reg[18]/P0001  & n16369 ;
  assign n16372 = ~n16370 & ~n16371 ;
  assign n16373 = decrypt_pad & ~\u2_uk_K_r6_reg[54]/NET0131  ;
  assign n16374 = ~decrypt_pad & ~\u2_uk_K_r6_reg[47]/NET0131  ;
  assign n16375 = ~n16373 & ~n16374 ;
  assign n16376 = \u2_R6_reg[4]/NET0131  & ~n16375 ;
  assign n16377 = ~\u2_R6_reg[4]/NET0131  & n16375 ;
  assign n16378 = ~n16376 & ~n16377 ;
  assign n16406 = decrypt_pad & ~\u2_uk_K_r6_reg[19]/NET0131  ;
  assign n16407 = ~decrypt_pad & ~\u2_uk_K_r6_reg[12]/NET0131  ;
  assign n16408 = ~n16406 & ~n16407 ;
  assign n16409 = \u2_R6_reg[3]/NET0131  & ~n16408 ;
  assign n16410 = ~\u2_R6_reg[3]/NET0131  & n16408 ;
  assign n16411 = ~n16409 & ~n16410 ;
  assign n16379 = decrypt_pad & ~\u2_uk_K_r6_reg[10]/NET0131  ;
  assign n16380 = ~decrypt_pad & ~\u2_uk_K_r6_reg[3]/NET0131  ;
  assign n16381 = ~n16379 & ~n16380 ;
  assign n16382 = \u2_R6_reg[2]/NET0131  & ~n16381 ;
  assign n16383 = ~\u2_R6_reg[2]/NET0131  & n16381 ;
  assign n16384 = ~n16382 & ~n16383 ;
  assign n16392 = decrypt_pad & ~\u2_uk_K_r6_reg[25]/NET0131  ;
  assign n16393 = ~decrypt_pad & ~\u2_uk_K_r6_reg[18]/NET0131  ;
  assign n16394 = ~n16392 & ~n16393 ;
  assign n16395 = \u2_R6_reg[5]/NET0131  & ~n16394 ;
  assign n16396 = ~\u2_R6_reg[5]/NET0131  & n16394 ;
  assign n16397 = ~n16395 & ~n16396 ;
  assign n16385 = decrypt_pad & ~\u2_uk_K_r6_reg[27]/NET0131  ;
  assign n16386 = ~decrypt_pad & ~\u2_uk_K_r6_reg[20]/NET0131  ;
  assign n16387 = ~n16385 & ~n16386 ;
  assign n16388 = \u2_R6_reg[1]/NET0131  & ~n16387 ;
  assign n16389 = ~\u2_R6_reg[1]/NET0131  & n16387 ;
  assign n16390 = ~n16388 & ~n16389 ;
  assign n16399 = decrypt_pad & ~\u2_uk_K_r6_reg[6]/NET0131  ;
  assign n16400 = ~decrypt_pad & ~\u2_uk_K_r6_reg[24]/NET0131  ;
  assign n16401 = ~n16399 & ~n16400 ;
  assign n16402 = \u2_R6_reg[32]/NET0131  & ~n16401 ;
  assign n16403 = ~\u2_R6_reg[32]/NET0131  & n16401 ;
  assign n16404 = ~n16402 & ~n16403 ;
  assign n16413 = ~n16390 & n16404 ;
  assign n16414 = ~n16397 & n16413 ;
  assign n16415 = n16384 & n16414 ;
  assign n16416 = ~n16384 & ~n16404 ;
  assign n16417 = ~n16390 & n16397 ;
  assign n16418 = n16416 & ~n16417 ;
  assign n16419 = ~n16415 & ~n16418 ;
  assign n16420 = ~n16411 & ~n16419 ;
  assign n16421 = n16397 & ~n16404 ;
  assign n16422 = n16384 & n16411 ;
  assign n16423 = n16421 & n16422 ;
  assign n16424 = ~n16397 & n16416 ;
  assign n16425 = ~n16423 & ~n16424 ;
  assign n16426 = n16390 & ~n16425 ;
  assign n16391 = n16384 & n16390 ;
  assign n16398 = n16391 & ~n16397 ;
  assign n16405 = n16398 & n16404 ;
  assign n16412 = n16405 & n16411 ;
  assign n16427 = n16397 & n16404 ;
  assign n16428 = ~n16384 & n16411 ;
  assign n16429 = ~n16384 & ~n16390 ;
  assign n16430 = ~n16428 & ~n16429 ;
  assign n16431 = n16427 & ~n16430 ;
  assign n16432 = ~n16412 & ~n16431 ;
  assign n16433 = ~n16426 & n16432 ;
  assign n16434 = ~n16420 & n16433 ;
  assign n16435 = ~n16378 & ~n16434 ;
  assign n16443 = ~n16384 & ~n16397 ;
  assign n16444 = n16404 & ~n16443 ;
  assign n16445 = ~n16390 & ~n16424 ;
  assign n16446 = ~n16444 & n16445 ;
  assign n16437 = n16384 & ~n16404 ;
  assign n16438 = ~n16397 & n16437 ;
  assign n16439 = ~n16417 & ~n16438 ;
  assign n16440 = n16411 & ~n16439 ;
  assign n16436 = n16421 & n16428 ;
  assign n16441 = n16390 & n16404 ;
  assign n16442 = ~n16411 & n16441 ;
  assign n16447 = ~n16436 & ~n16442 ;
  assign n16448 = ~n16440 & n16447 ;
  assign n16449 = ~n16446 & n16448 ;
  assign n16450 = n16378 & ~n16449 ;
  assign n16451 = ~n16390 & n16411 ;
  assign n16452 = ~n16384 & n16404 ;
  assign n16453 = ~n16438 & ~n16452 ;
  assign n16454 = n16451 & ~n16453 ;
  assign n16457 = n16391 & n16397 ;
  assign n16458 = n16404 & n16457 ;
  assign n16455 = n16390 & n16443 ;
  assign n16456 = n16417 & n16437 ;
  assign n16459 = ~n16455 & ~n16456 ;
  assign n16460 = ~n16458 & n16459 ;
  assign n16461 = ~n16411 & ~n16460 ;
  assign n16462 = ~n16454 & ~n16461 ;
  assign n16463 = ~n16450 & n16462 ;
  assign n16464 = ~n16435 & n16463 ;
  assign n16465 = ~\u2_L6_reg[31]/NET0131  & ~n16464 ;
  assign n16466 = \u2_L6_reg[31]/NET0131  & n16464 ;
  assign n16467 = ~n16465 & ~n16466 ;
  assign n16474 = decrypt_pad & ~\u2_uk_K_r6_reg[21]/NET0131  ;
  assign n16475 = ~decrypt_pad & ~\u2_uk_K_r6_reg[14]/NET0131  ;
  assign n16476 = ~n16474 & ~n16475 ;
  assign n16477 = \u2_R6_reg[23]/NET0131  & ~n16476 ;
  assign n16478 = ~\u2_R6_reg[23]/NET0131  & n16476 ;
  assign n16479 = ~n16477 & ~n16478 ;
  assign n16480 = decrypt_pad & ~\u2_uk_K_r6_reg[8]/NET0131  ;
  assign n16481 = ~decrypt_pad & ~\u2_uk_K_r6_reg[1]/NET0131  ;
  assign n16482 = ~n16480 & ~n16481 ;
  assign n16483 = \u2_R6_reg[22]/NET0131  & ~n16482 ;
  assign n16484 = ~\u2_R6_reg[22]/NET0131  & n16482 ;
  assign n16485 = ~n16483 & ~n16484 ;
  assign n16487 = decrypt_pad & ~\u2_uk_K_r6_reg[2]/NET0131  ;
  assign n16488 = ~decrypt_pad & ~\u2_uk_K_r6_reg[50]/NET0131  ;
  assign n16489 = ~n16487 & ~n16488 ;
  assign n16490 = \u2_R6_reg[20]/NET0131  & ~n16489 ;
  assign n16491 = ~\u2_R6_reg[20]/NET0131  & n16489 ;
  assign n16492 = ~n16490 & ~n16491 ;
  assign n16506 = decrypt_pad & ~\u2_uk_K_r6_reg[42]/NET0131  ;
  assign n16507 = ~decrypt_pad & ~\u2_uk_K_r6_reg[35]/NET0131  ;
  assign n16508 = ~n16506 & ~n16507 ;
  assign n16509 = \u2_R6_reg[25]/NET0131  & ~n16508 ;
  assign n16510 = ~\u2_R6_reg[25]/NET0131  & n16508 ;
  assign n16511 = ~n16509 & ~n16510 ;
  assign n16512 = n16492 & ~n16511 ;
  assign n16494 = decrypt_pad & ~\u2_uk_K_r6_reg[45]/NET0131  ;
  assign n16495 = ~decrypt_pad & ~\u2_uk_K_r6_reg[38]/NET0131  ;
  assign n16496 = ~n16494 & ~n16495 ;
  assign n16497 = \u2_R6_reg[21]/NET0131  & ~n16496 ;
  assign n16498 = ~\u2_R6_reg[21]/NET0131  & n16496 ;
  assign n16499 = ~n16497 & ~n16498 ;
  assign n16521 = ~n16492 & ~n16499 ;
  assign n16549 = ~n16512 & ~n16521 ;
  assign n16550 = n16485 & n16549 ;
  assign n16551 = n16499 & n16511 ;
  assign n16552 = ~n16492 & n16551 ;
  assign n16518 = n16492 & n16511 ;
  assign n16519 = ~n16499 & n16518 ;
  assign n16553 = ~n16485 & ~n16519 ;
  assign n16554 = ~n16552 & n16553 ;
  assign n16555 = ~n16550 & ~n16554 ;
  assign n16556 = ~n16479 & ~n16555 ;
  assign n16468 = decrypt_pad & ~\u2_uk_K_r6_reg[23]/P0001  ;
  assign n16469 = ~decrypt_pad & ~\u2_uk_K_r6_reg[16]/NET0131  ;
  assign n16470 = ~n16468 & ~n16469 ;
  assign n16471 = \u2_R6_reg[24]/NET0131  & ~n16470 ;
  assign n16472 = ~\u2_R6_reg[24]/NET0131  & n16470 ;
  assign n16473 = ~n16471 & ~n16472 ;
  assign n16500 = n16485 & ~n16492 ;
  assign n16501 = n16499 & n16500 ;
  assign n16546 = n16479 & ~n16501 ;
  assign n16543 = ~n16485 & ~n16499 ;
  assign n16544 = n16512 & n16543 ;
  assign n16545 = n16499 & n16518 ;
  assign n16547 = ~n16544 & ~n16545 ;
  assign n16548 = n16546 & n16547 ;
  assign n16557 = n16473 & ~n16548 ;
  assign n16558 = ~n16556 & n16557 ;
  assign n16502 = ~n16485 & n16499 ;
  assign n16524 = n16502 & ~n16511 ;
  assign n16525 = n16492 & n16524 ;
  assign n16520 = n16485 & n16519 ;
  assign n16522 = n16511 & n16521 ;
  assign n16523 = n16479 & n16522 ;
  assign n16528 = ~n16520 & ~n16523 ;
  assign n16529 = ~n16525 & n16528 ;
  assign n16503 = n16492 & n16502 ;
  assign n16504 = ~n16501 & ~n16503 ;
  assign n16505 = ~n16479 & ~n16504 ;
  assign n16515 = n16492 & ~n16499 ;
  assign n16516 = n16479 & n16485 ;
  assign n16517 = n16515 & n16516 ;
  assign n16486 = n16479 & ~n16485 ;
  assign n16493 = n16486 & ~n16492 ;
  assign n16513 = ~n16479 & ~n16485 ;
  assign n16514 = n16512 & n16513 ;
  assign n16526 = ~n16493 & ~n16514 ;
  assign n16527 = ~n16517 & n16526 ;
  assign n16530 = ~n16505 & n16527 ;
  assign n16531 = n16529 & n16530 ;
  assign n16532 = ~n16473 & ~n16531 ;
  assign n16537 = n16499 & n16512 ;
  assign n16538 = ~n16479 & n16537 ;
  assign n16539 = ~n16523 & ~n16538 ;
  assign n16540 = ~n16485 & ~n16539 ;
  assign n16533 = n16485 & n16518 ;
  assign n16534 = ~n16492 & n16524 ;
  assign n16535 = ~n16533 & ~n16534 ;
  assign n16536 = n16479 & ~n16535 ;
  assign n16541 = ~n16511 & n16521 ;
  assign n16542 = n16513 & n16541 ;
  assign n16559 = ~n16536 & ~n16542 ;
  assign n16560 = ~n16540 & n16559 ;
  assign n16561 = ~n16532 & n16560 ;
  assign n16562 = ~n16558 & n16561 ;
  assign n16563 = \u2_L6_reg[11]/NET0131  & ~n16562 ;
  assign n16564 = ~\u2_L6_reg[11]/NET0131  & n16562 ;
  assign n16565 = ~n16563 & ~n16564 ;
  assign n16578 = decrypt_pad & ~\u2_uk_K_r6_reg[14]/NET0131  ;
  assign n16579 = ~decrypt_pad & ~\u2_uk_K_r6_reg[7]/NET0131  ;
  assign n16580 = ~n16578 & ~n16579 ;
  assign n16581 = \u2_R6_reg[24]/NET0131  & ~n16580 ;
  assign n16582 = ~\u2_R6_reg[24]/NET0131  & n16580 ;
  assign n16583 = ~n16581 & ~n16582 ;
  assign n16601 = decrypt_pad & ~\u2_uk_K_r6_reg[43]/NET0131  ;
  assign n16602 = ~decrypt_pad & ~\u2_uk_K_r6_reg[36]/NET0131  ;
  assign n16603 = ~n16601 & ~n16602 ;
  assign n16604 = \u2_R6_reg[27]/NET0131  & ~n16603 ;
  assign n16605 = ~\u2_R6_reg[27]/NET0131  & n16603 ;
  assign n16606 = ~n16604 & ~n16605 ;
  assign n16620 = n16583 & ~n16606 ;
  assign n16572 = decrypt_pad & ~\u2_uk_K_r6_reg[49]/NET0131  ;
  assign n16573 = ~decrypt_pad & ~\u2_uk_K_r6_reg[42]/NET0131  ;
  assign n16574 = ~n16572 & ~n16573 ;
  assign n16575 = \u2_R6_reg[25]/NET0131  & ~n16574 ;
  assign n16576 = ~\u2_R6_reg[25]/NET0131  & n16574 ;
  assign n16577 = ~n16575 & ~n16576 ;
  assign n16585 = decrypt_pad & ~\u2_uk_K_r6_reg[38]/NET0131  ;
  assign n16586 = ~decrypt_pad & ~\u2_uk_K_r6_reg[31]/NET0131  ;
  assign n16587 = ~n16585 & ~n16586 ;
  assign n16588 = \u2_R6_reg[26]/NET0131  & ~n16587 ;
  assign n16589 = ~\u2_R6_reg[26]/NET0131  & n16587 ;
  assign n16590 = ~n16588 & ~n16589 ;
  assign n16623 = n16583 & ~n16590 ;
  assign n16591 = decrypt_pad & ~\u2_uk_K_r6_reg[22]/NET0131  ;
  assign n16592 = ~decrypt_pad & ~\u2_uk_K_r6_reg[15]/NET0131  ;
  assign n16593 = ~n16591 & ~n16592 ;
  assign n16594 = \u2_R6_reg[29]/NET0131  & ~n16593 ;
  assign n16595 = ~\u2_R6_reg[29]/NET0131  & n16593 ;
  assign n16596 = ~n16594 & ~n16595 ;
  assign n16598 = n16590 & ~n16596 ;
  assign n16624 = n16598 & ~n16606 ;
  assign n16625 = ~n16623 & ~n16624 ;
  assign n16626 = ~n16577 & ~n16625 ;
  assign n16627 = ~n16620 & ~n16626 ;
  assign n16566 = decrypt_pad & ~\u2_uk_K_r6_reg[30]/P0001  ;
  assign n16567 = ~decrypt_pad & ~\u2_uk_K_r6_reg[23]/P0001  ;
  assign n16568 = ~n16566 & ~n16567 ;
  assign n16569 = \u2_R6_reg[28]/NET0131  & ~n16568 ;
  assign n16570 = ~\u2_R6_reg[28]/NET0131  & n16568 ;
  assign n16571 = ~n16569 & ~n16570 ;
  assign n16597 = ~n16590 & n16596 ;
  assign n16607 = ~n16577 & n16590 ;
  assign n16621 = ~n16597 & ~n16607 ;
  assign n16622 = n16620 & ~n16621 ;
  assign n16628 = ~n16571 & ~n16622 ;
  assign n16629 = ~n16627 & n16628 ;
  assign n16613 = n16577 & n16597 ;
  assign n16614 = ~n16607 & ~n16613 ;
  assign n16615 = n16583 & n16606 ;
  assign n16616 = ~n16614 & n16615 ;
  assign n16584 = ~n16577 & ~n16583 ;
  assign n16599 = ~n16597 & ~n16598 ;
  assign n16600 = n16584 & n16599 ;
  assign n16608 = n16577 & n16583 ;
  assign n16609 = ~n16584 & ~n16608 ;
  assign n16610 = n16596 & ~n16606 ;
  assign n16611 = ~n16607 & n16610 ;
  assign n16612 = n16609 & n16611 ;
  assign n16617 = ~n16600 & ~n16612 ;
  assign n16618 = ~n16616 & n16617 ;
  assign n16619 = n16571 & ~n16618 ;
  assign n16630 = ~n16583 & n16590 ;
  assign n16631 = ~n16577 & ~n16596 ;
  assign n16633 = n16577 & n16596 ;
  assign n16634 = ~n16631 & ~n16633 ;
  assign n16635 = n16630 & ~n16634 ;
  assign n16632 = ~n16630 & ~n16631 ;
  assign n16636 = n16606 & ~n16632 ;
  assign n16637 = ~n16635 & n16636 ;
  assign n16639 = n16577 & ~n16606 ;
  assign n16640 = ~n16571 & n16596 ;
  assign n16641 = ~n16639 & ~n16640 ;
  assign n16638 = ~n16623 & ~n16630 ;
  assign n16642 = ~n16577 & n16606 ;
  assign n16643 = n16638 & ~n16642 ;
  assign n16644 = ~n16641 & n16643 ;
  assign n16645 = ~n16637 & ~n16644 ;
  assign n16646 = ~n16619 & n16645 ;
  assign n16647 = ~n16629 & n16646 ;
  assign n16648 = ~\u2_L6_reg[22]/NET0131  & ~n16647 ;
  assign n16649 = \u2_L6_reg[22]/NET0131  & n16647 ;
  assign n16650 = ~n16648 & ~n16649 ;
  assign n16667 = ~n16397 & ~n16404 ;
  assign n16668 = ~n16427 & ~n16667 ;
  assign n16669 = ~n16390 & ~n16668 ;
  assign n16670 = ~n16424 & ~n16669 ;
  assign n16671 = ~n16411 & ~n16670 ;
  assign n16672 = n16397 & n16441 ;
  assign n16673 = ~n16414 & ~n16672 ;
  assign n16674 = n16411 & ~n16673 ;
  assign n16675 = ~n16405 & ~n16456 ;
  assign n16676 = ~n16674 & n16675 ;
  assign n16677 = ~n16671 & n16676 ;
  assign n16678 = ~n16378 & ~n16677 ;
  assign n16651 = n16390 & n16421 ;
  assign n16652 = ~n16384 & n16651 ;
  assign n16653 = n16398 & ~n16404 ;
  assign n16654 = ~n16652 & ~n16653 ;
  assign n16655 = n16411 & ~n16654 ;
  assign n16657 = ~n16404 & ~n16429 ;
  assign n16658 = n16427 & n16429 ;
  assign n16659 = ~n16657 & ~n16658 ;
  assign n16660 = n16411 & ~n16659 ;
  assign n16661 = ~n16411 & ~n16452 ;
  assign n16662 = ~n16657 & n16661 ;
  assign n16656 = n16404 & n16455 ;
  assign n16663 = ~n16457 & ~n16656 ;
  assign n16664 = ~n16662 & n16663 ;
  assign n16665 = ~n16660 & n16664 ;
  assign n16666 = n16378 & ~n16665 ;
  assign n16679 = ~n16655 & ~n16666 ;
  assign n16680 = ~n16678 & n16679 ;
  assign n16681 = ~\u2_L6_reg[17]/NET0131  & ~n16680 ;
  assign n16682 = \u2_L6_reg[17]/NET0131  & n16680 ;
  assign n16683 = ~n16681 & ~n16682 ;
  assign n16697 = decrypt_pad & ~\u2_uk_K_r6_reg[48]/NET0131  ;
  assign n16698 = ~decrypt_pad & ~\u2_uk_K_r6_reg[41]/NET0131  ;
  assign n16699 = ~n16697 & ~n16698 ;
  assign n16700 = \u2_R6_reg[15]/NET0131  & ~n16699 ;
  assign n16701 = ~\u2_R6_reg[15]/NET0131  & n16699 ;
  assign n16702 = ~n16700 & ~n16701 ;
  assign n16711 = decrypt_pad & ~\u2_uk_K_r6_reg[40]/NET0131  ;
  assign n16712 = ~decrypt_pad & ~\u2_uk_K_r6_reg[33]/NET0131  ;
  assign n16713 = ~n16711 & ~n16712 ;
  assign n16714 = \u2_R6_reg[14]/NET0131  & ~n16713 ;
  assign n16715 = ~\u2_R6_reg[14]/NET0131  & n16713 ;
  assign n16716 = ~n16714 & ~n16715 ;
  assign n16726 = ~n16702 & ~n16716 ;
  assign n16690 = decrypt_pad & ~\u2_uk_K_r6_reg[20]/NET0131  ;
  assign n16691 = ~decrypt_pad & ~\u2_uk_K_r6_reg[13]/NET0131  ;
  assign n16692 = ~n16690 & ~n16691 ;
  assign n16693 = \u2_R6_reg[12]/NET0131  & ~n16692 ;
  assign n16694 = ~\u2_R6_reg[12]/NET0131  & n16692 ;
  assign n16695 = ~n16693 & ~n16694 ;
  assign n16704 = decrypt_pad & ~\u2_uk_K_r6_reg[39]/NET0131  ;
  assign n16705 = ~decrypt_pad & ~\u2_uk_K_r6_reg[32]/NET0131  ;
  assign n16706 = ~n16704 & ~n16705 ;
  assign n16707 = \u2_R6_reg[13]/NET0131  & ~n16706 ;
  assign n16708 = ~\u2_R6_reg[13]/NET0131  & n16706 ;
  assign n16709 = ~n16707 & ~n16708 ;
  assign n16727 = n16695 & ~n16709 ;
  assign n16728 = ~n16695 & n16709 ;
  assign n16729 = ~n16727 & ~n16728 ;
  assign n16730 = n16726 & ~n16729 ;
  assign n16684 = decrypt_pad & ~\u2_uk_K_r6_reg[4]/NET0131  ;
  assign n16685 = ~decrypt_pad & ~\u2_uk_K_r6_reg[54]/NET0131  ;
  assign n16686 = ~n16684 & ~n16685 ;
  assign n16687 = \u2_R6_reg[17]/NET0131  & ~n16686 ;
  assign n16688 = ~\u2_R6_reg[17]/NET0131  & n16686 ;
  assign n16689 = ~n16687 & ~n16688 ;
  assign n16696 = n16689 & ~n16695 ;
  assign n16703 = n16696 & n16702 ;
  assign n16710 = n16703 & ~n16709 ;
  assign n16723 = n16695 & n16702 ;
  assign n16724 = ~n16689 & n16709 ;
  assign n16725 = n16723 & n16724 ;
  assign n16731 = decrypt_pad & ~\u2_uk_K_r6_reg[24]/NET0131  ;
  assign n16732 = ~decrypt_pad & ~\u2_uk_K_r6_reg[17]/NET0131  ;
  assign n16733 = ~n16731 & ~n16732 ;
  assign n16734 = \u2_R6_reg[16]/NET0131  & ~n16733 ;
  assign n16735 = ~\u2_R6_reg[16]/NET0131  & n16733 ;
  assign n16736 = ~n16734 & ~n16735 ;
  assign n16741 = ~n16725 & n16736 ;
  assign n16742 = ~n16710 & n16741 ;
  assign n16743 = ~n16730 & n16742 ;
  assign n16717 = n16696 & n16709 ;
  assign n16718 = ~n16716 & n16717 ;
  assign n16719 = n16689 & n16695 ;
  assign n16720 = n16716 & n16719 ;
  assign n16721 = n16709 & n16720 ;
  assign n16722 = ~n16718 & ~n16721 ;
  assign n16737 = ~n16709 & n16716 ;
  assign n16738 = ~n16695 & n16737 ;
  assign n16739 = ~n16702 & n16738 ;
  assign n16740 = ~n16689 & n16739 ;
  assign n16744 = n16722 & ~n16740 ;
  assign n16745 = n16743 & n16744 ;
  assign n16755 = n16709 & n16719 ;
  assign n16750 = ~n16689 & ~n16709 ;
  assign n16756 = ~n16695 & n16750 ;
  assign n16757 = n16702 & ~n16756 ;
  assign n16758 = ~n16755 & n16757 ;
  assign n16760 = ~n16689 & n16695 ;
  assign n16761 = n16716 & n16760 ;
  assign n16759 = n16689 & ~n16709 ;
  assign n16762 = ~n16702 & ~n16759 ;
  assign n16763 = ~n16761 & n16762 ;
  assign n16764 = ~n16758 & ~n16763 ;
  assign n16753 = n16702 & n16716 ;
  assign n16754 = n16728 & n16753 ;
  assign n16751 = ~n16695 & ~n16716 ;
  assign n16752 = n16750 & n16751 ;
  assign n16765 = ~n16736 & ~n16752 ;
  assign n16766 = ~n16754 & n16765 ;
  assign n16746 = ~n16716 & n16727 ;
  assign n16747 = n16689 & n16746 ;
  assign n16748 = ~n16689 & n16728 ;
  assign n16749 = n16716 & n16748 ;
  assign n16767 = ~n16747 & ~n16749 ;
  assign n16768 = n16766 & n16767 ;
  assign n16769 = ~n16764 & n16768 ;
  assign n16770 = ~n16745 & ~n16769 ;
  assign n16771 = ~n16702 & ~n16718 ;
  assign n16772 = ~n16709 & n16761 ;
  assign n16773 = n16702 & ~n16772 ;
  assign n16774 = n16709 & ~n16716 ;
  assign n16775 = n16760 & n16774 ;
  assign n16776 = ~n16752 & ~n16775 ;
  assign n16777 = n16773 & n16776 ;
  assign n16778 = ~n16771 & ~n16777 ;
  assign n16779 = ~n16770 & ~n16778 ;
  assign n16780 = ~\u2_L6_reg[20]/NET0131  & ~n16779 ;
  assign n16781 = \u2_L6_reg[20]/NET0131  & n16779 ;
  assign n16782 = ~n16780 & ~n16781 ;
  assign n16806 = ~n16499 & n16512 ;
  assign n16807 = ~n16545 & ~n16806 ;
  assign n16808 = ~n16501 & ~n16543 ;
  assign n16809 = ~n16511 & ~n16808 ;
  assign n16810 = n16807 & ~n16809 ;
  assign n16811 = n16479 & ~n16810 ;
  assign n16783 = n16485 & n16537 ;
  assign n16803 = ~n16485 & n16549 ;
  assign n16804 = ~n16783 & ~n16803 ;
  assign n16805 = ~n16479 & ~n16804 ;
  assign n16812 = n16485 & n16522 ;
  assign n16813 = ~n16805 & ~n16812 ;
  assign n16814 = ~n16811 & n16813 ;
  assign n16815 = ~n16473 & ~n16814 ;
  assign n16784 = ~n16485 & ~n16492 ;
  assign n16785 = n16499 & n16784 ;
  assign n16786 = ~n16552 & ~n16785 ;
  assign n16787 = ~n16783 & n16786 ;
  assign n16788 = n16479 & ~n16787 ;
  assign n16789 = ~n16492 & ~n16511 ;
  assign n16793 = n16485 & n16789 ;
  assign n16794 = n16511 & n16784 ;
  assign n16795 = ~n16793 & ~n16794 ;
  assign n16796 = ~n16499 & ~n16795 ;
  assign n16790 = ~n16502 & n16789 ;
  assign n16791 = ~n16533 & ~n16790 ;
  assign n16792 = ~n16479 & ~n16791 ;
  assign n16797 = ~n16514 & ~n16520 ;
  assign n16798 = ~n16792 & n16797 ;
  assign n16799 = ~n16796 & n16798 ;
  assign n16800 = ~n16788 & n16799 ;
  assign n16801 = n16473 & ~n16800 ;
  assign n16802 = n16486 & n16551 ;
  assign n16816 = ~n16544 & ~n16802 ;
  assign n16817 = ~n16801 & n16816 ;
  assign n16818 = ~n16815 & n16817 ;
  assign n16819 = \u2_L6_reg[29]/NET0131  & ~n16818 ;
  assign n16820 = ~\u2_L6_reg[29]/NET0131  & n16818 ;
  assign n16821 = ~n16819 & ~n16820 ;
  assign n16822 = decrypt_pad & ~\u2_uk_K_r6_reg[55]/P0001  ;
  assign n16823 = ~decrypt_pad & ~\u2_uk_K_r6_reg[48]/NET0131  ;
  assign n16824 = ~n16822 & ~n16823 ;
  assign n16825 = \u2_R6_reg[8]/NET0131  & ~n16824 ;
  assign n16826 = ~\u2_R6_reg[8]/NET0131  & n16824 ;
  assign n16827 = ~n16825 & ~n16826 ;
  assign n16828 = decrypt_pad & ~\u2_uk_K_r6_reg[47]/NET0131  ;
  assign n16829 = ~decrypt_pad & ~\u2_uk_K_r6_reg[40]/NET0131  ;
  assign n16830 = ~n16828 & ~n16829 ;
  assign n16831 = \u2_R6_reg[5]/NET0131  & ~n16830 ;
  assign n16832 = ~\u2_R6_reg[5]/NET0131  & n16830 ;
  assign n16833 = ~n16831 & ~n16832 ;
  assign n16834 = decrypt_pad & ~\u2_uk_K_r6_reg[3]/NET0131  ;
  assign n16835 = ~decrypt_pad & ~\u2_uk_K_r6_reg[53]/NET0131  ;
  assign n16836 = ~n16834 & ~n16835 ;
  assign n16837 = \u2_R6_reg[9]/NET0131  & ~n16836 ;
  assign n16838 = ~\u2_R6_reg[9]/NET0131  & n16836 ;
  assign n16839 = ~n16837 & ~n16838 ;
  assign n16840 = n16833 & ~n16839 ;
  assign n16841 = ~n16833 & n16839 ;
  assign n16842 = decrypt_pad & ~\u2_uk_K_r6_reg[11]/NET0131  ;
  assign n16843 = ~decrypt_pad & ~\u2_uk_K_r6_reg[4]/NET0131  ;
  assign n16844 = ~n16842 & ~n16843 ;
  assign n16845 = \u2_R6_reg[4]/NET0131  & ~n16844 ;
  assign n16846 = ~\u2_R6_reg[4]/NET0131  & n16844 ;
  assign n16847 = ~n16845 & ~n16846 ;
  assign n16848 = n16841 & ~n16847 ;
  assign n16849 = ~n16840 & ~n16848 ;
  assign n16850 = decrypt_pad & ~\u2_uk_K_r6_reg[13]/NET0131  ;
  assign n16851 = ~decrypt_pad & ~\u2_uk_K_r6_reg[6]/NET0131  ;
  assign n16852 = ~n16850 & ~n16851 ;
  assign n16853 = \u2_R6_reg[6]/NET0131  & ~n16852 ;
  assign n16854 = ~\u2_R6_reg[6]/NET0131  & n16852 ;
  assign n16855 = ~n16853 & ~n16854 ;
  assign n16856 = ~n16849 & ~n16855 ;
  assign n16857 = decrypt_pad & ~\u2_uk_K_r6_reg[32]/NET0131  ;
  assign n16858 = ~decrypt_pad & ~\u2_uk_K_r6_reg[25]/NET0131  ;
  assign n16859 = ~n16857 & ~n16858 ;
  assign n16860 = \u2_R6_reg[7]/NET0131  & ~n16859 ;
  assign n16861 = ~\u2_R6_reg[7]/NET0131  & n16859 ;
  assign n16862 = ~n16860 & ~n16861 ;
  assign n16863 = ~n16833 & n16855 ;
  assign n16864 = n16839 & n16847 ;
  assign n16865 = n16863 & n16864 ;
  assign n16866 = n16862 & n16865 ;
  assign n16880 = ~n16856 & ~n16866 ;
  assign n16867 = n16847 & n16855 ;
  assign n16868 = ~n16841 & n16867 ;
  assign n16869 = ~n16848 & ~n16868 ;
  assign n16870 = ~n16862 & ~n16869 ;
  assign n16874 = n16833 & ~n16855 ;
  assign n16875 = ~n16855 & n16862 ;
  assign n16876 = ~n16874 & ~n16875 ;
  assign n16871 = n16839 & ~n16847 ;
  assign n16872 = n16833 & ~n16871 ;
  assign n16873 = ~n16839 & ~n16855 ;
  assign n16877 = ~n16863 & ~n16873 ;
  assign n16878 = ~n16872 & n16877 ;
  assign n16879 = n16876 & n16878 ;
  assign n16881 = ~n16870 & ~n16879 ;
  assign n16882 = n16880 & n16881 ;
  assign n16883 = ~n16827 & ~n16882 ;
  assign n16896 = ~n16839 & ~n16847 ;
  assign n16900 = ~n16865 & ~n16896 ;
  assign n16901 = n16827 & ~n16900 ;
  assign n16902 = ~n16863 & n16871 ;
  assign n16903 = ~n16901 & ~n16902 ;
  assign n16904 = ~n16862 & ~n16874 ;
  assign n16905 = ~n16903 & n16904 ;
  assign n16890 = ~n16855 & n16864 ;
  assign n16891 = n16833 & n16890 ;
  assign n16884 = ~n16839 & n16847 ;
  assign n16885 = ~n16833 & n16884 ;
  assign n16886 = ~n16855 & n16885 ;
  assign n16887 = ~n16847 & n16855 ;
  assign n16888 = n16833 & n16862 ;
  assign n16889 = ~n16887 & n16888 ;
  assign n16892 = ~n16886 & ~n16889 ;
  assign n16893 = ~n16891 & n16892 ;
  assign n16894 = n16827 & ~n16893 ;
  assign n16897 = ~n16874 & ~n16896 ;
  assign n16895 = ~n16847 & ~n16863 ;
  assign n16898 = n16862 & ~n16895 ;
  assign n16899 = ~n16897 & n16898 ;
  assign n16906 = ~n16894 & ~n16899 ;
  assign n16907 = ~n16905 & n16906 ;
  assign n16908 = ~n16883 & n16907 ;
  assign n16909 = \u2_L6_reg[2]/NET0131  & n16908 ;
  assign n16910 = ~\u2_L6_reg[2]/NET0131  & ~n16908 ;
  assign n16911 = ~n16909 & ~n16910 ;
  assign n16916 = ~n16537 & ~n16794 ;
  assign n16917 = ~n16520 & n16916 ;
  assign n16918 = n16479 & ~n16917 ;
  assign n16912 = n16499 & n16789 ;
  assign n16913 = ~n16812 & ~n16912 ;
  assign n16914 = ~n16479 & ~n16913 ;
  assign n16915 = n16513 & n16518 ;
  assign n16919 = ~n16544 & ~n16915 ;
  assign n16920 = ~n16914 & n16919 ;
  assign n16921 = ~n16918 & n16920 ;
  assign n16922 = ~n16473 & ~n16921 ;
  assign n16930 = ~n16524 & ~n16784 ;
  assign n16931 = ~n16479 & ~n16930 ;
  assign n16932 = n16485 & n16551 ;
  assign n16933 = n16486 & n16518 ;
  assign n16934 = ~n16932 & ~n16933 ;
  assign n16935 = ~n16534 & n16934 ;
  assign n16936 = ~n16931 & n16935 ;
  assign n16937 = n16473 & ~n16936 ;
  assign n16923 = ~n16541 & ~n16552 ;
  assign n16924 = ~n16537 & n16923 ;
  assign n16925 = n16516 & ~n16924 ;
  assign n16926 = n16485 & n16807 ;
  assign n16927 = ~n16485 & ~n16789 ;
  assign n16928 = ~n16479 & ~n16927 ;
  assign n16929 = ~n16926 & n16928 ;
  assign n16938 = ~n16925 & ~n16929 ;
  assign n16939 = ~n16937 & n16938 ;
  assign n16940 = ~n16922 & n16939 ;
  assign n16941 = ~\u2_L6_reg[4]/NET0131  & ~n16940 ;
  assign n16942 = \u2_L6_reg[4]/NET0131  & n16940 ;
  assign n16943 = ~n16941 & ~n16942 ;
  assign n16944 = decrypt_pad & ~\u2_uk_K_r6_reg[50]/NET0131  ;
  assign n16945 = ~decrypt_pad & ~\u2_uk_K_r6_reg[43]/NET0131  ;
  assign n16946 = ~n16944 & ~n16945 ;
  assign n16947 = \u2_R6_reg[32]/NET0131  & ~n16946 ;
  assign n16948 = ~\u2_R6_reg[32]/NET0131  & n16946 ;
  assign n16949 = ~n16947 & ~n16948 ;
  assign n16983 = decrypt_pad & ~\u2_uk_K_r6_reg[44]/NET0131  ;
  assign n16984 = ~decrypt_pad & ~\u2_uk_K_r6_reg[37]/NET0131  ;
  assign n16985 = ~n16983 & ~n16984 ;
  assign n16986 = \u2_R6_reg[31]/P0001  & ~n16985 ;
  assign n16987 = ~\u2_R6_reg[31]/P0001  & n16985 ;
  assign n16988 = ~n16986 & ~n16987 ;
  assign n16950 = decrypt_pad & ~\u2_uk_K_r6_reg[1]/NET0131  ;
  assign n16951 = ~decrypt_pad & ~\u2_uk_K_r6_reg[49]/NET0131  ;
  assign n16952 = ~n16950 & ~n16951 ;
  assign n16953 = \u2_R6_reg[30]/NET0131  & ~n16952 ;
  assign n16954 = ~\u2_R6_reg[30]/NET0131  & n16952 ;
  assign n16955 = ~n16953 & ~n16954 ;
  assign n16963 = decrypt_pad & ~\u2_uk_K_r6_reg[28]/NET0131  ;
  assign n16964 = ~decrypt_pad & ~\u2_uk_K_r6_reg[21]/NET0131  ;
  assign n16965 = ~n16963 & ~n16964 ;
  assign n16966 = \u2_R6_reg[28]/NET0131  & ~n16965 ;
  assign n16967 = ~\u2_R6_reg[28]/NET0131  & n16965 ;
  assign n16968 = ~n16966 & ~n16967 ;
  assign n16990 = ~n16955 & n16968 ;
  assign n16956 = decrypt_pad & ~\u2_uk_K_r6_reg[0]/NET0131  ;
  assign n16957 = ~decrypt_pad & ~\u2_uk_K_r6_reg[52]/NET0131  ;
  assign n16958 = ~n16956 & ~n16957 ;
  assign n16959 = \u2_R6_reg[29]/NET0131  & ~n16958 ;
  assign n16960 = ~\u2_R6_reg[29]/NET0131  & n16958 ;
  assign n16961 = ~n16959 & ~n16960 ;
  assign n16969 = decrypt_pad & ~\u2_uk_K_r6_reg[16]/NET0131  ;
  assign n16970 = ~decrypt_pad & ~\u2_uk_K_r6_reg[9]/NET0131  ;
  assign n16971 = ~n16969 & ~n16970 ;
  assign n16972 = \u2_R6_reg[1]/NET0131  & ~n16971 ;
  assign n16973 = ~\u2_R6_reg[1]/NET0131  & n16971 ;
  assign n16974 = ~n16972 & ~n16973 ;
  assign n16980 = ~n16961 & n16974 ;
  assign n16991 = n16955 & ~n16968 ;
  assign n16992 = ~n16974 & ~n16991 ;
  assign n16993 = ~n16980 & ~n16992 ;
  assign n16994 = ~n16990 & ~n16993 ;
  assign n16995 = ~n16988 & ~n16994 ;
  assign n16977 = ~n16961 & ~n16974 ;
  assign n16978 = n16955 & n16977 ;
  assign n16979 = n16968 & n16978 ;
  assign n16981 = ~n16968 & n16980 ;
  assign n16982 = ~n16979 & ~n16981 ;
  assign n16989 = ~n16982 & n16988 ;
  assign n16962 = n16955 & n16961 ;
  assign n16975 = n16968 & n16974 ;
  assign n16976 = n16962 & n16975 ;
  assign n16996 = n16968 & ~n16974 ;
  assign n16997 = ~n16955 & n16961 ;
  assign n16998 = n16996 & n16997 ;
  assign n16999 = ~n16976 & ~n16998 ;
  assign n17000 = ~n16989 & n16999 ;
  assign n17001 = ~n16995 & n17000 ;
  assign n17002 = ~n16949 & ~n17001 ;
  assign n17015 = n16961 & ~n16974 ;
  assign n17016 = ~n16990 & ~n17015 ;
  assign n17017 = n16949 & ~n16998 ;
  assign n17018 = ~n17016 & n17017 ;
  assign n17011 = ~n16968 & n16977 ;
  assign n17012 = ~n16955 & n17011 ;
  assign n17004 = n16962 & ~n16968 ;
  assign n17013 = ~n16974 & n17004 ;
  assign n17014 = ~n17012 & ~n17013 ;
  assign n17006 = ~n16990 & ~n16991 ;
  assign n17019 = n16980 & ~n17006 ;
  assign n17020 = n17014 & ~n17019 ;
  assign n17021 = ~n17018 & n17020 ;
  assign n17022 = n16988 & ~n17021 ;
  assign n17003 = ~n16988 & n16998 ;
  assign n17005 = n16974 & n17004 ;
  assign n17007 = ~n16961 & ~n16988 ;
  assign n17008 = n17006 & n17007 ;
  assign n17009 = ~n17005 & ~n17008 ;
  assign n17010 = n16949 & ~n17009 ;
  assign n17023 = ~n17003 & ~n17010 ;
  assign n17024 = ~n17022 & n17023 ;
  assign n17025 = ~n17002 & n17024 ;
  assign n17026 = \u2_L6_reg[5]/NET0131  & ~n17025 ;
  assign n17027 = ~\u2_L6_reg[5]/NET0131  & n17025 ;
  assign n17028 = ~n17026 & ~n17027 ;
  assign n17042 = ~n16747 & ~n16748 ;
  assign n17043 = n16702 & ~n17042 ;
  assign n17040 = n16689 & n16738 ;
  assign n17041 = ~n16721 & ~n17040 ;
  assign n17044 = n16689 & n16774 ;
  assign n17045 = ~n16760 & ~n17044 ;
  assign n17031 = n16695 & n16774 ;
  assign n17046 = ~n16702 & ~n17031 ;
  assign n17047 = ~n17045 & n17046 ;
  assign n17048 = n17041 & ~n17047 ;
  assign n17049 = ~n17043 & n17048 ;
  assign n17050 = n16736 & ~n17049 ;
  assign n17029 = ~n16703 & ~n16756 ;
  assign n17030 = ~n16753 & ~n17029 ;
  assign n17033 = ~n16737 & ~n16750 ;
  assign n17034 = n16723 & ~n17033 ;
  assign n17032 = n16719 & n16726 ;
  assign n17035 = ~n17031 & ~n17032 ;
  assign n17036 = ~n16749 & n17035 ;
  assign n17037 = ~n17034 & n17036 ;
  assign n17038 = ~n17030 & n17037 ;
  assign n17039 = ~n16736 & ~n17038 ;
  assign n17052 = ~n16752 & n17041 ;
  assign n17053 = ~n16702 & ~n17052 ;
  assign n17051 = ~n16716 & n16725 ;
  assign n17054 = ~n16754 & ~n17051 ;
  assign n17055 = ~n17053 & n17054 ;
  assign n17056 = ~n17039 & n17055 ;
  assign n17057 = ~n17050 & n17056 ;
  assign n17058 = ~\u2_L6_reg[10]/NET0131  & ~n17057 ;
  assign n17059 = \u2_L6_reg[10]/NET0131  & n17057 ;
  assign n17060 = ~n17058 & ~n17059 ;
  assign n17061 = ~n16583 & n16596 ;
  assign n17065 = n16606 & ~n16630 ;
  assign n17066 = ~n17061 & n17065 ;
  assign n17067 = ~n16609 & n17066 ;
  assign n17064 = ~n16599 & n16609 ;
  assign n17062 = n16607 & n17061 ;
  assign n17063 = ~n16606 & n17062 ;
  assign n17068 = n16571 & ~n17063 ;
  assign n17069 = ~n17064 & n17068 ;
  assign n17070 = ~n17067 & n17069 ;
  assign n17075 = ~n16577 & ~n16590 ;
  assign n17076 = n16583 & ~n16596 ;
  assign n17077 = ~n17061 & ~n17076 ;
  assign n17078 = ~n17075 & n17077 ;
  assign n17079 = n16577 & n16590 ;
  assign n17080 = ~n16623 & ~n17079 ;
  assign n17081 = n17078 & n17080 ;
  assign n17071 = ~n16590 & ~n16631 ;
  assign n17072 = n16590 & n16606 ;
  assign n17073 = n16583 & ~n17072 ;
  assign n17074 = ~n17071 & n17073 ;
  assign n17085 = ~n16571 & ~n17074 ;
  assign n17082 = ~n16642 & ~n17079 ;
  assign n17083 = n17061 & ~n17082 ;
  assign n17084 = ~n16606 & ~n16634 ;
  assign n17086 = ~n17083 & ~n17084 ;
  assign n17087 = n17085 & n17086 ;
  assign n17088 = ~n17081 & n17087 ;
  assign n17089 = ~n17070 & ~n17088 ;
  assign n17090 = \u2_L6_reg[12]/NET0131  & n17089 ;
  assign n17091 = ~\u2_L6_reg[12]/NET0131  & ~n17089 ;
  assign n17092 = ~n17090 & ~n17091 ;
  assign n17093 = n16840 & n16867 ;
  assign n17094 = ~n16891 & ~n17093 ;
  assign n17095 = n16848 & n16855 ;
  assign n17096 = n16840 & ~n16847 ;
  assign n17097 = ~n16886 & ~n17096 ;
  assign n17098 = ~n17095 & n17097 ;
  assign n17099 = ~n16827 & ~n17098 ;
  assign n17100 = n17094 & ~n17099 ;
  assign n17101 = ~n16862 & ~n17100 ;
  assign n17105 = ~n16833 & ~n16871 ;
  assign n17106 = ~n16884 & ~n17105 ;
  assign n17107 = ~n16874 & n16884 ;
  assign n17108 = n16862 & ~n17107 ;
  assign n17109 = ~n17106 & n17108 ;
  assign n17103 = ~n16840 & n16862 ;
  assign n17104 = n16867 & n17103 ;
  assign n17102 = n16871 & ~n16876 ;
  assign n17110 = ~n16827 & ~n17102 ;
  assign n17111 = ~n17104 & n17110 ;
  assign n17112 = ~n17109 & n17111 ;
  assign n17119 = ~n16855 & n17096 ;
  assign n17120 = n16827 & ~n17119 ;
  assign n17121 = ~n16879 & n17120 ;
  assign n17117 = ~n16873 & n17105 ;
  assign n17118 = ~n16862 & n17117 ;
  assign n17113 = ~n16833 & n16873 ;
  assign n17114 = n16855 & n16871 ;
  assign n17115 = ~n17113 & ~n17114 ;
  assign n17116 = n16862 & ~n17115 ;
  assign n17122 = n17094 & ~n17116 ;
  assign n17123 = ~n17118 & n17122 ;
  assign n17124 = n17121 & n17123 ;
  assign n17125 = ~n17112 & ~n17124 ;
  assign n17126 = ~n17101 & ~n17125 ;
  assign n17127 = ~\u2_L6_reg[13]/NET0131  & n17126 ;
  assign n17128 = \u2_L6_reg[13]/NET0131  & ~n17126 ;
  assign n17129 = ~n17127 & ~n17128 ;
  assign n17190 = decrypt_pad & ~\u2_uk_K_r6_reg[35]/NET0131  ;
  assign n17191 = ~decrypt_pad & ~\u2_uk_K_r6_reg[28]/NET0131  ;
  assign n17192 = ~n17190 & ~n17191 ;
  assign n17193 = \u2_R6_reg[20]/NET0131  & ~n17192 ;
  assign n17194 = ~\u2_R6_reg[20]/NET0131  & n17192 ;
  assign n17195 = ~n17193 & ~n17194 ;
  assign n17155 = decrypt_pad & ~\u2_uk_K_r6_reg[51]/NET0131  ;
  assign n17156 = ~decrypt_pad & ~\u2_uk_K_r6_reg[44]/NET0131  ;
  assign n17157 = ~n17155 & ~n17156 ;
  assign n17158 = \u2_R6_reg[19]/NET0131  & ~n17157 ;
  assign n17159 = ~\u2_R6_reg[19]/NET0131  & n17157 ;
  assign n17160 = ~n17158 & ~n17159 ;
  assign n17130 = decrypt_pad & ~\u2_uk_K_r6_reg[52]/NET0131  ;
  assign n17131 = ~decrypt_pad & ~\u2_uk_K_r6_reg[45]/NET0131  ;
  assign n17132 = ~n17130 & ~n17131 ;
  assign n17133 = \u2_R6_reg[16]/NET0131  & ~n17132 ;
  assign n17134 = ~\u2_R6_reg[16]/NET0131  & n17132 ;
  assign n17135 = ~n17133 & ~n17134 ;
  assign n17143 = decrypt_pad & ~\u2_uk_K_r6_reg[15]/NET0131  ;
  assign n17144 = ~decrypt_pad & ~\u2_uk_K_r6_reg[8]/NET0131  ;
  assign n17145 = ~n17143 & ~n17144 ;
  assign n17146 = \u2_R6_reg[17]/NET0131  & ~n17145 ;
  assign n17147 = ~\u2_R6_reg[17]/NET0131  & n17145 ;
  assign n17148 = ~n17146 & ~n17147 ;
  assign n17136 = decrypt_pad & ~\u2_uk_K_r6_reg[36]/NET0131  ;
  assign n17137 = ~decrypt_pad & ~\u2_uk_K_r6_reg[29]/NET0131  ;
  assign n17138 = ~n17136 & ~n17137 ;
  assign n17139 = \u2_R6_reg[21]/NET0131  & ~n17138 ;
  assign n17140 = ~\u2_R6_reg[21]/NET0131  & n17138 ;
  assign n17141 = ~n17139 & ~n17140 ;
  assign n17163 = decrypt_pad & ~\u2_uk_K_r6_reg[9]/NET0131  ;
  assign n17164 = ~decrypt_pad & ~\u2_uk_K_r6_reg[2]/NET0131  ;
  assign n17165 = ~n17163 & ~n17164 ;
  assign n17166 = \u2_R6_reg[18]/NET0131  & ~n17165 ;
  assign n17167 = ~\u2_R6_reg[18]/NET0131  & n17165 ;
  assign n17168 = ~n17166 & ~n17167 ;
  assign n17197 = n17141 & ~n17168 ;
  assign n17198 = n17148 & n17197 ;
  assign n17199 = n17135 & n17198 ;
  assign n17142 = n17135 & ~n17141 ;
  assign n17171 = ~n17148 & ~n17168 ;
  assign n17201 = n17142 & n17171 ;
  assign n17178 = ~n17135 & n17141 ;
  assign n17179 = ~n17148 & n17178 ;
  assign n17172 = n17148 & n17168 ;
  assign n17200 = ~n17141 & n17172 ;
  assign n17202 = ~n17179 & ~n17200 ;
  assign n17203 = ~n17201 & n17202 ;
  assign n17204 = ~n17199 & n17203 ;
  assign n17205 = ~n17160 & ~n17204 ;
  assign n17152 = ~n17135 & n17148 ;
  assign n17206 = n17152 & ~n17168 ;
  assign n17207 = ~n17152 & ~n17197 ;
  assign n17208 = ~n17142 & ~n17178 ;
  assign n17209 = n17207 & n17208 ;
  assign n17210 = ~n17206 & ~n17209 ;
  assign n17211 = n17160 & ~n17210 ;
  assign n17212 = ~n17142 & ~n17197 ;
  assign n17150 = ~n17135 & ~n17148 ;
  assign n17213 = ~n17150 & ~n17172 ;
  assign n17214 = n17212 & n17213 ;
  assign n17215 = ~n17211 & ~n17214 ;
  assign n17216 = ~n17205 & n17215 ;
  assign n17217 = ~n17195 & ~n17216 ;
  assign n17149 = n17142 & n17148 ;
  assign n17151 = ~n17141 & n17150 ;
  assign n17153 = n17141 & n17152 ;
  assign n17154 = ~n17151 & ~n17153 ;
  assign n17161 = ~n17154 & ~n17160 ;
  assign n17162 = ~n17149 & ~n17161 ;
  assign n17169 = ~n17162 & ~n17168 ;
  assign n17183 = ~n17149 & ~n17179 ;
  assign n17170 = n17135 & n17141 ;
  assign n17180 = ~n17168 & n17170 ;
  assign n17181 = ~n17135 & n17168 ;
  assign n17182 = n17141 & n17181 ;
  assign n17184 = ~n17180 & ~n17182 ;
  assign n17185 = n17183 & n17184 ;
  assign n17186 = n17160 & ~n17185 ;
  assign n17173 = ~n17160 & n17172 ;
  assign n17174 = ~n17171 & ~n17173 ;
  assign n17175 = n17170 & ~n17174 ;
  assign n17176 = ~n17148 & n17168 ;
  assign n17177 = n17142 & n17176 ;
  assign n17187 = ~n17175 & ~n17177 ;
  assign n17188 = ~n17186 & n17187 ;
  assign n17189 = ~n17169 & n17188 ;
  assign n17196 = ~n17189 & n17195 ;
  assign n17218 = ~n17148 & n17182 ;
  assign n17219 = ~n17200 & ~n17218 ;
  assign n17220 = ~n17135 & ~n17219 ;
  assign n17221 = ~n17160 & n17220 ;
  assign n17222 = n17149 & ~n17168 ;
  assign n17223 = n17151 & n17168 ;
  assign n17224 = ~n17222 & ~n17223 ;
  assign n17225 = n17160 & ~n17224 ;
  assign n17226 = ~n17221 & ~n17225 ;
  assign n17227 = ~n17196 & n17226 ;
  assign n17228 = ~n17217 & n17227 ;
  assign n17229 = ~\u2_L6_reg[14]/NET0131  & ~n17228 ;
  assign n17230 = \u2_L6_reg[14]/NET0131  & n17228 ;
  assign n17231 = ~n17229 & ~n17230 ;
  assign n17232 = ~n16968 & n16974 ;
  assign n17233 = n16961 & ~n16991 ;
  assign n17234 = ~n17232 & n17233 ;
  assign n17235 = ~n16981 & ~n17234 ;
  assign n17236 = n16988 & ~n17235 ;
  assign n17237 = n16977 & n16990 ;
  assign n17238 = ~n17236 & ~n17237 ;
  assign n17239 = ~n16949 & ~n17238 ;
  assign n17240 = n16968 & n16997 ;
  assign n17244 = n16955 & ~n16988 ;
  assign n17245 = n16980 & n17244 ;
  assign n17246 = ~n17240 & ~n17245 ;
  assign n17247 = ~n17013 & n17246 ;
  assign n17241 = n16988 & n17011 ;
  assign n17242 = ~n16961 & n16975 ;
  assign n17243 = n16955 & n17242 ;
  assign n17248 = ~n17241 & ~n17243 ;
  assign n17249 = n17247 & n17248 ;
  assign n17250 = n16949 & ~n17249 ;
  assign n17252 = ~n16961 & n16968 ;
  assign n17253 = n16949 & ~n16955 ;
  assign n17254 = n17252 & ~n17253 ;
  assign n17251 = n16997 & n17232 ;
  assign n17255 = ~n16988 & ~n17251 ;
  assign n17256 = ~n17254 & n17255 ;
  assign n17257 = n17014 & n17256 ;
  assign n17258 = ~n16955 & ~n16961 ;
  assign n17259 = ~n16968 & n17258 ;
  assign n17260 = n16974 & n17259 ;
  assign n17261 = n16988 & ~n17005 ;
  assign n17262 = ~n17260 & n17261 ;
  assign n17263 = ~n17257 & ~n17262 ;
  assign n17264 = ~n17250 & ~n17263 ;
  assign n17265 = ~n17239 & n17264 ;
  assign n17266 = ~\u2_L6_reg[15]/NET0131  & ~n17265 ;
  assign n17267 = \u2_L6_reg[15]/NET0131  & n17265 ;
  assign n17268 = ~n17266 & ~n17267 ;
  assign n17271 = n16492 & ~n16502 ;
  assign n17272 = ~n16912 & ~n17271 ;
  assign n17273 = n16479 & ~n17272 ;
  assign n17270 = ~n16479 & ~n16923 ;
  assign n17269 = n16485 & n16545 ;
  assign n17274 = ~n16473 & ~n17269 ;
  assign n17275 = ~n17270 & n17274 ;
  assign n17276 = ~n17273 & n17275 ;
  assign n17279 = n16485 & n16552 ;
  assign n17280 = ~n16479 & n16515 ;
  assign n17281 = n16473 & ~n16524 ;
  assign n17282 = ~n17280 & n17281 ;
  assign n17283 = ~n17279 & n17282 ;
  assign n17277 = ~n16503 & ~n16522 ;
  assign n17278 = n16479 & ~n17277 ;
  assign n17284 = ~n16796 & ~n17278 ;
  assign n17285 = n17283 & n17284 ;
  assign n17286 = ~n17276 & ~n17285 ;
  assign n17287 = n16513 & n16519 ;
  assign n17288 = ~n16540 & ~n17287 ;
  assign n17289 = ~n17286 & n17288 ;
  assign n17290 = ~\u2_L6_reg[19]/NET0131  & ~n17289 ;
  assign n17291 = \u2_L6_reg[19]/NET0131  & n17289 ;
  assign n17292 = ~n17290 & ~n17291 ;
  assign n17306 = ~n16689 & ~n16716 ;
  assign n17307 = ~n16759 & ~n17306 ;
  assign n17308 = n16695 & ~n17307 ;
  assign n17309 = ~n16702 & ~n17308 ;
  assign n17310 = ~n16695 & n17306 ;
  assign n17311 = n16773 & ~n17310 ;
  assign n17312 = ~n17309 & ~n17311 ;
  assign n17313 = n16722 & ~n16775 ;
  assign n17314 = ~n17312 & n17313 ;
  assign n17315 = ~n16736 & ~n17314 ;
  assign n17300 = ~n16760 & n16774 ;
  assign n17301 = ~n16717 & ~n17300 ;
  assign n17302 = ~n16702 & ~n17301 ;
  assign n17295 = n16709 & n16761 ;
  assign n17303 = ~n16738 & ~n17295 ;
  assign n17304 = ~n17302 & n17303 ;
  assign n17305 = n16736 & ~n17304 ;
  assign n17293 = ~n16749 & n17041 ;
  assign n17294 = n16702 & ~n17293 ;
  assign n17297 = ~n16746 & ~n16759 ;
  assign n17298 = n16702 & n16736 ;
  assign n17299 = ~n17297 & n17298 ;
  assign n17296 = ~n16702 & n17295 ;
  assign n17316 = ~n16740 & ~n17296 ;
  assign n17317 = ~n17299 & n17316 ;
  assign n17318 = ~n17294 & n17317 ;
  assign n17319 = ~n17305 & n17318 ;
  assign n17320 = ~n17315 & n17319 ;
  assign n17321 = ~\u2_L6_reg[1]/NET0131  & ~n17320 ;
  assign n17322 = \u2_L6_reg[1]/NET0131  & n17320 ;
  assign n17323 = ~n17321 & ~n17322 ;
  assign n17327 = ~n16980 & n16990 ;
  assign n17328 = ~n16988 & ~n17327 ;
  assign n17329 = ~n17243 & n17328 ;
  assign n17330 = n16988 & ~n17259 ;
  assign n17333 = n16962 & n16968 ;
  assign n17331 = n16974 & n17258 ;
  assign n17332 = n16961 & n17232 ;
  assign n17334 = ~n17331 & ~n17332 ;
  assign n17335 = ~n17333 & n17334 ;
  assign n17336 = n17330 & n17335 ;
  assign n17337 = ~n17329 & ~n17336 ;
  assign n17324 = n16961 & n16996 ;
  assign n17325 = ~n17011 & ~n17324 ;
  assign n17326 = n16955 & ~n17325 ;
  assign n17338 = n16949 & ~n17260 ;
  assign n17339 = ~n17326 & n17338 ;
  assign n17340 = ~n17337 & n17339 ;
  assign n17342 = n16974 & ~n17006 ;
  assign n17343 = ~n16988 & ~n17342 ;
  assign n17344 = n16955 & n17252 ;
  assign n17345 = ~n17324 & ~n17344 ;
  assign n17346 = n17330 & n17345 ;
  assign n17347 = ~n17343 & ~n17346 ;
  assign n17349 = ~n16968 & ~n16988 ;
  assign n17350 = n17015 & n17349 ;
  assign n17351 = ~n16979 & ~n17350 ;
  assign n17348 = n16974 & n17240 ;
  assign n17341 = ~n16949 & ~n17004 ;
  assign n17352 = ~n17012 & n17341 ;
  assign n17353 = ~n17348 & n17352 ;
  assign n17354 = n17351 & n17353 ;
  assign n17355 = ~n17347 & n17354 ;
  assign n17356 = ~n17340 & ~n17355 ;
  assign n17357 = ~\u2_L6_reg[21]/NET0131  & n17356 ;
  assign n17358 = \u2_L6_reg[21]/NET0131  & ~n17356 ;
  assign n17359 = ~n17357 & ~n17358 ;
  assign n17360 = n16390 & n16667 ;
  assign n17361 = ~n16417 & ~n17360 ;
  assign n17362 = ~n16404 & ~n17361 ;
  assign n17363 = ~n16415 & ~n17362 ;
  assign n17364 = n16378 & ~n17363 ;
  assign n17365 = n16421 & n16429 ;
  assign n17366 = ~n16458 & ~n17365 ;
  assign n17367 = ~n16656 & n17366 ;
  assign n17368 = ~n17364 & n17367 ;
  assign n17369 = ~n16411 & ~n17368 ;
  assign n17383 = ~n16405 & ~n16651 ;
  assign n17384 = n16411 & ~n17383 ;
  assign n17382 = n16438 & n16451 ;
  assign n17385 = ~n16658 & ~n17382 ;
  assign n17386 = ~n17384 & n17385 ;
  assign n17387 = n16378 & ~n17386 ;
  assign n17370 = ~n16413 & ~n17360 ;
  assign n17371 = n16428 & ~n17370 ;
  assign n17373 = n16384 & ~n16411 ;
  assign n17374 = n16427 & n17373 ;
  assign n17372 = ~n16390 & n16443 ;
  assign n17377 = ~n16457 & ~n17372 ;
  assign n17378 = ~n17374 & n17377 ;
  assign n17375 = n16411 & n17360 ;
  assign n17376 = ~n16423 & ~n16442 ;
  assign n17379 = ~n17375 & n17376 ;
  assign n17380 = n17378 & n17379 ;
  assign n17381 = ~n16378 & ~n17380 ;
  assign n17388 = ~n17371 & ~n17381 ;
  assign n17389 = ~n17387 & n17388 ;
  assign n17390 = ~n17369 & n17389 ;
  assign n17391 = \u2_L6_reg[23]/NET0131  & ~n17390 ;
  assign n17392 = ~\u2_L6_reg[23]/NET0131  & n17390 ;
  assign n17393 = ~n17391 & ~n17392 ;
  assign n17414 = ~n17171 & ~n17181 ;
  assign n17415 = ~n17141 & ~n17414 ;
  assign n17413 = n17148 & n17170 ;
  assign n17416 = ~n17150 & ~n17413 ;
  assign n17417 = ~n17415 & n17416 ;
  assign n17418 = n17160 & ~n17417 ;
  assign n17394 = ~n17148 & n17170 ;
  assign n17419 = ~n17206 & ~n17394 ;
  assign n17420 = ~n17160 & ~n17419 ;
  assign n17406 = n17149 & n17168 ;
  assign n17421 = ~n17198 & ~n17406 ;
  assign n17422 = ~n17420 & n17421 ;
  assign n17423 = ~n17418 & n17422 ;
  assign n17424 = n17195 & ~n17423 ;
  assign n17395 = ~n17160 & ~n17394 ;
  assign n17400 = n17181 & n17395 ;
  assign n17398 = ~n17141 & ~n17168 ;
  assign n17399 = n17160 & n17398 ;
  assign n17401 = n17148 & ~n17182 ;
  assign n17402 = ~n17399 & n17401 ;
  assign n17403 = ~n17400 & n17402 ;
  assign n17396 = ~n17181 & n17395 ;
  assign n17397 = ~n17148 & ~n17396 ;
  assign n17404 = ~n17195 & ~n17397 ;
  assign n17405 = ~n17403 & n17404 ;
  assign n17407 = ~n17223 & ~n17406 ;
  assign n17408 = n17171 & n17178 ;
  assign n17409 = n17407 & ~n17408 ;
  assign n17410 = n17160 & ~n17409 ;
  assign n17411 = n17135 & ~n17160 ;
  assign n17412 = n17176 & n17411 ;
  assign n17425 = ~n17199 & ~n17412 ;
  assign n17426 = ~n17410 & n17425 ;
  assign n17427 = ~n17405 & n17426 ;
  assign n17428 = ~n17424 & n17427 ;
  assign n17429 = ~\u2_L6_reg[25]/NET0131  & ~n17428 ;
  assign n17430 = \u2_L6_reg[25]/NET0131  & n17428 ;
  assign n17431 = ~n17429 & ~n17430 ;
  assign n17440 = n16751 & n16759 ;
  assign n17441 = ~n16702 & ~n16720 ;
  assign n17442 = ~n17440 & n17441 ;
  assign n17443 = ~n16757 & ~n17442 ;
  assign n17445 = ~n16703 & ~n16717 ;
  assign n17446 = n16716 & ~n17445 ;
  assign n17444 = n16728 & n17306 ;
  assign n17447 = n16736 & ~n17444 ;
  assign n17448 = ~n17295 & n17447 ;
  assign n17449 = ~n17446 & n17448 ;
  assign n17450 = ~n17443 & n17449 ;
  assign n17453 = ~n16702 & n16750 ;
  assign n17454 = ~n16725 & ~n16736 ;
  assign n17455 = ~n17453 & n17454 ;
  assign n17451 = ~n16696 & n16709 ;
  assign n17452 = n16753 & n17451 ;
  assign n17456 = ~n16718 & ~n16739 ;
  assign n17457 = ~n17452 & n17456 ;
  assign n17458 = n17455 & n17457 ;
  assign n17459 = ~n17450 & ~n17458 ;
  assign n17432 = n16727 & ~n16736 ;
  assign n17433 = ~n16689 & ~n16729 ;
  assign n17434 = ~n16755 & ~n17433 ;
  assign n17435 = ~n16702 & ~n17434 ;
  assign n17436 = ~n17432 & ~n17435 ;
  assign n17437 = ~n16716 & ~n17436 ;
  assign n17438 = ~n16718 & ~n16747 ;
  assign n17439 = n16702 & ~n17438 ;
  assign n17460 = ~n17437 & ~n17439 ;
  assign n17461 = ~n17459 & n17460 ;
  assign n17462 = ~\u2_L6_reg[26]/NET0131  & ~n17461 ;
  assign n17463 = \u2_L6_reg[26]/NET0131  & n17461 ;
  assign n17464 = ~n17462 & ~n17463 ;
  assign n17467 = n16833 & n16871 ;
  assign n17468 = ~n16855 & n16896 ;
  assign n17469 = ~n17467 & ~n17468 ;
  assign n17470 = n16862 & n17469 ;
  assign n17474 = n16847 & ~n17117 ;
  assign n17471 = ~n16847 & n16863 ;
  assign n17472 = ~n16862 & ~n17093 ;
  assign n17473 = ~n17471 & n17472 ;
  assign n17475 = ~n16848 & n17473 ;
  assign n17476 = ~n17474 & n17475 ;
  assign n17477 = ~n17470 & ~n17476 ;
  assign n17465 = n16855 & ~n16885 ;
  assign n17466 = ~n17106 & n17465 ;
  assign n17478 = ~n16827 & ~n17466 ;
  assign n17479 = ~n17477 & n17478 ;
  assign n17483 = n17469 & n17473 ;
  assign n17484 = ~n16839 & ~n16887 ;
  assign n17485 = n16872 & ~n17484 ;
  assign n17486 = n16862 & ~n16885 ;
  assign n17487 = ~n17485 & n17486 ;
  assign n17488 = ~n17483 & ~n17487 ;
  assign n17480 = ~n16841 & ~n16862 ;
  assign n17481 = n16847 & ~n16855 ;
  assign n17482 = ~n17480 & n17481 ;
  assign n17489 = n16827 & ~n17095 ;
  assign n17490 = ~n17482 & n17489 ;
  assign n17491 = ~n17488 & n17490 ;
  assign n17492 = ~n17479 & ~n17491 ;
  assign n17493 = ~\u2_L6_reg[28]/NET0131  & n17492 ;
  assign n17494 = \u2_L6_reg[28]/NET0131  & ~n17492 ;
  assign n17495 = ~n17493 & ~n17494 ;
  assign n17507 = n17160 & ~n17201 ;
  assign n17508 = ~n17413 & n17507 ;
  assign n17509 = ~n17176 & n17178 ;
  assign n17510 = n17395 & ~n17509 ;
  assign n17511 = ~n17508 & ~n17510 ;
  assign n17512 = ~n17206 & n17407 ;
  assign n17513 = ~n17511 & n17512 ;
  assign n17514 = ~n17195 & ~n17513 ;
  assign n17497 = n17150 & n17398 ;
  assign n17498 = ~n17394 & ~n17497 ;
  assign n17499 = n17160 & ~n17498 ;
  assign n17500 = ~n17168 & n17411 ;
  assign n17501 = ~n17499 & ~n17500 ;
  assign n17502 = ~n17220 & n17501 ;
  assign n17503 = n17195 & ~n17502 ;
  assign n17496 = ~n17141 & n17412 ;
  assign n17504 = n17152 & n17197 ;
  assign n17505 = n17219 & ~n17504 ;
  assign n17506 = n17160 & ~n17505 ;
  assign n17515 = ~n17496 & ~n17506 ;
  assign n17516 = ~n17503 & n17515 ;
  assign n17517 = ~n17514 & n17516 ;
  assign n17518 = ~\u2_L6_reg[8]/NET0131  & ~n17517 ;
  assign n17519 = \u2_L6_reg[8]/NET0131  & n17517 ;
  assign n17520 = ~n17518 & ~n17519 ;
  assign n17523 = ~n17259 & ~n17324 ;
  assign n17524 = ~n17332 & n17523 ;
  assign n17525 = ~n16988 & ~n17524 ;
  assign n17521 = n16988 & ~n16996 ;
  assign n17522 = n17234 & n17521 ;
  assign n17526 = ~n16979 & ~n17331 ;
  assign n17527 = ~n17005 & n17526 ;
  assign n17528 = ~n17522 & n17527 ;
  assign n17529 = ~n17525 & n17528 ;
  assign n17530 = n16949 & ~n17529 ;
  assign n17531 = n16974 & ~n16997 ;
  assign n17532 = ~n16974 & n16997 ;
  assign n17533 = ~n17531 & ~n17532 ;
  assign n17534 = n17341 & n17533 ;
  assign n17535 = ~n16978 & ~n17534 ;
  assign n17536 = n16988 & ~n17535 ;
  assign n17538 = n16980 & n16991 ;
  assign n17537 = n16975 & n17244 ;
  assign n17539 = ~n17350 & ~n17537 ;
  assign n17540 = ~n17538 & n17539 ;
  assign n17541 = ~n16949 & ~n17540 ;
  assign n17542 = ~n17015 & ~n17242 ;
  assign n17543 = ~n16988 & ~n17006 ;
  assign n17544 = ~n17542 & n17543 ;
  assign n17545 = ~n17541 & ~n17544 ;
  assign n17546 = ~n17536 & n17545 ;
  assign n17547 = ~n17530 & n17546 ;
  assign n17548 = ~\u2_L6_reg[27]/NET0131  & ~n17547 ;
  assign n17549 = \u2_L6_reg[27]/NET0131  & n17547 ;
  assign n17550 = ~n17548 & ~n17549 ;
  assign n17554 = n17075 & ~n17077 ;
  assign n17555 = n16609 & n17078 ;
  assign n17556 = ~n17554 & ~n17555 ;
  assign n17557 = ~n16606 & ~n17556 ;
  assign n17551 = ~n16577 & ~n16606 ;
  assign n17552 = n16583 & ~n17551 ;
  assign n17553 = n16598 & n17552 ;
  assign n17558 = n16584 & ~n16596 ;
  assign n17559 = ~n16613 & ~n17558 ;
  assign n17560 = n16606 & ~n17559 ;
  assign n17561 = ~n17553 & ~n17560 ;
  assign n17562 = ~n17557 & n17561 ;
  assign n17563 = n16571 & ~n17562 ;
  assign n17566 = ~n16590 & n17076 ;
  assign n17567 = n17084 & ~n17566 ;
  assign n17568 = n17077 & n17079 ;
  assign n17569 = ~n16598 & ~n16633 ;
  assign n17570 = n17552 & n17569 ;
  assign n17571 = ~n17568 & ~n17570 ;
  assign n17572 = ~n17567 & n17571 ;
  assign n17573 = ~n16571 & ~n17572 ;
  assign n17564 = n16571 & ~n16606 ;
  assign n17565 = n17062 & ~n17564 ;
  assign n17574 = n16639 & ~n17076 ;
  assign n17575 = ~n16638 & n17574 ;
  assign n17576 = ~n17565 & ~n17575 ;
  assign n17577 = ~n17573 & n17576 ;
  assign n17578 = ~n17563 & n17577 ;
  assign n17579 = \u2_L6_reg[32]/NET0131  & n17578 ;
  assign n17580 = ~\u2_L6_reg[32]/NET0131  & ~n17578 ;
  assign n17581 = ~n17579 & ~n17580 ;
  assign n17582 = ~n17142 & n17176 ;
  assign n17583 = ~n17195 & ~n17582 ;
  assign n17584 = ~n17212 & ~n17394 ;
  assign n17585 = n17583 & n17584 ;
  assign n17586 = ~n17177 & n17195 ;
  assign n17587 = ~n17153 & ~n17199 ;
  assign n17588 = n17586 & n17587 ;
  assign n17589 = ~n17585 & ~n17588 ;
  assign n17590 = n17168 & n17394 ;
  assign n17591 = ~n17160 & ~n17497 ;
  assign n17592 = ~n17222 & n17591 ;
  assign n17593 = ~n17590 & n17592 ;
  assign n17594 = ~n17589 & n17593 ;
  assign n17595 = ~n17178 & ~n17207 ;
  assign n17596 = n17586 & ~n17595 ;
  assign n17597 = ~n17168 & n17178 ;
  assign n17598 = ~n17149 & ~n17597 ;
  assign n17599 = n17583 & n17598 ;
  assign n17600 = ~n17596 & ~n17599 ;
  assign n17601 = ~n17218 & n17507 ;
  assign n17602 = ~n17600 & n17601 ;
  assign n17603 = ~n17594 & ~n17602 ;
  assign n17604 = ~\u2_L6_reg[3]/NET0131  & n17603 ;
  assign n17605 = \u2_L6_reg[3]/NET0131  & ~n17603 ;
  assign n17606 = ~n17604 & ~n17605 ;
  assign n17607 = decrypt_pad & ~\u2_uk_K_r6_reg[46]/NET0131  ;
  assign n17608 = ~decrypt_pad & ~\u2_uk_K_r6_reg[39]/NET0131  ;
  assign n17609 = ~n17607 & ~n17608 ;
  assign n17610 = \u2_R6_reg[13]/NET0131  & ~n17609 ;
  assign n17611 = ~\u2_R6_reg[13]/NET0131  & n17609 ;
  assign n17612 = ~n17610 & ~n17611 ;
  assign n17620 = decrypt_pad & ~\u2_uk_K_r6_reg[41]/NET0131  ;
  assign n17621 = ~decrypt_pad & ~\u2_uk_K_r6_reg[34]/NET0131  ;
  assign n17622 = ~n17620 & ~n17621 ;
  assign n17623 = \u2_R6_reg[9]/NET0131  & ~n17622 ;
  assign n17624 = ~\u2_R6_reg[9]/NET0131  & n17622 ;
  assign n17625 = ~n17623 & ~n17624 ;
  assign n17634 = ~n17612 & n17625 ;
  assign n17635 = decrypt_pad & ~\u2_uk_K_r6_reg[18]/NET0131  ;
  assign n17636 = ~decrypt_pad & ~\u2_uk_K_r6_reg[11]/NET0131  ;
  assign n17637 = ~n17635 & ~n17636 ;
  assign n17638 = \u2_R6_reg[11]/NET0131  & ~n17637 ;
  assign n17639 = ~\u2_R6_reg[11]/NET0131  & n17637 ;
  assign n17640 = ~n17638 & ~n17639 ;
  assign n17641 = ~n17634 & ~n17640 ;
  assign n17626 = decrypt_pad & ~\u2_uk_K_r6_reg[17]/NET0131  ;
  assign n17627 = ~decrypt_pad & ~\u2_uk_K_r6_reg[10]/NET0131  ;
  assign n17628 = ~n17626 & ~n17627 ;
  assign n17629 = \u2_R6_reg[10]/NET0131  & ~n17628 ;
  assign n17630 = ~\u2_R6_reg[10]/NET0131  & n17628 ;
  assign n17631 = ~n17629 & ~n17630 ;
  assign n17642 = n17625 & ~n17631 ;
  assign n17613 = decrypt_pad & ~\u2_uk_K_r6_reg[12]/NET0131  ;
  assign n17614 = ~decrypt_pad & ~\u2_uk_K_r6_reg[5]/NET0131  ;
  assign n17615 = ~n17613 & ~n17614 ;
  assign n17616 = \u2_R6_reg[8]/NET0131  & ~n17615 ;
  assign n17617 = ~\u2_R6_reg[8]/NET0131  & n17615 ;
  assign n17618 = ~n17616 & ~n17617 ;
  assign n17643 = n17612 & ~n17625 ;
  assign n17644 = n17618 & ~n17643 ;
  assign n17645 = ~n17642 & ~n17644 ;
  assign n17646 = n17641 & ~n17645 ;
  assign n17619 = ~n17612 & ~n17618 ;
  assign n17632 = n17625 & n17631 ;
  assign n17633 = n17619 & n17632 ;
  assign n17647 = decrypt_pad & ~\u2_uk_K_r6_reg[33]/NET0131  ;
  assign n17648 = ~decrypt_pad & ~\u2_uk_K_r6_reg[26]/NET0131  ;
  assign n17649 = ~n17647 & ~n17648 ;
  assign n17650 = \u2_R6_reg[12]/NET0131  & ~n17649 ;
  assign n17651 = ~\u2_R6_reg[12]/NET0131  & n17649 ;
  assign n17652 = ~n17650 & ~n17651 ;
  assign n17653 = ~n17633 & n17652 ;
  assign n17654 = ~n17646 & n17653 ;
  assign n17659 = n17612 & n17618 ;
  assign n17660 = ~n17619 & ~n17659 ;
  assign n17661 = ~n17625 & ~n17631 ;
  assign n17664 = ~n17660 & ~n17661 ;
  assign n17665 = ~n17632 & n17664 ;
  assign n17667 = n17618 & n17631 ;
  assign n17668 = n17634 & n17667 ;
  assign n17658 = ~n17618 & n17640 ;
  assign n17666 = n17642 & n17658 ;
  assign n17669 = ~n17652 & ~n17666 ;
  assign n17670 = ~n17668 & n17669 ;
  assign n17655 = n17612 & ~n17618 ;
  assign n17656 = n17632 & n17655 ;
  assign n17657 = ~n17640 & n17656 ;
  assign n17662 = ~n17658 & n17661 ;
  assign n17663 = n17660 & n17662 ;
  assign n17671 = ~n17657 & ~n17663 ;
  assign n17672 = n17670 & n17671 ;
  assign n17673 = ~n17665 & n17672 ;
  assign n17674 = ~n17654 & ~n17673 ;
  assign n17676 = ~n17618 & ~n17631 ;
  assign n17677 = n17618 & ~n17625 ;
  assign n17678 = ~n17676 & ~n17677 ;
  assign n17679 = n17660 & n17678 ;
  assign n17680 = ~n17643 & ~n17679 ;
  assign n17681 = n17652 & ~n17680 ;
  assign n17675 = n17631 & n17643 ;
  assign n17682 = n17619 & ~n17631 ;
  assign n17683 = ~n17625 & n17682 ;
  assign n17684 = ~n17675 & ~n17683 ;
  assign n17685 = ~n17681 & n17684 ;
  assign n17686 = n17640 & ~n17685 ;
  assign n17687 = ~n17674 & ~n17686 ;
  assign n17688 = ~\u2_L6_reg[6]/NET0131  & ~n17687 ;
  assign n17689 = \u2_L6_reg[6]/NET0131  & n17687 ;
  assign n17690 = ~n17688 & ~n17689 ;
  assign n17692 = ~n16598 & n17077 ;
  assign n17693 = ~n17079 & ~n17692 ;
  assign n17691 = ~n16571 & n16606 ;
  assign n17694 = ~n17568 & n17691 ;
  assign n17695 = ~n17693 & n17694 ;
  assign n17696 = ~n17077 & ~n17079 ;
  assign n17697 = ~n16631 & ~n17568 ;
  assign n17698 = ~n17696 & n17697 ;
  assign n17699 = ~n17564 & ~n17691 ;
  assign n17700 = ~n17698 & n17699 ;
  assign n17701 = ~n17695 & ~n17700 ;
  assign n17702 = n16590 & n17558 ;
  assign n17703 = ~n17701 & ~n17702 ;
  assign n17704 = n16577 & ~n17692 ;
  assign n17705 = ~n16577 & n16638 ;
  assign n17706 = n17564 & ~n17705 ;
  assign n17707 = ~n17704 & n17706 ;
  assign n17708 = ~n17703 & ~n17707 ;
  assign n17709 = ~\u2_L6_reg[7]/NET0131  & n17708 ;
  assign n17710 = \u2_L6_reg[7]/NET0131  & ~n17708 ;
  assign n17711 = ~n17709 & ~n17710 ;
  assign n17727 = n16673 & ~n17362 ;
  assign n17728 = n16384 & ~n17727 ;
  assign n17719 = n16390 & ~n16421 ;
  assign n17720 = ~n16417 & ~n17719 ;
  assign n17726 = n16428 & n17720 ;
  assign n17729 = ~n16656 & ~n17726 ;
  assign n17730 = ~n17728 & n17729 ;
  assign n17731 = n16378 & ~n17730 ;
  assign n17712 = ~n16384 & n16672 ;
  assign n17713 = n16384 & n16651 ;
  assign n17714 = ~n17712 & ~n17713 ;
  assign n17715 = ~n16411 & ~n17714 ;
  assign n17717 = ~n16398 & n17361 ;
  assign n17718 = n16411 & ~n17717 ;
  assign n17721 = ~n16411 & n17720 ;
  assign n17716 = n16384 & n16669 ;
  assign n17722 = ~n17712 & ~n17716 ;
  assign n17723 = ~n17721 & n17722 ;
  assign n17724 = ~n17718 & n17723 ;
  assign n17725 = ~n16378 & ~n17724 ;
  assign n17732 = ~n17715 & ~n17725 ;
  assign n17733 = ~n17731 & n17732 ;
  assign n17734 = ~\u2_L6_reg[9]/NET0131  & ~n17733 ;
  assign n17735 = \u2_L6_reg[9]/NET0131  & n17733 ;
  assign n17736 = ~n17734 & ~n17735 ;
  assign n17739 = n17625 & ~n17659 ;
  assign n17740 = ~n17625 & n17659 ;
  assign n17741 = ~n17739 & ~n17740 ;
  assign n17742 = ~n17619 & n17741 ;
  assign n17743 = n17634 & n17658 ;
  assign n17744 = ~n17742 & ~n17743 ;
  assign n17745 = ~n17631 & ~n17744 ;
  assign n17746 = ~n17640 & ~n17667 ;
  assign n17747 = ~n17612 & ~n17676 ;
  assign n17748 = n17746 & n17747 ;
  assign n17749 = ~n17656 & ~n17748 ;
  assign n17750 = ~n17745 & n17749 ;
  assign n17751 = n17652 & ~n17750 ;
  assign n17752 = ~n17619 & n17640 ;
  assign n17753 = ~n17741 & n17752 ;
  assign n17754 = n17640 & ~n17683 ;
  assign n17755 = ~n17625 & ~n17655 ;
  assign n17756 = ~n17739 & ~n17755 ;
  assign n17757 = ~n17682 & ~n17756 ;
  assign n17758 = ~n17754 & ~n17757 ;
  assign n17759 = ~n17753 & ~n17758 ;
  assign n17760 = ~n17652 & ~n17759 ;
  assign n17737 = ~n17640 & n17667 ;
  assign n17738 = ~n17625 & n17737 ;
  assign n17761 = n17619 & n17631 ;
  assign n17762 = ~n17625 & n17761 ;
  assign n17763 = ~n17668 & ~n17762 ;
  assign n17764 = n17640 & ~n17763 ;
  assign n17765 = ~n17738 & ~n17764 ;
  assign n17766 = ~n17760 & n17765 ;
  assign n17767 = ~n17751 & n17766 ;
  assign n17768 = ~\u2_L6_reg[16]/NET0131  & ~n17767 ;
  assign n17769 = \u2_L6_reg[16]/NET0131  & n17767 ;
  assign n17770 = ~n17768 & ~n17769 ;
  assign n17774 = ~n16885 & ~n16890 ;
  assign n17775 = ~n16862 & ~n17774 ;
  assign n17772 = n16863 & n16896 ;
  assign n17773 = ~n16849 & n16862 ;
  assign n17776 = ~n17772 & ~n17773 ;
  assign n17777 = ~n17775 & n17776 ;
  assign n17778 = n16827 & ~n17777 ;
  assign n17780 = ~n16874 & ~n16888 ;
  assign n17781 = n16895 & n17780 ;
  assign n17782 = ~n16865 & ~n17093 ;
  assign n17779 = n16864 & n16888 ;
  assign n17783 = ~n17113 & ~n17779 ;
  assign n17784 = n17782 & n17783 ;
  assign n17785 = ~n17781 & n17784 ;
  assign n17786 = ~n16827 & ~n17785 ;
  assign n17771 = ~n16862 & n17467 ;
  assign n17787 = n16839 & n16867 ;
  assign n17788 = ~n17119 & ~n17787 ;
  assign n17789 = n16862 & ~n17788 ;
  assign n17790 = ~n17771 & ~n17789 ;
  assign n17791 = ~n17786 & n17790 ;
  assign n17792 = ~n17778 & n17791 ;
  assign n17793 = ~\u2_L6_reg[18]/P0001  & ~n17792 ;
  assign n17794 = \u2_L6_reg[18]/P0001  & n17792 ;
  assign n17795 = ~n17793 & ~n17794 ;
  assign n17803 = ~n17631 & n17655 ;
  assign n17804 = ~n17761 & ~n17803 ;
  assign n17805 = n17631 & n17677 ;
  assign n17802 = n17619 & n17625 ;
  assign n17806 = n17640 & ~n17802 ;
  assign n17807 = ~n17805 & n17806 ;
  assign n17808 = n17804 & n17807 ;
  assign n17811 = ~n17660 & n17661 ;
  assign n17809 = ~n17631 & ~n17634 ;
  assign n17810 = n17660 & ~n17809 ;
  assign n17812 = ~n17640 & ~n17810 ;
  assign n17813 = ~n17811 & n17812 ;
  assign n17814 = ~n17808 & ~n17813 ;
  assign n17815 = ~n17652 & ~n17814 ;
  assign n17816 = ~n17640 & n17664 ;
  assign n17820 = n17652 & ~n17663 ;
  assign n17817 = n17631 & ~n17677 ;
  assign n17818 = n17752 & n17817 ;
  assign n17798 = ~n17631 & n17640 ;
  assign n17819 = n17755 & n17798 ;
  assign n17821 = ~n17818 & ~n17819 ;
  assign n17822 = n17820 & n17821 ;
  assign n17823 = ~n17816 & n17822 ;
  assign n17824 = ~n17815 & ~n17823 ;
  assign n17796 = n17612 & n17625 ;
  assign n17797 = ~n17677 & ~n17796 ;
  assign n17799 = ~n17659 & n17798 ;
  assign n17800 = ~n17797 & n17799 ;
  assign n17801 = n17737 & n17796 ;
  assign n17825 = ~n17800 & ~n17801 ;
  assign n17826 = ~n17824 & n17825 ;
  assign n17827 = ~\u2_L6_reg[24]/NET0131  & ~n17826 ;
  assign n17828 = \u2_L6_reg[24]/NET0131  & n17826 ;
  assign n17829 = ~n17827 & ~n17828 ;
  assign n17846 = ~n17634 & n17667 ;
  assign n17841 = ~n17612 & ~n17631 ;
  assign n17845 = n17625 & n17841 ;
  assign n17847 = ~n17652 & ~n17845 ;
  assign n17848 = ~n17846 & n17847 ;
  assign n17842 = n17677 & n17841 ;
  assign n17843 = n17652 & ~n17842 ;
  assign n17844 = n17804 & n17843 ;
  assign n17849 = n17640 & ~n17844 ;
  assign n17850 = ~n17848 & n17849 ;
  assign n17831 = ~n17667 & ~n17802 ;
  assign n17832 = ~n17640 & ~n17831 ;
  assign n17830 = n17631 & n17739 ;
  assign n17833 = n17652 & ~n17830 ;
  assign n17834 = ~n17832 & n17833 ;
  assign n17837 = ~n17652 & ~n17811 ;
  assign n17835 = ~n17618 & n17675 ;
  assign n17836 = n17746 & ~n17797 ;
  assign n17838 = ~n17835 & ~n17836 ;
  assign n17839 = n17837 & n17838 ;
  assign n17840 = ~n17834 & ~n17839 ;
  assign n17851 = n17640 & ~n17740 ;
  assign n17852 = n17631 & ~n17641 ;
  assign n17853 = ~n17851 & n17852 ;
  assign n17854 = ~n17840 & ~n17853 ;
  assign n17855 = ~n17850 & n17854 ;
  assign n17856 = \u2_L6_reg[30]/NET0131  & ~n17855 ;
  assign n17857 = ~\u2_L6_reg[30]/NET0131  & n17855 ;
  assign n17858 = ~n17856 & ~n17857 ;
  assign n17882 = decrypt_pad & ~\u2_uk_K_r5_reg[44]/NET0131  ;
  assign n17883 = ~decrypt_pad & ~\u2_uk_K_r5_reg[9]/P0001  ;
  assign n17884 = ~n17882 & ~n17883 ;
  assign n17885 = \u2_R5_reg[28]/NET0131  & ~n17884 ;
  assign n17886 = ~\u2_R5_reg[28]/NET0131  & n17884 ;
  assign n17887 = ~n17885 & ~n17886 ;
  assign n17902 = decrypt_pad & ~\u2_uk_K_r5_reg[2]/NET0131  ;
  assign n17903 = ~decrypt_pad & ~\u2_uk_K_r5_reg[22]/NET0131  ;
  assign n17904 = ~n17902 & ~n17903 ;
  assign n17905 = \u2_R5_reg[27]/NET0131  & ~n17904 ;
  assign n17906 = ~\u2_R5_reg[27]/NET0131  & n17904 ;
  assign n17907 = ~n17905 & ~n17906 ;
  assign n17872 = decrypt_pad & ~\u2_uk_K_r5_reg[52]/NET0131  ;
  assign n17873 = ~decrypt_pad & ~\u2_uk_K_r5_reg[44]/NET0131  ;
  assign n17874 = ~n17872 & ~n17873 ;
  assign n17875 = \u2_R5_reg[26]/NET0131  & ~n17874 ;
  assign n17876 = ~\u2_R5_reg[26]/NET0131  & n17874 ;
  assign n17877 = ~n17875 & ~n17876 ;
  assign n17859 = decrypt_pad & ~\u2_uk_K_r5_reg[28]/NET0131  ;
  assign n17860 = ~decrypt_pad & ~\u2_uk_K_r5_reg[52]/NET0131  ;
  assign n17861 = ~n17859 & ~n17860 ;
  assign n17862 = \u2_R5_reg[24]/NET0131  & ~n17861 ;
  assign n17863 = ~\u2_R5_reg[24]/NET0131  & n17861 ;
  assign n17864 = ~n17862 & ~n17863 ;
  assign n17888 = decrypt_pad & ~\u2_uk_K_r5_reg[36]/NET0131  ;
  assign n17889 = ~decrypt_pad & ~\u2_uk_K_r5_reg[1]/NET0131  ;
  assign n17890 = ~n17888 & ~n17889 ;
  assign n17891 = \u2_R5_reg[29]/NET0131  & ~n17890 ;
  assign n17892 = ~\u2_R5_reg[29]/NET0131  & n17890 ;
  assign n17893 = ~n17891 & ~n17892 ;
  assign n17894 = n17864 & n17893 ;
  assign n17865 = decrypt_pad & ~\u2_uk_K_r5_reg[8]/NET0131  ;
  assign n17866 = ~decrypt_pad & ~\u2_uk_K_r5_reg[28]/NET0131  ;
  assign n17867 = ~n17865 & ~n17866 ;
  assign n17868 = \u2_R5_reg[25]/NET0131  & ~n17867 ;
  assign n17869 = ~\u2_R5_reg[25]/NET0131  & n17867 ;
  assign n17870 = ~n17868 & ~n17869 ;
  assign n17924 = ~n17864 & ~n17893 ;
  assign n17934 = ~n17870 & n17924 ;
  assign n17935 = ~n17894 & ~n17934 ;
  assign n17936 = n17877 & ~n17935 ;
  assign n17937 = n17864 & ~n17893 ;
  assign n17938 = n17870 & n17937 ;
  assign n17939 = ~n17936 & ~n17938 ;
  assign n17940 = ~n17907 & ~n17939 ;
  assign n17909 = ~n17864 & n17893 ;
  assign n17930 = ~n17907 & n17909 ;
  assign n17920 = n17864 & n17907 ;
  assign n17931 = ~n17870 & n17920 ;
  assign n17932 = ~n17930 & ~n17931 ;
  assign n17933 = ~n17877 & ~n17932 ;
  assign n17871 = n17864 & n17870 ;
  assign n17878 = n17871 & n17877 ;
  assign n17879 = n17870 & ~n17877 ;
  assign n17880 = ~n17864 & n17879 ;
  assign n17881 = ~n17878 & ~n17880 ;
  assign n17929 = ~n17881 & n17893 ;
  assign n17941 = ~n17877 & n17937 ;
  assign n17942 = ~n17870 & n17941 ;
  assign n17943 = ~n17929 & ~n17942 ;
  assign n17944 = ~n17933 & n17943 ;
  assign n17945 = ~n17940 & n17944 ;
  assign n17946 = ~n17887 & ~n17945 ;
  assign n17910 = ~n17870 & n17877 ;
  assign n17897 = n17870 & n17893 ;
  assign n17921 = ~n17877 & n17897 ;
  assign n17922 = ~n17910 & ~n17921 ;
  assign n17923 = n17920 & ~n17922 ;
  assign n17911 = n17909 & n17910 ;
  assign n17895 = ~n17870 & ~n17877 ;
  assign n17925 = n17895 & n17924 ;
  assign n17926 = ~n17911 & ~n17925 ;
  assign n17927 = ~n17923 & n17926 ;
  assign n17928 = n17887 & ~n17927 ;
  assign n17896 = n17894 & n17895 ;
  assign n17898 = ~n17864 & n17897 ;
  assign n17899 = ~n17896 & ~n17898 ;
  assign n17900 = n17887 & ~n17899 ;
  assign n17901 = n17881 & ~n17900 ;
  assign n17908 = ~n17901 & ~n17907 ;
  assign n17912 = ~n17864 & n17877 ;
  assign n17913 = n17870 & n17912 ;
  assign n17914 = ~n17893 & n17913 ;
  assign n17915 = ~n17911 & ~n17914 ;
  assign n17916 = ~n17870 & ~n17893 ;
  assign n17917 = ~n17912 & n17916 ;
  assign n17918 = n17915 & ~n17917 ;
  assign n17919 = n17907 & ~n17918 ;
  assign n17947 = ~n17908 & ~n17919 ;
  assign n17948 = ~n17928 & n17947 ;
  assign n17949 = ~n17946 & n17948 ;
  assign n17950 = ~\u2_L5_reg[22]/NET0131  & ~n17949 ;
  assign n17951 = \u2_L5_reg[22]/NET0131  & n17949 ;
  assign n17952 = ~n17950 & ~n17951 ;
  assign n17953 = decrypt_pad & ~\u2_uk_K_r5_reg[11]/NET0131  ;
  assign n17954 = ~decrypt_pad & ~\u2_uk_K_r5_reg[33]/NET0131  ;
  assign n17955 = ~n17953 & ~n17954 ;
  assign n17956 = \u2_R5_reg[4]/NET0131  & ~n17955 ;
  assign n17957 = ~\u2_R5_reg[4]/NET0131  & n17955 ;
  assign n17958 = ~n17956 & ~n17957 ;
  assign n17959 = decrypt_pad & ~\u2_uk_K_r5_reg[33]/NET0131  ;
  assign n17960 = ~decrypt_pad & ~\u2_uk_K_r5_reg[55]/NET0131  ;
  assign n17961 = ~n17959 & ~n17960 ;
  assign n17962 = \u2_R5_reg[3]/NET0131  & ~n17961 ;
  assign n17963 = ~\u2_R5_reg[3]/NET0131  & n17961 ;
  assign n17964 = ~n17962 & ~n17963 ;
  assign n17972 = decrypt_pad & ~\u2_uk_K_r5_reg[41]/NET0131  ;
  assign n17973 = ~decrypt_pad & ~\u2_uk_K_r5_reg[6]/NET0131  ;
  assign n17974 = ~n17972 & ~n17973 ;
  assign n17975 = \u2_R5_reg[1]/NET0131  & ~n17974 ;
  assign n17976 = ~\u2_R5_reg[1]/NET0131  & n17974 ;
  assign n17977 = ~n17975 & ~n17976 ;
  assign n17978 = decrypt_pad & ~\u2_uk_K_r5_reg[39]/NET0131  ;
  assign n17979 = ~decrypt_pad & ~\u2_uk_K_r5_reg[4]/NET0131  ;
  assign n17980 = ~n17978 & ~n17979 ;
  assign n17981 = \u2_R5_reg[5]/NET0131  & ~n17980 ;
  assign n17982 = ~\u2_R5_reg[5]/NET0131  & n17980 ;
  assign n17983 = ~n17981 & ~n17982 ;
  assign n17998 = ~n17977 & n17983 ;
  assign n17965 = decrypt_pad & ~\u2_uk_K_r5_reg[24]/NET0131  ;
  assign n17966 = ~decrypt_pad & ~\u2_uk_K_r5_reg[46]/NET0131  ;
  assign n17967 = ~n17965 & ~n17966 ;
  assign n17968 = \u2_R5_reg[2]/NET0131  & ~n17967 ;
  assign n17969 = ~\u2_R5_reg[2]/NET0131  & n17967 ;
  assign n17970 = ~n17968 & ~n17969 ;
  assign n17984 = decrypt_pad & ~\u2_uk_K_r5_reg[20]/NET0131  ;
  assign n17985 = ~decrypt_pad & ~\u2_uk_K_r5_reg[10]/NET0131  ;
  assign n17986 = ~n17984 & ~n17985 ;
  assign n17987 = \u2_R5_reg[32]/NET0131  & ~n17986 ;
  assign n17988 = ~\u2_R5_reg[32]/NET0131  & n17986 ;
  assign n17989 = ~n17987 & ~n17988 ;
  assign n17991 = ~n17983 & ~n17989 ;
  assign n18027 = n17970 & n17991 ;
  assign n18028 = ~n17998 & ~n18027 ;
  assign n18029 = n17964 & ~n18028 ;
  assign n18019 = n17983 & ~n17989 ;
  assign n18012 = n17964 & ~n17970 ;
  assign n18032 = n17977 & ~n18012 ;
  assign n18033 = n18019 & ~n18032 ;
  assign n18003 = ~n17964 & n17989 ;
  assign n18004 = n17977 & ~n18003 ;
  assign n17999 = ~n17970 & ~n17989 ;
  assign n18011 = ~n17977 & n17989 ;
  assign n18030 = ~n17999 & ~n18011 ;
  assign n18031 = ~n18004 & n18030 ;
  assign n18034 = ~n17970 & n17989 ;
  assign n18035 = ~n17977 & ~n17983 ;
  assign n18036 = n18034 & n18035 ;
  assign n18037 = ~n18031 & ~n18036 ;
  assign n18038 = ~n18033 & n18037 ;
  assign n18039 = ~n18029 & n18038 ;
  assign n18040 = n17958 & ~n18039 ;
  assign n18005 = ~n17998 & ~n18004 ;
  assign n17990 = n17983 & n17989 ;
  assign n17992 = ~n17990 & ~n17991 ;
  assign n18006 = ~n17970 & ~n17992 ;
  assign n18007 = ~n18005 & n18006 ;
  assign n17971 = n17964 & n17970 ;
  assign n17993 = n17977 & n17992 ;
  assign n17994 = n17971 & n17993 ;
  assign n17995 = n17970 & ~n17977 ;
  assign n17996 = ~n17983 & n17989 ;
  assign n17997 = n17995 & n17996 ;
  assign n18000 = ~n17998 & n17999 ;
  assign n18001 = ~n17997 & ~n18000 ;
  assign n18002 = ~n17964 & ~n18001 ;
  assign n18008 = ~n17994 & ~n18002 ;
  assign n18009 = ~n18007 & n18008 ;
  assign n18010 = ~n17958 & ~n18009 ;
  assign n18020 = ~n17977 & n18019 ;
  assign n18021 = n17970 & n18020 ;
  assign n18016 = n17970 & n17977 ;
  assign n18017 = n17983 & n18016 ;
  assign n18018 = n17989 & n18017 ;
  assign n18022 = ~n17970 & n17977 ;
  assign n18023 = ~n17983 & n18022 ;
  assign n18024 = ~n18018 & ~n18023 ;
  assign n18025 = ~n18021 & n18024 ;
  assign n18026 = ~n17964 & ~n18025 ;
  assign n18013 = n18011 & n18012 ;
  assign n18014 = n17964 & n17991 ;
  assign n18015 = n17995 & n18014 ;
  assign n18041 = ~n18013 & ~n18015 ;
  assign n18042 = ~n18026 & n18041 ;
  assign n18043 = ~n18010 & n18042 ;
  assign n18044 = ~n18040 & n18043 ;
  assign n18045 = ~\u2_L5_reg[31]/NET0131  & ~n18044 ;
  assign n18046 = \u2_L5_reg[31]/NET0131  & n18044 ;
  assign n18047 = ~n18045 & ~n18046 ;
  assign n18099 = decrypt_pad & ~\u2_uk_K_r5_reg[37]/P0001  ;
  assign n18100 = ~decrypt_pad & ~\u2_uk_K_r5_reg[2]/NET0131  ;
  assign n18101 = ~n18099 & ~n18100 ;
  assign n18102 = \u2_R5_reg[24]/NET0131  & ~n18101 ;
  assign n18103 = ~\u2_R5_reg[24]/NET0131  & n18101 ;
  assign n18104 = ~n18102 & ~n18103 ;
  assign n18054 = decrypt_pad & ~\u2_uk_K_r5_reg[16]/NET0131  ;
  assign n18055 = ~decrypt_pad & ~\u2_uk_K_r5_reg[36]/NET0131  ;
  assign n18056 = ~n18054 & ~n18055 ;
  assign n18057 = \u2_R5_reg[20]/NET0131  & ~n18056 ;
  assign n18058 = ~\u2_R5_reg[20]/NET0131  & n18056 ;
  assign n18059 = ~n18057 & ~n18058 ;
  assign n18067 = decrypt_pad & ~\u2_uk_K_r5_reg[22]/NET0131  ;
  assign n18068 = ~decrypt_pad & ~\u2_uk_K_r5_reg[42]/NET0131  ;
  assign n18069 = ~n18067 & ~n18068 ;
  assign n18070 = \u2_R5_reg[22]/NET0131  & ~n18069 ;
  assign n18071 = ~\u2_R5_reg[22]/NET0131  & n18069 ;
  assign n18072 = ~n18070 & ~n18071 ;
  assign n18073 = decrypt_pad & ~\u2_uk_K_r5_reg[0]/NET0131  ;
  assign n18074 = ~decrypt_pad & ~\u2_uk_K_r5_reg[51]/NET0131  ;
  assign n18075 = ~n18073 & ~n18074 ;
  assign n18076 = \u2_R5_reg[21]/NET0131  & ~n18075 ;
  assign n18077 = ~\u2_R5_reg[21]/NET0131  & n18075 ;
  assign n18078 = ~n18076 & ~n18077 ;
  assign n18108 = ~n18072 & n18078 ;
  assign n18124 = n18059 & n18108 ;
  assign n18048 = decrypt_pad & ~\u2_uk_K_r5_reg[35]/NET0131  ;
  assign n18049 = ~decrypt_pad & ~\u2_uk_K_r5_reg[0]/NET0131  ;
  assign n18050 = ~n18048 & ~n18049 ;
  assign n18051 = \u2_R5_reg[23]/NET0131  & ~n18050 ;
  assign n18052 = ~\u2_R5_reg[23]/NET0131  & n18050 ;
  assign n18053 = ~n18051 & ~n18052 ;
  assign n18081 = ~n18059 & n18078 ;
  assign n18082 = n18072 & n18081 ;
  assign n18125 = ~n18053 & ~n18082 ;
  assign n18126 = ~n18124 & n18125 ;
  assign n18060 = decrypt_pad & ~\u2_uk_K_r5_reg[1]/NET0131  ;
  assign n18061 = ~decrypt_pad & ~\u2_uk_K_r5_reg[21]/NET0131  ;
  assign n18062 = ~n18060 & ~n18061 ;
  assign n18063 = \u2_R5_reg[25]/NET0131  & ~n18062 ;
  assign n18064 = ~\u2_R5_reg[25]/NET0131  & n18062 ;
  assign n18065 = ~n18063 & ~n18064 ;
  assign n18116 = n18065 & ~n18078 ;
  assign n18117 = ~n18059 & n18116 ;
  assign n18118 = n18053 & ~n18117 ;
  assign n18127 = n18072 & ~n18078 ;
  assign n18128 = n18059 & n18127 ;
  assign n18129 = ~n18059 & ~n18072 ;
  assign n18130 = ~n18128 & ~n18129 ;
  assign n18131 = n18118 & n18130 ;
  assign n18132 = ~n18126 & ~n18131 ;
  assign n18083 = n18059 & n18065 ;
  assign n18094 = ~n18078 & n18083 ;
  assign n18121 = n18072 & n18094 ;
  assign n18066 = n18059 & ~n18065 ;
  assign n18088 = ~n18053 & ~n18072 ;
  assign n18122 = ~n18088 & ~n18108 ;
  assign n18123 = n18066 & ~n18122 ;
  assign n18133 = ~n18121 & ~n18123 ;
  assign n18134 = ~n18132 & n18133 ;
  assign n18135 = ~n18104 & ~n18134 ;
  assign n18084 = n18078 & n18083 ;
  assign n18079 = ~n18072 & ~n18078 ;
  assign n18080 = n18066 & n18079 ;
  assign n18085 = ~n18080 & ~n18082 ;
  assign n18086 = ~n18084 & n18085 ;
  assign n18087 = n18053 & ~n18086 ;
  assign n18089 = ~n18081 & ~n18083 ;
  assign n18090 = ~n18053 & n18089 ;
  assign n18091 = ~n18088 & ~n18090 ;
  assign n18092 = n18065 & n18078 ;
  assign n18093 = ~n18059 & n18092 ;
  assign n18095 = ~n18072 & ~n18093 ;
  assign n18096 = ~n18094 & n18095 ;
  assign n18097 = ~n18091 & ~n18096 ;
  assign n18098 = ~n18087 & ~n18097 ;
  assign n18105 = ~n18098 & n18104 ;
  assign n18114 = n18066 & n18078 ;
  assign n18115 = ~n18053 & ~n18114 ;
  assign n18119 = ~n18072 & ~n18115 ;
  assign n18120 = ~n18118 & n18119 ;
  assign n18109 = ~n18083 & ~n18108 ;
  assign n18106 = ~n18059 & ~n18065 ;
  assign n18107 = ~n18072 & ~n18106 ;
  assign n18110 = n18053 & ~n18107 ;
  assign n18111 = ~n18109 & n18110 ;
  assign n18112 = ~n18078 & n18106 ;
  assign n18113 = n18088 & n18112 ;
  assign n18136 = ~n18111 & ~n18113 ;
  assign n18137 = ~n18120 & n18136 ;
  assign n18138 = ~n18105 & n18137 ;
  assign n18139 = ~n18135 & n18138 ;
  assign n18140 = \u2_L5_reg[11]/NET0131  & ~n18139 ;
  assign n18141 = ~\u2_L5_reg[11]/NET0131  & n18139 ;
  assign n18142 = ~n18140 & ~n18141 ;
  assign n18156 = decrypt_pad & ~\u2_uk_K_r5_reg[54]/NET0131  ;
  assign n18157 = ~decrypt_pad & ~\u2_uk_K_r5_reg[19]/NET0131  ;
  assign n18158 = ~n18156 & ~n18157 ;
  assign n18159 = \u2_R5_reg[14]/NET0131  & ~n18158 ;
  assign n18160 = ~\u2_R5_reg[14]/NET0131  & n18158 ;
  assign n18161 = ~n18159 & ~n18160 ;
  assign n18149 = decrypt_pad & ~\u2_uk_K_r5_reg[34]/NET0131  ;
  assign n18150 = ~decrypt_pad & ~\u2_uk_K_r5_reg[24]/NET0131  ;
  assign n18151 = ~n18149 & ~n18150 ;
  assign n18152 = \u2_R5_reg[12]/NET0131  & ~n18151 ;
  assign n18153 = ~\u2_R5_reg[12]/NET0131  & n18151 ;
  assign n18154 = ~n18152 & ~n18153 ;
  assign n18163 = decrypt_pad & ~\u2_uk_K_r5_reg[18]/NET0131  ;
  assign n18164 = ~decrypt_pad & ~\u2_uk_K_r5_reg[40]/NET0131  ;
  assign n18165 = ~n18163 & ~n18164 ;
  assign n18166 = \u2_R5_reg[17]/NET0131  & ~n18165 ;
  assign n18167 = ~\u2_R5_reg[17]/NET0131  & n18165 ;
  assign n18168 = ~n18166 & ~n18167 ;
  assign n18177 = n18154 & ~n18168 ;
  assign n18178 = n18161 & n18177 ;
  assign n18170 = decrypt_pad & ~\u2_uk_K_r5_reg[5]/NET0131  ;
  assign n18171 = ~decrypt_pad & ~\u2_uk_K_r5_reg[27]/NET0131  ;
  assign n18172 = ~n18170 & ~n18171 ;
  assign n18173 = \u2_R5_reg[15]/NET0131  & ~n18172 ;
  assign n18174 = ~\u2_R5_reg[15]/NET0131  & n18172 ;
  assign n18175 = ~n18173 & ~n18174 ;
  assign n18143 = decrypt_pad & ~\u2_uk_K_r5_reg[53]/NET0131  ;
  assign n18144 = ~decrypt_pad & ~\u2_uk_K_r5_reg[18]/NET0131  ;
  assign n18145 = ~n18143 & ~n18144 ;
  assign n18146 = \u2_R5_reg[13]/NET0131  & ~n18145 ;
  assign n18147 = ~\u2_R5_reg[13]/NET0131  & n18145 ;
  assign n18148 = ~n18146 & ~n18147 ;
  assign n18176 = ~n18148 & n18168 ;
  assign n18179 = ~n18175 & ~n18176 ;
  assign n18180 = ~n18178 & n18179 ;
  assign n18183 = ~n18148 & ~n18168 ;
  assign n18184 = ~n18154 & n18183 ;
  assign n18181 = n18148 & n18154 ;
  assign n18182 = n18168 & n18181 ;
  assign n18185 = n18175 & ~n18182 ;
  assign n18186 = ~n18184 & n18185 ;
  assign n18187 = ~n18180 & ~n18186 ;
  assign n18155 = ~n18148 & n18154 ;
  assign n18162 = n18155 & ~n18161 ;
  assign n18169 = n18162 & n18168 ;
  assign n18188 = decrypt_pad & ~\u2_uk_K_r5_reg[13]/P0001  ;
  assign n18189 = ~decrypt_pad & ~\u2_uk_K_r5_reg[3]/NET0131  ;
  assign n18190 = ~n18188 & ~n18189 ;
  assign n18191 = \u2_R5_reg[16]/NET0131  & ~n18190 ;
  assign n18192 = ~\u2_R5_reg[16]/NET0131  & n18190 ;
  assign n18193 = ~n18191 & ~n18192 ;
  assign n18201 = ~n18169 & ~n18193 ;
  assign n18200 = ~n18161 & n18184 ;
  assign n18194 = n18161 & n18175 ;
  assign n18195 = n18148 & n18194 ;
  assign n18196 = ~n18154 & n18195 ;
  assign n18197 = n18148 & ~n18154 ;
  assign n18198 = ~n18168 & n18197 ;
  assign n18199 = n18161 & n18198 ;
  assign n18202 = ~n18196 & ~n18199 ;
  assign n18203 = ~n18200 & n18202 ;
  assign n18204 = n18201 & n18203 ;
  assign n18205 = ~n18187 & n18204 ;
  assign n18213 = ~n18155 & ~n18197 ;
  assign n18214 = ~n18161 & ~n18213 ;
  assign n18215 = n18161 & n18184 ;
  assign n18216 = ~n18214 & ~n18215 ;
  assign n18217 = ~n18175 & ~n18216 ;
  assign n18206 = n18161 & n18182 ;
  assign n18207 = ~n18154 & n18168 ;
  assign n18208 = n18148 & n18207 ;
  assign n18209 = ~n18161 & n18208 ;
  assign n18210 = ~n18206 & ~n18209 ;
  assign n18218 = ~n18148 & n18175 ;
  assign n18219 = n18207 & n18218 ;
  assign n18211 = ~n18168 & n18175 ;
  assign n18212 = n18181 & n18211 ;
  assign n18220 = n18193 & ~n18212 ;
  assign n18221 = ~n18219 & n18220 ;
  assign n18222 = n18210 & n18221 ;
  assign n18223 = ~n18217 & n18222 ;
  assign n18224 = ~n18205 & ~n18223 ;
  assign n18225 = ~n18175 & n18209 ;
  assign n18226 = ~n18148 & n18161 ;
  assign n18227 = n18148 & ~n18161 ;
  assign n18228 = ~n18226 & ~n18227 ;
  assign n18229 = n18177 & ~n18228 ;
  assign n18230 = ~n18200 & ~n18229 ;
  assign n18231 = n18175 & ~n18230 ;
  assign n18232 = ~n18225 & ~n18231 ;
  assign n18233 = ~n18224 & n18232 ;
  assign n18234 = ~\u2_L5_reg[20]/NET0131  & ~n18233 ;
  assign n18235 = \u2_L5_reg[20]/NET0131  & n18233 ;
  assign n18236 = ~n18234 & ~n18235 ;
  assign n18271 = decrypt_pad & ~\u2_uk_K_r5_reg[9]/P0001  ;
  assign n18272 = ~decrypt_pad & ~\u2_uk_K_r5_reg[29]/NET0131  ;
  assign n18273 = ~n18271 & ~n18272 ;
  assign n18274 = \u2_R5_reg[32]/NET0131  & ~n18273 ;
  assign n18275 = ~\u2_R5_reg[32]/NET0131  & n18273 ;
  assign n18276 = ~n18274 & ~n18275 ;
  assign n18243 = decrypt_pad & ~\u2_uk_K_r5_reg[42]/NET0131  ;
  assign n18244 = ~decrypt_pad & ~\u2_uk_K_r5_reg[7]/NET0131  ;
  assign n18245 = ~n18243 & ~n18244 ;
  assign n18246 = \u2_R5_reg[28]/NET0131  & ~n18245 ;
  assign n18247 = ~\u2_R5_reg[28]/NET0131  & n18245 ;
  assign n18248 = ~n18246 & ~n18247 ;
  assign n18249 = decrypt_pad & ~\u2_uk_K_r5_reg[15]/NET0131  ;
  assign n18250 = ~decrypt_pad & ~\u2_uk_K_r5_reg[35]/NET0131  ;
  assign n18251 = ~n18249 & ~n18250 ;
  assign n18252 = \u2_R5_reg[30]/NET0131  & ~n18251 ;
  assign n18253 = ~\u2_R5_reg[30]/NET0131  & n18251 ;
  assign n18254 = ~n18252 & ~n18253 ;
  assign n18255 = n18248 & ~n18254 ;
  assign n18256 = decrypt_pad & ~\u2_uk_K_r5_reg[14]/NET0131  ;
  assign n18257 = ~decrypt_pad & ~\u2_uk_K_r5_reg[38]/NET0131  ;
  assign n18258 = ~n18256 & ~n18257 ;
  assign n18259 = \u2_R5_reg[29]/NET0131  & ~n18258 ;
  assign n18260 = ~\u2_R5_reg[29]/NET0131  & n18258 ;
  assign n18261 = ~n18259 & ~n18260 ;
  assign n18262 = decrypt_pad & ~\u2_uk_K_r5_reg[30]/NET0131  ;
  assign n18263 = ~decrypt_pad & ~\u2_uk_K_r5_reg[50]/NET0131  ;
  assign n18264 = ~n18262 & ~n18263 ;
  assign n18265 = \u2_R5_reg[1]/NET0131  & ~n18264 ;
  assign n18266 = ~\u2_R5_reg[1]/NET0131  & n18264 ;
  assign n18267 = ~n18265 & ~n18266 ;
  assign n18268 = n18261 & ~n18267 ;
  assign n18303 = ~n18255 & ~n18268 ;
  assign n18237 = decrypt_pad & ~\u2_uk_K_r5_reg[31]/NET0131  ;
  assign n18238 = ~decrypt_pad & ~\u2_uk_K_r5_reg[23]/NET0131  ;
  assign n18239 = ~n18237 & ~n18238 ;
  assign n18240 = \u2_R5_reg[31]/P0001  & ~n18239 ;
  assign n18241 = ~\u2_R5_reg[31]/P0001  & n18239 ;
  assign n18242 = ~n18240 & ~n18241 ;
  assign n18269 = n18255 & n18268 ;
  assign n18304 = n18242 & ~n18269 ;
  assign n18305 = ~n18303 & n18304 ;
  assign n18284 = n18248 & ~n18261 ;
  assign n18296 = n18254 & n18284 ;
  assign n18297 = ~n18254 & ~n18261 ;
  assign n18298 = ~n18248 & n18297 ;
  assign n18299 = ~n18296 & ~n18298 ;
  assign n18300 = ~n18242 & ~n18299 ;
  assign n18288 = ~n18248 & n18254 ;
  assign n18301 = n18261 & n18288 ;
  assign n18302 = n18267 & n18301 ;
  assign n18306 = ~n18300 & ~n18302 ;
  assign n18307 = ~n18305 & n18306 ;
  assign n18308 = n18276 & ~n18307 ;
  assign n18282 = ~n18261 & n18267 ;
  assign n18289 = ~n18267 & ~n18288 ;
  assign n18290 = ~n18282 & ~n18289 ;
  assign n18291 = ~n18255 & ~n18290 ;
  assign n18292 = ~n18242 & ~n18291 ;
  assign n18277 = n18248 & n18261 ;
  assign n18278 = n18254 & ~n18267 ;
  assign n18279 = ~n18254 & n18267 ;
  assign n18280 = ~n18278 & ~n18279 ;
  assign n18281 = n18277 & n18280 ;
  assign n18283 = ~n18248 & n18282 ;
  assign n18285 = n18278 & n18284 ;
  assign n18286 = ~n18283 & ~n18285 ;
  assign n18287 = n18242 & ~n18286 ;
  assign n18293 = ~n18281 & ~n18287 ;
  assign n18294 = ~n18292 & n18293 ;
  assign n18295 = ~n18276 & ~n18294 ;
  assign n18270 = ~n18242 & n18269 ;
  assign n18311 = ~n18254 & n18261 ;
  assign n18312 = n18248 & ~n18267 ;
  assign n18313 = ~n18311 & ~n18312 ;
  assign n18314 = ~n18303 & n18313 ;
  assign n18309 = ~n18267 & n18298 ;
  assign n18310 = n18282 & n18288 ;
  assign n18315 = ~n18309 & ~n18310 ;
  assign n18316 = ~n18314 & n18315 ;
  assign n18317 = n18242 & ~n18316 ;
  assign n18318 = ~n18270 & ~n18317 ;
  assign n18319 = ~n18295 & n18318 ;
  assign n18320 = ~n18308 & n18319 ;
  assign n18321 = \u2_L5_reg[5]/NET0131  & ~n18320 ;
  assign n18322 = ~\u2_L5_reg[5]/NET0131  & n18320 ;
  assign n18323 = ~n18321 & ~n18322 ;
  assign n18329 = ~n18169 & ~n18198 ;
  assign n18330 = n18175 & ~n18329 ;
  assign n18324 = n18207 & n18226 ;
  assign n18325 = ~n18206 & ~n18324 ;
  assign n18326 = n18177 & ~n18227 ;
  assign n18327 = ~n18209 & ~n18326 ;
  assign n18328 = ~n18175 & ~n18327 ;
  assign n18331 = n18325 & ~n18328 ;
  assign n18332 = ~n18330 & n18331 ;
  assign n18333 = n18193 & ~n18332 ;
  assign n18337 = ~n18161 & n18168 ;
  assign n18338 = n18175 & n18337 ;
  assign n18339 = ~n18218 & ~n18337 ;
  assign n18340 = ~n18338 & ~n18339 ;
  assign n18341 = ~n18227 & ~n18340 ;
  assign n18342 = n18154 & ~n18341 ;
  assign n18343 = n18175 & n18207 ;
  assign n18344 = ~n18184 & ~n18343 ;
  assign n18345 = ~n18194 & ~n18344 ;
  assign n18346 = ~n18199 & ~n18345 ;
  assign n18347 = ~n18342 & n18346 ;
  assign n18348 = ~n18193 & ~n18347 ;
  assign n18334 = ~n18200 & n18325 ;
  assign n18335 = ~n18175 & ~n18334 ;
  assign n18336 = ~n18161 & n18212 ;
  assign n18349 = ~n18196 & ~n18336 ;
  assign n18350 = ~n18335 & n18349 ;
  assign n18351 = ~n18348 & n18350 ;
  assign n18352 = ~n18333 & n18351 ;
  assign n18353 = ~\u2_L5_reg[10]/NET0131  & ~n18352 ;
  assign n18354 = \u2_L5_reg[10]/NET0131  & n18352 ;
  assign n18355 = ~n18353 & ~n18354 ;
  assign n18358 = n17880 & n17893 ;
  assign n18357 = ~n17907 & n17911 ;
  assign n18363 = ~n17914 & ~n18357 ;
  assign n18364 = ~n18358 & n18363 ;
  assign n18359 = ~n17871 & ~n17925 ;
  assign n18360 = n17907 & ~n18359 ;
  assign n18356 = n17910 & n17937 ;
  assign n18361 = n17887 & ~n17896 ;
  assign n18362 = ~n18356 & n18361 ;
  assign n18365 = ~n18360 & n18362 ;
  assign n18366 = n18364 & n18365 ;
  assign n18372 = n17864 & ~n17907 ;
  assign n18373 = ~n17909 & ~n17937 ;
  assign n18374 = ~n17870 & n18373 ;
  assign n18375 = ~n18372 & ~n18374 ;
  assign n18376 = n17877 & ~n18375 ;
  assign n18367 = n17879 & n17924 ;
  assign n18379 = ~n17887 & ~n18367 ;
  assign n18380 = ~n17942 & n18379 ;
  assign n18368 = ~n17864 & ~n17879 ;
  assign n18369 = ~n17870 & ~n17907 ;
  assign n18370 = n17893 & ~n18369 ;
  assign n18371 = n18368 & n18370 ;
  assign n18377 = ~n17897 & ~n17916 ;
  assign n18378 = ~n17907 & ~n18377 ;
  assign n18381 = ~n18371 & ~n18378 ;
  assign n18382 = n18380 & n18381 ;
  assign n18383 = ~n18376 & n18382 ;
  assign n18384 = ~n18366 & ~n18383 ;
  assign n18385 = \u2_L5_reg[12]/NET0131  & n18384 ;
  assign n18386 = ~\u2_L5_reg[12]/NET0131  & ~n18384 ;
  assign n18387 = ~n18385 & ~n18386 ;
  assign n18388 = decrypt_pad & ~\u2_uk_K_r5_reg[38]/NET0131  ;
  assign n18389 = ~decrypt_pad & ~\u2_uk_K_r5_reg[30]/NET0131  ;
  assign n18390 = ~n18388 & ~n18389 ;
  assign n18391 = \u2_R5_reg[19]/NET0131  & ~n18390 ;
  assign n18392 = ~\u2_R5_reg[19]/NET0131  & n18390 ;
  assign n18393 = ~n18391 & ~n18392 ;
  assign n18394 = decrypt_pad & ~\u2_uk_K_r5_reg[23]/NET0131  ;
  assign n18395 = ~decrypt_pad & ~\u2_uk_K_r5_reg[43]/NET0131  ;
  assign n18396 = ~n18394 & ~n18395 ;
  assign n18397 = \u2_R5_reg[18]/NET0131  & ~n18396 ;
  assign n18398 = ~\u2_R5_reg[18]/NET0131  & n18396 ;
  assign n18399 = ~n18397 & ~n18398 ;
  assign n18400 = decrypt_pad & ~\u2_uk_K_r5_reg[29]/NET0131  ;
  assign n18401 = ~decrypt_pad & ~\u2_uk_K_r5_reg[49]/NET0131  ;
  assign n18402 = ~n18400 & ~n18401 ;
  assign n18403 = \u2_R5_reg[17]/NET0131  & ~n18402 ;
  assign n18404 = ~\u2_R5_reg[17]/NET0131  & n18402 ;
  assign n18405 = ~n18403 & ~n18404 ;
  assign n18407 = decrypt_pad & ~\u2_uk_K_r5_reg[7]/NET0131  ;
  assign n18408 = ~decrypt_pad & ~\u2_uk_K_r5_reg[31]/NET0131  ;
  assign n18409 = ~n18407 & ~n18408 ;
  assign n18410 = \u2_R5_reg[16]/NET0131  & ~n18409 ;
  assign n18411 = ~\u2_R5_reg[16]/NET0131  & n18409 ;
  assign n18412 = ~n18410 & ~n18411 ;
  assign n18414 = decrypt_pad & ~\u2_uk_K_r5_reg[50]/NET0131  ;
  assign n18415 = ~decrypt_pad & ~\u2_uk_K_r5_reg[15]/NET0131  ;
  assign n18416 = ~n18414 & ~n18415 ;
  assign n18417 = \u2_R5_reg[21]/NET0131  & ~n18416 ;
  assign n18418 = ~\u2_R5_reg[21]/NET0131  & n18416 ;
  assign n18419 = ~n18417 & ~n18418 ;
  assign n18420 = n18412 & ~n18419 ;
  assign n18431 = ~n18405 & n18420 ;
  assign n18432 = ~n18399 & n18431 ;
  assign n18406 = ~n18399 & n18405 ;
  assign n18433 = n18412 & n18419 ;
  assign n18434 = n18406 & n18433 ;
  assign n18423 = n18405 & ~n18419 ;
  assign n18428 = n18399 & n18423 ;
  assign n18429 = ~n18412 & n18419 ;
  assign n18430 = ~n18405 & n18429 ;
  assign n18435 = ~n18428 & ~n18430 ;
  assign n18436 = ~n18434 & n18435 ;
  assign n18437 = ~n18432 & n18436 ;
  assign n18438 = ~n18393 & ~n18437 ;
  assign n18413 = n18406 & ~n18412 ;
  assign n18421 = n18399 & n18412 ;
  assign n18422 = n18419 & ~n18421 ;
  assign n18424 = ~n18420 & ~n18423 ;
  assign n18425 = ~n18422 & n18424 ;
  assign n18426 = ~n18413 & ~n18425 ;
  assign n18427 = n18393 & ~n18426 ;
  assign n18439 = ~n18399 & n18419 ;
  assign n18440 = ~n18420 & ~n18439 ;
  assign n18441 = ~n18405 & ~n18412 ;
  assign n18442 = n18399 & n18405 ;
  assign n18443 = ~n18441 & ~n18442 ;
  assign n18444 = n18440 & n18443 ;
  assign n18445 = ~n18427 & ~n18444 ;
  assign n18446 = ~n18438 & n18445 ;
  assign n18447 = decrypt_pad & ~\u2_uk_K_r5_reg[49]/NET0131  ;
  assign n18448 = ~decrypt_pad & ~\u2_uk_K_r5_reg[14]/NET0131  ;
  assign n18449 = ~n18447 & ~n18448 ;
  assign n18450 = \u2_R5_reg[20]/NET0131  & ~n18449 ;
  assign n18451 = ~\u2_R5_reg[20]/NET0131  & n18449 ;
  assign n18452 = ~n18450 & ~n18451 ;
  assign n18453 = ~n18446 & ~n18452 ;
  assign n18457 = ~n18413 & n18422 ;
  assign n18458 = n18412 & n18423 ;
  assign n18459 = ~n18457 & ~n18458 ;
  assign n18460 = n18393 & ~n18459 ;
  assign n18461 = n18405 & n18429 ;
  assign n18462 = ~n18419 & n18441 ;
  assign n18463 = ~n18461 & ~n18462 ;
  assign n18464 = ~n18393 & ~n18399 ;
  assign n18465 = ~n18463 & n18464 ;
  assign n18454 = n18399 & ~n18405 ;
  assign n18455 = ~n18406 & ~n18454 ;
  assign n18456 = n18420 & ~n18455 ;
  assign n18466 = n18393 & n18399 ;
  assign n18467 = n18433 & ~n18466 ;
  assign n18468 = n18455 & n18467 ;
  assign n18469 = ~n18456 & ~n18468 ;
  assign n18470 = ~n18465 & n18469 ;
  assign n18471 = ~n18460 & n18470 ;
  assign n18472 = n18452 & ~n18471 ;
  assign n18473 = n18399 & n18462 ;
  assign n18474 = ~n18399 & n18458 ;
  assign n18475 = ~n18473 & ~n18474 ;
  assign n18476 = n18393 & ~n18475 ;
  assign n18477 = n18399 & n18430 ;
  assign n18478 = ~n18412 & n18428 ;
  assign n18479 = ~n18477 & ~n18478 ;
  assign n18480 = ~n18393 & ~n18479 ;
  assign n18481 = ~n18476 & ~n18480 ;
  assign n18482 = ~n18472 & n18481 ;
  assign n18483 = ~n18453 & n18482 ;
  assign n18484 = ~\u2_L5_reg[14]/NET0131  & ~n18483 ;
  assign n18485 = \u2_L5_reg[14]/NET0131  & n18483 ;
  assign n18486 = ~n18484 & ~n18485 ;
  assign n18487 = ~n18267 & n18311 ;
  assign n18488 = ~n18277 & ~n18487 ;
  assign n18489 = ~n18283 & n18488 ;
  assign n18490 = n18242 & ~n18489 ;
  assign n18491 = n18297 & n18312 ;
  assign n18492 = ~n18490 & ~n18491 ;
  assign n18493 = ~n18276 & ~n18492 ;
  assign n18495 = n18267 & n18296 ;
  assign n18494 = ~n18254 & n18277 ;
  assign n18496 = ~n18242 & n18254 ;
  assign n18497 = n18282 & n18496 ;
  assign n18502 = ~n18494 & ~n18497 ;
  assign n18498 = ~n18248 & ~n18267 ;
  assign n18499 = n18242 & ~n18261 ;
  assign n18500 = n18498 & n18499 ;
  assign n18501 = n18268 & n18288 ;
  assign n18503 = ~n18500 & ~n18501 ;
  assign n18504 = n18502 & n18503 ;
  assign n18505 = ~n18495 & n18504 ;
  assign n18506 = n18276 & ~n18505 ;
  assign n18507 = ~n18248 & n18261 ;
  assign n18508 = ~n18280 & n18507 ;
  assign n18509 = ~n18254 & n18276 ;
  assign n18510 = n18284 & ~n18509 ;
  assign n18511 = ~n18242 & ~n18510 ;
  assign n18512 = ~n18309 & n18511 ;
  assign n18513 = ~n18508 & n18512 ;
  assign n18514 = ~n18254 & n18283 ;
  assign n18515 = n18242 & ~n18302 ;
  assign n18516 = ~n18514 & n18515 ;
  assign n18517 = ~n18513 & ~n18516 ;
  assign n18518 = ~n18506 & ~n18517 ;
  assign n18519 = ~n18493 & n18518 ;
  assign n18520 = ~\u2_L5_reg[15]/NET0131  & ~n18519 ;
  assign n18521 = \u2_L5_reg[15]/NET0131  & n18519 ;
  assign n18522 = ~n18520 & ~n18521 ;
  assign n18523 = ~n17977 & ~n17992 ;
  assign n18524 = ~n17970 & n17991 ;
  assign n18525 = ~n18523 & ~n18524 ;
  assign n18526 = ~n17964 & ~n18525 ;
  assign n18528 = n17964 & ~n17998 ;
  assign n18529 = n17977 & ~n17983 ;
  assign n18530 = n17989 & ~n18529 ;
  assign n18531 = n18528 & n18530 ;
  assign n18527 = n17996 & n18016 ;
  assign n18532 = ~n18021 & ~n18527 ;
  assign n18533 = ~n18531 & n18532 ;
  assign n18534 = ~n18526 & n18533 ;
  assign n18535 = ~n17958 & ~n18534 ;
  assign n18537 = ~n17970 & ~n17977 ;
  assign n18538 = ~n17989 & ~n18537 ;
  assign n18539 = n17990 & n18537 ;
  assign n18540 = ~n18538 & ~n18539 ;
  assign n18541 = n17964 & ~n18540 ;
  assign n18542 = ~n17964 & ~n18034 ;
  assign n18543 = ~n18538 & n18542 ;
  assign n18536 = n17996 & n18022 ;
  assign n18544 = ~n18017 & ~n18536 ;
  assign n18545 = ~n18543 & n18544 ;
  assign n18546 = ~n18541 & n18545 ;
  assign n18547 = n17958 & ~n18546 ;
  assign n18548 = ~n17970 & n18019 ;
  assign n18549 = ~n18027 & ~n18548 ;
  assign n18550 = n17964 & n17977 ;
  assign n18551 = ~n18549 & n18550 ;
  assign n18552 = ~n18547 & ~n18551 ;
  assign n18553 = ~n18535 & n18552 ;
  assign n18554 = ~\u2_L5_reg[17]/NET0131  & ~n18553 ;
  assign n18555 = \u2_L5_reg[17]/NET0131  & n18553 ;
  assign n18556 = ~n18554 & ~n18555 ;
  assign n18557 = ~n18162 & ~n18176 ;
  assign n18558 = n18193 & ~n18557 ;
  assign n18559 = n18175 & ~n18199 ;
  assign n18560 = n18325 & n18559 ;
  assign n18561 = ~n18558 & n18560 ;
  assign n18562 = n18148 & n18178 ;
  assign n18563 = ~n18175 & ~n18215 ;
  assign n18564 = ~n18562 & n18563 ;
  assign n18565 = ~n18561 & ~n18564 ;
  assign n18571 = ~n18161 & ~n18168 ;
  assign n18572 = ~n18176 & ~n18571 ;
  assign n18573 = n18154 & ~n18218 ;
  assign n18574 = ~n18572 & n18573 ;
  assign n18566 = n18154 & ~n18161 ;
  assign n18567 = ~n18154 & n18161 ;
  assign n18568 = ~n18566 & ~n18567 ;
  assign n18569 = ~n18181 & n18211 ;
  assign n18570 = n18568 & n18569 ;
  assign n18575 = ~n18193 & ~n18570 ;
  assign n18576 = ~n18574 & n18575 ;
  assign n18577 = n18210 & n18576 ;
  assign n18579 = ~n18177 & n18227 ;
  assign n18580 = ~n18208 & ~n18579 ;
  assign n18581 = ~n18175 & ~n18580 ;
  assign n18578 = ~n18154 & n18226 ;
  assign n18582 = n18193 & ~n18578 ;
  assign n18583 = ~n18562 & n18582 ;
  assign n18584 = ~n18581 & n18583 ;
  assign n18585 = ~n18577 & ~n18584 ;
  assign n18586 = ~n18565 & ~n18585 ;
  assign n18587 = ~\u2_L5_reg[1]/NET0131  & ~n18586 ;
  assign n18588 = \u2_L5_reg[1]/NET0131  & n18586 ;
  assign n18589 = ~n18587 & ~n18588 ;
  assign n18596 = n18261 & ~n18498 ;
  assign n18597 = ~n18255 & n18596 ;
  assign n18598 = ~n18254 & n18282 ;
  assign n18599 = ~n18597 & ~n18598 ;
  assign n18600 = n18242 & ~n18599 ;
  assign n18590 = ~n18254 & n18312 ;
  assign n18591 = ~n18495 & ~n18590 ;
  assign n18592 = ~n18242 & ~n18591 ;
  assign n18593 = ~n18267 & ~n18507 ;
  assign n18594 = n18254 & ~n18284 ;
  assign n18595 = n18593 & n18594 ;
  assign n18601 = n18276 & ~n18514 ;
  assign n18602 = ~n18595 & n18601 ;
  assign n18603 = ~n18592 & n18602 ;
  assign n18604 = ~n18600 & n18603 ;
  assign n18611 = n18248 & n18267 ;
  assign n18612 = ~n18254 & ~n18499 ;
  assign n18613 = n18611 & n18612 ;
  assign n18616 = ~n18276 & ~n18301 ;
  assign n18605 = ~n18242 & n18267 ;
  assign n18606 = n18288 & n18605 ;
  assign n18614 = ~n18242 & ~n18248 ;
  assign n18615 = n18268 & n18614 ;
  assign n18617 = ~n18606 & ~n18615 ;
  assign n18618 = n18616 & n18617 ;
  assign n18619 = ~n18613 & n18618 ;
  assign n18607 = n18261 & n18312 ;
  assign n18608 = ~n18296 & ~n18607 ;
  assign n18609 = n18242 & ~n18608 ;
  assign n18610 = ~n18267 & ~n18299 ;
  assign n18620 = ~n18609 & ~n18610 ;
  assign n18621 = n18619 & n18620 ;
  assign n18622 = ~n18604 & ~n18621 ;
  assign n18623 = n18494 & n18605 ;
  assign n18624 = n18242 & n18298 ;
  assign n18625 = ~n18623 & ~n18624 ;
  assign n18626 = ~n18622 & n18625 ;
  assign n18627 = ~\u2_L5_reg[21]/NET0131  & ~n18626 ;
  assign n18628 = \u2_L5_reg[21]/NET0131  & n18626 ;
  assign n18629 = ~n18627 & ~n18628 ;
  assign n18632 = ~n18406 & ~n18419 ;
  assign n18633 = ~n18421 & n18632 ;
  assign n18631 = n18405 & n18433 ;
  assign n18634 = ~n18441 & ~n18631 ;
  assign n18635 = ~n18633 & n18634 ;
  assign n18636 = n18393 & ~n18635 ;
  assign n18637 = ~n18405 & n18433 ;
  assign n18638 = ~n18413 & ~n18637 ;
  assign n18639 = ~n18393 & ~n18638 ;
  assign n18630 = n18405 & n18439 ;
  assign n18640 = n18421 & n18423 ;
  assign n18641 = ~n18630 & ~n18640 ;
  assign n18642 = ~n18639 & n18641 ;
  assign n18643 = ~n18636 & n18642 ;
  assign n18644 = n18452 & ~n18643 ;
  assign n18656 = ~n18473 & ~n18640 ;
  assign n18657 = ~n18399 & n18430 ;
  assign n18658 = n18656 & ~n18657 ;
  assign n18659 = n18393 & ~n18658 ;
  assign n18650 = n18393 & ~n18423 ;
  assign n18649 = ~n18393 & ~n18441 ;
  assign n18651 = ~n18399 & ~n18649 ;
  assign n18652 = ~n18650 & n18651 ;
  assign n18645 = ~n18393 & n18431 ;
  assign n18646 = n18393 & ~n18419 ;
  assign n18647 = ~n18412 & n18442 ;
  assign n18648 = ~n18646 & n18647 ;
  assign n18653 = ~n18645 & ~n18648 ;
  assign n18654 = ~n18652 & n18653 ;
  assign n18655 = ~n18452 & ~n18654 ;
  assign n18660 = ~n18393 & n18412 ;
  assign n18661 = n18454 & n18660 ;
  assign n18662 = ~n18434 & ~n18661 ;
  assign n18663 = ~n18655 & n18662 ;
  assign n18664 = ~n18659 & n18663 ;
  assign n18665 = ~n18644 & n18664 ;
  assign n18666 = ~\u2_L5_reg[25]/NET0131  & ~n18665 ;
  assign n18667 = \u2_L5_reg[25]/NET0131  & n18665 ;
  assign n18668 = ~n18666 & ~n18667 ;
  assign n18677 = ~n18208 & ~n18343 ;
  assign n18678 = n18161 & ~n18677 ;
  assign n18679 = n18197 & n18571 ;
  assign n18683 = ~n18562 & ~n18679 ;
  assign n18676 = n18175 & n18184 ;
  assign n18680 = n18168 & ~n18175 ;
  assign n18681 = ~n18197 & n18680 ;
  assign n18682 = n18568 & n18681 ;
  assign n18684 = ~n18676 & ~n18682 ;
  assign n18685 = n18683 & n18684 ;
  assign n18686 = ~n18678 & n18685 ;
  assign n18687 = n18193 & ~n18686 ;
  assign n18669 = ~n18183 & ~n18578 ;
  assign n18670 = ~n18193 & ~n18669 ;
  assign n18671 = ~n18168 & ~n18213 ;
  assign n18672 = ~n18182 & ~n18671 ;
  assign n18673 = ~n18161 & ~n18672 ;
  assign n18674 = ~n18670 & ~n18673 ;
  assign n18675 = ~n18175 & ~n18674 ;
  assign n18688 = ~n18213 & n18338 ;
  assign n18689 = n18195 & ~n18207 ;
  assign n18690 = ~n18162 & ~n18212 ;
  assign n18691 = ~n18209 & n18690 ;
  assign n18692 = ~n18689 & n18691 ;
  assign n18693 = ~n18193 & ~n18692 ;
  assign n18694 = ~n18688 & ~n18693 ;
  assign n18695 = ~n18675 & n18694 ;
  assign n18696 = ~n18687 & n18695 ;
  assign n18697 = ~\u2_L5_reg[26]/NET0131  & ~n18696 ;
  assign n18698 = \u2_L5_reg[26]/NET0131  & n18696 ;
  assign n18699 = ~n18697 & ~n18698 ;
  assign n18700 = decrypt_pad & ~\u2_uk_K_r5_reg[12]/NET0131  ;
  assign n18701 = ~decrypt_pad & ~\u2_uk_K_r5_reg[34]/NET0131  ;
  assign n18702 = ~n18700 & ~n18701 ;
  assign n18703 = \u2_R5_reg[8]/NET0131  & ~n18702 ;
  assign n18704 = ~\u2_R5_reg[8]/NET0131  & n18702 ;
  assign n18705 = ~n18703 & ~n18704 ;
  assign n18706 = decrypt_pad & ~\u2_uk_K_r5_reg[25]/NET0131  ;
  assign n18707 = ~decrypt_pad & ~\u2_uk_K_r5_reg[47]/NET0131  ;
  assign n18708 = ~n18706 & ~n18707 ;
  assign n18709 = \u2_R5_reg[4]/NET0131  & ~n18708 ;
  assign n18710 = ~\u2_R5_reg[4]/NET0131  & n18708 ;
  assign n18711 = ~n18709 & ~n18710 ;
  assign n18712 = decrypt_pad & ~\u2_uk_K_r5_reg[17]/NET0131  ;
  assign n18713 = ~decrypt_pad & ~\u2_uk_K_r5_reg[39]/NET0131  ;
  assign n18714 = ~n18712 & ~n18713 ;
  assign n18715 = \u2_R5_reg[9]/NET0131  & ~n18714 ;
  assign n18716 = ~\u2_R5_reg[9]/NET0131  & n18714 ;
  assign n18717 = ~n18715 & ~n18716 ;
  assign n18718 = n18711 & n18717 ;
  assign n18719 = decrypt_pad & ~\u2_uk_K_r5_reg[4]/NET0131  ;
  assign n18720 = ~decrypt_pad & ~\u2_uk_K_r5_reg[26]/NET0131  ;
  assign n18721 = ~n18719 & ~n18720 ;
  assign n18722 = \u2_R5_reg[5]/NET0131  & ~n18721 ;
  assign n18723 = ~\u2_R5_reg[5]/NET0131  & n18721 ;
  assign n18724 = ~n18722 & ~n18723 ;
  assign n18725 = n18717 & ~n18724 ;
  assign n18726 = ~n18717 & n18724 ;
  assign n18727 = ~n18725 & ~n18726 ;
  assign n18728 = ~n18718 & ~n18727 ;
  assign n18729 = decrypt_pad & ~\u2_uk_K_r5_reg[27]/NET0131  ;
  assign n18730 = ~decrypt_pad & ~\u2_uk_K_r5_reg[17]/NET0131  ;
  assign n18731 = ~n18729 & ~n18730 ;
  assign n18732 = \u2_R5_reg[6]/NET0131  & ~n18731 ;
  assign n18733 = ~\u2_R5_reg[6]/NET0131  & n18731 ;
  assign n18734 = ~n18732 & ~n18733 ;
  assign n18735 = n18728 & ~n18734 ;
  assign n18736 = decrypt_pad & ~\u2_uk_K_r5_reg[46]/NET0131  ;
  assign n18737 = ~decrypt_pad & ~\u2_uk_K_r5_reg[11]/NET0131  ;
  assign n18738 = ~n18736 & ~n18737 ;
  assign n18739 = \u2_R5_reg[7]/NET0131  & ~n18738 ;
  assign n18740 = ~\u2_R5_reg[7]/NET0131  & n18738 ;
  assign n18741 = ~n18739 & ~n18740 ;
  assign n18742 = n18711 & n18734 ;
  assign n18743 = n18725 & n18742 ;
  assign n18744 = n18741 & n18743 ;
  assign n18761 = ~n18735 & ~n18744 ;
  assign n18745 = n18724 & ~n18734 ;
  assign n18746 = n18717 & ~n18734 ;
  assign n18747 = ~n18741 & n18746 ;
  assign n18748 = ~n18711 & n18717 ;
  assign n18749 = n18724 & n18748 ;
  assign n18750 = ~n18747 & ~n18749 ;
  assign n18751 = ~n18745 & ~n18750 ;
  assign n18753 = ~n18711 & ~n18717 ;
  assign n18754 = ~n18718 & ~n18753 ;
  assign n18755 = ~n18724 & ~n18754 ;
  assign n18752 = n18711 & ~n18734 ;
  assign n18756 = ~n18724 & ~n18741 ;
  assign n18757 = n18711 & ~n18741 ;
  assign n18758 = ~n18756 & ~n18757 ;
  assign n18759 = ~n18752 & ~n18758 ;
  assign n18760 = ~n18755 & n18759 ;
  assign n18762 = ~n18751 & ~n18760 ;
  assign n18763 = n18761 & n18762 ;
  assign n18764 = ~n18705 & ~n18763 ;
  assign n18778 = ~n18743 & ~n18753 ;
  assign n18779 = n18705 & ~n18778 ;
  assign n18780 = ~n18724 & n18734 ;
  assign n18781 = n18748 & ~n18780 ;
  assign n18782 = ~n18779 & ~n18781 ;
  assign n18783 = ~n18741 & ~n18745 ;
  assign n18784 = ~n18782 & n18783 ;
  assign n18765 = ~n18717 & ~n18724 ;
  assign n18766 = ~n18711 & n18734 ;
  assign n18767 = n18765 & n18766 ;
  assign n18768 = n18711 & n18745 ;
  assign n18769 = ~n18767 & ~n18768 ;
  assign n18770 = n18741 & ~n18769 ;
  assign n18774 = n18717 & n18768 ;
  assign n18771 = n18752 & n18765 ;
  assign n18772 = n18724 & n18741 ;
  assign n18773 = ~n18766 & n18772 ;
  assign n18775 = ~n18771 & ~n18773 ;
  assign n18776 = ~n18774 & n18775 ;
  assign n18777 = n18705 & ~n18776 ;
  assign n18785 = ~n18770 & ~n18777 ;
  assign n18786 = ~n18784 & n18785 ;
  assign n18787 = ~n18764 & n18786 ;
  assign n18788 = \u2_L5_reg[2]/NET0131  & n18787 ;
  assign n18789 = ~\u2_L5_reg[2]/NET0131  & ~n18787 ;
  assign n18790 = ~n18788 & ~n18789 ;
  assign n18807 = n18066 & ~n18078 ;
  assign n18808 = ~n18084 & ~n18807 ;
  assign n18809 = ~n18079 & ~n18082 ;
  assign n18810 = ~n18065 & ~n18809 ;
  assign n18811 = n18808 & ~n18810 ;
  assign n18812 = n18053 & ~n18811 ;
  assign n18791 = n18072 & n18114 ;
  assign n18798 = ~n18072 & ~n18089 ;
  assign n18813 = ~n18791 & ~n18798 ;
  assign n18814 = ~n18053 & ~n18813 ;
  assign n18815 = n18072 & n18117 ;
  assign n18816 = ~n18814 & ~n18815 ;
  assign n18817 = ~n18812 & n18816 ;
  assign n18818 = ~n18104 & ~n18817 ;
  assign n18792 = n18078 & n18129 ;
  assign n18793 = ~n18093 & ~n18792 ;
  assign n18794 = ~n18791 & n18793 ;
  assign n18795 = n18053 & ~n18794 ;
  assign n18799 = n18053 & ~n18116 ;
  assign n18800 = ~n18127 & n18799 ;
  assign n18796 = n18072 & ~n18083 ;
  assign n18797 = ~n18106 & n18796 ;
  assign n18801 = ~n18797 & ~n18798 ;
  assign n18802 = ~n18800 & n18801 ;
  assign n18803 = ~n18795 & ~n18802 ;
  assign n18804 = n18104 & ~n18803 ;
  assign n18805 = n18053 & n18065 ;
  assign n18806 = n18108 & n18805 ;
  assign n18819 = ~n18080 & ~n18806 ;
  assign n18820 = ~n18804 & n18819 ;
  assign n18821 = ~n18818 & n18820 ;
  assign n18822 = \u2_L5_reg[29]/NET0131  & ~n18821 ;
  assign n18823 = ~\u2_L5_reg[29]/NET0131  & n18821 ;
  assign n18824 = ~n18822 & ~n18823 ;
  assign n18825 = n18711 & n18726 ;
  assign n18826 = n18734 & n18825 ;
  assign n18827 = ~n18711 & n18780 ;
  assign n18828 = ~n18826 & ~n18827 ;
  assign n18829 = ~n18741 & ~n18828 ;
  assign n18838 = ~n18755 & ~n18825 ;
  assign n18839 = n18734 & ~n18838 ;
  assign n18830 = ~n18711 & ~n18725 ;
  assign n18831 = ~n18717 & n18734 ;
  assign n18832 = ~n18718 & ~n18831 ;
  assign n18833 = ~n18724 & ~n18832 ;
  assign n18834 = ~n18741 & ~n18833 ;
  assign n18835 = ~n18830 & n18834 ;
  assign n18836 = n18830 & ~n18831 ;
  assign n18837 = n18741 & n18836 ;
  assign n18840 = ~n18705 & ~n18837 ;
  assign n18841 = ~n18835 & n18840 ;
  assign n18842 = ~n18839 & n18841 ;
  assign n18844 = ~n18725 & ~n18741 ;
  assign n18845 = n18752 & ~n18844 ;
  assign n18843 = n18717 & n18827 ;
  assign n18851 = n18705 & ~n18843 ;
  assign n18852 = ~n18845 & n18851 ;
  assign n18847 = ~n18727 & ~n18766 ;
  assign n18846 = ~n18711 & ~n18726 ;
  assign n18848 = n18741 & ~n18846 ;
  assign n18849 = ~n18847 & n18848 ;
  assign n18850 = ~n18741 & n18836 ;
  assign n18853 = ~n18849 & ~n18850 ;
  assign n18854 = n18852 & n18853 ;
  assign n18855 = ~n18842 & ~n18854 ;
  assign n18856 = ~n18829 & ~n18855 ;
  assign n18857 = ~\u2_L5_reg[28]/NET0131  & ~n18856 ;
  assign n18858 = \u2_L5_reg[28]/NET0131  & n18856 ;
  assign n18859 = ~n18857 & ~n18858 ;
  assign n18863 = n18065 & n18129 ;
  assign n18864 = ~n18114 & ~n18863 ;
  assign n18865 = ~n18121 & n18864 ;
  assign n18866 = n18053 & ~n18865 ;
  assign n18860 = n18078 & n18106 ;
  assign n18861 = ~n18815 & ~n18860 ;
  assign n18862 = ~n18053 & ~n18861 ;
  assign n18867 = n18083 & n18088 ;
  assign n18868 = ~n18080 & ~n18867 ;
  assign n18869 = ~n18862 & n18868 ;
  assign n18870 = ~n18866 & n18869 ;
  assign n18871 = ~n18104 & ~n18870 ;
  assign n18875 = n18053 & n18083 ;
  assign n18876 = ~n18860 & ~n18875 ;
  assign n18877 = ~n18072 & ~n18876 ;
  assign n18872 = ~n18065 & n18108 ;
  assign n18873 = ~n18129 & ~n18872 ;
  assign n18874 = ~n18053 & ~n18873 ;
  assign n18878 = n18072 & n18092 ;
  assign n18879 = ~n18874 & ~n18878 ;
  assign n18880 = ~n18877 & n18879 ;
  assign n18881 = n18104 & ~n18880 ;
  assign n18882 = n18072 & n18808 ;
  assign n18883 = ~n18053 & ~n18107 ;
  assign n18884 = ~n18882 & n18883 ;
  assign n18885 = ~n18093 & ~n18112 ;
  assign n18886 = ~n18114 & n18885 ;
  assign n18887 = n18053 & n18072 ;
  assign n18888 = ~n18886 & n18887 ;
  assign n18889 = ~n18884 & ~n18888 ;
  assign n18890 = ~n18881 & n18889 ;
  assign n18891 = ~n18871 & n18890 ;
  assign n18892 = ~\u2_L5_reg[4]/NET0131  & ~n18891 ;
  assign n18893 = \u2_L5_reg[4]/NET0131  & n18891 ;
  assign n18894 = ~n18892 & ~n18893 ;
  assign n18914 = n18717 & n18766 ;
  assign n18913 = ~n18734 & n18765 ;
  assign n18915 = n18741 & ~n18913 ;
  assign n18916 = ~n18914 & n18915 ;
  assign n18917 = ~n18834 & ~n18916 ;
  assign n18912 = n18745 & ~n18754 ;
  assign n18918 = ~n18826 & ~n18912 ;
  assign n18919 = ~n18751 & n18918 ;
  assign n18920 = ~n18917 & n18919 ;
  assign n18921 = n18705 & ~n18920 ;
  assign n18895 = ~n18734 & n18825 ;
  assign n18896 = ~n18755 & ~n18895 ;
  assign n18897 = n18741 & ~n18896 ;
  assign n18898 = ~n18726 & n18741 ;
  assign n18899 = n18742 & n18898 ;
  assign n18900 = ~n18711 & n18746 ;
  assign n18901 = ~n18756 & n18900 ;
  assign n18902 = ~n18899 & ~n18901 ;
  assign n18903 = ~n18897 & n18902 ;
  assign n18904 = ~n18705 & ~n18903 ;
  assign n18905 = ~n18711 & n18726 ;
  assign n18906 = ~n18771 & ~n18905 ;
  assign n18907 = ~n18843 & n18906 ;
  assign n18908 = ~n18705 & ~n18907 ;
  assign n18909 = ~n18774 & ~n18826 ;
  assign n18910 = ~n18908 & n18909 ;
  assign n18911 = ~n18741 & ~n18910 ;
  assign n18922 = ~n18904 & ~n18911 ;
  assign n18923 = ~n18921 & n18922 ;
  assign n18924 = ~\u2_L5_reg[13]/NET0131  & n18923 ;
  assign n18925 = \u2_L5_reg[13]/NET0131  & ~n18923 ;
  assign n18926 = ~n18924 & ~n18925 ;
  assign n18927 = ~n18053 & n18059 ;
  assign n18928 = ~n18863 & ~n18927 ;
  assign n18929 = ~n18078 & ~n18928 ;
  assign n18933 = n18104 & ~n18872 ;
  assign n18934 = ~n18929 & n18933 ;
  assign n18930 = n18072 & ~n18885 ;
  assign n18931 = ~n18117 & ~n18124 ;
  assign n18932 = n18053 & ~n18931 ;
  assign n18935 = ~n18930 & ~n18932 ;
  assign n18936 = n18934 & n18935 ;
  assign n18939 = n18059 & ~n18108 ;
  assign n18940 = ~n18860 & ~n18939 ;
  assign n18941 = n18053 & ~n18940 ;
  assign n18938 = ~n18053 & ~n18885 ;
  assign n18937 = n18072 & n18084 ;
  assign n18942 = ~n18104 & ~n18937 ;
  assign n18943 = ~n18938 & n18942 ;
  assign n18944 = ~n18941 & n18943 ;
  assign n18945 = ~n18936 & ~n18944 ;
  assign n18946 = ~n18078 & n18867 ;
  assign n18947 = ~n18120 & ~n18946 ;
  assign n18948 = ~n18945 & n18947 ;
  assign n18949 = ~\u2_L5_reg[19]/NET0131  & ~n18948 ;
  assign n18950 = \u2_L5_reg[19]/NET0131  & n18948 ;
  assign n18951 = ~n18949 & ~n18950 ;
  assign n18953 = n17977 & n17991 ;
  assign n18972 = ~n17997 & ~n18020 ;
  assign n18973 = ~n18953 & n18972 ;
  assign n18974 = n17958 & ~n18973 ;
  assign n18975 = ~n18018 & ~n18536 ;
  assign n18976 = ~n18974 & n18975 ;
  assign n18977 = ~n17964 & ~n18976 ;
  assign n18967 = n17964 & ~n18034 ;
  assign n18968 = n17993 & n18967 ;
  assign n18969 = ~n18015 & ~n18539 ;
  assign n18970 = ~n18968 & n18969 ;
  assign n18971 = n17958 & ~n18970 ;
  assign n18954 = n17964 & ~n18011 ;
  assign n18955 = ~n18953 & n18954 ;
  assign n18952 = ~n17964 & ~n18020 ;
  assign n18956 = ~n17970 & ~n18952 ;
  assign n18957 = ~n18955 & n18956 ;
  assign n18960 = n18003 & ~n18537 ;
  assign n18961 = ~n18014 & ~n18960 ;
  assign n18962 = ~n18035 & ~n18961 ;
  assign n18959 = ~n17983 & n18537 ;
  assign n18958 = n17971 & n18019 ;
  assign n18963 = ~n18017 & ~n18958 ;
  assign n18964 = ~n18959 & n18963 ;
  assign n18965 = ~n18962 & n18964 ;
  assign n18966 = ~n17958 & ~n18965 ;
  assign n18978 = ~n18957 & ~n18966 ;
  assign n18979 = ~n18971 & n18978 ;
  assign n18980 = ~n18977 & n18979 ;
  assign n18981 = \u2_L5_reg[23]/NET0131  & ~n18980 ;
  assign n18982 = ~\u2_L5_reg[23]/NET0131  & n18980 ;
  assign n18983 = ~n18981 & ~n18982 ;
  assign n18996 = ~n18298 & ~n18596 ;
  assign n18997 = ~n18242 & ~n18611 ;
  assign n18998 = ~n18996 & n18997 ;
  assign n18994 = n18242 & ~n18312 ;
  assign n18995 = ~n18488 & n18994 ;
  assign n18999 = ~n18285 & ~n18598 ;
  assign n19000 = ~n18302 & n18999 ;
  assign n19001 = ~n18995 & n19000 ;
  assign n19002 = ~n18998 & n19001 ;
  assign n19003 = n18276 & ~n19002 ;
  assign n18985 = ~n18311 & ~n18593 ;
  assign n18986 = n18242 & ~n18487 ;
  assign n18987 = ~n18985 & n18986 ;
  assign n18984 = n18496 & n18611 ;
  assign n18988 = ~n18310 & ~n18615 ;
  assign n18989 = ~n18984 & n18988 ;
  assign n18990 = ~n18987 & n18989 ;
  assign n18991 = ~n18276 & ~n18990 ;
  assign n18992 = ~n18242 & n18314 ;
  assign n18993 = n18278 & n18499 ;
  assign n19004 = ~n18270 & ~n18993 ;
  assign n19005 = ~n18992 & n19004 ;
  assign n19006 = ~n18991 & n19005 ;
  assign n19007 = ~n19003 & n19006 ;
  assign n19008 = ~\u2_L5_reg[27]/NET0131  & ~n19007 ;
  assign n19009 = \u2_L5_reg[27]/NET0131  & n19007 ;
  assign n19010 = ~n19008 & ~n19009 ;
  assign n19013 = ~n17895 & ~n17924 ;
  assign n19014 = ~n18374 & ~n19013 ;
  assign n19015 = ~n17870 & n17894 ;
  assign n19016 = n17877 & n19015 ;
  assign n19017 = ~n19014 & ~n19016 ;
  assign n19018 = ~n17907 & ~n19017 ;
  assign n19011 = n17877 & n17937 ;
  assign n19012 = ~n18369 & n19011 ;
  assign n19019 = ~n17921 & ~n17934 ;
  assign n19020 = n17907 & ~n19019 ;
  assign n19021 = ~n19012 & ~n19020 ;
  assign n19022 = ~n19018 & n19021 ;
  assign n19023 = n17887 & ~n19022 ;
  assign n19024 = n17879 & n17937 ;
  assign n19028 = n17878 & n17893 ;
  assign n19029 = ~n19024 & ~n19028 ;
  assign n19030 = n17915 & n19029 ;
  assign n19025 = ~n17941 & ~n19015 ;
  assign n19026 = n17907 & ~n19025 ;
  assign n19027 = ~n17941 & n18378 ;
  assign n19031 = ~n19026 & ~n19027 ;
  assign n19032 = n19030 & n19031 ;
  assign n19033 = ~n17887 & ~n19032 ;
  assign n19034 = n17907 & n17911 ;
  assign n19035 = n17879 & n17894 ;
  assign n19036 = ~n17913 & ~n19035 ;
  assign n19037 = ~n17907 & ~n19036 ;
  assign n19038 = ~n19034 & ~n19037 ;
  assign n19039 = ~n19033 & n19038 ;
  assign n19040 = ~n19023 & n19039 ;
  assign n19041 = \u2_L5_reg[32]/NET0131  & n19040 ;
  assign n19042 = ~\u2_L5_reg[32]/NET0131  & ~n19040 ;
  assign n19043 = ~n19041 & ~n19042 ;
  assign n19077 = decrypt_pad & ~\u2_uk_K_r5_reg[47]/NET0131  ;
  assign n19078 = ~decrypt_pad & ~\u2_uk_K_r5_reg[12]/NET0131  ;
  assign n19079 = ~n19077 & ~n19078 ;
  assign n19080 = \u2_R5_reg[12]/NET0131  & ~n19079 ;
  assign n19081 = ~\u2_R5_reg[12]/NET0131  & n19079 ;
  assign n19082 = ~n19080 & ~n19081 ;
  assign n19044 = decrypt_pad & ~\u2_uk_K_r5_reg[3]/NET0131  ;
  assign n19045 = ~decrypt_pad & ~\u2_uk_K_r5_reg[25]/NET0131  ;
  assign n19046 = ~n19044 & ~n19045 ;
  assign n19047 = \u2_R5_reg[13]/NET0131  & ~n19046 ;
  assign n19048 = ~\u2_R5_reg[13]/NET0131  & n19046 ;
  assign n19049 = ~n19047 & ~n19048 ;
  assign n19057 = decrypt_pad & ~\u2_uk_K_r5_reg[26]/NET0131  ;
  assign n19058 = ~decrypt_pad & ~\u2_uk_K_r5_reg[48]/NET0131  ;
  assign n19059 = ~n19057 & ~n19058 ;
  assign n19060 = \u2_R5_reg[8]/NET0131  & ~n19059 ;
  assign n19061 = ~\u2_R5_reg[8]/NET0131  & n19059 ;
  assign n19062 = ~n19060 & ~n19061 ;
  assign n19064 = ~n19049 & ~n19062 ;
  assign n19065 = n19049 & n19062 ;
  assign n19066 = ~n19064 & ~n19065 ;
  assign n19050 = decrypt_pad & ~\u2_uk_K_r5_reg[55]/NET0131  ;
  assign n19051 = ~decrypt_pad & ~\u2_uk_K_r5_reg[20]/NET0131  ;
  assign n19052 = ~n19050 & ~n19051 ;
  assign n19053 = \u2_R5_reg[9]/NET0131  & ~n19052 ;
  assign n19054 = ~\u2_R5_reg[9]/NET0131  & n19052 ;
  assign n19055 = ~n19053 & ~n19054 ;
  assign n19067 = decrypt_pad & ~\u2_uk_K_r5_reg[6]/NET0131  ;
  assign n19068 = ~decrypt_pad & ~\u2_uk_K_r5_reg[53]/NET0131  ;
  assign n19069 = ~n19067 & ~n19068 ;
  assign n19070 = \u2_R5_reg[10]/NET0131  & ~n19069 ;
  assign n19071 = ~\u2_R5_reg[10]/NET0131  & n19069 ;
  assign n19072 = ~n19070 & ~n19071 ;
  assign n19118 = ~n19055 & n19072 ;
  assign n19119 = ~n19066 & n19118 ;
  assign n19107 = n19049 & ~n19062 ;
  assign n19108 = n19055 & n19107 ;
  assign n19089 = decrypt_pad & ~\u2_uk_K_r5_reg[32]/NET0131  ;
  assign n19090 = ~decrypt_pad & ~\u2_uk_K_r5_reg[54]/NET0131  ;
  assign n19091 = ~n19089 & ~n19090 ;
  assign n19092 = \u2_R5_reg[11]/NET0131  & ~n19091 ;
  assign n19093 = ~\u2_R5_reg[11]/NET0131  & n19091 ;
  assign n19094 = ~n19092 & ~n19093 ;
  assign n19109 = n19072 & ~n19094 ;
  assign n19110 = n19108 & n19109 ;
  assign n19115 = ~n19049 & n19055 ;
  assign n19116 = n19072 & n19115 ;
  assign n19117 = n19062 & n19116 ;
  assign n19120 = ~n19110 & ~n19117 ;
  assign n19121 = ~n19119 & n19120 ;
  assign n19100 = n19055 & ~n19072 ;
  assign n19111 = n19049 & n19094 ;
  assign n19112 = n19066 & ~n19111 ;
  assign n19113 = n19100 & ~n19112 ;
  assign n19084 = ~n19055 & ~n19072 ;
  assign n19114 = n19084 & n19112 ;
  assign n19122 = ~n19113 & ~n19114 ;
  assign n19123 = n19121 & n19122 ;
  assign n19124 = ~n19082 & ~n19123 ;
  assign n19056 = n19049 & ~n19055 ;
  assign n19063 = ~n19055 & n19062 ;
  assign n19073 = ~n19062 & ~n19072 ;
  assign n19074 = ~n19063 & ~n19073 ;
  assign n19075 = n19066 & n19074 ;
  assign n19076 = ~n19056 & ~n19075 ;
  assign n19083 = ~n19076 & n19082 ;
  assign n19085 = n19064 & n19084 ;
  assign n19086 = n19056 & n19072 ;
  assign n19087 = ~n19085 & ~n19086 ;
  assign n19088 = ~n19083 & n19087 ;
  assign n19095 = ~n19088 & n19094 ;
  assign n19096 = n19072 & n19082 ;
  assign n19097 = n19055 & n19064 ;
  assign n19098 = n19096 & n19097 ;
  assign n19099 = n19082 & ~n19094 ;
  assign n19101 = n19049 & n19100 ;
  assign n19102 = ~n19049 & n19063 ;
  assign n19103 = n19055 & n19065 ;
  assign n19104 = ~n19102 & ~n19103 ;
  assign n19105 = ~n19101 & n19104 ;
  assign n19106 = n19099 & ~n19105 ;
  assign n19125 = ~n19098 & ~n19106 ;
  assign n19126 = ~n19095 & n19125 ;
  assign n19127 = ~n19124 & n19126 ;
  assign n19128 = ~\u2_L5_reg[6]/NET0131  & ~n19127 ;
  assign n19129 = \u2_L5_reg[6]/NET0131  & n19127 ;
  assign n19130 = ~n19128 & ~n19129 ;
  assign n19136 = ~n17877 & n18373 ;
  assign n19137 = ~n17916 & n19136 ;
  assign n19134 = n17870 & ~n18373 ;
  assign n19135 = n17877 & n19134 ;
  assign n19131 = n17912 & n17916 ;
  assign n19132 = ~n17887 & n17907 ;
  assign n19133 = n17887 & ~n17907 ;
  assign n19138 = ~n19132 & ~n19133 ;
  assign n19139 = ~n19131 & n19138 ;
  assign n19140 = ~n19135 & n19139 ;
  assign n19141 = ~n19137 & n19140 ;
  assign n19142 = ~n17910 & n18368 ;
  assign n19143 = ~n19011 & n19133 ;
  assign n19144 = ~n19134 & n19143 ;
  assign n19145 = ~n19142 & n19144 ;
  assign n19146 = ~n19141 & ~n19145 ;
  assign n19147 = ~n19016 & ~n19146 ;
  assign n19148 = ~n19015 & ~n19136 ;
  assign n19149 = ~n19135 & n19148 ;
  assign n19150 = ~n19131 & n19132 ;
  assign n19151 = ~n19149 & n19150 ;
  assign n19152 = ~n19147 & ~n19151 ;
  assign n19153 = ~\u2_L5_reg[7]/NET0131  & n19152 ;
  assign n19154 = \u2_L5_reg[7]/NET0131  & ~n19152 ;
  assign n19155 = ~n19153 & ~n19154 ;
  assign n19167 = ~n18432 & ~n18631 ;
  assign n19168 = n18393 & ~n19167 ;
  assign n19169 = n18429 & ~n18454 ;
  assign n19170 = ~n18637 & ~n19169 ;
  assign n19171 = ~n18393 & ~n19170 ;
  assign n19172 = ~n18413 & n18656 ;
  assign n19173 = ~n19171 & n19172 ;
  assign n19174 = ~n19168 & n19173 ;
  assign n19175 = ~n18452 & ~n19174 ;
  assign n19160 = ~n18399 & n18462 ;
  assign n19161 = ~n18637 & ~n19160 ;
  assign n19162 = n18393 & ~n19161 ;
  assign n19163 = ~n18399 & n18660 ;
  assign n19164 = n18479 & ~n19163 ;
  assign n19165 = ~n19162 & n19164 ;
  assign n19166 = n18452 & ~n19165 ;
  assign n19156 = n18429 & ~n18455 ;
  assign n19157 = ~n18428 & ~n19156 ;
  assign n19158 = n18393 & ~n19157 ;
  assign n19159 = n18399 & n18645 ;
  assign n19176 = ~n19158 & ~n19159 ;
  assign n19177 = ~n19166 & n19176 ;
  assign n19178 = ~n19175 & n19177 ;
  assign n19179 = ~\u2_L5_reg[8]/NET0131  & ~n19178 ;
  assign n19180 = \u2_L5_reg[8]/NET0131  & n19178 ;
  assign n19181 = ~n19179 & ~n19180 ;
  assign n19182 = n19072 & ~n19108 ;
  assign n19184 = n19094 & n19097 ;
  assign n19183 = n19056 & ~n19062 ;
  assign n19185 = ~n19072 & ~n19183 ;
  assign n19186 = n19104 & n19185 ;
  assign n19187 = ~n19184 & n19186 ;
  assign n19188 = ~n19182 & ~n19187 ;
  assign n19189 = n19064 & n19072 ;
  assign n19190 = ~n19055 & n19189 ;
  assign n19191 = n19094 & ~n19117 ;
  assign n19192 = ~n19190 & n19191 ;
  assign n19193 = n19062 & n19072 ;
  assign n19194 = ~n19049 & ~n19073 ;
  assign n19195 = ~n19193 & n19194 ;
  assign n19196 = ~n19192 & n19195 ;
  assign n19197 = ~n19188 & ~n19196 ;
  assign n19198 = n19082 & ~n19197 ;
  assign n19199 = ~n19055 & n19193 ;
  assign n19200 = ~n19094 & ~n19199 ;
  assign n19201 = ~n19192 & ~n19200 ;
  assign n19206 = n19064 & ~n19072 ;
  assign n19207 = ~n19103 & ~n19183 ;
  assign n19208 = ~n19206 & n19207 ;
  assign n19209 = ~n19094 & ~n19208 ;
  assign n19203 = ~n19064 & n19094 ;
  assign n19202 = ~n19055 & ~n19065 ;
  assign n19204 = ~n19103 & ~n19202 ;
  assign n19205 = n19203 & n19204 ;
  assign n19210 = ~n19085 & ~n19205 ;
  assign n19211 = ~n19209 & n19210 ;
  assign n19212 = ~n19082 & ~n19211 ;
  assign n19213 = ~n19201 & ~n19212 ;
  assign n19214 = ~n19198 & n19213 ;
  assign n19215 = ~\u2_L5_reg[16]/NET0131  & ~n19214 ;
  assign n19216 = \u2_L5_reg[16]/NET0131  & n19214 ;
  assign n19217 = ~n19215 & ~n19216 ;
  assign n19227 = ~n19072 & n19094 ;
  assign n19238 = ~n19055 & ~n19107 ;
  assign n19239 = n19227 & n19238 ;
  assign n19234 = ~n19084 & ~n19094 ;
  assign n19235 = ~n19066 & n19234 ;
  assign n19236 = ~n19063 & n19072 ;
  assign n19237 = n19203 & n19236 ;
  assign n19240 = ~n19235 & ~n19237 ;
  assign n19241 = ~n19239 & n19240 ;
  assign n19242 = ~n19114 & n19241 ;
  assign n19243 = n19082 & ~n19242 ;
  assign n19218 = n19049 & n19073 ;
  assign n19219 = ~n19189 & ~n19218 ;
  assign n19220 = ~n19097 & ~n19199 ;
  assign n19221 = n19219 & n19220 ;
  assign n19222 = n19094 & ~n19221 ;
  assign n19223 = ~n19049 & n19199 ;
  assign n19224 = ~n19222 & ~n19223 ;
  assign n19225 = ~n19082 & ~n19224 ;
  assign n19230 = ~n19066 & n19084 ;
  assign n19231 = ~n19075 & ~n19230 ;
  assign n19232 = ~n19082 & ~n19094 ;
  assign n19233 = ~n19231 & n19232 ;
  assign n19226 = n19103 & n19109 ;
  assign n19228 = ~n19102 & ~n19108 ;
  assign n19229 = n19227 & ~n19228 ;
  assign n19244 = ~n19226 & ~n19229 ;
  assign n19245 = ~n19233 & n19244 ;
  assign n19246 = ~n19225 & n19245 ;
  assign n19247 = ~n19243 & n19246 ;
  assign n19248 = ~\u2_L5_reg[24]/NET0131  & ~n19247 ;
  assign n19249 = \u2_L5_reg[24]/NET0131  & n19247 ;
  assign n19250 = ~n19248 & ~n19249 ;
  assign n19252 = ~n19072 & n19102 ;
  assign n19253 = n19219 & ~n19252 ;
  assign n19254 = n19082 & ~n19253 ;
  assign n19255 = ~n19115 & ~n19193 ;
  assign n19256 = ~n19082 & ~n19116 ;
  assign n19257 = ~n19255 & n19256 ;
  assign n19258 = ~n19254 & ~n19257 ;
  assign n19259 = n19094 & ~n19258 ;
  assign n19263 = n19072 & n19183 ;
  assign n19260 = ~n19055 & ~n19062 ;
  assign n19261 = ~n19094 & ~n19260 ;
  assign n19262 = n19255 & n19261 ;
  assign n19264 = ~n19230 & ~n19262 ;
  assign n19265 = ~n19263 & n19264 ;
  assign n19266 = ~n19082 & ~n19265 ;
  assign n19267 = ~n19097 & ~n19193 ;
  assign n19268 = n19099 & ~n19267 ;
  assign n19270 = n19055 & ~n19065 ;
  assign n19271 = n19096 & n19270 ;
  assign n19251 = n19109 & n19115 ;
  assign n19269 = n19111 & n19199 ;
  assign n19272 = ~n19251 & ~n19269 ;
  assign n19273 = ~n19271 & n19272 ;
  assign n19274 = ~n19268 & n19273 ;
  assign n19275 = ~n19266 & n19274 ;
  assign n19276 = ~n19259 & n19275 ;
  assign n19277 = \u2_L5_reg[30]/NET0131  & ~n19276 ;
  assign n19278 = ~\u2_L5_reg[30]/NET0131  & n19276 ;
  assign n19279 = ~n19277 & ~n19278 ;
  assign n19283 = ~n18399 & n18429 ;
  assign n19284 = ~n18458 & ~n19283 ;
  assign n19285 = n18393 & ~n19284 ;
  assign n19280 = n18393 & ~n18454 ;
  assign n19281 = ~n18440 & ~n18637 ;
  assign n19282 = ~n19280 & ~n19281 ;
  assign n19286 = ~n18452 & ~n19282 ;
  assign n19287 = ~n19285 & n19286 ;
  assign n19290 = n18412 & ~n18439 ;
  assign n19289 = ~n18412 & ~n18423 ;
  assign n19291 = n18393 & ~n19289 ;
  assign n19292 = ~n19290 & n19291 ;
  assign n19293 = ~n18393 & n18461 ;
  assign n19288 = n18399 & n18431 ;
  assign n19294 = ~n18434 & n18452 ;
  assign n19295 = ~n19288 & n19294 ;
  assign n19296 = ~n19293 & n19295 ;
  assign n19297 = ~n19292 & n19296 ;
  assign n19298 = ~n19287 & ~n19297 ;
  assign n19299 = n18433 & n18454 ;
  assign n19300 = ~n18393 & ~n19299 ;
  assign n19301 = ~n18474 & n19300 ;
  assign n19302 = ~n19160 & n19301 ;
  assign n19303 = n18393 & ~n18432 ;
  assign n19304 = ~n18477 & n19303 ;
  assign n19305 = ~n19302 & ~n19304 ;
  assign n19306 = ~n19298 & ~n19305 ;
  assign n19307 = ~\u2_L5_reg[3]/NET0131  & ~n19306 ;
  assign n19308 = \u2_L5_reg[3]/NET0131  & n19306 ;
  assign n19309 = ~n19307 & ~n19308 ;
  assign n19311 = n17977 & n18019 ;
  assign n19315 = ~n18035 & ~n19311 ;
  assign n19322 = ~n17964 & n19315 ;
  assign n19323 = ~n18034 & n18529 ;
  assign n19324 = n18528 & ~n19323 ;
  assign n19325 = ~n19322 & ~n19324 ;
  assign n19310 = n17990 & n18022 ;
  assign n19326 = n17970 & n18523 ;
  assign n19327 = ~n19310 & ~n19326 ;
  assign n19328 = ~n19325 & n19327 ;
  assign n19329 = ~n17958 & ~n19328 ;
  assign n19312 = n17970 & n19311 ;
  assign n19313 = ~n19310 & ~n19312 ;
  assign n19314 = ~n17964 & ~n19313 ;
  assign n19317 = n17970 & ~n17993 ;
  assign n19318 = ~n18523 & n19317 ;
  assign n19316 = n18012 & ~n19315 ;
  assign n19319 = ~n18536 & ~n19316 ;
  assign n19320 = ~n19318 & n19319 ;
  assign n19321 = n17958 & ~n19320 ;
  assign n19330 = ~n19314 & ~n19321 ;
  assign n19331 = ~n19329 & n19330 ;
  assign n19332 = ~\u2_L5_reg[9]/NET0131  & ~n19331 ;
  assign n19333 = \u2_L5_reg[9]/NET0131  & n19331 ;
  assign n19334 = ~n19332 & ~n19333 ;
  assign n19349 = n18705 & n18728 ;
  assign n19338 = ~n18711 & ~n18745 ;
  assign n19350 = ~n18746 & ~n18754 ;
  assign n19351 = ~n19338 & n19350 ;
  assign n19352 = ~n19349 & ~n19351 ;
  assign n19353 = n18741 & ~n19352 ;
  assign n19335 = ~n18741 & n18749 ;
  assign n19340 = ~n18705 & ~n18913 ;
  assign n19341 = ~n18826 & n19340 ;
  assign n19336 = ~n18772 & ~n18780 ;
  assign n19337 = n18718 & ~n19336 ;
  assign n19339 = n19336 & n19338 ;
  assign n19342 = ~n19337 & ~n19339 ;
  assign n19343 = n19341 & n19342 ;
  assign n19344 = ~n18746 & ~n18765 ;
  assign n19345 = n18757 & ~n19344 ;
  assign n19346 = n18705 & ~n18767 ;
  assign n19347 = ~n19345 & n19346 ;
  assign n19348 = ~n19343 & ~n19347 ;
  assign n19354 = ~n19335 & ~n19348 ;
  assign n19355 = ~n19353 & n19354 ;
  assign n19356 = ~\u2_L5_reg[18]/NET0131  & ~n19355 ;
  assign n19357 = \u2_L5_reg[18]/NET0131  & n19355 ;
  assign n19358 = ~n19356 & ~n19357 ;
  assign n19365 = decrypt_pad & ~\u2_uk_K_r4_reg[53]/NET0131  ;
  assign n19366 = ~decrypt_pad & ~\u2_uk_K_r4_reg[47]/NET0131  ;
  assign n19367 = ~n19365 & ~n19366 ;
  assign n19368 = \u2_R4_reg[5]/NET0131  & ~n19367 ;
  assign n19369 = ~\u2_R4_reg[5]/NET0131  & n19367 ;
  assign n19370 = ~n19368 & ~n19369 ;
  assign n19384 = decrypt_pad & ~\u2_uk_K_r4_reg[34]/NET0131  ;
  assign n19385 = ~decrypt_pad & ~\u2_uk_K_r4_reg[53]/NET0131  ;
  assign n19386 = ~n19384 & ~n19385 ;
  assign n19387 = \u2_R4_reg[32]/NET0131  & ~n19386 ;
  assign n19388 = ~\u2_R4_reg[32]/NET0131  & n19386 ;
  assign n19389 = ~n19387 & ~n19388 ;
  assign n19421 = ~n19370 & ~n19389 ;
  assign n19371 = decrypt_pad & ~\u2_uk_K_r4_reg[55]/NET0131  ;
  assign n19372 = ~decrypt_pad & ~\u2_uk_K_r4_reg[17]/NET0131  ;
  assign n19373 = ~n19371 & ~n19372 ;
  assign n19374 = \u2_R4_reg[1]/NET0131  & ~n19373 ;
  assign n19375 = ~\u2_R4_reg[1]/NET0131  & n19373 ;
  assign n19376 = ~n19374 & ~n19375 ;
  assign n19359 = decrypt_pad & ~\u2_uk_K_r4_reg[47]/NET0131  ;
  assign n19360 = ~decrypt_pad & ~\u2_uk_K_r4_reg[41]/NET0131  ;
  assign n19361 = ~n19359 & ~n19360 ;
  assign n19362 = \u2_R4_reg[3]/NET0131  & ~n19361 ;
  assign n19363 = ~\u2_R4_reg[3]/NET0131  & n19361 ;
  assign n19364 = ~n19362 & ~n19363 ;
  assign n19378 = decrypt_pad & ~\u2_uk_K_r4_reg[13]/NET0131  ;
  assign n19379 = ~decrypt_pad & ~\u2_uk_K_r4_reg[32]/NET0131  ;
  assign n19380 = ~n19378 & ~n19379 ;
  assign n19381 = \u2_R4_reg[2]/NET0131  & ~n19380 ;
  assign n19382 = ~\u2_R4_reg[2]/NET0131  & n19380 ;
  assign n19383 = ~n19381 & ~n19382 ;
  assign n19425 = n19364 & ~n19383 ;
  assign n19426 = n19376 & ~n19425 ;
  assign n19427 = ~n19389 & ~n19426 ;
  assign n19414 = ~n19376 & ~n19383 ;
  assign n19428 = ~n19370 & n19414 ;
  assign n19429 = ~n19427 & ~n19428 ;
  assign n19430 = ~n19421 & ~n19429 ;
  assign n19377 = n19370 & ~n19376 ;
  assign n19422 = n19383 & n19421 ;
  assign n19423 = ~n19377 & ~n19422 ;
  assign n19424 = n19364 & ~n19423 ;
  assign n19390 = n19383 & ~n19389 ;
  assign n19431 = ~n19376 & n19390 ;
  assign n19398 = decrypt_pad & ~\u2_uk_K_r4_reg[25]/NET0131  ;
  assign n19399 = ~decrypt_pad & ~\u2_uk_K_r4_reg[19]/NET0131  ;
  assign n19400 = ~n19398 & ~n19399 ;
  assign n19401 = \u2_R4_reg[4]/NET0131  & ~n19400 ;
  assign n19402 = ~\u2_R4_reg[4]/NET0131  & n19400 ;
  assign n19403 = ~n19401 & ~n19402 ;
  assign n19419 = ~n19364 & n19389 ;
  assign n19420 = n19376 & n19419 ;
  assign n19432 = n19403 & ~n19420 ;
  assign n19433 = ~n19431 & n19432 ;
  assign n19434 = ~n19424 & n19433 ;
  assign n19435 = ~n19430 & n19434 ;
  assign n19417 = n19364 & n19390 ;
  assign n19436 = n19370 & n19417 ;
  assign n19437 = ~n19383 & n19421 ;
  assign n19438 = ~n19436 & ~n19437 ;
  assign n19439 = n19376 & ~n19438 ;
  assign n19407 = n19370 & n19389 ;
  assign n19443 = ~n19414 & ~n19425 ;
  assign n19444 = n19407 & ~n19443 ;
  assign n19415 = n19364 & n19389 ;
  assign n19440 = n19376 & n19383 ;
  assign n19441 = ~n19370 & n19440 ;
  assign n19442 = n19415 & n19441 ;
  assign n19445 = ~n19403 & ~n19442 ;
  assign n19446 = ~n19444 & n19445 ;
  assign n19447 = ~n19439 & n19446 ;
  assign n19448 = ~n19435 & ~n19447 ;
  assign n19392 = ~n19370 & ~n19376 ;
  assign n19393 = n19389 & n19392 ;
  assign n19394 = n19383 & n19393 ;
  assign n19395 = ~n19383 & ~n19389 ;
  assign n19396 = ~n19377 & n19395 ;
  assign n19397 = ~n19394 & ~n19396 ;
  assign n19404 = ~n19397 & ~n19403 ;
  assign n19408 = n19376 & n19407 ;
  assign n19409 = n19383 & n19408 ;
  assign n19391 = n19377 & n19390 ;
  assign n19405 = n19376 & ~n19383 ;
  assign n19406 = ~n19370 & n19405 ;
  assign n19410 = ~n19391 & ~n19406 ;
  assign n19411 = ~n19409 & n19410 ;
  assign n19412 = ~n19404 & n19411 ;
  assign n19413 = ~n19364 & ~n19412 ;
  assign n19416 = n19414 & n19415 ;
  assign n19418 = n19392 & n19417 ;
  assign n19449 = ~n19416 & ~n19418 ;
  assign n19450 = ~n19413 & n19449 ;
  assign n19451 = ~n19448 & n19450 ;
  assign n19452 = ~\u2_L4_reg[31]/NET0131  & ~n19451 ;
  assign n19453 = \u2_L4_reg[31]/NET0131  & n19451 ;
  assign n19454 = ~n19452 & ~n19453 ;
  assign n19506 = decrypt_pad & ~\u2_uk_K_r4_reg[51]/NET0131  ;
  assign n19507 = ~decrypt_pad & ~\u2_uk_K_r4_reg[43]/NET0131  ;
  assign n19508 = ~n19506 & ~n19507 ;
  assign n19509 = \u2_R4_reg[24]/NET0131  & ~n19508 ;
  assign n19510 = ~\u2_R4_reg[24]/NET0131  & n19508 ;
  assign n19511 = ~n19509 & ~n19510 ;
  assign n19461 = decrypt_pad & ~\u2_uk_K_r4_reg[30]/NET0131  ;
  assign n19462 = ~decrypt_pad & ~\u2_uk_K_r4_reg[22]/NET0131  ;
  assign n19463 = ~n19461 & ~n19462 ;
  assign n19464 = \u2_R4_reg[20]/NET0131  & ~n19463 ;
  assign n19465 = ~\u2_R4_reg[20]/NET0131  & n19463 ;
  assign n19466 = ~n19464 & ~n19465 ;
  assign n19474 = decrypt_pad & ~\u2_uk_K_r4_reg[36]/NET0131  ;
  assign n19475 = ~decrypt_pad & ~\u2_uk_K_r4_reg[28]/NET0131  ;
  assign n19476 = ~n19474 & ~n19475 ;
  assign n19477 = \u2_R4_reg[22]/NET0131  & ~n19476 ;
  assign n19478 = ~\u2_R4_reg[22]/NET0131  & n19476 ;
  assign n19479 = ~n19477 & ~n19478 ;
  assign n19480 = decrypt_pad & ~\u2_uk_K_r4_reg[14]/NET0131  ;
  assign n19481 = ~decrypt_pad & ~\u2_uk_K_r4_reg[37]/NET0131  ;
  assign n19482 = ~n19480 & ~n19481 ;
  assign n19483 = \u2_R4_reg[21]/NET0131  & ~n19482 ;
  assign n19484 = ~\u2_R4_reg[21]/NET0131  & n19482 ;
  assign n19485 = ~n19483 & ~n19484 ;
  assign n19515 = ~n19479 & n19485 ;
  assign n19531 = n19466 & n19515 ;
  assign n19455 = decrypt_pad & ~\u2_uk_K_r4_reg[49]/NET0131  ;
  assign n19456 = ~decrypt_pad & ~\u2_uk_K_r4_reg[45]/NET0131  ;
  assign n19457 = ~n19455 & ~n19456 ;
  assign n19458 = \u2_R4_reg[23]/NET0131  & ~n19457 ;
  assign n19459 = ~\u2_R4_reg[23]/NET0131  & n19457 ;
  assign n19460 = ~n19458 & ~n19459 ;
  assign n19488 = ~n19466 & n19485 ;
  assign n19489 = n19479 & n19488 ;
  assign n19532 = ~n19460 & ~n19489 ;
  assign n19533 = ~n19531 & n19532 ;
  assign n19467 = decrypt_pad & ~\u2_uk_K_r4_reg[15]/NET0131  ;
  assign n19468 = ~decrypt_pad & ~\u2_uk_K_r4_reg[7]/NET0131  ;
  assign n19469 = ~n19467 & ~n19468 ;
  assign n19470 = \u2_R4_reg[25]/NET0131  & ~n19469 ;
  assign n19471 = ~\u2_R4_reg[25]/NET0131  & n19469 ;
  assign n19472 = ~n19470 & ~n19471 ;
  assign n19523 = n19472 & ~n19485 ;
  assign n19524 = ~n19466 & n19523 ;
  assign n19525 = n19460 & ~n19524 ;
  assign n19534 = n19479 & ~n19485 ;
  assign n19535 = n19466 & n19534 ;
  assign n19536 = ~n19466 & ~n19479 ;
  assign n19537 = ~n19535 & ~n19536 ;
  assign n19538 = n19525 & n19537 ;
  assign n19539 = ~n19533 & ~n19538 ;
  assign n19490 = n19466 & n19472 ;
  assign n19501 = ~n19485 & n19490 ;
  assign n19528 = n19479 & n19501 ;
  assign n19473 = n19466 & ~n19472 ;
  assign n19495 = ~n19460 & ~n19479 ;
  assign n19529 = ~n19495 & ~n19515 ;
  assign n19530 = n19473 & ~n19529 ;
  assign n19540 = ~n19528 & ~n19530 ;
  assign n19541 = ~n19539 & n19540 ;
  assign n19542 = ~n19511 & ~n19541 ;
  assign n19491 = n19485 & n19490 ;
  assign n19486 = ~n19479 & ~n19485 ;
  assign n19487 = n19473 & n19486 ;
  assign n19492 = ~n19487 & ~n19489 ;
  assign n19493 = ~n19491 & n19492 ;
  assign n19494 = n19460 & ~n19493 ;
  assign n19496 = ~n19488 & ~n19490 ;
  assign n19497 = ~n19460 & n19496 ;
  assign n19498 = ~n19495 & ~n19497 ;
  assign n19499 = n19472 & n19485 ;
  assign n19500 = ~n19466 & n19499 ;
  assign n19502 = ~n19479 & ~n19500 ;
  assign n19503 = ~n19501 & n19502 ;
  assign n19504 = ~n19498 & ~n19503 ;
  assign n19505 = ~n19494 & ~n19504 ;
  assign n19512 = ~n19505 & n19511 ;
  assign n19521 = n19473 & n19485 ;
  assign n19522 = ~n19460 & ~n19521 ;
  assign n19526 = ~n19479 & ~n19522 ;
  assign n19527 = ~n19525 & n19526 ;
  assign n19516 = ~n19490 & ~n19515 ;
  assign n19513 = ~n19466 & ~n19472 ;
  assign n19514 = ~n19479 & ~n19513 ;
  assign n19517 = n19460 & ~n19514 ;
  assign n19518 = ~n19516 & n19517 ;
  assign n19519 = ~n19485 & n19513 ;
  assign n19520 = n19495 & n19519 ;
  assign n19543 = ~n19518 & ~n19520 ;
  assign n19544 = ~n19527 & n19543 ;
  assign n19545 = ~n19512 & n19544 ;
  assign n19546 = ~n19542 & n19545 ;
  assign n19547 = \u2_L4_reg[11]/NET0131  & ~n19546 ;
  assign n19548 = ~\u2_L4_reg[11]/NET0131  & n19546 ;
  assign n19549 = ~n19547 & ~n19548 ;
  assign n19550 = decrypt_pad & ~\u2_uk_K_r4_reg[31]/P0001  ;
  assign n19551 = ~decrypt_pad & ~\u2_uk_K_r4_reg[50]/NET0131  ;
  assign n19552 = ~n19550 & ~n19551 ;
  assign n19553 = \u2_R4_reg[28]/NET0131  & ~n19552 ;
  assign n19554 = ~\u2_R4_reg[28]/NET0131  & n19552 ;
  assign n19555 = ~n19553 & ~n19554 ;
  assign n19556 = decrypt_pad & ~\u2_uk_K_r4_reg[16]/NET0131  ;
  assign n19557 = ~decrypt_pad & ~\u2_uk_K_r4_reg[8]/NET0131  ;
  assign n19558 = ~n19556 & ~n19557 ;
  assign n19559 = \u2_R4_reg[27]/NET0131  & ~n19558 ;
  assign n19560 = ~\u2_R4_reg[27]/NET0131  & n19558 ;
  assign n19561 = ~n19559 & ~n19560 ;
  assign n19562 = decrypt_pad & ~\u2_uk_K_r4_reg[22]/NET0131  ;
  assign n19563 = ~decrypt_pad & ~\u2_uk_K_r4_reg[14]/NET0131  ;
  assign n19564 = ~n19562 & ~n19563 ;
  assign n19565 = \u2_R4_reg[25]/NET0131  & ~n19564 ;
  assign n19566 = ~\u2_R4_reg[25]/NET0131  & n19564 ;
  assign n19567 = ~n19565 & ~n19566 ;
  assign n19568 = decrypt_pad & ~\u2_uk_K_r4_reg[7]/NET0131  ;
  assign n19569 = ~decrypt_pad & ~\u2_uk_K_r4_reg[30]/NET0131  ;
  assign n19570 = ~n19568 & ~n19569 ;
  assign n19571 = \u2_R4_reg[26]/NET0131  & ~n19570 ;
  assign n19572 = ~\u2_R4_reg[26]/NET0131  & n19570 ;
  assign n19573 = ~n19571 & ~n19572 ;
  assign n19574 = ~n19567 & ~n19573 ;
  assign n19575 = decrypt_pad & ~\u2_uk_K_r4_reg[42]/NET0131  ;
  assign n19576 = ~decrypt_pad & ~\u2_uk_K_r4_reg[38]/NET0131  ;
  assign n19577 = ~n19575 & ~n19576 ;
  assign n19578 = \u2_R4_reg[24]/NET0131  & ~n19577 ;
  assign n19579 = ~\u2_R4_reg[24]/NET0131  & n19577 ;
  assign n19580 = ~n19578 & ~n19579 ;
  assign n19581 = n19574 & n19580 ;
  assign n19584 = decrypt_pad & ~\u2_uk_K_r4_reg[50]/NET0131  ;
  assign n19585 = ~decrypt_pad & ~\u2_uk_K_r4_reg[42]/NET0131  ;
  assign n19586 = ~n19584 & ~n19585 ;
  assign n19587 = \u2_R4_reg[29]/NET0131  & ~n19586 ;
  assign n19588 = ~\u2_R4_reg[29]/NET0131  & n19586 ;
  assign n19589 = ~n19587 & ~n19588 ;
  assign n19618 = n19581 & n19589 ;
  assign n19602 = ~n19580 & n19589 ;
  assign n19619 = n19567 & n19602 ;
  assign n19620 = ~n19618 & ~n19619 ;
  assign n19621 = ~n19561 & ~n19620 ;
  assign n19583 = n19567 & n19573 ;
  assign n19622 = ~n19574 & ~n19583 ;
  assign n19590 = ~n19573 & ~n19589 ;
  assign n19623 = n19561 & n19580 ;
  assign n19624 = ~n19590 & n19623 ;
  assign n19625 = n19622 & n19624 ;
  assign n19603 = ~n19567 & n19573 ;
  assign n19604 = n19602 & n19603 ;
  assign n19600 = ~n19580 & ~n19589 ;
  assign n19617 = n19574 & n19600 ;
  assign n19626 = ~n19604 & ~n19617 ;
  assign n19627 = ~n19625 & n19626 ;
  assign n19628 = ~n19621 & n19627 ;
  assign n19629 = n19555 & ~n19628 ;
  assign n19593 = ~n19567 & ~n19589 ;
  assign n19594 = n19573 & ~n19580 ;
  assign n19605 = n19593 & ~n19594 ;
  assign n19601 = n19583 & n19600 ;
  assign n19606 = ~n19601 & ~n19604 ;
  assign n19607 = ~n19605 & n19606 ;
  assign n19608 = n19561 & ~n19607 ;
  assign n19591 = ~n19583 & ~n19590 ;
  assign n19592 = n19580 & ~n19591 ;
  assign n19595 = n19593 & n19594 ;
  assign n19596 = ~n19561 & ~n19595 ;
  assign n19597 = ~n19592 & n19596 ;
  assign n19582 = n19561 & ~n19581 ;
  assign n19598 = ~n19555 & ~n19582 ;
  assign n19599 = ~n19597 & n19598 ;
  assign n19611 = ~n19561 & n19567 ;
  assign n19612 = ~n19555 & n19589 ;
  assign n19613 = ~n19611 & ~n19612 ;
  assign n19609 = ~n19573 & n19580 ;
  assign n19610 = ~n19594 & ~n19609 ;
  assign n19614 = n19561 & ~n19567 ;
  assign n19615 = n19610 & ~n19614 ;
  assign n19616 = ~n19613 & n19615 ;
  assign n19630 = ~n19599 & ~n19616 ;
  assign n19631 = ~n19608 & n19630 ;
  assign n19632 = ~n19629 & n19631 ;
  assign n19633 = ~\u2_L4_reg[22]/NET0131  & ~n19632 ;
  assign n19634 = \u2_L4_reg[22]/NET0131  & n19632 ;
  assign n19635 = ~n19633 & ~n19634 ;
  assign n19637 = n19370 & n19405 ;
  assign n19638 = ~n19441 & ~n19637 ;
  assign n19639 = ~n19389 & ~n19638 ;
  assign n19636 = ~n19393 & ~n19408 ;
  assign n19640 = n19364 & n19636 ;
  assign n19641 = ~n19639 & n19640 ;
  assign n19642 = ~n19407 & ~n19421 ;
  assign n19643 = ~n19376 & ~n19642 ;
  assign n19644 = ~n19364 & ~n19437 ;
  assign n19645 = ~n19643 & n19644 ;
  assign n19646 = ~n19641 & ~n19645 ;
  assign n19647 = ~n19431 & ~n19441 ;
  assign n19648 = ~n19421 & ~n19647 ;
  assign n19649 = ~n19403 & ~n19648 ;
  assign n19650 = ~n19646 & n19649 ;
  assign n19651 = n19407 & n19414 ;
  assign n19652 = ~n19389 & ~n19414 ;
  assign n19653 = ~n19651 & ~n19652 ;
  assign n19654 = n19364 & ~n19653 ;
  assign n19655 = n19389 & n19406 ;
  assign n19656 = ~n19364 & ~n19389 ;
  assign n19657 = n19414 & n19656 ;
  assign n19660 = n19403 & ~n19657 ;
  assign n19658 = n19370 & n19440 ;
  assign n19659 = n19383 & n19419 ;
  assign n19661 = ~n19658 & ~n19659 ;
  assign n19662 = n19660 & n19661 ;
  assign n19663 = ~n19655 & n19662 ;
  assign n19664 = ~n19654 & n19663 ;
  assign n19665 = ~n19650 & ~n19664 ;
  assign n19666 = ~\u2_L4_reg[17]/NET0131  & n19665 ;
  assign n19667 = \u2_L4_reg[17]/NET0131  & ~n19665 ;
  assign n19668 = ~n19666 & ~n19667 ;
  assign n19669 = decrypt_pad & ~\u2_uk_K_r4_reg[10]/NET0131  ;
  assign n19670 = ~decrypt_pad & ~\u2_uk_K_r4_reg[4]/NET0131  ;
  assign n19671 = ~n19669 & ~n19670 ;
  assign n19672 = \u2_R4_reg[13]/NET0131  & ~n19671 ;
  assign n19673 = ~\u2_R4_reg[13]/NET0131  & n19671 ;
  assign n19674 = ~n19672 & ~n19673 ;
  assign n19675 = decrypt_pad & ~\u2_uk_K_r4_reg[48]/NET0131  ;
  assign n19676 = ~decrypt_pad & ~\u2_uk_K_r4_reg[10]/NET0131  ;
  assign n19677 = ~n19675 & ~n19676 ;
  assign n19678 = \u2_R4_reg[12]/NET0131  & ~n19677 ;
  assign n19679 = ~\u2_R4_reg[12]/NET0131  & n19677 ;
  assign n19680 = ~n19678 & ~n19679 ;
  assign n19681 = decrypt_pad & ~\u2_uk_K_r4_reg[32]/NET0131  ;
  assign n19682 = ~decrypt_pad & ~\u2_uk_K_r4_reg[26]/NET0131  ;
  assign n19683 = ~n19681 & ~n19682 ;
  assign n19684 = \u2_R4_reg[17]/NET0131  & ~n19683 ;
  assign n19685 = ~\u2_R4_reg[17]/NET0131  & n19683 ;
  assign n19686 = ~n19684 & ~n19685 ;
  assign n19687 = ~n19680 & n19686 ;
  assign n19688 = decrypt_pad & ~\u2_uk_K_r4_reg[19]/NET0131  ;
  assign n19689 = ~decrypt_pad & ~\u2_uk_K_r4_reg[13]/NET0131  ;
  assign n19690 = ~n19688 & ~n19689 ;
  assign n19691 = \u2_R4_reg[15]/NET0131  & ~n19690 ;
  assign n19692 = ~\u2_R4_reg[15]/NET0131  & n19690 ;
  assign n19693 = ~n19691 & ~n19692 ;
  assign n19694 = n19687 & n19693 ;
  assign n19695 = ~n19674 & n19694 ;
  assign n19696 = decrypt_pad & ~\u2_uk_K_r4_reg[27]/P0001  ;
  assign n19697 = ~decrypt_pad & ~\u2_uk_K_r4_reg[46]/NET0131  ;
  assign n19698 = ~n19696 & ~n19697 ;
  assign n19699 = \u2_R4_reg[16]/NET0131  & ~n19698 ;
  assign n19700 = ~\u2_R4_reg[16]/NET0131  & n19698 ;
  assign n19701 = ~n19699 & ~n19700 ;
  assign n19726 = ~n19695 & n19701 ;
  assign n19715 = n19680 & ~n19686 ;
  assign n19716 = n19674 & n19715 ;
  assign n19717 = n19693 & n19716 ;
  assign n19702 = n19674 & ~n19680 ;
  assign n19718 = ~n19674 & n19680 ;
  assign n19719 = ~n19702 & ~n19718 ;
  assign n19703 = decrypt_pad & ~\u2_uk_K_r4_reg[11]/NET0131  ;
  assign n19704 = ~decrypt_pad & ~\u2_uk_K_r4_reg[5]/NET0131  ;
  assign n19705 = ~n19703 & ~n19704 ;
  assign n19706 = \u2_R4_reg[14]/NET0131  & ~n19705 ;
  assign n19707 = ~\u2_R4_reg[14]/NET0131  & n19705 ;
  assign n19708 = ~n19706 & ~n19707 ;
  assign n19720 = ~n19693 & ~n19708 ;
  assign n19721 = ~n19719 & n19720 ;
  assign n19727 = ~n19717 & ~n19721 ;
  assign n19728 = n19726 & n19727 ;
  assign n19709 = n19686 & ~n19708 ;
  assign n19710 = n19702 & n19709 ;
  assign n19711 = n19680 & n19686 ;
  assign n19712 = n19708 & n19711 ;
  assign n19713 = n19674 & n19712 ;
  assign n19714 = ~n19710 & ~n19713 ;
  assign n19722 = ~n19674 & ~n19686 ;
  assign n19723 = ~n19680 & n19722 ;
  assign n19724 = n19708 & n19723 ;
  assign n19725 = ~n19693 & n19724 ;
  assign n19729 = n19714 & ~n19725 ;
  assign n19730 = n19728 & n19729 ;
  assign n19739 = n19674 & n19711 ;
  assign n19740 = n19693 & ~n19723 ;
  assign n19741 = ~n19739 & n19740 ;
  assign n19742 = n19708 & n19715 ;
  assign n19743 = ~n19674 & n19686 ;
  assign n19744 = ~n19693 & ~n19743 ;
  assign n19745 = ~n19742 & n19744 ;
  assign n19746 = ~n19741 & ~n19745 ;
  assign n19737 = n19693 & n19708 ;
  assign n19738 = n19702 & n19737 ;
  assign n19733 = ~n19680 & ~n19708 ;
  assign n19734 = n19722 & n19733 ;
  assign n19747 = ~n19701 & ~n19734 ;
  assign n19748 = ~n19738 & n19747 ;
  assign n19731 = ~n19686 & n19702 ;
  assign n19732 = n19708 & n19731 ;
  assign n19735 = ~n19708 & n19718 ;
  assign n19736 = n19686 & n19735 ;
  assign n19749 = ~n19732 & ~n19736 ;
  assign n19750 = n19748 & n19749 ;
  assign n19751 = ~n19746 & n19750 ;
  assign n19752 = ~n19730 & ~n19751 ;
  assign n19753 = ~n19693 & ~n19710 ;
  assign n19754 = ~n19674 & n19708 ;
  assign n19755 = n19715 & n19754 ;
  assign n19756 = n19693 & ~n19755 ;
  assign n19757 = n19674 & ~n19708 ;
  assign n19758 = n19715 & n19757 ;
  assign n19759 = ~n19734 & ~n19758 ;
  assign n19760 = n19756 & n19759 ;
  assign n19761 = ~n19753 & ~n19760 ;
  assign n19762 = ~n19752 & ~n19761 ;
  assign n19763 = ~\u2_L4_reg[20]/NET0131  & ~n19762 ;
  assign n19764 = \u2_L4_reg[20]/NET0131  & n19762 ;
  assign n19765 = ~n19763 & ~n19764 ;
  assign n19782 = n19473 & ~n19485 ;
  assign n19783 = ~n19491 & ~n19782 ;
  assign n19784 = ~n19486 & ~n19489 ;
  assign n19785 = ~n19472 & ~n19784 ;
  assign n19786 = n19783 & ~n19785 ;
  assign n19787 = n19460 & ~n19786 ;
  assign n19766 = n19479 & n19521 ;
  assign n19773 = ~n19479 & ~n19496 ;
  assign n19788 = ~n19766 & ~n19773 ;
  assign n19789 = ~n19460 & ~n19788 ;
  assign n19790 = n19479 & n19524 ;
  assign n19791 = ~n19789 & ~n19790 ;
  assign n19792 = ~n19787 & n19791 ;
  assign n19793 = ~n19511 & ~n19792 ;
  assign n19767 = n19485 & n19536 ;
  assign n19768 = ~n19500 & ~n19767 ;
  assign n19769 = ~n19766 & n19768 ;
  assign n19770 = n19460 & ~n19769 ;
  assign n19774 = n19460 & ~n19523 ;
  assign n19775 = ~n19534 & n19774 ;
  assign n19771 = n19479 & ~n19490 ;
  assign n19772 = ~n19513 & n19771 ;
  assign n19776 = ~n19772 & ~n19773 ;
  assign n19777 = ~n19775 & n19776 ;
  assign n19778 = ~n19770 & ~n19777 ;
  assign n19779 = n19511 & ~n19778 ;
  assign n19780 = n19460 & n19472 ;
  assign n19781 = n19515 & n19780 ;
  assign n19794 = ~n19487 & ~n19781 ;
  assign n19795 = ~n19779 & n19794 ;
  assign n19796 = ~n19793 & n19795 ;
  assign n19797 = \u2_L4_reg[29]/NET0131  & ~n19796 ;
  assign n19798 = ~\u2_L4_reg[29]/NET0131  & n19796 ;
  assign n19799 = ~n19797 & ~n19798 ;
  assign n19800 = decrypt_pad & ~\u2_uk_K_r4_reg[26]/NET0131  ;
  assign n19801 = ~decrypt_pad & ~\u2_uk_K_r4_reg[20]/NET0131  ;
  assign n19802 = ~n19800 & ~n19801 ;
  assign n19803 = \u2_R4_reg[8]/NET0131  & ~n19802 ;
  assign n19804 = ~\u2_R4_reg[8]/NET0131  & n19802 ;
  assign n19805 = ~n19803 & ~n19804 ;
  assign n19806 = decrypt_pad & ~\u2_uk_K_r4_reg[18]/NET0131  ;
  assign n19807 = ~decrypt_pad & ~\u2_uk_K_r4_reg[12]/NET0131  ;
  assign n19808 = ~n19806 & ~n19807 ;
  assign n19809 = \u2_R4_reg[5]/NET0131  & ~n19808 ;
  assign n19810 = ~\u2_R4_reg[5]/NET0131  & n19808 ;
  assign n19811 = ~n19809 & ~n19810 ;
  assign n19812 = decrypt_pad & ~\u2_uk_K_r4_reg[6]/NET0131  ;
  assign n19813 = ~decrypt_pad & ~\u2_uk_K_r4_reg[25]/NET0131  ;
  assign n19814 = ~n19812 & ~n19813 ;
  assign n19815 = \u2_R4_reg[9]/NET0131  & ~n19814 ;
  assign n19816 = ~\u2_R4_reg[9]/NET0131  & n19814 ;
  assign n19817 = ~n19815 & ~n19816 ;
  assign n19818 = n19811 & ~n19817 ;
  assign n19819 = ~n19811 & n19817 ;
  assign n19820 = decrypt_pad & ~\u2_uk_K_r4_reg[39]/NET0131  ;
  assign n19821 = ~decrypt_pad & ~\u2_uk_K_r4_reg[33]/NET0131  ;
  assign n19822 = ~n19820 & ~n19821 ;
  assign n19823 = \u2_R4_reg[4]/NET0131  & ~n19822 ;
  assign n19824 = ~\u2_R4_reg[4]/NET0131  & n19822 ;
  assign n19825 = ~n19823 & ~n19824 ;
  assign n19826 = n19819 & ~n19825 ;
  assign n19827 = ~n19818 & ~n19826 ;
  assign n19828 = decrypt_pad & ~\u2_uk_K_r4_reg[41]/NET0131  ;
  assign n19829 = ~decrypt_pad & ~\u2_uk_K_r4_reg[3]/NET0131  ;
  assign n19830 = ~n19828 & ~n19829 ;
  assign n19831 = \u2_R4_reg[6]/NET0131  & ~n19830 ;
  assign n19832 = ~\u2_R4_reg[6]/NET0131  & n19830 ;
  assign n19833 = ~n19831 & ~n19832 ;
  assign n19834 = ~n19827 & ~n19833 ;
  assign n19835 = decrypt_pad & ~\u2_uk_K_r4_reg[3]/NET0131  ;
  assign n19836 = ~decrypt_pad & ~\u2_uk_K_r4_reg[54]/NET0131  ;
  assign n19837 = ~n19835 & ~n19836 ;
  assign n19838 = \u2_R4_reg[7]/NET0131  & ~n19837 ;
  assign n19839 = ~\u2_R4_reg[7]/NET0131  & n19837 ;
  assign n19840 = ~n19838 & ~n19839 ;
  assign n19841 = ~n19811 & n19833 ;
  assign n19842 = n19817 & n19825 ;
  assign n19843 = n19841 & n19842 ;
  assign n19844 = n19840 & n19843 ;
  assign n19858 = ~n19834 & ~n19844 ;
  assign n19845 = n19825 & n19833 ;
  assign n19846 = ~n19819 & n19845 ;
  assign n19847 = ~n19826 & ~n19846 ;
  assign n19848 = ~n19840 & ~n19847 ;
  assign n19852 = n19811 & ~n19833 ;
  assign n19853 = ~n19833 & n19840 ;
  assign n19854 = ~n19852 & ~n19853 ;
  assign n19849 = n19817 & ~n19825 ;
  assign n19850 = n19811 & ~n19849 ;
  assign n19851 = ~n19817 & ~n19833 ;
  assign n19855 = ~n19841 & ~n19851 ;
  assign n19856 = ~n19850 & n19855 ;
  assign n19857 = n19854 & n19856 ;
  assign n19859 = ~n19848 & ~n19857 ;
  assign n19860 = n19858 & n19859 ;
  assign n19861 = ~n19805 & ~n19860 ;
  assign n19874 = ~n19817 & ~n19825 ;
  assign n19878 = ~n19843 & ~n19874 ;
  assign n19879 = n19805 & ~n19878 ;
  assign n19880 = ~n19841 & n19849 ;
  assign n19881 = ~n19879 & ~n19880 ;
  assign n19882 = ~n19840 & ~n19852 ;
  assign n19883 = ~n19881 & n19882 ;
  assign n19868 = ~n19833 & n19842 ;
  assign n19869 = n19811 & n19868 ;
  assign n19862 = ~n19817 & n19825 ;
  assign n19863 = ~n19811 & n19862 ;
  assign n19864 = ~n19833 & n19863 ;
  assign n19865 = ~n19825 & n19833 ;
  assign n19866 = n19811 & n19840 ;
  assign n19867 = ~n19865 & n19866 ;
  assign n19870 = ~n19864 & ~n19867 ;
  assign n19871 = ~n19869 & n19870 ;
  assign n19872 = n19805 & ~n19871 ;
  assign n19875 = ~n19852 & ~n19874 ;
  assign n19873 = ~n19825 & ~n19841 ;
  assign n19876 = n19840 & ~n19873 ;
  assign n19877 = ~n19875 & n19876 ;
  assign n19884 = ~n19872 & ~n19877 ;
  assign n19885 = ~n19883 & n19884 ;
  assign n19886 = ~n19861 & n19885 ;
  assign n19887 = \u2_L4_reg[2]/NET0131  & n19886 ;
  assign n19888 = ~\u2_L4_reg[2]/NET0131  & ~n19886 ;
  assign n19889 = ~n19887 & ~n19888 ;
  assign n19893 = n19472 & n19536 ;
  assign n19894 = ~n19521 & ~n19893 ;
  assign n19895 = ~n19528 & n19894 ;
  assign n19896 = n19460 & ~n19895 ;
  assign n19890 = n19485 & n19513 ;
  assign n19891 = ~n19790 & ~n19890 ;
  assign n19892 = ~n19460 & ~n19891 ;
  assign n19897 = n19490 & n19495 ;
  assign n19898 = ~n19487 & ~n19897 ;
  assign n19899 = ~n19892 & n19898 ;
  assign n19900 = ~n19896 & n19899 ;
  assign n19901 = ~n19511 & ~n19900 ;
  assign n19905 = n19460 & n19490 ;
  assign n19906 = ~n19890 & ~n19905 ;
  assign n19907 = ~n19479 & ~n19906 ;
  assign n19902 = ~n19472 & n19515 ;
  assign n19903 = ~n19536 & ~n19902 ;
  assign n19904 = ~n19460 & ~n19903 ;
  assign n19908 = n19479 & n19499 ;
  assign n19909 = ~n19904 & ~n19908 ;
  assign n19910 = ~n19907 & n19909 ;
  assign n19911 = n19511 & ~n19910 ;
  assign n19912 = n19479 & n19783 ;
  assign n19913 = ~n19460 & ~n19514 ;
  assign n19914 = ~n19912 & n19913 ;
  assign n19915 = ~n19500 & ~n19519 ;
  assign n19916 = ~n19521 & n19915 ;
  assign n19917 = n19460 & n19479 ;
  assign n19918 = ~n19916 & n19917 ;
  assign n19919 = ~n19914 & ~n19918 ;
  assign n19920 = ~n19911 & n19919 ;
  assign n19921 = ~n19901 & n19920 ;
  assign n19922 = ~\u2_L4_reg[4]/NET0131  & ~n19921 ;
  assign n19923 = \u2_L4_reg[4]/NET0131  & n19921 ;
  assign n19924 = ~n19922 & ~n19923 ;
  assign n19925 = decrypt_pad & ~\u2_uk_K_r4_reg[23]/NET0131  ;
  assign n19926 = ~decrypt_pad & ~\u2_uk_K_r4_reg[15]/NET0131  ;
  assign n19927 = ~n19925 & ~n19926 ;
  assign n19928 = \u2_R4_reg[32]/NET0131  & ~n19927 ;
  assign n19929 = ~\u2_R4_reg[32]/NET0131  & n19927 ;
  assign n19930 = ~n19928 & ~n19929 ;
  assign n19969 = decrypt_pad & ~\u2_uk_K_r4_reg[45]/NET0131  ;
  assign n19970 = ~decrypt_pad & ~\u2_uk_K_r4_reg[9]/NET0131  ;
  assign n19971 = ~n19969 & ~n19970 ;
  assign n19972 = \u2_R4_reg[31]/P0001  & ~n19971 ;
  assign n19973 = ~\u2_R4_reg[31]/P0001  & n19971 ;
  assign n19974 = ~n19972 & ~n19973 ;
  assign n19944 = decrypt_pad & ~\u2_uk_K_r4_reg[1]/NET0131  ;
  assign n19945 = ~decrypt_pad & ~\u2_uk_K_r4_reg[52]/NET0131  ;
  assign n19946 = ~n19944 & ~n19945 ;
  assign n19947 = \u2_R4_reg[28]/NET0131  & ~n19946 ;
  assign n19948 = ~\u2_R4_reg[28]/NET0131  & n19946 ;
  assign n19949 = ~n19947 & ~n19948 ;
  assign n19931 = decrypt_pad & ~\u2_uk_K_r4_reg[28]/NET0131  ;
  assign n19932 = ~decrypt_pad & ~\u2_uk_K_r4_reg[51]/NET0131  ;
  assign n19933 = ~n19931 & ~n19932 ;
  assign n19934 = \u2_R4_reg[29]/NET0131  & ~n19933 ;
  assign n19935 = ~\u2_R4_reg[29]/NET0131  & n19933 ;
  assign n19936 = ~n19934 & ~n19935 ;
  assign n19937 = decrypt_pad & ~\u2_uk_K_r4_reg[44]/NET0131  ;
  assign n19938 = ~decrypt_pad & ~\u2_uk_K_r4_reg[36]/NET0131  ;
  assign n19939 = ~n19937 & ~n19938 ;
  assign n19940 = \u2_R4_reg[1]/NET0131  & ~n19939 ;
  assign n19941 = ~\u2_R4_reg[1]/NET0131  & n19939 ;
  assign n19942 = ~n19940 & ~n19941 ;
  assign n19977 = ~n19936 & n19942 ;
  assign n19978 = ~n19949 & n19977 ;
  assign n19950 = decrypt_pad & ~\u2_uk_K_r4_reg[29]/NET0131  ;
  assign n19951 = ~decrypt_pad & ~\u2_uk_K_r4_reg[21]/NET0131  ;
  assign n19952 = ~n19950 & ~n19951 ;
  assign n19953 = \u2_R4_reg[30]/NET0131  & ~n19952 ;
  assign n19954 = ~\u2_R4_reg[30]/NET0131  & n19952 ;
  assign n19955 = ~n19953 & ~n19954 ;
  assign n19998 = ~n19936 & ~n19942 ;
  assign n19999 = n19955 & n19998 ;
  assign n20000 = n19949 & n19999 ;
  assign n20001 = ~n19978 & ~n20000 ;
  assign n20002 = n19974 & ~n20001 ;
  assign n19943 = n19936 & n19942 ;
  assign n19984 = n19949 & ~n19955 ;
  assign n19956 = ~n19949 & n19955 ;
  assign n19992 = ~n19942 & n19956 ;
  assign n19993 = ~n19984 & ~n19992 ;
  assign n19994 = ~n19943 & n19993 ;
  assign n19995 = ~n19974 & ~n19994 ;
  assign n19965 = n19936 & n19949 ;
  assign n19966 = ~n19955 & n19965 ;
  assign n19967 = ~n19942 & n19966 ;
  assign n19996 = n19955 & n19965 ;
  assign n19997 = n19942 & n19996 ;
  assign n20003 = ~n19967 & ~n19997 ;
  assign n20004 = ~n19995 & n20003 ;
  assign n20005 = ~n20002 & n20004 ;
  assign n20006 = ~n19930 & ~n20005 ;
  assign n19980 = n19936 & ~n19955 ;
  assign n19981 = ~n19942 & n19949 ;
  assign n19982 = ~n19980 & ~n19981 ;
  assign n19983 = ~n19930 & ~n19982 ;
  assign n19985 = n19936 & ~n19942 ;
  assign n19986 = ~n19984 & ~n19985 ;
  assign n19987 = ~n19967 & ~n19986 ;
  assign n19988 = ~n19983 & n19987 ;
  assign n19961 = ~n19949 & ~n19955 ;
  assign n19962 = ~n19936 & n19961 ;
  assign n19976 = ~n19942 & n19962 ;
  assign n19979 = n19955 & n19978 ;
  assign n19989 = ~n19976 & ~n19979 ;
  assign n19990 = ~n19988 & n19989 ;
  assign n19991 = n19974 & ~n19990 ;
  assign n19957 = n19943 & n19956 ;
  assign n19958 = n19930 & n19957 ;
  assign n19959 = ~n19936 & n19949 ;
  assign n19960 = n19955 & n19959 ;
  assign n19963 = ~n19960 & ~n19962 ;
  assign n19964 = n19930 & ~n19963 ;
  assign n19968 = ~n19964 & ~n19967 ;
  assign n19975 = ~n19968 & ~n19974 ;
  assign n20007 = ~n19958 & ~n19975 ;
  assign n20008 = ~n19991 & n20007 ;
  assign n20009 = ~n20006 & n20008 ;
  assign n20010 = \u2_L4_reg[5]/NET0131  & ~n20009 ;
  assign n20011 = ~\u2_L4_reg[5]/NET0131  & n20009 ;
  assign n20012 = ~n20010 & ~n20011 ;
  assign n20029 = ~n19731 & ~n19736 ;
  assign n20030 = n19693 & ~n20029 ;
  assign n20025 = n19687 & n19754 ;
  assign n20026 = ~n19713 & ~n20025 ;
  assign n20031 = n19686 & n19757 ;
  assign n20032 = ~n19715 & ~n20031 ;
  assign n20016 = n19680 & n19757 ;
  assign n20033 = ~n19693 & ~n20016 ;
  assign n20034 = ~n20032 & n20033 ;
  assign n20035 = n20026 & ~n20034 ;
  assign n20036 = ~n20030 & n20035 ;
  assign n20037 = n19701 & ~n20036 ;
  assign n20013 = ~n19694 & ~n19723 ;
  assign n20014 = ~n19737 & ~n20013 ;
  assign n20017 = n19693 & ~n19709 ;
  assign n20018 = n19718 & n20017 ;
  assign n20015 = n19711 & n19720 ;
  assign n20019 = ~n20015 & ~n20016 ;
  assign n20020 = ~n19732 & n20019 ;
  assign n20021 = ~n20018 & n20020 ;
  assign n20022 = ~n20014 & n20021 ;
  assign n20023 = ~n19701 & ~n20022 ;
  assign n20027 = ~n19734 & n20026 ;
  assign n20028 = ~n19693 & ~n20027 ;
  assign n20024 = ~n19708 & n19717 ;
  assign n20038 = ~n19738 & ~n20024 ;
  assign n20039 = ~n20028 & n20038 ;
  assign n20040 = ~n20023 & n20039 ;
  assign n20041 = ~n20037 & n20040 ;
  assign n20042 = ~\u2_L4_reg[10]/NET0131  & ~n20041 ;
  assign n20043 = \u2_L4_reg[10]/NET0131  & n20041 ;
  assign n20044 = ~n20042 & ~n20043 ;
  assign n20054 = n19600 & n19622 ;
  assign n20052 = ~n19583 & ~n19614 ;
  assign n20053 = n19602 & ~n20052 ;
  assign n20055 = n19580 & n19589 ;
  assign n20056 = n19603 & n20055 ;
  assign n20057 = ~n20053 & ~n20056 ;
  assign n20058 = ~n20054 & n20057 ;
  assign n20045 = ~n19555 & ~n19581 ;
  assign n20046 = ~n19612 & ~n20045 ;
  assign n20047 = n19573 & n19580 ;
  assign n20048 = n19567 & n19589 ;
  assign n20049 = ~n19593 & ~n20048 ;
  assign n20050 = ~n20047 & n20049 ;
  assign n20051 = ~n19561 & ~n20050 ;
  assign n20059 = ~n20046 & ~n20051 ;
  assign n20060 = n20058 & n20059 ;
  assign n20063 = ~n19561 & ~n19604 ;
  assign n20064 = n19567 & n19580 ;
  assign n20065 = n19561 & ~n20064 ;
  assign n20066 = ~n19617 & n20065 ;
  assign n20067 = ~n20063 & ~n20066 ;
  assign n20061 = n19610 & n19622 ;
  assign n20062 = ~n20049 & n20061 ;
  assign n20068 = n19555 & ~n19601 ;
  assign n20069 = ~n19618 & n20068 ;
  assign n20070 = ~n20062 & n20069 ;
  assign n20071 = ~n20067 & n20070 ;
  assign n20072 = ~n20060 & ~n20071 ;
  assign n20073 = \u2_L4_reg[12]/NET0131  & n20072 ;
  assign n20074 = ~\u2_L4_reg[12]/NET0131  & ~n20072 ;
  assign n20075 = ~n20073 & ~n20074 ;
  assign n20076 = n19818 & n19845 ;
  assign n20077 = ~n19869 & ~n20076 ;
  assign n20078 = n19826 & n19833 ;
  assign n20079 = n19818 & ~n19825 ;
  assign n20080 = ~n19864 & ~n20079 ;
  assign n20081 = ~n20078 & n20080 ;
  assign n20082 = ~n19805 & ~n20081 ;
  assign n20083 = n20077 & ~n20082 ;
  assign n20084 = ~n19840 & ~n20083 ;
  assign n20088 = ~n19811 & ~n19849 ;
  assign n20089 = ~n19862 & ~n20088 ;
  assign n20090 = ~n19852 & n19862 ;
  assign n20091 = n19840 & ~n20090 ;
  assign n20092 = ~n20089 & n20091 ;
  assign n20086 = ~n19818 & n19840 ;
  assign n20087 = n19845 & n20086 ;
  assign n20085 = n19849 & ~n19854 ;
  assign n20093 = ~n19805 & ~n20085 ;
  assign n20094 = ~n20087 & n20093 ;
  assign n20095 = ~n20092 & n20094 ;
  assign n20102 = ~n19833 & n20079 ;
  assign n20103 = n19805 & ~n20102 ;
  assign n20104 = ~n19857 & n20103 ;
  assign n20100 = ~n19851 & n20088 ;
  assign n20101 = ~n19840 & n20100 ;
  assign n20096 = ~n19811 & n19851 ;
  assign n20097 = n19833 & n19849 ;
  assign n20098 = ~n20096 & ~n20097 ;
  assign n20099 = n19840 & ~n20098 ;
  assign n20105 = n20077 & ~n20099 ;
  assign n20106 = ~n20101 & n20105 ;
  assign n20107 = n20104 & n20106 ;
  assign n20108 = ~n20095 & ~n20107 ;
  assign n20109 = ~n20084 & ~n20108 ;
  assign n20110 = ~\u2_L4_reg[13]/NET0131  & n20109 ;
  assign n20111 = \u2_L4_reg[13]/NET0131  & ~n20109 ;
  assign n20112 = ~n20110 & ~n20111 ;
  assign n20114 = n19936 & ~n19993 ;
  assign n20115 = ~n19949 & n19998 ;
  assign n20116 = n19974 & n20115 ;
  assign n20113 = n19942 & n19960 ;
  assign n20117 = n19955 & ~n19974 ;
  assign n20118 = n19977 & n20117 ;
  assign n20119 = n19930 & ~n20118 ;
  assign n20120 = ~n20113 & n20119 ;
  assign n20121 = ~n20116 & n20120 ;
  assign n20122 = ~n20114 & n20121 ;
  assign n20124 = ~n19955 & n19985 ;
  assign n20125 = ~n19965 & ~n20124 ;
  assign n20126 = ~n19978 & n20125 ;
  assign n20127 = n19974 & ~n20126 ;
  assign n20123 = n19984 & n19998 ;
  assign n20128 = ~n19930 & ~n20123 ;
  assign n20129 = ~n20127 & n20128 ;
  assign n20130 = ~n20122 & ~n20129 ;
  assign n20132 = n19961 & ~n19977 ;
  assign n20133 = ~n19985 & n20132 ;
  assign n20134 = n19930 & ~n19955 ;
  assign n20135 = n19959 & ~n20134 ;
  assign n20131 = n19956 & n19985 ;
  assign n20136 = ~n19974 & ~n20131 ;
  assign n20137 = ~n20135 & n20136 ;
  assign n20138 = ~n20133 & n20137 ;
  assign n20139 = ~n19955 & n19977 ;
  assign n20140 = ~n19949 & n20139 ;
  assign n20141 = ~n19957 & n19974 ;
  assign n20142 = ~n20140 & n20141 ;
  assign n20143 = ~n20138 & ~n20142 ;
  assign n20144 = ~n20130 & ~n20143 ;
  assign n20145 = ~\u2_L4_reg[15]/NET0131  & ~n20144 ;
  assign n20146 = \u2_L4_reg[15]/NET0131  & n20144 ;
  assign n20147 = ~n20145 & ~n20146 ;
  assign n20209 = decrypt_pad & ~\u2_uk_K_r4_reg[8]/NET0131  ;
  assign n20210 = ~decrypt_pad & ~\u2_uk_K_r4_reg[0]/P0001  ;
  assign n20211 = ~n20209 & ~n20210 ;
  assign n20212 = \u2_R4_reg[20]/NET0131  & ~n20211 ;
  assign n20213 = ~\u2_R4_reg[20]/NET0131  & n20211 ;
  assign n20214 = ~n20212 & ~n20213 ;
  assign n20148 = decrypt_pad & ~\u2_uk_K_r4_reg[52]/NET0131  ;
  assign n20149 = ~decrypt_pad & ~\u2_uk_K_r4_reg[16]/NET0131  ;
  assign n20150 = ~n20148 & ~n20149 ;
  assign n20151 = \u2_R4_reg[19]/NET0131  & ~n20150 ;
  assign n20152 = ~\u2_R4_reg[19]/NET0131  & n20150 ;
  assign n20153 = ~n20151 & ~n20152 ;
  assign n20174 = decrypt_pad & ~\u2_uk_K_r4_reg[37]/NET0131  ;
  assign n20175 = ~decrypt_pad & ~\u2_uk_K_r4_reg[29]/NET0131  ;
  assign n20176 = ~n20174 & ~n20175 ;
  assign n20177 = \u2_R4_reg[18]/NET0131  & ~n20176 ;
  assign n20178 = ~\u2_R4_reg[18]/NET0131  & n20176 ;
  assign n20179 = ~n20177 & ~n20178 ;
  assign n20154 = decrypt_pad & ~\u2_uk_K_r4_reg[9]/NET0131  ;
  assign n20155 = ~decrypt_pad & ~\u2_uk_K_r4_reg[1]/NET0131  ;
  assign n20156 = ~n20154 & ~n20155 ;
  assign n20157 = \u2_R4_reg[21]/NET0131  & ~n20156 ;
  assign n20158 = ~\u2_R4_reg[21]/NET0131  & n20156 ;
  assign n20159 = ~n20157 & ~n20158 ;
  assign n20160 = decrypt_pad & ~\u2_uk_K_r4_reg[21]/NET0131  ;
  assign n20161 = ~decrypt_pad & ~\u2_uk_K_r4_reg[44]/NET0131  ;
  assign n20162 = ~n20160 & ~n20161 ;
  assign n20163 = \u2_R4_reg[16]/NET0131  & ~n20162 ;
  assign n20164 = ~\u2_R4_reg[16]/NET0131  & n20162 ;
  assign n20165 = ~n20163 & ~n20164 ;
  assign n20166 = ~n20159 & n20165 ;
  assign n20167 = decrypt_pad & ~\u2_uk_K_r4_reg[43]/NET0131  ;
  assign n20168 = ~decrypt_pad & ~\u2_uk_K_r4_reg[35]/NET0131  ;
  assign n20169 = ~n20167 & ~n20168 ;
  assign n20170 = \u2_R4_reg[17]/NET0131  & ~n20169 ;
  assign n20171 = ~\u2_R4_reg[17]/NET0131  & n20169 ;
  assign n20172 = ~n20170 & ~n20171 ;
  assign n20194 = n20166 & ~n20172 ;
  assign n20226 = ~n20179 & n20194 ;
  assign n20181 = n20172 & ~n20179 ;
  assign n20200 = n20159 & n20165 ;
  assign n20229 = n20181 & n20200 ;
  assign n20188 = ~n20165 & ~n20172 ;
  assign n20225 = n20159 & n20188 ;
  assign n20227 = ~n20159 & n20172 ;
  assign n20228 = n20179 & n20227 ;
  assign n20230 = ~n20225 & ~n20228 ;
  assign n20231 = ~n20229 & n20230 ;
  assign n20232 = ~n20226 & n20231 ;
  assign n20233 = ~n20153 & ~n20232 ;
  assign n20197 = n20159 & ~n20179 ;
  assign n20216 = ~n20166 & ~n20197 ;
  assign n20196 = n20165 & ~n20172 ;
  assign n20217 = ~n20181 & ~n20196 ;
  assign n20218 = n20216 & ~n20217 ;
  assign n20219 = ~n20165 & n20172 ;
  assign n20190 = n20159 & ~n20165 ;
  assign n20220 = ~n20190 & n20216 ;
  assign n20221 = ~n20219 & ~n20220 ;
  assign n20222 = n20179 & n20219 ;
  assign n20223 = n20153 & ~n20222 ;
  assign n20224 = ~n20221 & n20223 ;
  assign n20234 = ~n20218 & ~n20224 ;
  assign n20235 = ~n20233 & n20234 ;
  assign n20236 = ~n20214 & ~n20235 ;
  assign n20173 = n20166 & n20172 ;
  assign n20182 = ~n20165 & n20181 ;
  assign n20180 = n20165 & n20179 ;
  assign n20183 = n20159 & ~n20180 ;
  assign n20184 = ~n20182 & n20183 ;
  assign n20185 = ~n20173 & ~n20184 ;
  assign n20186 = n20153 & ~n20185 ;
  assign n20187 = ~n20153 & ~n20179 ;
  assign n20189 = ~n20159 & n20188 ;
  assign n20191 = n20172 & n20190 ;
  assign n20192 = ~n20189 & ~n20191 ;
  assign n20193 = n20187 & ~n20192 ;
  assign n20195 = n20179 & n20194 ;
  assign n20198 = n20196 & n20197 ;
  assign n20204 = ~n20195 & ~n20198 ;
  assign n20199 = ~n20153 & n20179 ;
  assign n20201 = n20172 & n20200 ;
  assign n20202 = n20199 & n20201 ;
  assign n20203 = n20173 & ~n20179 ;
  assign n20205 = ~n20202 & ~n20203 ;
  assign n20206 = n20204 & n20205 ;
  assign n20207 = ~n20193 & n20206 ;
  assign n20208 = ~n20186 & n20207 ;
  assign n20215 = ~n20208 & n20214 ;
  assign n20237 = ~n20172 & n20179 ;
  assign n20238 = n20190 & n20237 ;
  assign n20239 = ~n20228 & ~n20238 ;
  assign n20240 = ~n20165 & ~n20239 ;
  assign n20241 = ~n20153 & n20240 ;
  assign n20242 = n20179 & n20189 ;
  assign n20243 = ~n20203 & ~n20242 ;
  assign n20244 = n20153 & ~n20243 ;
  assign n20245 = ~n20241 & ~n20244 ;
  assign n20246 = ~n20215 & n20245 ;
  assign n20247 = ~n20236 & n20246 ;
  assign n20248 = ~\u2_L4_reg[14]/NET0131  & ~n20247 ;
  assign n20249 = \u2_L4_reg[14]/NET0131  & n20247 ;
  assign n20250 = ~n20248 & ~n20249 ;
  assign n20251 = ~n19460 & n19466 ;
  assign n20252 = ~n19893 & ~n20251 ;
  assign n20253 = ~n19485 & ~n20252 ;
  assign n20257 = n19511 & ~n19902 ;
  assign n20258 = ~n20253 & n20257 ;
  assign n20254 = n19479 & ~n19915 ;
  assign n20255 = ~n19524 & ~n19531 ;
  assign n20256 = n19460 & ~n20255 ;
  assign n20259 = ~n20254 & ~n20256 ;
  assign n20260 = n20258 & n20259 ;
  assign n20263 = n19466 & ~n19515 ;
  assign n20264 = ~n19890 & ~n20263 ;
  assign n20265 = n19460 & ~n20264 ;
  assign n20262 = ~n19460 & ~n19915 ;
  assign n20261 = n19479 & n19491 ;
  assign n20266 = ~n19511 & ~n20261 ;
  assign n20267 = ~n20262 & n20266 ;
  assign n20268 = ~n20265 & n20267 ;
  assign n20269 = ~n20260 & ~n20268 ;
  assign n20270 = ~n19485 & n19897 ;
  assign n20271 = ~n19527 & ~n20270 ;
  assign n20272 = ~n20269 & n20271 ;
  assign n20273 = ~\u2_L4_reg[19]/NET0131  & ~n20272 ;
  assign n20274 = \u2_L4_reg[19]/NET0131  & n20272 ;
  assign n20275 = ~n20273 & ~n20274 ;
  assign n20297 = ~n19735 & ~n19743 ;
  assign n20298 = n19701 & ~n20297 ;
  assign n20299 = ~n19732 & n20026 ;
  assign n20300 = ~n20298 & n20299 ;
  assign n20301 = n19693 & ~n20300 ;
  assign n20287 = ~n19686 & ~n19708 ;
  assign n20288 = ~n19743 & ~n20287 ;
  assign n20289 = n19680 & ~n20288 ;
  assign n20290 = ~n19693 & ~n20289 ;
  assign n20291 = ~n19680 & n20287 ;
  assign n20292 = n19756 & ~n20291 ;
  assign n20293 = ~n20290 & ~n20292 ;
  assign n20294 = n19714 & ~n19758 ;
  assign n20295 = ~n20293 & n20294 ;
  assign n20296 = ~n19701 & ~n20295 ;
  assign n20277 = ~n19715 & n19757 ;
  assign n20278 = n19674 & n19687 ;
  assign n20279 = ~n20277 & ~n20278 ;
  assign n20280 = ~n19693 & ~n20279 ;
  assign n20276 = ~n19680 & n19754 ;
  assign n20281 = n19708 & n19716 ;
  assign n20282 = ~n20276 & ~n20281 ;
  assign n20283 = ~n20280 & n20282 ;
  assign n20284 = n19701 & ~n20283 ;
  assign n20285 = ~n19724 & ~n20281 ;
  assign n20286 = ~n19693 & ~n20285 ;
  assign n20302 = ~n20284 & ~n20286 ;
  assign n20303 = ~n20296 & n20302 ;
  assign n20304 = ~n20301 & n20303 ;
  assign n20305 = ~\u2_L4_reg[1]/NET0131  & ~n20304 ;
  assign n20306 = \u2_L4_reg[1]/NET0131  & n20304 ;
  assign n20307 = ~n20305 & ~n20306 ;
  assign n20311 = ~n19942 & n19984 ;
  assign n20312 = ~n19974 & ~n20311 ;
  assign n20313 = ~n20113 & n20312 ;
  assign n20315 = n19974 & ~n19996 ;
  assign n20314 = n19943 & ~n19949 ;
  assign n20316 = ~n20139 & ~n20314 ;
  assign n20317 = n20315 & n20316 ;
  assign n20318 = ~n20313 & ~n20317 ;
  assign n20319 = ~n19942 & n19965 ;
  assign n20320 = ~n20115 & ~n20319 ;
  assign n20321 = n19955 & ~n20320 ;
  assign n20322 = n19930 & ~n20140 ;
  assign n20323 = ~n20321 & n20322 ;
  assign n20324 = ~n20318 & n20323 ;
  assign n20309 = n19942 & ~n19974 ;
  assign n20329 = ~n19943 & ~n20309 ;
  assign n20330 = n19984 & ~n20329 ;
  assign n20325 = ~n19936 & ~n20309 ;
  assign n20326 = n19956 & ~n20325 ;
  assign n20335 = ~n20000 & ~n20326 ;
  assign n20336 = ~n20330 & n20335 ;
  assign n20327 = ~n19960 & ~n20319 ;
  assign n20328 = n19974 & ~n20327 ;
  assign n20331 = ~n19949 & ~n19974 ;
  assign n20332 = n19985 & n20331 ;
  assign n20333 = ~n19930 & ~n20332 ;
  assign n20334 = ~n19976 & n20333 ;
  assign n20337 = ~n20328 & n20334 ;
  assign n20338 = n20336 & n20337 ;
  assign n20339 = ~n20324 & ~n20338 ;
  assign n20308 = n19962 & n19974 ;
  assign n20310 = n19966 & n20309 ;
  assign n20340 = ~n20308 & ~n20310 ;
  assign n20341 = ~n20339 & n20340 ;
  assign n20342 = ~\u2_L4_reg[21]/NET0131  & ~n20341 ;
  assign n20343 = \u2_L4_reg[21]/NET0131  & n20341 ;
  assign n20344 = ~n20342 & ~n20343 ;
  assign n20357 = n19403 & ~n19651 ;
  assign n20358 = ~n19418 & n20357 ;
  assign n20354 = n19370 & n19376 ;
  assign n20355 = ~n19389 & n20354 ;
  assign n20356 = n19364 & n20355 ;
  assign n20359 = ~n19442 & ~n20356 ;
  assign n20360 = n20358 & n20359 ;
  assign n20361 = ~n19417 & ~n19659 ;
  assign n20362 = n19370 & ~n20361 ;
  assign n20345 = n19376 & n19421 ;
  assign n20363 = n19364 & n20345 ;
  assign n20364 = ~n19403 & ~n19420 ;
  assign n20365 = ~n19428 & ~n19658 ;
  assign n20366 = n20364 & n20365 ;
  assign n20367 = ~n20363 & n20366 ;
  assign n20368 = ~n20362 & n20367 ;
  assign n20369 = ~n20360 & ~n20368 ;
  assign n20346 = n19377 & ~n19389 ;
  assign n20347 = ~n20345 & ~n20346 ;
  assign n20348 = ~n19394 & n20347 ;
  assign n20349 = n19403 & ~n20348 ;
  assign n20350 = n19377 & n19395 ;
  assign n20351 = ~n19655 & ~n20350 ;
  assign n20352 = ~n20349 & n20351 ;
  assign n20353 = ~n19364 & ~n20352 ;
  assign n20370 = ~n19364 & n19409 ;
  assign n20371 = n19425 & n20345 ;
  assign n20372 = ~n19416 & ~n20371 ;
  assign n20373 = ~n20370 & n20372 ;
  assign n20374 = ~n20353 & n20373 ;
  assign n20375 = ~n20369 & n20374 ;
  assign n20376 = \u2_L4_reg[23]/NET0131  & ~n20375 ;
  assign n20377 = ~\u2_L4_reg[23]/NET0131  & n20375 ;
  assign n20378 = ~n20376 & ~n20377 ;
  assign n20383 = n19733 & n19743 ;
  assign n20384 = ~n19693 & ~n19712 ;
  assign n20385 = ~n20383 & n20384 ;
  assign n20386 = ~n19740 & ~n20385 ;
  assign n20379 = ~n19708 & n19731 ;
  assign n20380 = ~n19694 & ~n19716 ;
  assign n20381 = ~n20278 & n20380 ;
  assign n20382 = n19708 & ~n20381 ;
  assign n20387 = ~n20379 & ~n20382 ;
  assign n20388 = ~n20386 & n20387 ;
  assign n20389 = n19701 & ~n20388 ;
  assign n20390 = ~n19686 & ~n19719 ;
  assign n20391 = ~n19739 & ~n20390 ;
  assign n20392 = ~n19693 & ~n20391 ;
  assign n20393 = ~n19718 & ~n20278 ;
  assign n20394 = n19686 & n19693 ;
  assign n20395 = n19701 & ~n20394 ;
  assign n20396 = ~n20393 & ~n20395 ;
  assign n20397 = ~n20392 & ~n20396 ;
  assign n20398 = ~n19708 & ~n20397 ;
  assign n20399 = ~n19722 & ~n20276 ;
  assign n20400 = ~n19693 & ~n20399 ;
  assign n20401 = n19674 & ~n19687 ;
  assign n20402 = n19737 & n20401 ;
  assign n20403 = ~n19717 & ~n20402 ;
  assign n20404 = ~n20400 & n20403 ;
  assign n20405 = ~n19701 & ~n20404 ;
  assign n20406 = ~n20398 & ~n20405 ;
  assign n20407 = ~n20389 & n20406 ;
  assign n20408 = ~\u2_L4_reg[26]/NET0131  & ~n20407 ;
  assign n20409 = \u2_L4_reg[26]/NET0131  & n20407 ;
  assign n20410 = ~n20408 & ~n20409 ;
  assign n20411 = ~n20172 & n20200 ;
  assign n20412 = ~n20153 & ~n20411 ;
  assign n20413 = ~n20182 & n20412 ;
  assign n20414 = ~n20159 & ~n20180 ;
  assign n20415 = ~n20181 & n20414 ;
  assign n20416 = n20153 & ~n20188 ;
  assign n20417 = ~n20201 & n20416 ;
  assign n20418 = ~n20415 & n20417 ;
  assign n20419 = ~n20413 & ~n20418 ;
  assign n20420 = n20165 & n20228 ;
  assign n20421 = n20172 & n20197 ;
  assign n20422 = n20214 & ~n20421 ;
  assign n20423 = ~n20420 & n20422 ;
  assign n20424 = ~n20419 & n20423 ;
  assign n20429 = n20153 & ~n20227 ;
  assign n20428 = ~n20153 & ~n20188 ;
  assign n20430 = ~n20179 & ~n20428 ;
  assign n20431 = ~n20429 & n20430 ;
  assign n20425 = n20153 & ~n20159 ;
  assign n20426 = ~n20194 & ~n20222 ;
  assign n20427 = ~n20425 & ~n20426 ;
  assign n20432 = ~n20214 & ~n20427 ;
  assign n20433 = ~n20431 & n20432 ;
  assign n20434 = ~n20424 & ~n20433 ;
  assign n20435 = ~n20242 & ~n20420 ;
  assign n20436 = n20188 & n20197 ;
  assign n20437 = n20435 & ~n20436 ;
  assign n20438 = n20153 & ~n20437 ;
  assign n20439 = n20196 & n20199 ;
  assign n20440 = ~n20229 & ~n20439 ;
  assign n20441 = ~n20438 & n20440 ;
  assign n20442 = ~n20434 & n20441 ;
  assign n20443 = ~\u2_L4_reg[25]/NET0131  & ~n20442 ;
  assign n20444 = \u2_L4_reg[25]/NET0131  & n20442 ;
  assign n20445 = ~n20443 & ~n20444 ;
  assign n20448 = n19811 & n19849 ;
  assign n20449 = ~n19833 & n19874 ;
  assign n20450 = ~n20448 & ~n20449 ;
  assign n20451 = n19840 & n20450 ;
  assign n20455 = n19825 & ~n20100 ;
  assign n20452 = ~n19825 & n19841 ;
  assign n20453 = ~n19840 & ~n20076 ;
  assign n20454 = ~n20452 & n20453 ;
  assign n20456 = ~n19826 & n20454 ;
  assign n20457 = ~n20455 & n20456 ;
  assign n20458 = ~n20451 & ~n20457 ;
  assign n20446 = n19833 & ~n19863 ;
  assign n20447 = ~n20089 & n20446 ;
  assign n20459 = ~n19805 & ~n20447 ;
  assign n20460 = ~n20458 & n20459 ;
  assign n20464 = n20450 & n20454 ;
  assign n20465 = ~n19817 & ~n19865 ;
  assign n20466 = n19850 & ~n20465 ;
  assign n20467 = n19840 & ~n19863 ;
  assign n20468 = ~n20466 & n20467 ;
  assign n20469 = ~n20464 & ~n20468 ;
  assign n20461 = ~n19819 & ~n19840 ;
  assign n20462 = n19825 & ~n19833 ;
  assign n20463 = ~n20461 & n20462 ;
  assign n20470 = n19805 & ~n20078 ;
  assign n20471 = ~n20463 & n20470 ;
  assign n20472 = ~n20469 & n20471 ;
  assign n20473 = ~n20460 & ~n20472 ;
  assign n20474 = ~\u2_L4_reg[28]/NET0131  & n20473 ;
  assign n20475 = \u2_L4_reg[28]/NET0131  & ~n20473 ;
  assign n20476 = ~n20474 & ~n20475 ;
  assign n20477 = n20153 & ~n20226 ;
  assign n20478 = ~n20201 & n20477 ;
  assign n20479 = n20190 & ~n20237 ;
  assign n20480 = n20412 & ~n20479 ;
  assign n20481 = ~n20478 & ~n20480 ;
  assign n20482 = ~n20182 & n20435 ;
  assign n20483 = ~n20481 & n20482 ;
  assign n20484 = ~n20214 & ~n20483 ;
  assign n20485 = ~n20179 & n20189 ;
  assign n20486 = ~n20411 & ~n20485 ;
  assign n20487 = n20153 & ~n20486 ;
  assign n20488 = n20165 & n20187 ;
  assign n20489 = ~n20240 & ~n20488 ;
  assign n20490 = ~n20487 & n20489 ;
  assign n20491 = n20214 & ~n20490 ;
  assign n20492 = n20159 & n20182 ;
  assign n20493 = n20239 & ~n20492 ;
  assign n20494 = n20153 & ~n20493 ;
  assign n20495 = ~n20153 & n20195 ;
  assign n20496 = ~n20494 & ~n20495 ;
  assign n20497 = ~n20491 & n20496 ;
  assign n20498 = ~n20484 & n20497 ;
  assign n20499 = ~\u2_L4_reg[8]/NET0131  & ~n20498 ;
  assign n20500 = \u2_L4_reg[8]/NET0131  & n20498 ;
  assign n20501 = ~n20499 & ~n20500 ;
  assign n20502 = ~n19962 & ~n20314 ;
  assign n20503 = ~n20319 & n20502 ;
  assign n20504 = ~n19974 & ~n20503 ;
  assign n20505 = n19974 & ~n19981 ;
  assign n20506 = ~n20125 & n20505 ;
  assign n20507 = ~n19957 & ~n20139 ;
  assign n20508 = ~n20000 & n20507 ;
  assign n20509 = ~n20506 & n20508 ;
  assign n20510 = ~n20504 & n20509 ;
  assign n20511 = n19930 & ~n20510 ;
  assign n20518 = n19982 & ~n19998 ;
  assign n20519 = n19974 & ~n20124 ;
  assign n20520 = ~n20518 & n20519 ;
  assign n20516 = n19942 & n19949 ;
  assign n20517 = n20117 & n20516 ;
  assign n20521 = ~n20332 & ~n20517 ;
  assign n20522 = ~n19979 & n20521 ;
  assign n20523 = ~n20520 & n20522 ;
  assign n20524 = ~n19930 & ~n20523 ;
  assign n20512 = n19974 & n19999 ;
  assign n20513 = n19982 & ~n19986 ;
  assign n20514 = ~n19967 & ~n20513 ;
  assign n20515 = ~n19974 & ~n20514 ;
  assign n20525 = ~n20512 & ~n20515 ;
  assign n20526 = ~n20524 & n20525 ;
  assign n20527 = ~n20511 & n20526 ;
  assign n20528 = ~\u2_L4_reg[27]/NET0131  & ~n20527 ;
  assign n20529 = \u2_L4_reg[27]/NET0131  & n20527 ;
  assign n20530 = ~n20528 & ~n20529 ;
  assign n20541 = ~n19600 & ~n20055 ;
  assign n20543 = ~n19574 & n20049 ;
  assign n20544 = ~n20541 & ~n20543 ;
  assign n20542 = ~n19574 & n20541 ;
  assign n20545 = ~n19561 & ~n20542 ;
  assign n20546 = ~n20544 & n20545 ;
  assign n20533 = ~n19573 & n20048 ;
  assign n20534 = ~n19580 & n19593 ;
  assign n20535 = ~n20533 & ~n20534 ;
  assign n20536 = n19561 & ~n20535 ;
  assign n20538 = ~n19561 & ~n19567 ;
  assign n20537 = n19573 & ~n19589 ;
  assign n20539 = n19580 & n20537 ;
  assign n20540 = ~n20538 & n20539 ;
  assign n20547 = ~n20536 & ~n20540 ;
  assign n20548 = ~n20546 & n20547 ;
  assign n20549 = n19555 & ~n20548 ;
  assign n20550 = n20045 & ~n20049 ;
  assign n20551 = n19580 & ~n20048 ;
  assign n20552 = ~n19603 & ~n19610 ;
  assign n20553 = ~n20551 & n20552 ;
  assign n20554 = ~n20550 & ~n20553 ;
  assign n20555 = ~n19561 & ~n20554 ;
  assign n20531 = n19555 & ~n19561 ;
  assign n20532 = n19604 & ~n20531 ;
  assign n20556 = n19583 & ~n20541 ;
  assign n20557 = ~n20537 & ~n20538 ;
  assign n20558 = n20551 & n20557 ;
  assign n20559 = ~n20556 & ~n20558 ;
  assign n20560 = ~n19555 & ~n20559 ;
  assign n20561 = ~n20532 & ~n20560 ;
  assign n20562 = ~n20555 & n20561 ;
  assign n20563 = ~n20549 & n20562 ;
  assign n20564 = \u2_L4_reg[32]/NET0131  & n20563 ;
  assign n20565 = ~\u2_L4_reg[32]/NET0131  & ~n20563 ;
  assign n20566 = ~n20564 & ~n20565 ;
  assign n20571 = n20214 & ~n20229 ;
  assign n20572 = ~n20195 & n20571 ;
  assign n20567 = ~n20153 & n20191 ;
  assign n20568 = ~n20197 & ~n20219 ;
  assign n20569 = n20153 & ~n20190 ;
  assign n20570 = ~n20568 & n20569 ;
  assign n20573 = ~n20567 & ~n20570 ;
  assign n20574 = n20572 & n20573 ;
  assign n20578 = ~n20165 & n20197 ;
  assign n20579 = ~n20173 & ~n20578 ;
  assign n20580 = n20153 & ~n20579 ;
  assign n20575 = n20153 & ~n20237 ;
  assign n20576 = ~n20198 & ~n20216 ;
  assign n20577 = ~n20575 & ~n20576 ;
  assign n20581 = ~n20214 & ~n20577 ;
  assign n20582 = ~n20580 & n20581 ;
  assign n20583 = ~n20574 & ~n20582 ;
  assign n20584 = ~n20238 & n20477 ;
  assign n20585 = ~n20187 & ~n20412 ;
  assign n20586 = ~n20203 & ~n20485 ;
  assign n20587 = ~n20585 & n20586 ;
  assign n20588 = ~n20584 & ~n20587 ;
  assign n20589 = ~n20583 & ~n20588 ;
  assign n20590 = ~\u2_L4_reg[3]/NET0131  & ~n20589 ;
  assign n20591 = \u2_L4_reg[3]/NET0131  & n20589 ;
  assign n20592 = ~n20590 & ~n20591 ;
  assign n20619 = decrypt_pad & ~\u2_uk_K_r4_reg[46]/NET0131  ;
  assign n20620 = ~decrypt_pad & ~\u2_uk_K_r4_reg[40]/NET0131  ;
  assign n20621 = ~n20619 & ~n20620 ;
  assign n20622 = \u2_R4_reg[11]/NET0131  & ~n20621 ;
  assign n20623 = ~\u2_R4_reg[11]/NET0131  & n20621 ;
  assign n20624 = ~n20622 & ~n20623 ;
  assign n20593 = decrypt_pad & ~\u2_uk_K_r4_reg[4]/NET0131  ;
  assign n20594 = ~decrypt_pad & ~\u2_uk_K_r4_reg[55]/NET0131  ;
  assign n20595 = ~n20593 & ~n20594 ;
  assign n20596 = \u2_R4_reg[12]/NET0131  & ~n20595 ;
  assign n20597 = ~\u2_R4_reg[12]/NET0131  & n20595 ;
  assign n20598 = ~n20596 & ~n20597 ;
  assign n20599 = decrypt_pad & ~\u2_uk_K_r4_reg[17]/NET0131  ;
  assign n20600 = ~decrypt_pad & ~\u2_uk_K_r4_reg[11]/NET0131  ;
  assign n20601 = ~n20599 & ~n20600 ;
  assign n20602 = \u2_R4_reg[13]/NET0131  & ~n20601 ;
  assign n20603 = ~\u2_R4_reg[13]/NET0131  & n20601 ;
  assign n20604 = ~n20602 & ~n20603 ;
  assign n20612 = decrypt_pad & ~\u2_uk_K_r4_reg[12]/NET0131  ;
  assign n20613 = ~decrypt_pad & ~\u2_uk_K_r4_reg[6]/NET0131  ;
  assign n20614 = ~n20612 & ~n20613 ;
  assign n20615 = \u2_R4_reg[9]/NET0131  & ~n20614 ;
  assign n20616 = ~\u2_R4_reg[9]/NET0131  & n20614 ;
  assign n20617 = ~n20615 & ~n20616 ;
  assign n20655 = n20604 & ~n20617 ;
  assign n20605 = decrypt_pad & ~\u2_uk_K_r4_reg[40]/NET0131  ;
  assign n20606 = ~decrypt_pad & ~\u2_uk_K_r4_reg[34]/NET0131  ;
  assign n20607 = ~n20605 & ~n20606 ;
  assign n20608 = \u2_R4_reg[8]/NET0131  & ~n20607 ;
  assign n20609 = ~\u2_R4_reg[8]/NET0131  & n20607 ;
  assign n20610 = ~n20608 & ~n20609 ;
  assign n20611 = n20604 & ~n20610 ;
  assign n20625 = decrypt_pad & ~\u2_uk_K_r4_reg[20]/NET0131  ;
  assign n20626 = ~decrypt_pad & ~\u2_uk_K_r4_reg[39]/NET0131  ;
  assign n20627 = ~n20625 & ~n20626 ;
  assign n20628 = \u2_R4_reg[10]/NET0131  & ~n20627 ;
  assign n20629 = ~\u2_R4_reg[10]/NET0131  & n20627 ;
  assign n20630 = ~n20628 & ~n20629 ;
  assign n20663 = n20611 & n20630 ;
  assign n20664 = ~n20604 & n20610 ;
  assign n20665 = n20617 & n20664 ;
  assign n20666 = ~n20663 & ~n20665 ;
  assign n20667 = ~n20655 & n20666 ;
  assign n20668 = n20598 & ~n20667 ;
  assign n20635 = ~n20604 & ~n20610 ;
  assign n20661 = ~n20630 & n20635 ;
  assign n20662 = ~n20617 & n20661 ;
  assign n20642 = ~n20617 & n20630 ;
  assign n20669 = n20604 & n20642 ;
  assign n20670 = ~n20662 & ~n20669 ;
  assign n20671 = ~n20668 & n20670 ;
  assign n20672 = n20624 & ~n20671 ;
  assign n20636 = n20604 & n20610 ;
  assign n20637 = ~n20635 & ~n20636 ;
  assign n20643 = ~n20637 & n20642 ;
  assign n20618 = n20611 & n20617 ;
  assign n20631 = ~n20624 & n20630 ;
  assign n20632 = n20618 & n20631 ;
  assign n20644 = n20610 & n20630 ;
  assign n20645 = ~n20604 & n20617 ;
  assign n20646 = n20644 & n20645 ;
  assign n20647 = ~n20632 & ~n20646 ;
  assign n20648 = ~n20643 & n20647 ;
  assign n20633 = ~n20617 & ~n20630 ;
  assign n20634 = n20604 & n20624 ;
  assign n20638 = ~n20634 & n20637 ;
  assign n20639 = n20633 & n20638 ;
  assign n20640 = n20617 & ~n20630 ;
  assign n20641 = ~n20638 & n20640 ;
  assign n20649 = ~n20639 & ~n20641 ;
  assign n20650 = n20648 & n20649 ;
  assign n20651 = ~n20598 & ~n20650 ;
  assign n20652 = n20598 & n20630 ;
  assign n20653 = n20617 & n20635 ;
  assign n20654 = n20652 & n20653 ;
  assign n20656 = ~n20610 & ~n20640 ;
  assign n20657 = n20598 & ~n20624 ;
  assign n20658 = ~n20645 & ~n20655 ;
  assign n20659 = n20657 & n20658 ;
  assign n20660 = ~n20656 & n20659 ;
  assign n20673 = ~n20654 & ~n20660 ;
  assign n20674 = ~n20651 & n20673 ;
  assign n20675 = ~n20672 & n20674 ;
  assign n20676 = ~\u2_L4_reg[6]/NET0131  & ~n20675 ;
  assign n20677 = \u2_L4_reg[6]/NET0131  & n20675 ;
  assign n20678 = ~n20676 & ~n20677 ;
  assign n20680 = ~n19583 & n20541 ;
  assign n20681 = ~n19573 & ~n19593 ;
  assign n20682 = ~n20541 & ~n20681 ;
  assign n20683 = ~n20680 & ~n20682 ;
  assign n20679 = ~n19555 & n19561 ;
  assign n20684 = ~n20531 & ~n20679 ;
  assign n20685 = ~n20056 & n20684 ;
  assign n20686 = ~n20683 & n20685 ;
  assign n20687 = n19573 & ~n19602 ;
  assign n20688 = ~n20551 & n20687 ;
  assign n20689 = n20679 & ~n20680 ;
  assign n20690 = ~n20688 & n20689 ;
  assign n20691 = ~n20686 & ~n20690 ;
  assign n20692 = ~n19595 & ~n20691 ;
  assign n20694 = ~n19567 & ~n20047 ;
  assign n20695 = n20541 & ~n20694 ;
  assign n20693 = ~n19580 & ~n19622 ;
  assign n20696 = ~n20056 & n20531 ;
  assign n20697 = ~n20693 & n20696 ;
  assign n20698 = ~n20695 & n20697 ;
  assign n20699 = ~n20692 & ~n20698 ;
  assign n20700 = ~\u2_L4_reg[7]/NET0131  & n20699 ;
  assign n20701 = \u2_L4_reg[7]/NET0131  & ~n20699 ;
  assign n20702 = ~n20700 & ~n20701 ;
  assign n20717 = n19636 & n20347 ;
  assign n20718 = n19383 & ~n20717 ;
  assign n20708 = ~n19392 & ~n20355 ;
  assign n20719 = n19425 & ~n20708 ;
  assign n20720 = ~n19655 & ~n20719 ;
  assign n20721 = ~n20718 & n20720 ;
  assign n20722 = n19403 & ~n20721 ;
  assign n20703 = ~n19383 & n19408 ;
  assign n20704 = n19383 & n20355 ;
  assign n20705 = ~n20703 & ~n20704 ;
  assign n20706 = ~n19364 & ~n20705 ;
  assign n20709 = ~n19364 & n20708 ;
  assign n20710 = n19364 & ~n19377 ;
  assign n20711 = ~n19441 & n20710 ;
  assign n20712 = ~n20345 & n20711 ;
  assign n20713 = ~n20709 & ~n20712 ;
  assign n20707 = n19383 & n19643 ;
  assign n20714 = ~n20703 & ~n20707 ;
  assign n20715 = ~n20713 & n20714 ;
  assign n20716 = ~n19403 & ~n20715 ;
  assign n20723 = ~n20706 & ~n20716 ;
  assign n20724 = ~n20722 & n20723 ;
  assign n20725 = ~\u2_L4_reg[9]/NET0131  & ~n20724 ;
  assign n20726 = \u2_L4_reg[9]/NET0131  & n20724 ;
  assign n20727 = ~n20725 & ~n20726 ;
  assign n20732 = ~n20617 & ~n20636 ;
  assign n20731 = n20617 & n20636 ;
  assign n20733 = ~n20635 & ~n20731 ;
  assign n20734 = ~n20732 & n20733 ;
  assign n20729 = n20617 & n20624 ;
  assign n20730 = n20635 & ~n20729 ;
  assign n20735 = ~n20630 & ~n20730 ;
  assign n20736 = ~n20734 & n20735 ;
  assign n20737 = n20630 & n20635 ;
  assign n20738 = ~n20630 & n20664 ;
  assign n20739 = ~n20737 & ~n20738 ;
  assign n20740 = ~n20624 & ~n20739 ;
  assign n20728 = n20618 & n20630 ;
  assign n20741 = n20598 & ~n20728 ;
  assign n20742 = ~n20740 & n20741 ;
  assign n20743 = ~n20736 & n20742 ;
  assign n20745 = ~n20610 & n20655 ;
  assign n20746 = ~n20661 & ~n20731 ;
  assign n20747 = ~n20745 & n20746 ;
  assign n20748 = ~n20624 & ~n20747 ;
  assign n20744 = n20624 & n20734 ;
  assign n20749 = ~n20598 & ~n20662 ;
  assign n20750 = ~n20744 & n20749 ;
  assign n20751 = ~n20748 & n20750 ;
  assign n20752 = ~n20743 & ~n20751 ;
  assign n20753 = ~n20617 & n20644 ;
  assign n20754 = ~n20624 & n20753 ;
  assign n20755 = ~n20617 & n20737 ;
  assign n20756 = ~n20646 & ~n20755 ;
  assign n20757 = n20624 & ~n20756 ;
  assign n20758 = ~n20754 & ~n20757 ;
  assign n20759 = ~n20752 & n20758 ;
  assign n20760 = ~\u2_L4_reg[16]/NET0131  & ~n20759 ;
  assign n20761 = \u2_L4_reg[16]/NET0131  & n20759 ;
  assign n20762 = ~n20760 & ~n20761 ;
  assign n20766 = ~n19863 & ~n19868 ;
  assign n20767 = ~n19840 & ~n20766 ;
  assign n20764 = n19841 & n19874 ;
  assign n20765 = ~n19827 & n19840 ;
  assign n20768 = ~n20764 & ~n20765 ;
  assign n20769 = ~n20767 & n20768 ;
  assign n20770 = n19805 & ~n20769 ;
  assign n20772 = ~n19852 & ~n19866 ;
  assign n20773 = n19873 & n20772 ;
  assign n20774 = ~n19843 & ~n20076 ;
  assign n20771 = n19842 & n19866 ;
  assign n20775 = ~n20096 & ~n20771 ;
  assign n20776 = n20774 & n20775 ;
  assign n20777 = ~n20773 & n20776 ;
  assign n20778 = ~n19805 & ~n20777 ;
  assign n20763 = ~n19840 & n20448 ;
  assign n20779 = n19817 & n19845 ;
  assign n20780 = ~n20102 & ~n20779 ;
  assign n20781 = n19840 & ~n20780 ;
  assign n20782 = ~n20763 & ~n20781 ;
  assign n20783 = ~n20778 & n20782 ;
  assign n20784 = ~n20770 & n20783 ;
  assign n20785 = ~\u2_L4_reg[18]/P0001  & ~n20784 ;
  assign n20786 = \u2_L4_reg[18]/P0001  & n20784 ;
  assign n20787 = ~n20785 & ~n20786 ;
  assign n20789 = n20611 & ~n20630 ;
  assign n20790 = ~n20737 & ~n20789 ;
  assign n20791 = ~n20653 & ~n20753 ;
  assign n20792 = n20790 & n20791 ;
  assign n20793 = n20624 & ~n20792 ;
  assign n20794 = n20642 & n20664 ;
  assign n20795 = ~n20793 & ~n20794 ;
  assign n20796 = ~n20598 & ~n20795 ;
  assign n20805 = ~n20633 & ~n20664 ;
  assign n20806 = ~n20624 & ~n20805 ;
  assign n20807 = n20624 & ~n20633 ;
  assign n20808 = ~n20611 & ~n20807 ;
  assign n20809 = ~n20806 & n20808 ;
  assign n20810 = ~n20639 & ~n20809 ;
  assign n20811 = n20598 & ~n20810 ;
  assign n20798 = n20617 & n20644 ;
  assign n20799 = ~n20663 & ~n20798 ;
  assign n20800 = n20598 & ~n20799 ;
  assign n20797 = n20633 & n20664 ;
  assign n20801 = n20617 & n20789 ;
  assign n20802 = ~n20797 & ~n20801 ;
  assign n20803 = ~n20800 & n20802 ;
  assign n20804 = n20624 & ~n20803 ;
  assign n20788 = n20631 & n20731 ;
  assign n20812 = n20633 & ~n20637 ;
  assign n20813 = n20666 & ~n20812 ;
  assign n20814 = ~n20598 & ~n20624 ;
  assign n20815 = ~n20813 & n20814 ;
  assign n20816 = ~n20788 & ~n20815 ;
  assign n20817 = ~n20804 & n20816 ;
  assign n20818 = ~n20811 & n20817 ;
  assign n20819 = ~n20796 & n20818 ;
  assign n20820 = ~\u2_L4_reg[24]/NET0131  & ~n20819 ;
  assign n20821 = \u2_L4_reg[24]/NET0131  & n20819 ;
  assign n20822 = ~n20820 & ~n20821 ;
  assign n20823 = n20644 & ~n20645 ;
  assign n20824 = ~n20604 & n20640 ;
  assign n20825 = ~n20823 & ~n20824 ;
  assign n20826 = n20624 & ~n20825 ;
  assign n20828 = ~n20617 & ~n20664 ;
  assign n20829 = n20624 & ~n20828 ;
  assign n20830 = ~n20611 & n20630 ;
  assign n20827 = n20611 & n20633 ;
  assign n20831 = ~n20645 & ~n20827 ;
  assign n20832 = ~n20830 & n20831 ;
  assign n20833 = ~n20829 & n20832 ;
  assign n20834 = ~n20826 & ~n20833 ;
  assign n20835 = ~n20598 & ~n20834 ;
  assign n20842 = n20790 & ~n20797 ;
  assign n20843 = n20598 & n20624 ;
  assign n20844 = ~n20842 & n20843 ;
  assign n20836 = ~n20644 & ~n20653 ;
  assign n20837 = n20657 & ~n20836 ;
  assign n20840 = n20617 & ~n20636 ;
  assign n20841 = n20652 & n20840 ;
  assign n20838 = n20634 & n20753 ;
  assign n20839 = n20631 & n20645 ;
  assign n20845 = ~n20838 & ~n20839 ;
  assign n20846 = ~n20841 & n20845 ;
  assign n20847 = ~n20837 & n20846 ;
  assign n20848 = ~n20844 & n20847 ;
  assign n20849 = ~n20835 & n20848 ;
  assign n20850 = \u2_L4_reg[30]/NET0131  & ~n20849 ;
  assign n20851 = ~\u2_L4_reg[30]/NET0131  & n20849 ;
  assign n20852 = ~n20850 & ~n20851 ;
  assign n20853 = decrypt_pad & ~\u2_uk_K_r3_reg[30]/NET0131  ;
  assign n20854 = ~decrypt_pad & ~\u2_uk_K_r3_reg[49]/NET0131  ;
  assign n20855 = ~n20853 & ~n20854 ;
  assign n20856 = \u2_R3_reg[27]/NET0131  & ~n20855 ;
  assign n20857 = ~\u2_R3_reg[27]/NET0131  & n20855 ;
  assign n20858 = ~n20856 & ~n20857 ;
  assign n20865 = decrypt_pad & ~\u2_uk_K_r3_reg[36]/NET0131  ;
  assign n20866 = ~decrypt_pad & ~\u2_uk_K_r3_reg[0]/NET0131  ;
  assign n20867 = ~n20865 & ~n20866 ;
  assign n20868 = \u2_R3_reg[25]/NET0131  & ~n20867 ;
  assign n20869 = ~\u2_R3_reg[25]/NET0131  & n20867 ;
  assign n20870 = ~n20868 & ~n20869 ;
  assign n20859 = decrypt_pad & ~\u2_uk_K_r3_reg[21]/NET0131  ;
  assign n20860 = ~decrypt_pad & ~\u2_uk_K_r3_reg[16]/NET0131  ;
  assign n20861 = ~n20859 & ~n20860 ;
  assign n20862 = \u2_R3_reg[26]/NET0131  & ~n20861 ;
  assign n20863 = ~\u2_R3_reg[26]/NET0131  & n20861 ;
  assign n20864 = ~n20862 & ~n20863 ;
  assign n20872 = decrypt_pad & ~\u2_uk_K_r3_reg[1]/NET0131  ;
  assign n20873 = ~decrypt_pad & ~\u2_uk_K_r3_reg[51]/NET0131  ;
  assign n20874 = ~n20872 & ~n20873 ;
  assign n20875 = \u2_R3_reg[24]/NET0131  & ~n20874 ;
  assign n20876 = ~\u2_R3_reg[24]/NET0131  & n20874 ;
  assign n20877 = ~n20875 & ~n20876 ;
  assign n20878 = decrypt_pad & ~\u2_uk_K_r3_reg[9]/NET0131  ;
  assign n20879 = ~decrypt_pad & ~\u2_uk_K_r3_reg[28]/NET0131  ;
  assign n20880 = ~n20878 & ~n20879 ;
  assign n20881 = \u2_R3_reg[29]/NET0131  & ~n20880 ;
  assign n20882 = ~\u2_R3_reg[29]/NET0131  & n20880 ;
  assign n20883 = ~n20881 & ~n20882 ;
  assign n20890 = ~n20877 & ~n20883 ;
  assign n20891 = n20864 & n20890 ;
  assign n20892 = ~n20870 & n20891 ;
  assign n20871 = n20864 & ~n20870 ;
  assign n20884 = n20877 & ~n20883 ;
  assign n20885 = ~n20871 & n20884 ;
  assign n20886 = ~n20864 & ~n20877 ;
  assign n20887 = n20864 & n20877 ;
  assign n20888 = ~n20886 & ~n20887 ;
  assign n20889 = n20883 & ~n20888 ;
  assign n20893 = ~n20885 & ~n20889 ;
  assign n20894 = ~n20892 & n20893 ;
  assign n20895 = ~n20858 & ~n20894 ;
  assign n20896 = ~n20864 & ~n20870 ;
  assign n20897 = n20858 & n20877 ;
  assign n20898 = n20896 & n20897 ;
  assign n20899 = n20870 & n20883 ;
  assign n20900 = ~n20888 & n20899 ;
  assign n20901 = ~n20898 & ~n20900 ;
  assign n20902 = ~n20895 & n20901 ;
  assign n20903 = decrypt_pad & ~\u2_uk_K_r3_reg[45]/P0001  ;
  assign n20904 = ~decrypt_pad & ~\u2_uk_K_r3_reg[36]/NET0131  ;
  assign n20905 = ~n20903 & ~n20904 ;
  assign n20906 = \u2_R3_reg[28]/NET0131  & ~n20905 ;
  assign n20907 = ~\u2_R3_reg[28]/NET0131  & n20905 ;
  assign n20908 = ~n20906 & ~n20907 ;
  assign n20909 = ~n20902 & ~n20908 ;
  assign n20925 = n20877 & n20883 ;
  assign n20926 = n20896 & n20925 ;
  assign n20912 = ~n20877 & n20883 ;
  assign n20927 = n20870 & n20912 ;
  assign n20928 = ~n20926 & ~n20927 ;
  assign n20929 = ~n20858 & ~n20928 ;
  assign n20930 = n20864 & n20870 ;
  assign n20931 = ~n20896 & ~n20930 ;
  assign n20920 = ~n20864 & ~n20883 ;
  assign n20932 = n20897 & ~n20920 ;
  assign n20933 = n20931 & n20932 ;
  assign n20913 = n20871 & n20912 ;
  assign n20923 = ~n20870 & ~n20877 ;
  assign n20924 = n20920 & n20923 ;
  assign n20934 = ~n20913 & ~n20924 ;
  assign n20935 = ~n20933 & n20934 ;
  assign n20936 = ~n20929 & n20935 ;
  assign n20937 = n20908 & ~n20936 ;
  assign n20914 = n20870 & n20891 ;
  assign n20915 = ~n20913 & ~n20914 ;
  assign n20916 = ~n20870 & ~n20883 ;
  assign n20917 = n20877 & n20916 ;
  assign n20918 = n20915 & ~n20917 ;
  assign n20919 = n20858 & ~n20918 ;
  assign n20910 = ~n20858 & n20870 ;
  assign n20911 = ~n20888 & n20910 ;
  assign n20921 = n20858 & ~n20870 ;
  assign n20922 = n20920 & n20921 ;
  assign n20938 = ~n20911 & ~n20922 ;
  assign n20939 = ~n20919 & n20938 ;
  assign n20940 = ~n20937 & n20939 ;
  assign n20941 = ~n20909 & n20940 ;
  assign n20942 = ~\u2_L3_reg[22]/NET0131  & ~n20941 ;
  assign n20943 = \u2_L3_reg[22]/NET0131  & n20941 ;
  assign n20944 = ~n20942 & ~n20943 ;
  assign n20945 = decrypt_pad & ~\u2_uk_K_r3_reg[39]/NET0131  ;
  assign n20946 = ~decrypt_pad & ~\u2_uk_K_r3_reg[5]/NET0131  ;
  assign n20947 = ~n20945 & ~n20946 ;
  assign n20948 = \u2_R3_reg[4]/NET0131  & ~n20947 ;
  assign n20949 = ~\u2_R3_reg[4]/NET0131  & n20947 ;
  assign n20950 = ~n20948 & ~n20949 ;
  assign n20978 = decrypt_pad & ~\u2_uk_K_r3_reg[4]/NET0131  ;
  assign n20979 = ~decrypt_pad & ~\u2_uk_K_r3_reg[27]/NET0131  ;
  assign n20980 = ~n20978 & ~n20979 ;
  assign n20981 = \u2_R3_reg[3]/NET0131  & ~n20980 ;
  assign n20982 = ~\u2_R3_reg[3]/NET0131  & n20980 ;
  assign n20983 = ~n20981 & ~n20982 ;
  assign n20951 = decrypt_pad & ~\u2_uk_K_r3_reg[27]/NET0131  ;
  assign n20952 = ~decrypt_pad & ~\u2_uk_K_r3_reg[18]/NET0131  ;
  assign n20953 = ~n20951 & ~n20952 ;
  assign n20954 = \u2_R3_reg[2]/NET0131  & ~n20953 ;
  assign n20955 = ~\u2_R3_reg[2]/NET0131  & n20953 ;
  assign n20956 = ~n20954 & ~n20955 ;
  assign n20971 = decrypt_pad & ~\u2_uk_K_r3_reg[48]/NET0131  ;
  assign n20972 = ~decrypt_pad & ~\u2_uk_K_r3_reg[39]/NET0131  ;
  assign n20973 = ~n20971 & ~n20972 ;
  assign n20974 = \u2_R3_reg[32]/NET0131  & ~n20973 ;
  assign n20975 = ~\u2_R3_reg[32]/NET0131  & n20973 ;
  assign n20976 = ~n20974 & ~n20975 ;
  assign n20957 = decrypt_pad & ~\u2_uk_K_r3_reg[12]/NET0131  ;
  assign n20958 = ~decrypt_pad & ~\u2_uk_K_r3_reg[3]/NET0131  ;
  assign n20959 = ~n20957 & ~n20958 ;
  assign n20960 = \u2_R3_reg[1]/NET0131  & ~n20959 ;
  assign n20961 = ~\u2_R3_reg[1]/NET0131  & n20959 ;
  assign n20962 = ~n20960 & ~n20961 ;
  assign n20964 = decrypt_pad & ~\u2_uk_K_r3_reg[10]/NET0131  ;
  assign n20965 = ~decrypt_pad & ~\u2_uk_K_r3_reg[33]/NET0131  ;
  assign n20966 = ~n20964 & ~n20965 ;
  assign n20967 = \u2_R3_reg[5]/NET0131  & ~n20966 ;
  assign n20968 = ~\u2_R3_reg[5]/NET0131  & n20966 ;
  assign n20969 = ~n20967 & ~n20968 ;
  assign n20985 = ~n20962 & ~n20969 ;
  assign n20986 = n20976 & n20985 ;
  assign n20987 = n20956 & n20986 ;
  assign n20988 = ~n20962 & n20969 ;
  assign n20989 = ~n20956 & ~n20976 ;
  assign n20990 = ~n20988 & n20989 ;
  assign n20991 = ~n20987 & ~n20990 ;
  assign n20992 = ~n20983 & ~n20991 ;
  assign n20993 = n20969 & ~n20976 ;
  assign n20994 = n20956 & n20983 ;
  assign n20995 = n20993 & n20994 ;
  assign n20996 = ~n20969 & ~n20976 ;
  assign n20997 = ~n20956 & n20996 ;
  assign n20998 = ~n20995 & ~n20997 ;
  assign n20999 = n20962 & ~n20998 ;
  assign n20963 = n20956 & n20962 ;
  assign n20970 = n20963 & ~n20969 ;
  assign n20977 = n20970 & n20976 ;
  assign n20984 = n20977 & n20983 ;
  assign n21000 = n20969 & n20976 ;
  assign n21001 = ~n20956 & n20983 ;
  assign n21002 = ~n20956 & ~n20962 ;
  assign n21003 = ~n21001 & ~n21002 ;
  assign n21004 = n21000 & ~n21003 ;
  assign n21005 = ~n20984 & ~n21004 ;
  assign n21006 = ~n20999 & n21005 ;
  assign n21007 = ~n20992 & n21006 ;
  assign n21008 = ~n20950 & ~n21007 ;
  assign n21010 = n20956 & n20996 ;
  assign n21011 = ~n20988 & ~n21010 ;
  assign n21012 = n20983 & ~n21011 ;
  assign n21018 = n20962 & ~n21001 ;
  assign n21019 = n20993 & ~n21018 ;
  assign n21009 = ~n20956 & n20986 ;
  assign n21013 = ~n20962 & n20976 ;
  assign n21014 = n20956 & ~n20962 ;
  assign n21015 = n20976 & ~n20983 ;
  assign n21016 = ~n21014 & ~n21015 ;
  assign n21017 = ~n21013 & ~n21016 ;
  assign n21020 = ~n21009 & ~n21017 ;
  assign n21021 = ~n21019 & n21020 ;
  assign n21022 = ~n21012 & n21021 ;
  assign n21023 = n20950 & ~n21022 ;
  assign n21024 = ~n20962 & n20983 ;
  assign n21025 = ~n20956 & n20976 ;
  assign n21026 = ~n21010 & ~n21025 ;
  assign n21027 = n21024 & ~n21026 ;
  assign n21032 = ~n20962 & n20993 ;
  assign n21033 = n20956 & n21032 ;
  assign n21028 = n20963 & n20969 ;
  assign n21029 = n20976 & n21028 ;
  assign n21030 = ~n20956 & n20962 ;
  assign n21031 = ~n20969 & n21030 ;
  assign n21034 = ~n21029 & ~n21031 ;
  assign n21035 = ~n21033 & n21034 ;
  assign n21036 = ~n20983 & ~n21035 ;
  assign n21037 = ~n21027 & ~n21036 ;
  assign n21038 = ~n21023 & n21037 ;
  assign n21039 = ~n21008 & n21038 ;
  assign n21040 = ~\u2_L3_reg[31]/NET0131  & ~n21039 ;
  assign n21041 = \u2_L3_reg[31]/NET0131  & n21039 ;
  assign n21042 = ~n21040 & ~n21041 ;
  assign n21094 = decrypt_pad & ~\u2_uk_K_r3_reg[38]/NET0131  ;
  assign n21095 = ~decrypt_pad & ~\u2_uk_K_r3_reg[29]/NET0131  ;
  assign n21096 = ~n21094 & ~n21095 ;
  assign n21097 = \u2_R3_reg[24]/NET0131  & ~n21096 ;
  assign n21098 = ~\u2_R3_reg[24]/NET0131  & n21096 ;
  assign n21099 = ~n21097 & ~n21098 ;
  assign n21049 = decrypt_pad & ~\u2_uk_K_r3_reg[44]/NET0131  ;
  assign n21050 = ~decrypt_pad & ~\u2_uk_K_r3_reg[8]/NET0131  ;
  assign n21051 = ~n21049 & ~n21050 ;
  assign n21052 = \u2_R3_reg[20]/NET0131  & ~n21051 ;
  assign n21053 = ~\u2_R3_reg[20]/NET0131  & n21051 ;
  assign n21054 = ~n21052 & ~n21053 ;
  assign n21062 = decrypt_pad & ~\u2_uk_K_r3_reg[50]/NET0131  ;
  assign n21063 = ~decrypt_pad & ~\u2_uk_K_r3_reg[14]/NET0131  ;
  assign n21064 = ~n21062 & ~n21063 ;
  assign n21065 = \u2_R3_reg[22]/NET0131  & ~n21064 ;
  assign n21066 = ~\u2_R3_reg[22]/NET0131  & n21064 ;
  assign n21067 = ~n21065 & ~n21066 ;
  assign n21068 = decrypt_pad & ~\u2_uk_K_r3_reg[28]/NET0131  ;
  assign n21069 = ~decrypt_pad & ~\u2_uk_K_r3_reg[23]/NET0131  ;
  assign n21070 = ~n21068 & ~n21069 ;
  assign n21071 = \u2_R3_reg[21]/NET0131  & ~n21070 ;
  assign n21072 = ~\u2_R3_reg[21]/NET0131  & n21070 ;
  assign n21073 = ~n21071 & ~n21072 ;
  assign n21103 = ~n21067 & n21073 ;
  assign n21119 = n21054 & n21103 ;
  assign n21043 = decrypt_pad & ~\u2_uk_K_r3_reg[8]/NET0131  ;
  assign n21044 = ~decrypt_pad & ~\u2_uk_K_r3_reg[31]/NET0131  ;
  assign n21045 = ~n21043 & ~n21044 ;
  assign n21046 = \u2_R3_reg[23]/NET0131  & ~n21045 ;
  assign n21047 = ~\u2_R3_reg[23]/NET0131  & n21045 ;
  assign n21048 = ~n21046 & ~n21047 ;
  assign n21076 = ~n21054 & n21073 ;
  assign n21077 = n21067 & n21076 ;
  assign n21120 = ~n21048 & ~n21077 ;
  assign n21121 = ~n21119 & n21120 ;
  assign n21055 = decrypt_pad & ~\u2_uk_K_r3_reg[29]/NET0131  ;
  assign n21056 = ~decrypt_pad & ~\u2_uk_K_r3_reg[52]/NET0131  ;
  assign n21057 = ~n21055 & ~n21056 ;
  assign n21058 = \u2_R3_reg[25]/NET0131  & ~n21057 ;
  assign n21059 = ~\u2_R3_reg[25]/NET0131  & n21057 ;
  assign n21060 = ~n21058 & ~n21059 ;
  assign n21111 = n21060 & ~n21073 ;
  assign n21112 = ~n21054 & n21111 ;
  assign n21113 = n21048 & ~n21112 ;
  assign n21122 = n21067 & ~n21073 ;
  assign n21123 = n21054 & n21122 ;
  assign n21124 = ~n21054 & ~n21067 ;
  assign n21125 = ~n21123 & ~n21124 ;
  assign n21126 = n21113 & n21125 ;
  assign n21127 = ~n21121 & ~n21126 ;
  assign n21078 = n21054 & n21060 ;
  assign n21089 = ~n21073 & n21078 ;
  assign n21116 = n21067 & n21089 ;
  assign n21061 = n21054 & ~n21060 ;
  assign n21083 = ~n21048 & ~n21067 ;
  assign n21117 = ~n21083 & ~n21103 ;
  assign n21118 = n21061 & ~n21117 ;
  assign n21128 = ~n21116 & ~n21118 ;
  assign n21129 = ~n21127 & n21128 ;
  assign n21130 = ~n21099 & ~n21129 ;
  assign n21079 = n21073 & n21078 ;
  assign n21074 = ~n21067 & ~n21073 ;
  assign n21075 = n21061 & n21074 ;
  assign n21080 = ~n21075 & ~n21077 ;
  assign n21081 = ~n21079 & n21080 ;
  assign n21082 = n21048 & ~n21081 ;
  assign n21084 = ~n21076 & ~n21078 ;
  assign n21085 = ~n21048 & n21084 ;
  assign n21086 = ~n21083 & ~n21085 ;
  assign n21087 = n21060 & n21073 ;
  assign n21088 = ~n21054 & n21087 ;
  assign n21090 = ~n21067 & ~n21088 ;
  assign n21091 = ~n21089 & n21090 ;
  assign n21092 = ~n21086 & ~n21091 ;
  assign n21093 = ~n21082 & ~n21092 ;
  assign n21100 = ~n21093 & n21099 ;
  assign n21109 = n21061 & n21073 ;
  assign n21110 = ~n21048 & ~n21109 ;
  assign n21114 = ~n21067 & ~n21110 ;
  assign n21115 = ~n21113 & n21114 ;
  assign n21104 = ~n21078 & ~n21103 ;
  assign n21101 = ~n21054 & ~n21060 ;
  assign n21102 = ~n21067 & ~n21101 ;
  assign n21105 = n21048 & ~n21102 ;
  assign n21106 = ~n21104 & n21105 ;
  assign n21107 = ~n21073 & n21101 ;
  assign n21108 = n21083 & n21107 ;
  assign n21131 = ~n21106 & ~n21108 ;
  assign n21132 = ~n21115 & n21131 ;
  assign n21133 = ~n21100 & n21132 ;
  assign n21134 = ~n21130 & n21133 ;
  assign n21135 = \u2_L3_reg[11]/NET0131  & ~n21134 ;
  assign n21136 = ~\u2_L3_reg[11]/NET0131  & n21134 ;
  assign n21137 = ~n21135 & ~n21136 ;
  assign n21138 = decrypt_pad & ~\u2_uk_K_r3_reg[5]/NET0131  ;
  assign n21139 = ~decrypt_pad & ~\u2_uk_K_r3_reg[53]/NET0131  ;
  assign n21140 = ~n21138 & ~n21139 ;
  assign n21141 = \u2_R3_reg[12]/NET0131  & ~n21140 ;
  assign n21142 = ~\u2_R3_reg[12]/NET0131  & n21140 ;
  assign n21143 = ~n21141 & ~n21142 ;
  assign n21158 = decrypt_pad & ~\u2_uk_K_r3_reg[24]/NET0131  ;
  assign n21159 = ~decrypt_pad & ~\u2_uk_K_r3_reg[47]/NET0131  ;
  assign n21160 = ~n21158 & ~n21159 ;
  assign n21161 = \u2_R3_reg[13]/NET0131  & ~n21160 ;
  assign n21162 = ~\u2_R3_reg[13]/NET0131  & n21160 ;
  assign n21163 = ~n21161 & ~n21162 ;
  assign n21178 = ~n21143 & n21163 ;
  assign n21191 = n21143 & ~n21163 ;
  assign n21192 = ~n21178 & ~n21191 ;
  assign n21151 = decrypt_pad & ~\u2_uk_K_r3_reg[33]/NET0131  ;
  assign n21152 = ~decrypt_pad & ~\u2_uk_K_r3_reg[24]/NET0131  ;
  assign n21153 = ~n21151 & ~n21152 ;
  assign n21154 = \u2_R3_reg[15]/NET0131  & ~n21153 ;
  assign n21155 = ~\u2_R3_reg[15]/NET0131  & n21153 ;
  assign n21156 = ~n21154 & ~n21155 ;
  assign n21168 = decrypt_pad & ~\u2_uk_K_r3_reg[25]/NET0131  ;
  assign n21169 = ~decrypt_pad & ~\u2_uk_K_r3_reg[48]/NET0131  ;
  assign n21170 = ~n21168 & ~n21169 ;
  assign n21171 = \u2_R3_reg[14]/NET0131  & ~n21170 ;
  assign n21172 = ~\u2_R3_reg[14]/NET0131  & n21170 ;
  assign n21173 = ~n21171 & ~n21172 ;
  assign n21193 = ~n21156 & ~n21173 ;
  assign n21194 = ~n21192 & n21193 ;
  assign n21144 = decrypt_pad & ~\u2_uk_K_r3_reg[46]/NET0131  ;
  assign n21145 = ~decrypt_pad & ~\u2_uk_K_r3_reg[12]/NET0131  ;
  assign n21146 = ~n21144 & ~n21145 ;
  assign n21147 = \u2_R3_reg[17]/NET0131  & ~n21146 ;
  assign n21148 = ~\u2_R3_reg[17]/NET0131  & n21146 ;
  assign n21149 = ~n21147 & ~n21148 ;
  assign n21150 = ~n21143 & n21149 ;
  assign n21157 = n21150 & n21156 ;
  assign n21164 = n21157 & ~n21163 ;
  assign n21182 = n21143 & ~n21149 ;
  assign n21183 = n21156 & n21163 ;
  assign n21184 = n21182 & n21183 ;
  assign n21185 = decrypt_pad & ~\u2_uk_K_r3_reg[41]/NET0131  ;
  assign n21186 = ~decrypt_pad & ~\u2_uk_K_r3_reg[32]/NET0131  ;
  assign n21187 = ~n21185 & ~n21186 ;
  assign n21188 = \u2_R3_reg[16]/NET0131  & ~n21187 ;
  assign n21189 = ~\u2_R3_reg[16]/NET0131  & n21187 ;
  assign n21190 = ~n21188 & ~n21189 ;
  assign n21195 = ~n21184 & n21190 ;
  assign n21196 = ~n21164 & n21195 ;
  assign n21197 = ~n21194 & n21196 ;
  assign n21165 = ~n21143 & ~n21163 ;
  assign n21166 = ~n21149 & n21165 ;
  assign n21167 = ~n21156 & n21166 ;
  assign n21174 = n21167 & n21173 ;
  assign n21175 = n21143 & n21149 ;
  assign n21176 = n21163 & n21175 ;
  assign n21177 = n21173 & n21176 ;
  assign n21179 = n21149 & ~n21173 ;
  assign n21180 = n21178 & n21179 ;
  assign n21181 = ~n21177 & ~n21180 ;
  assign n21198 = ~n21174 & n21181 ;
  assign n21199 = n21197 & n21198 ;
  assign n21209 = ~n21173 & n21191 ;
  assign n21210 = n21149 & n21209 ;
  assign n21214 = n21175 & n21183 ;
  assign n21215 = ~n21190 & ~n21214 ;
  assign n21216 = ~n21210 & n21215 ;
  assign n21211 = n21156 & n21166 ;
  assign n21212 = n21173 & n21183 ;
  assign n21213 = ~n21143 & n21212 ;
  assign n21217 = ~n21211 & ~n21213 ;
  assign n21218 = n21216 & n21217 ;
  assign n21200 = n21173 & n21182 ;
  assign n21201 = n21149 & ~n21163 ;
  assign n21202 = ~n21200 & ~n21201 ;
  assign n21203 = ~n21156 & ~n21202 ;
  assign n21204 = ~n21149 & n21178 ;
  assign n21205 = n21173 & n21204 ;
  assign n21206 = ~n21149 & ~n21173 ;
  assign n21207 = n21165 & n21206 ;
  assign n21208 = ~n21205 & ~n21207 ;
  assign n21219 = ~n21203 & n21208 ;
  assign n21220 = n21218 & n21219 ;
  assign n21221 = ~n21199 & ~n21220 ;
  assign n21224 = ~n21163 & n21200 ;
  assign n21222 = n21163 & ~n21173 ;
  assign n21223 = n21182 & n21222 ;
  assign n21225 = ~n21207 & ~n21223 ;
  assign n21226 = ~n21224 & n21225 ;
  assign n21227 = n21156 & ~n21226 ;
  assign n21228 = n21149 & n21193 ;
  assign n21229 = n21178 & n21228 ;
  assign n21230 = ~n21227 & ~n21229 ;
  assign n21231 = ~n21221 & n21230 ;
  assign n21232 = ~\u2_L3_reg[20]/NET0131  & ~n21231 ;
  assign n21233 = \u2_L3_reg[20]/NET0131  & n21231 ;
  assign n21234 = ~n21232 & ~n21233 ;
  assign n21279 = decrypt_pad & ~\u2_uk_K_r3_reg[37]/NET0131  ;
  assign n21280 = ~decrypt_pad & ~\u2_uk_K_r3_reg[1]/NET0131  ;
  assign n21281 = ~n21279 & ~n21280 ;
  assign n21282 = \u2_R3_reg[32]/NET0131  & ~n21281 ;
  assign n21283 = ~\u2_R3_reg[32]/NET0131  & n21281 ;
  assign n21284 = ~n21282 & ~n21283 ;
  assign n21241 = decrypt_pad & ~\u2_uk_K_r3_reg[31]/NET0131  ;
  assign n21242 = ~decrypt_pad & ~\u2_uk_K_r3_reg[22]/NET0131  ;
  assign n21243 = ~n21241 & ~n21242 ;
  assign n21244 = \u2_R3_reg[1]/NET0131  & ~n21243 ;
  assign n21245 = ~\u2_R3_reg[1]/NET0131  & n21243 ;
  assign n21246 = ~n21244 & ~n21245 ;
  assign n21247 = decrypt_pad & ~\u2_uk_K_r3_reg[15]/NET0131  ;
  assign n21248 = ~decrypt_pad & ~\u2_uk_K_r3_reg[38]/NET0131  ;
  assign n21249 = ~n21247 & ~n21248 ;
  assign n21250 = \u2_R3_reg[28]/NET0131  & ~n21249 ;
  assign n21251 = ~\u2_R3_reg[28]/NET0131  & n21249 ;
  assign n21252 = ~n21250 & ~n21251 ;
  assign n21235 = decrypt_pad & ~\u2_uk_K_r3_reg[43]/NET0131  ;
  assign n21236 = ~decrypt_pad & ~\u2_uk_K_r3_reg[7]/NET0131  ;
  assign n21237 = ~n21235 & ~n21236 ;
  assign n21238 = \u2_R3_reg[30]/NET0131  & ~n21237 ;
  assign n21239 = ~\u2_R3_reg[30]/NET0131  & n21237 ;
  assign n21240 = ~n21238 & ~n21239 ;
  assign n21254 = decrypt_pad & ~\u2_uk_K_r3_reg[42]/NET0131  ;
  assign n21255 = ~decrypt_pad & ~\u2_uk_K_r3_reg[37]/NET0131  ;
  assign n21256 = ~n21254 & ~n21255 ;
  assign n21257 = \u2_R3_reg[29]/NET0131  & ~n21256 ;
  assign n21258 = ~\u2_R3_reg[29]/NET0131  & n21256 ;
  assign n21259 = ~n21257 & ~n21258 ;
  assign n21286 = n21240 & ~n21259 ;
  assign n21287 = n21252 & n21286 ;
  assign n21288 = ~n21246 & n21287 ;
  assign n21264 = decrypt_pad & ~\u2_uk_K_r3_reg[0]/NET0131  ;
  assign n21265 = ~decrypt_pad & ~\u2_uk_K_r3_reg[50]/NET0131  ;
  assign n21266 = ~n21264 & ~n21265 ;
  assign n21267 = \u2_R3_reg[31]/P0001  & ~n21266 ;
  assign n21268 = ~\u2_R3_reg[31]/P0001  & n21266 ;
  assign n21269 = ~n21267 & ~n21268 ;
  assign n21253 = n21246 & ~n21252 ;
  assign n21289 = n21253 & ~n21259 ;
  assign n21290 = n21269 & ~n21289 ;
  assign n21291 = ~n21288 & n21290 ;
  assign n21293 = ~n21246 & ~n21252 ;
  assign n21294 = n21240 & n21293 ;
  assign n21292 = n21246 & n21259 ;
  assign n21295 = ~n21269 & ~n21292 ;
  assign n21296 = ~n21294 & n21295 ;
  assign n21297 = ~n21291 & ~n21296 ;
  assign n21300 = n21240 & n21259 ;
  assign n21301 = n21246 & n21300 ;
  assign n21271 = ~n21246 & n21259 ;
  assign n21298 = ~n21240 & n21271 ;
  assign n21299 = ~n21240 & ~n21269 ;
  assign n21302 = ~n21298 & ~n21299 ;
  assign n21303 = ~n21301 & n21302 ;
  assign n21304 = n21252 & ~n21303 ;
  assign n21305 = ~n21297 & ~n21304 ;
  assign n21306 = ~n21284 & ~n21305 ;
  assign n21260 = n21253 & n21259 ;
  assign n21261 = n21240 & n21260 ;
  assign n21262 = ~n21240 & ~n21259 ;
  assign n21263 = ~n21252 & n21262 ;
  assign n21270 = ~n21263 & ~n21269 ;
  assign n21272 = ~n21240 & n21252 ;
  assign n21274 = n21271 & ~n21272 ;
  assign n21273 = ~n21271 & n21272 ;
  assign n21275 = n21269 & ~n21273 ;
  assign n21276 = ~n21274 & n21275 ;
  assign n21277 = ~n21270 & ~n21276 ;
  assign n21278 = ~n21261 & ~n21277 ;
  assign n21285 = ~n21278 & n21284 ;
  assign n21312 = ~n21252 & n21300 ;
  assign n21313 = ~n21246 & n21312 ;
  assign n21314 = ~n21246 & n21263 ;
  assign n21315 = ~n21313 & ~n21314 ;
  assign n21316 = n21246 & n21252 ;
  assign n21317 = n21262 & n21316 ;
  assign n21318 = n21240 & n21289 ;
  assign n21319 = ~n21317 & ~n21318 ;
  assign n21320 = n21315 & n21319 ;
  assign n21321 = n21269 & ~n21320 ;
  assign n21307 = ~n21269 & n21284 ;
  assign n21308 = n21287 & n21307 ;
  assign n21309 = n21252 & n21259 ;
  assign n21310 = ~n21246 & n21309 ;
  assign n21311 = n21299 & n21310 ;
  assign n21322 = ~n21308 & ~n21311 ;
  assign n21323 = ~n21321 & n21322 ;
  assign n21324 = ~n21285 & n21323 ;
  assign n21325 = ~n21306 & n21324 ;
  assign n21326 = \u2_L3_reg[5]/NET0131  & ~n21325 ;
  assign n21327 = ~\u2_L3_reg[5]/NET0131  & n21325 ;
  assign n21328 = ~n21326 & ~n21327 ;
  assign n21342 = n21156 & ~n21179 ;
  assign n21343 = n21191 & n21342 ;
  assign n21341 = n21157 & ~n21173 ;
  assign n21346 = ~n21167 & ~n21341 ;
  assign n21347 = ~n21343 & n21346 ;
  assign n21344 = ~n21222 & ~n21228 ;
  assign n21345 = n21143 & ~n21344 ;
  assign n21348 = n21208 & ~n21345 ;
  assign n21349 = n21347 & n21348 ;
  assign n21350 = ~n21190 & ~n21349 ;
  assign n21336 = ~n21204 & ~n21210 ;
  assign n21337 = n21156 & ~n21336 ;
  assign n21330 = n21165 & n21173 ;
  assign n21331 = n21149 & n21330 ;
  assign n21332 = ~n21177 & ~n21331 ;
  assign n21333 = n21182 & ~n21222 ;
  assign n21334 = ~n21180 & ~n21333 ;
  assign n21335 = ~n21156 & ~n21334 ;
  assign n21338 = n21332 & ~n21335 ;
  assign n21339 = ~n21337 & n21338 ;
  assign n21340 = n21190 & ~n21339 ;
  assign n21351 = ~n21207 & n21332 ;
  assign n21352 = ~n21156 & ~n21351 ;
  assign n21329 = n21156 & n21223 ;
  assign n21353 = ~n21213 & ~n21329 ;
  assign n21354 = ~n21352 & n21353 ;
  assign n21355 = ~n21340 & n21354 ;
  assign n21356 = ~n21350 & n21355 ;
  assign n21357 = ~\u2_L3_reg[10]/NET0131  & ~n21356 ;
  assign n21358 = \u2_L3_reg[10]/NET0131  & n21356 ;
  assign n21359 = ~n21357 & ~n21358 ;
  assign n21365 = n20871 & n20925 ;
  assign n21360 = ~n20858 & n20887 ;
  assign n21369 = ~n20908 & ~n21360 ;
  assign n21370 = ~n21365 & n21369 ;
  assign n21361 = ~n20921 & ~n20930 ;
  assign n21362 = n20912 & ~n21361 ;
  assign n21363 = ~n20899 & ~n20916 ;
  assign n21364 = ~n20858 & ~n21363 ;
  assign n21371 = ~n21362 & ~n21364 ;
  assign n21366 = n20888 & n20916 ;
  assign n21367 = n20870 & n20890 ;
  assign n21368 = ~n20864 & n21367 ;
  assign n21372 = ~n21366 & ~n21368 ;
  assign n21373 = n21371 & n21372 ;
  assign n21374 = n21370 & n21373 ;
  assign n21376 = n20864 & n20917 ;
  assign n21375 = ~n20858 & n20913 ;
  assign n21383 = ~n20914 & ~n21375 ;
  assign n21384 = ~n21376 & n21383 ;
  assign n21378 = n20870 & n20877 ;
  assign n21379 = ~n20924 & ~n21378 ;
  assign n21380 = n20858 & ~n21379 ;
  assign n21377 = n20886 & n20899 ;
  assign n21381 = n20908 & ~n20926 ;
  assign n21382 = ~n21377 & n21381 ;
  assign n21385 = ~n21380 & n21382 ;
  assign n21386 = n21384 & n21385 ;
  assign n21387 = ~n21374 & ~n21386 ;
  assign n21388 = \u2_L3_reg[12]/NET0131  & n21387 ;
  assign n21389 = ~\u2_L3_reg[12]/NET0131  & ~n21387 ;
  assign n21390 = ~n21388 & ~n21389 ;
  assign n21391 = decrypt_pad & ~\u2_uk_K_r3_reg[7]/NET0131  ;
  assign n21392 = ~decrypt_pad & ~\u2_uk_K_r3_reg[2]/NET0131  ;
  assign n21393 = ~n21391 & ~n21392 ;
  assign n21394 = \u2_R3_reg[19]/NET0131  & ~n21393 ;
  assign n21395 = ~\u2_R3_reg[19]/NET0131  & n21393 ;
  assign n21396 = ~n21394 & ~n21395 ;
  assign n21397 = decrypt_pad & ~\u2_uk_K_r3_reg[51]/NET0131  ;
  assign n21398 = ~decrypt_pad & ~\u2_uk_K_r3_reg[15]/NET0131  ;
  assign n21399 = ~n21397 & ~n21398 ;
  assign n21400 = \u2_R3_reg[18]/NET0131  & ~n21399 ;
  assign n21401 = ~\u2_R3_reg[18]/NET0131  & n21399 ;
  assign n21402 = ~n21400 & ~n21401 ;
  assign n21403 = decrypt_pad & ~\u2_uk_K_r3_reg[2]/NET0131  ;
  assign n21404 = ~decrypt_pad & ~\u2_uk_K_r3_reg[21]/NET0131  ;
  assign n21405 = ~n21403 & ~n21404 ;
  assign n21406 = \u2_R3_reg[17]/NET0131  & ~n21405 ;
  assign n21407 = ~\u2_R3_reg[17]/NET0131  & n21405 ;
  assign n21408 = ~n21406 & ~n21407 ;
  assign n21410 = decrypt_pad & ~\u2_uk_K_r3_reg[35]/NET0131  ;
  assign n21411 = ~decrypt_pad & ~\u2_uk_K_r3_reg[30]/NET0131  ;
  assign n21412 = ~n21410 & ~n21411 ;
  assign n21413 = \u2_R3_reg[16]/NET0131  & ~n21412 ;
  assign n21414 = ~\u2_R3_reg[16]/NET0131  & n21412 ;
  assign n21415 = ~n21413 & ~n21414 ;
  assign n21417 = decrypt_pad & ~\u2_uk_K_r3_reg[23]/NET0131  ;
  assign n21418 = ~decrypt_pad & ~\u2_uk_K_r3_reg[42]/NET0131  ;
  assign n21419 = ~n21417 & ~n21418 ;
  assign n21420 = \u2_R3_reg[21]/NET0131  & ~n21419 ;
  assign n21421 = ~\u2_R3_reg[21]/NET0131  & n21419 ;
  assign n21422 = ~n21420 & ~n21421 ;
  assign n21423 = n21415 & ~n21422 ;
  assign n21434 = ~n21408 & n21423 ;
  assign n21435 = ~n21402 & n21434 ;
  assign n21409 = ~n21402 & n21408 ;
  assign n21436 = n21415 & n21422 ;
  assign n21437 = n21409 & n21436 ;
  assign n21426 = n21408 & ~n21422 ;
  assign n21431 = n21402 & n21426 ;
  assign n21432 = ~n21415 & n21422 ;
  assign n21433 = ~n21408 & n21432 ;
  assign n21438 = ~n21431 & ~n21433 ;
  assign n21439 = ~n21437 & n21438 ;
  assign n21440 = ~n21435 & n21439 ;
  assign n21441 = ~n21396 & ~n21440 ;
  assign n21416 = n21409 & ~n21415 ;
  assign n21424 = n21402 & n21415 ;
  assign n21425 = n21422 & ~n21424 ;
  assign n21427 = ~n21423 & ~n21426 ;
  assign n21428 = ~n21425 & n21427 ;
  assign n21429 = ~n21416 & ~n21428 ;
  assign n21430 = n21396 & ~n21429 ;
  assign n21442 = ~n21402 & n21422 ;
  assign n21443 = ~n21423 & ~n21442 ;
  assign n21444 = ~n21408 & ~n21415 ;
  assign n21445 = n21402 & n21408 ;
  assign n21446 = ~n21444 & ~n21445 ;
  assign n21447 = n21443 & n21446 ;
  assign n21448 = ~n21430 & ~n21447 ;
  assign n21449 = ~n21441 & n21448 ;
  assign n21450 = decrypt_pad & ~\u2_uk_K_r3_reg[22]/NET0131  ;
  assign n21451 = ~decrypt_pad & ~\u2_uk_K_r3_reg[45]/P0001  ;
  assign n21452 = ~n21450 & ~n21451 ;
  assign n21453 = \u2_R3_reg[20]/NET0131  & ~n21452 ;
  assign n21454 = ~\u2_R3_reg[20]/NET0131  & n21452 ;
  assign n21455 = ~n21453 & ~n21454 ;
  assign n21456 = ~n21449 & ~n21455 ;
  assign n21460 = ~n21416 & n21425 ;
  assign n21461 = n21415 & n21426 ;
  assign n21462 = ~n21460 & ~n21461 ;
  assign n21463 = n21396 & ~n21462 ;
  assign n21464 = n21408 & n21432 ;
  assign n21465 = ~n21422 & n21444 ;
  assign n21466 = ~n21464 & ~n21465 ;
  assign n21467 = ~n21396 & ~n21402 ;
  assign n21468 = ~n21466 & n21467 ;
  assign n21457 = n21402 & ~n21408 ;
  assign n21458 = ~n21409 & ~n21457 ;
  assign n21459 = n21423 & ~n21458 ;
  assign n21469 = n21396 & n21402 ;
  assign n21470 = n21436 & ~n21469 ;
  assign n21471 = n21458 & n21470 ;
  assign n21472 = ~n21459 & ~n21471 ;
  assign n21473 = ~n21468 & n21472 ;
  assign n21474 = ~n21463 & n21473 ;
  assign n21475 = n21455 & ~n21474 ;
  assign n21476 = n21402 & n21465 ;
  assign n21477 = ~n21402 & n21461 ;
  assign n21478 = ~n21476 & ~n21477 ;
  assign n21479 = n21396 & ~n21478 ;
  assign n21480 = n21402 & n21433 ;
  assign n21481 = ~n21415 & n21431 ;
  assign n21482 = ~n21480 & ~n21481 ;
  assign n21483 = ~n21396 & ~n21482 ;
  assign n21484 = ~n21479 & ~n21483 ;
  assign n21485 = ~n21475 & n21484 ;
  assign n21486 = ~n21456 & n21485 ;
  assign n21487 = ~\u2_L3_reg[14]/NET0131  & ~n21486 ;
  assign n21488 = \u2_L3_reg[14]/NET0131  & n21486 ;
  assign n21489 = ~n21487 & ~n21488 ;
  assign n21506 = ~n20976 & ~n21002 ;
  assign n21507 = n21000 & n21002 ;
  assign n21508 = ~n21506 & ~n21507 ;
  assign n21509 = n20983 & ~n21508 ;
  assign n21510 = ~n20983 & ~n21025 ;
  assign n21511 = ~n21506 & n21510 ;
  assign n21505 = n20976 & n21031 ;
  assign n21512 = ~n21028 & ~n21505 ;
  assign n21513 = ~n21511 & n21512 ;
  assign n21514 = ~n21509 & n21513 ;
  assign n21515 = n20950 & ~n21514 ;
  assign n21490 = ~n20956 & n20993 ;
  assign n21491 = ~n21010 & ~n21490 ;
  assign n21492 = n20962 & ~n21491 ;
  assign n21493 = n20962 & n21000 ;
  assign n21494 = ~n20986 & ~n21493 ;
  assign n21495 = ~n20950 & ~n21494 ;
  assign n21496 = ~n21492 & ~n21495 ;
  assign n21497 = n20983 & ~n21496 ;
  assign n21499 = n20962 & ~n20997 ;
  assign n21498 = ~n20996 & ~n21000 ;
  assign n21500 = ~n20983 & ~n21498 ;
  assign n21501 = ~n21499 & n21500 ;
  assign n21502 = ~n20977 & ~n21033 ;
  assign n21503 = ~n21501 & n21502 ;
  assign n21504 = ~n20950 & ~n21503 ;
  assign n21516 = ~n21497 & ~n21504 ;
  assign n21517 = ~n21515 & n21516 ;
  assign n21518 = ~\u2_L3_reg[17]/NET0131  & ~n21517 ;
  assign n21519 = \u2_L3_reg[17]/NET0131  & n21517 ;
  assign n21520 = ~n21518 & ~n21519 ;
  assign n21521 = ~n21246 & n21272 ;
  assign n21522 = ~n21259 & n21521 ;
  assign n21523 = ~n21289 & ~n21309 ;
  assign n21524 = ~n21298 & n21523 ;
  assign n21525 = n21269 & ~n21524 ;
  assign n21526 = ~n21522 & ~n21525 ;
  assign n21527 = ~n21284 & ~n21526 ;
  assign n21538 = ~n21240 & n21260 ;
  assign n21539 = ~n21287 & ~n21538 ;
  assign n21540 = n21315 & n21539 ;
  assign n21541 = ~n21269 & ~n21540 ;
  assign n21528 = n21259 & n21272 ;
  assign n21534 = ~n21313 & ~n21528 ;
  assign n21529 = ~n21259 & n21293 ;
  assign n21530 = n21269 & n21529 ;
  assign n21531 = n21246 & n21286 ;
  assign n21532 = ~n21252 & n21269 ;
  assign n21533 = n21531 & ~n21532 ;
  assign n21535 = ~n21530 & ~n21533 ;
  assign n21536 = n21534 & n21535 ;
  assign n21537 = n21284 & ~n21536 ;
  assign n21542 = ~n21240 & n21289 ;
  assign n21543 = ~n21261 & ~n21542 ;
  assign n21544 = n21269 & ~n21543 ;
  assign n21545 = n21252 & ~n21259 ;
  assign n21546 = ~n21269 & ~n21284 ;
  assign n21547 = n21545 & n21546 ;
  assign n21548 = ~n21544 & ~n21547 ;
  assign n21549 = ~n21537 & n21548 ;
  assign n21550 = ~n21541 & n21549 ;
  assign n21551 = ~n21527 & n21550 ;
  assign n21552 = ~\u2_L3_reg[15]/NET0131  & ~n21551 ;
  assign n21553 = \u2_L3_reg[15]/NET0131  & n21551 ;
  assign n21554 = ~n21552 & ~n21553 ;
  assign n21569 = ~n21201 & ~n21206 ;
  assign n21570 = n21143 & ~n21569 ;
  assign n21571 = ~n21156 & ~n21570 ;
  assign n21572 = ~n21143 & n21206 ;
  assign n21573 = n21156 & ~n21572 ;
  assign n21574 = ~n21224 & n21573 ;
  assign n21575 = ~n21571 & ~n21574 ;
  assign n21576 = n21181 & ~n21223 ;
  assign n21577 = ~n21575 & n21576 ;
  assign n21578 = ~n21190 & ~n21577 ;
  assign n21562 = ~n21182 & n21222 ;
  assign n21563 = n21150 & n21163 ;
  assign n21564 = ~n21562 & ~n21563 ;
  assign n21565 = ~n21156 & ~n21564 ;
  assign n21560 = n21163 & n21200 ;
  assign n21566 = ~n21330 & ~n21560 ;
  assign n21567 = ~n21565 & n21566 ;
  assign n21568 = n21190 & ~n21567 ;
  assign n21555 = ~n21205 & n21332 ;
  assign n21556 = n21156 & ~n21555 ;
  assign n21561 = ~n21156 & n21560 ;
  assign n21557 = ~n21201 & ~n21209 ;
  assign n21558 = n21156 & n21190 ;
  assign n21559 = ~n21557 & n21558 ;
  assign n21579 = ~n21174 & ~n21559 ;
  assign n21580 = ~n21561 & n21579 ;
  assign n21581 = ~n21556 & n21580 ;
  assign n21582 = ~n21568 & n21581 ;
  assign n21583 = ~n21578 & n21582 ;
  assign n21584 = ~\u2_L3_reg[1]/NET0131  & ~n21583 ;
  assign n21585 = \u2_L3_reg[1]/NET0131  & n21583 ;
  assign n21586 = ~n21584 & ~n21585 ;
  assign n21612 = n21240 & n21309 ;
  assign n21611 = n21246 & n21262 ;
  assign n21613 = ~n21260 & ~n21611 ;
  assign n21614 = ~n21612 & n21613 ;
  assign n21615 = n21269 & ~n21614 ;
  assign n21606 = n21252 & n21531 ;
  assign n21607 = ~n21521 & ~n21606 ;
  assign n21608 = ~n21269 & ~n21607 ;
  assign n21609 = ~n21310 & ~n21529 ;
  assign n21610 = n21240 & ~n21609 ;
  assign n21616 = ~n21542 & ~n21610 ;
  assign n21617 = ~n21608 & n21616 ;
  assign n21618 = ~n21615 & n21617 ;
  assign n21619 = n21284 & ~n21618 ;
  assign n21593 = ~n21240 & n21259 ;
  assign n21594 = ~n21299 & ~n21593 ;
  assign n21595 = n21316 & ~n21594 ;
  assign n21598 = ~n21288 & ~n21314 ;
  assign n21599 = ~n21595 & n21598 ;
  assign n21587 = ~n21287 & ~n21310 ;
  assign n21588 = n21269 & ~n21587 ;
  assign n21591 = n21259 & ~n21269 ;
  assign n21592 = n21293 & n21591 ;
  assign n21589 = n21240 & ~n21269 ;
  assign n21590 = n21253 & n21589 ;
  assign n21596 = ~n21312 & ~n21590 ;
  assign n21597 = ~n21592 & n21596 ;
  assign n21600 = ~n21588 & n21597 ;
  assign n21601 = n21599 & n21600 ;
  assign n21602 = ~n21284 & ~n21601 ;
  assign n21603 = n21252 & n21292 ;
  assign n21604 = n21299 & n21603 ;
  assign n21605 = n21263 & n21269 ;
  assign n21620 = ~n21604 & ~n21605 ;
  assign n21621 = ~n21602 & n21620 ;
  assign n21622 = ~n21619 & n21621 ;
  assign n21623 = ~\u2_L3_reg[21]/NET0131  & ~n21622 ;
  assign n21624 = \u2_L3_reg[21]/NET0131  & n21622 ;
  assign n21625 = ~n21623 & ~n21624 ;
  assign n21644 = ~n21149 & ~n21163 ;
  assign n21645 = ~n21330 & ~n21644 ;
  assign n21646 = ~n21190 & ~n21645 ;
  assign n21647 = ~n21149 & ~n21192 ;
  assign n21648 = ~n21176 & ~n21647 ;
  assign n21649 = ~n21173 & ~n21648 ;
  assign n21650 = ~n21646 & ~n21649 ;
  assign n21651 = ~n21156 & ~n21650 ;
  assign n21632 = n21178 & n21206 ;
  assign n21633 = n21190 & ~n21632 ;
  assign n21634 = ~n21211 & n21633 ;
  assign n21635 = ~n21560 & n21634 ;
  assign n21626 = ~n21157 & ~n21563 ;
  assign n21627 = n21173 & ~n21626 ;
  assign n21628 = n21173 & n21175 ;
  assign n21629 = n21165 & n21179 ;
  assign n21630 = ~n21628 & ~n21629 ;
  assign n21631 = ~n21156 & ~n21630 ;
  assign n21636 = ~n21627 & ~n21631 ;
  assign n21637 = n21635 & n21636 ;
  assign n21638 = ~n21150 & n21212 ;
  assign n21639 = ~n21180 & ~n21190 ;
  assign n21640 = ~n21184 & ~n21209 ;
  assign n21641 = n21639 & n21640 ;
  assign n21642 = ~n21638 & n21641 ;
  assign n21643 = ~n21637 & ~n21642 ;
  assign n21652 = n21156 & n21179 ;
  assign n21653 = ~n21192 & n21652 ;
  assign n21654 = ~n21643 & ~n21653 ;
  assign n21655 = ~n21651 & n21654 ;
  assign n21656 = ~\u2_L3_reg[26]/NET0131  & ~n21655 ;
  assign n21657 = \u2_L3_reg[26]/NET0131  & n21655 ;
  assign n21658 = ~n21656 & ~n21657 ;
  assign n21675 = n21061 & ~n21073 ;
  assign n21676 = ~n21079 & ~n21675 ;
  assign n21677 = ~n21074 & ~n21077 ;
  assign n21678 = ~n21060 & ~n21677 ;
  assign n21679 = n21676 & ~n21678 ;
  assign n21680 = n21048 & ~n21679 ;
  assign n21659 = n21067 & n21109 ;
  assign n21666 = ~n21067 & ~n21084 ;
  assign n21681 = ~n21659 & ~n21666 ;
  assign n21682 = ~n21048 & ~n21681 ;
  assign n21683 = n21067 & n21112 ;
  assign n21684 = ~n21682 & ~n21683 ;
  assign n21685 = ~n21680 & n21684 ;
  assign n21686 = ~n21099 & ~n21685 ;
  assign n21660 = n21073 & n21124 ;
  assign n21661 = ~n21088 & ~n21660 ;
  assign n21662 = ~n21659 & n21661 ;
  assign n21663 = n21048 & ~n21662 ;
  assign n21667 = n21048 & ~n21111 ;
  assign n21668 = ~n21122 & n21667 ;
  assign n21664 = n21067 & ~n21078 ;
  assign n21665 = ~n21101 & n21664 ;
  assign n21669 = ~n21665 & ~n21666 ;
  assign n21670 = ~n21668 & n21669 ;
  assign n21671 = ~n21663 & ~n21670 ;
  assign n21672 = n21099 & ~n21671 ;
  assign n21673 = n21048 & n21060 ;
  assign n21674 = n21103 & n21673 ;
  assign n21687 = ~n21075 & ~n21674 ;
  assign n21688 = ~n21672 & n21687 ;
  assign n21689 = ~n21686 & n21688 ;
  assign n21690 = \u2_L3_reg[29]/NET0131  & ~n21689 ;
  assign n21691 = ~\u2_L3_reg[29]/NET0131  & n21689 ;
  assign n21692 = ~n21690 & ~n21691 ;
  assign n21695 = ~n21409 & ~n21422 ;
  assign n21696 = ~n21424 & n21695 ;
  assign n21694 = n21408 & n21436 ;
  assign n21697 = ~n21444 & ~n21694 ;
  assign n21698 = ~n21696 & n21697 ;
  assign n21699 = n21396 & ~n21698 ;
  assign n21700 = ~n21408 & n21436 ;
  assign n21701 = ~n21416 & ~n21700 ;
  assign n21702 = ~n21396 & ~n21701 ;
  assign n21693 = n21408 & n21442 ;
  assign n21703 = n21424 & n21426 ;
  assign n21704 = ~n21693 & ~n21703 ;
  assign n21705 = ~n21702 & n21704 ;
  assign n21706 = ~n21699 & n21705 ;
  assign n21707 = n21455 & ~n21706 ;
  assign n21719 = ~n21476 & ~n21703 ;
  assign n21720 = ~n21402 & n21433 ;
  assign n21721 = n21719 & ~n21720 ;
  assign n21722 = n21396 & ~n21721 ;
  assign n21713 = n21396 & ~n21426 ;
  assign n21712 = ~n21396 & ~n21444 ;
  assign n21714 = ~n21402 & ~n21712 ;
  assign n21715 = ~n21713 & n21714 ;
  assign n21708 = ~n21396 & n21434 ;
  assign n21709 = n21396 & ~n21422 ;
  assign n21710 = ~n21415 & n21445 ;
  assign n21711 = ~n21709 & n21710 ;
  assign n21716 = ~n21708 & ~n21711 ;
  assign n21717 = ~n21715 & n21716 ;
  assign n21718 = ~n21455 & ~n21717 ;
  assign n21723 = ~n21396 & n21415 ;
  assign n21724 = n21457 & n21723 ;
  assign n21725 = ~n21437 & ~n21724 ;
  assign n21726 = ~n21718 & n21725 ;
  assign n21727 = ~n21722 & n21726 ;
  assign n21728 = ~n21707 & n21727 ;
  assign n21729 = ~\u2_L3_reg[25]/NET0131  & ~n21728 ;
  assign n21730 = \u2_L3_reg[25]/NET0131  & n21728 ;
  assign n21731 = ~n21729 & ~n21730 ;
  assign n21732 = decrypt_pad & ~\u2_uk_K_r3_reg[40]/NET0131  ;
  assign n21733 = ~decrypt_pad & ~\u2_uk_K_r3_reg[6]/NET0131  ;
  assign n21734 = ~n21732 & ~n21733 ;
  assign n21735 = \u2_R3_reg[8]/NET0131  & ~n21734 ;
  assign n21736 = ~\u2_R3_reg[8]/NET0131  & n21734 ;
  assign n21737 = ~n21735 & ~n21736 ;
  assign n21738 = decrypt_pad & ~\u2_uk_K_r3_reg[32]/NET0131  ;
  assign n21739 = ~decrypt_pad & ~\u2_uk_K_r3_reg[55]/NET0131  ;
  assign n21740 = ~n21738 & ~n21739 ;
  assign n21741 = \u2_R3_reg[5]/NET0131  & ~n21740 ;
  assign n21742 = ~\u2_R3_reg[5]/NET0131  & n21740 ;
  assign n21743 = ~n21741 & ~n21742 ;
  assign n21744 = decrypt_pad & ~\u2_uk_K_r3_reg[20]/NET0131  ;
  assign n21745 = ~decrypt_pad & ~\u2_uk_K_r3_reg[11]/NET0131  ;
  assign n21746 = ~n21744 & ~n21745 ;
  assign n21747 = \u2_R3_reg[9]/NET0131  & ~n21746 ;
  assign n21748 = ~\u2_R3_reg[9]/NET0131  & n21746 ;
  assign n21749 = ~n21747 & ~n21748 ;
  assign n21750 = n21743 & ~n21749 ;
  assign n21751 = ~n21743 & n21749 ;
  assign n21752 = decrypt_pad & ~\u2_uk_K_r3_reg[53]/NET0131  ;
  assign n21753 = ~decrypt_pad & ~\u2_uk_K_r3_reg[19]/NET0131  ;
  assign n21754 = ~n21752 & ~n21753 ;
  assign n21755 = \u2_R3_reg[4]/NET0131  & ~n21754 ;
  assign n21756 = ~\u2_R3_reg[4]/NET0131  & n21754 ;
  assign n21757 = ~n21755 & ~n21756 ;
  assign n21758 = n21751 & ~n21757 ;
  assign n21759 = ~n21750 & ~n21758 ;
  assign n21760 = decrypt_pad & ~\u2_uk_K_r3_reg[55]/NET0131  ;
  assign n21761 = ~decrypt_pad & ~\u2_uk_K_r3_reg[46]/NET0131  ;
  assign n21762 = ~n21760 & ~n21761 ;
  assign n21763 = \u2_R3_reg[6]/NET0131  & ~n21762 ;
  assign n21764 = ~\u2_R3_reg[6]/NET0131  & n21762 ;
  assign n21765 = ~n21763 & ~n21764 ;
  assign n21766 = ~n21759 & ~n21765 ;
  assign n21767 = decrypt_pad & ~\u2_uk_K_r3_reg[17]/NET0131  ;
  assign n21768 = ~decrypt_pad & ~\u2_uk_K_r3_reg[40]/NET0131  ;
  assign n21769 = ~n21767 & ~n21768 ;
  assign n21770 = \u2_R3_reg[7]/NET0131  & ~n21769 ;
  assign n21771 = ~\u2_R3_reg[7]/NET0131  & n21769 ;
  assign n21772 = ~n21770 & ~n21771 ;
  assign n21773 = ~n21743 & n21765 ;
  assign n21774 = n21749 & n21757 ;
  assign n21775 = n21773 & n21774 ;
  assign n21776 = n21772 & n21775 ;
  assign n21790 = ~n21766 & ~n21776 ;
  assign n21777 = n21757 & n21765 ;
  assign n21778 = ~n21751 & n21777 ;
  assign n21779 = ~n21758 & ~n21778 ;
  assign n21780 = ~n21772 & ~n21779 ;
  assign n21784 = n21743 & ~n21765 ;
  assign n21785 = ~n21765 & n21772 ;
  assign n21786 = ~n21784 & ~n21785 ;
  assign n21781 = n21749 & ~n21757 ;
  assign n21782 = n21743 & ~n21781 ;
  assign n21783 = ~n21749 & ~n21765 ;
  assign n21787 = ~n21773 & ~n21783 ;
  assign n21788 = ~n21782 & n21787 ;
  assign n21789 = n21786 & n21788 ;
  assign n21791 = ~n21780 & ~n21789 ;
  assign n21792 = n21790 & n21791 ;
  assign n21793 = ~n21737 & ~n21792 ;
  assign n21806 = ~n21749 & ~n21757 ;
  assign n21810 = ~n21775 & ~n21806 ;
  assign n21811 = n21737 & ~n21810 ;
  assign n21812 = ~n21773 & n21781 ;
  assign n21813 = ~n21811 & ~n21812 ;
  assign n21814 = ~n21772 & ~n21784 ;
  assign n21815 = ~n21813 & n21814 ;
  assign n21800 = ~n21765 & n21774 ;
  assign n21801 = n21743 & n21800 ;
  assign n21794 = ~n21749 & n21757 ;
  assign n21795 = ~n21743 & n21794 ;
  assign n21796 = ~n21765 & n21795 ;
  assign n21797 = ~n21757 & n21765 ;
  assign n21798 = n21743 & n21772 ;
  assign n21799 = ~n21797 & n21798 ;
  assign n21802 = ~n21796 & ~n21799 ;
  assign n21803 = ~n21801 & n21802 ;
  assign n21804 = n21737 & ~n21803 ;
  assign n21807 = ~n21784 & ~n21806 ;
  assign n21805 = ~n21757 & ~n21773 ;
  assign n21808 = n21772 & ~n21805 ;
  assign n21809 = ~n21807 & n21808 ;
  assign n21816 = ~n21804 & ~n21809 ;
  assign n21817 = ~n21815 & n21816 ;
  assign n21818 = ~n21793 & n21817 ;
  assign n21819 = \u2_L3_reg[2]/NET0131  & n21818 ;
  assign n21820 = ~\u2_L3_reg[2]/NET0131  & ~n21818 ;
  assign n21821 = ~n21819 & ~n21820 ;
  assign n21825 = n21060 & n21124 ;
  assign n21826 = ~n21109 & ~n21825 ;
  assign n21827 = ~n21116 & n21826 ;
  assign n21828 = n21048 & ~n21827 ;
  assign n21822 = n21073 & n21101 ;
  assign n21823 = ~n21683 & ~n21822 ;
  assign n21824 = ~n21048 & ~n21823 ;
  assign n21829 = n21078 & n21083 ;
  assign n21830 = ~n21075 & ~n21829 ;
  assign n21831 = ~n21824 & n21830 ;
  assign n21832 = ~n21828 & n21831 ;
  assign n21833 = ~n21099 & ~n21832 ;
  assign n21837 = n21048 & n21078 ;
  assign n21838 = ~n21822 & ~n21837 ;
  assign n21839 = ~n21067 & ~n21838 ;
  assign n21834 = ~n21060 & n21103 ;
  assign n21835 = ~n21124 & ~n21834 ;
  assign n21836 = ~n21048 & ~n21835 ;
  assign n21840 = n21067 & n21087 ;
  assign n21841 = ~n21836 & ~n21840 ;
  assign n21842 = ~n21839 & n21841 ;
  assign n21843 = n21099 & ~n21842 ;
  assign n21844 = n21067 & n21676 ;
  assign n21845 = ~n21048 & ~n21102 ;
  assign n21846 = ~n21844 & n21845 ;
  assign n21847 = ~n21088 & ~n21107 ;
  assign n21848 = ~n21109 & n21847 ;
  assign n21849 = n21048 & n21067 ;
  assign n21850 = ~n21848 & n21849 ;
  assign n21851 = ~n21846 & ~n21850 ;
  assign n21852 = ~n21843 & n21851 ;
  assign n21853 = ~n21833 & n21852 ;
  assign n21854 = ~\u2_L3_reg[4]/NET0131  & ~n21853 ;
  assign n21855 = \u2_L3_reg[4]/NET0131  & n21853 ;
  assign n21856 = ~n21854 & ~n21855 ;
  assign n21857 = n21750 & n21777 ;
  assign n21858 = ~n21801 & ~n21857 ;
  assign n21859 = n21758 & n21765 ;
  assign n21860 = n21750 & ~n21757 ;
  assign n21861 = ~n21796 & ~n21860 ;
  assign n21862 = ~n21859 & n21861 ;
  assign n21863 = ~n21737 & ~n21862 ;
  assign n21864 = n21858 & ~n21863 ;
  assign n21865 = ~n21772 & ~n21864 ;
  assign n21869 = ~n21743 & ~n21781 ;
  assign n21870 = ~n21794 & ~n21869 ;
  assign n21871 = ~n21784 & n21794 ;
  assign n21872 = n21772 & ~n21871 ;
  assign n21873 = ~n21870 & n21872 ;
  assign n21867 = ~n21750 & n21772 ;
  assign n21868 = n21777 & n21867 ;
  assign n21866 = n21781 & ~n21786 ;
  assign n21874 = ~n21737 & ~n21866 ;
  assign n21875 = ~n21868 & n21874 ;
  assign n21876 = ~n21873 & n21875 ;
  assign n21883 = ~n21765 & n21860 ;
  assign n21884 = n21737 & ~n21883 ;
  assign n21885 = ~n21789 & n21884 ;
  assign n21881 = ~n21783 & n21869 ;
  assign n21882 = ~n21772 & n21881 ;
  assign n21877 = ~n21743 & n21783 ;
  assign n21878 = n21765 & n21781 ;
  assign n21879 = ~n21877 & ~n21878 ;
  assign n21880 = n21772 & ~n21879 ;
  assign n21886 = n21858 & ~n21880 ;
  assign n21887 = ~n21882 & n21886 ;
  assign n21888 = n21885 & n21887 ;
  assign n21889 = ~n21876 & ~n21888 ;
  assign n21890 = ~n21865 & ~n21889 ;
  assign n21891 = ~\u2_L3_reg[13]/NET0131  & n21890 ;
  assign n21892 = \u2_L3_reg[13]/NET0131  & ~n21890 ;
  assign n21893 = ~n21891 & ~n21892 ;
  assign n21894 = ~n21048 & n21054 ;
  assign n21895 = ~n21825 & ~n21894 ;
  assign n21896 = ~n21073 & ~n21895 ;
  assign n21900 = n21099 & ~n21834 ;
  assign n21901 = ~n21896 & n21900 ;
  assign n21897 = n21067 & ~n21847 ;
  assign n21898 = ~n21112 & ~n21119 ;
  assign n21899 = n21048 & ~n21898 ;
  assign n21902 = ~n21897 & ~n21899 ;
  assign n21903 = n21901 & n21902 ;
  assign n21906 = n21054 & ~n21103 ;
  assign n21907 = ~n21822 & ~n21906 ;
  assign n21908 = n21048 & ~n21907 ;
  assign n21905 = ~n21048 & ~n21847 ;
  assign n21904 = n21067 & n21079 ;
  assign n21909 = ~n21099 & ~n21904 ;
  assign n21910 = ~n21905 & n21909 ;
  assign n21911 = ~n21908 & n21910 ;
  assign n21912 = ~n21903 & ~n21911 ;
  assign n21913 = ~n21073 & n21829 ;
  assign n21914 = ~n21115 & ~n21913 ;
  assign n21915 = ~n21912 & n21914 ;
  assign n21916 = ~\u2_L3_reg[19]/NET0131  & ~n21915 ;
  assign n21917 = \u2_L3_reg[19]/NET0131  & n21915 ;
  assign n21918 = ~n21916 & ~n21917 ;
  assign n21940 = n20962 & n20993 ;
  assign n21941 = ~n20977 & ~n21940 ;
  assign n21942 = n20983 & ~n21941 ;
  assign n21939 = n21010 & n21024 ;
  assign n21943 = ~n21507 & ~n21939 ;
  assign n21944 = ~n21942 & n21943 ;
  assign n21945 = n20950 & ~n21944 ;
  assign n21935 = ~n20962 & n21490 ;
  assign n21936 = ~n21029 & ~n21505 ;
  assign n21937 = ~n21935 & n21936 ;
  assign n21938 = ~n20983 & ~n21937 ;
  assign n21921 = ~n20969 & n21002 ;
  assign n21924 = ~n20995 & ~n21028 ;
  assign n21925 = ~n21921 & n21924 ;
  assign n21919 = n20962 & n20996 ;
  assign n21920 = n20983 & n21919 ;
  assign n21922 = ~n20985 & ~n21002 ;
  assign n21923 = n21015 & n21922 ;
  assign n21926 = ~n21920 & ~n21923 ;
  assign n21927 = n21925 & n21926 ;
  assign n21928 = ~n20950 & ~n21927 ;
  assign n21929 = ~n21013 & ~n21919 ;
  assign n21930 = n21001 & ~n21929 ;
  assign n21931 = ~n21032 & ~n21919 ;
  assign n21932 = ~n20987 & n21931 ;
  assign n21933 = n20950 & ~n20983 ;
  assign n21934 = ~n21932 & n21933 ;
  assign n21946 = ~n21930 & ~n21934 ;
  assign n21947 = ~n21928 & n21946 ;
  assign n21948 = ~n21938 & n21947 ;
  assign n21949 = ~n21945 & n21948 ;
  assign n21950 = \u2_L3_reg[23]/NET0131  & ~n21949 ;
  assign n21951 = ~\u2_L3_reg[23]/NET0131  & n21949 ;
  assign n21952 = ~n21950 & ~n21951 ;
  assign n21966 = ~n21260 & ~n21310 ;
  assign n21967 = n21270 & n21966 ;
  assign n21968 = n21293 & n21593 ;
  assign n21969 = n21269 & ~n21603 ;
  assign n21970 = ~n21968 & n21969 ;
  assign n21971 = ~n21967 & ~n21970 ;
  assign n21972 = ~n21261 & ~n21611 ;
  assign n21973 = ~n21288 & n21972 ;
  assign n21974 = ~n21971 & n21973 ;
  assign n21975 = n21284 & ~n21974 ;
  assign n21955 = n21269 & ~n21298 ;
  assign n21954 = n21246 & ~n21593 ;
  assign n21956 = ~n21312 & ~n21954 ;
  assign n21957 = n21955 & n21956 ;
  assign n21953 = n21316 & n21589 ;
  assign n21958 = ~n21592 & ~n21953 ;
  assign n21959 = ~n21318 & n21958 ;
  assign n21960 = ~n21957 & n21959 ;
  assign n21961 = ~n21284 & ~n21960 ;
  assign n21964 = ~n21313 & ~n21317 ;
  assign n21965 = ~n21269 & ~n21964 ;
  assign n21962 = ~n21246 & n21269 ;
  assign n21963 = n21286 & n21962 ;
  assign n21976 = ~n21311 & ~n21963 ;
  assign n21977 = ~n21965 & n21976 ;
  assign n21978 = ~n21961 & n21977 ;
  assign n21979 = ~n21975 & n21978 ;
  assign n21980 = ~\u2_L3_reg[27]/NET0131  & ~n21979 ;
  assign n21981 = \u2_L3_reg[27]/NET0131  & n21979 ;
  assign n21982 = ~n21980 & ~n21981 ;
  assign n21985 = n21743 & n21781 ;
  assign n21986 = ~n21765 & n21806 ;
  assign n21987 = ~n21985 & ~n21986 ;
  assign n21988 = n21772 & n21987 ;
  assign n21992 = n21757 & ~n21881 ;
  assign n21989 = ~n21757 & n21773 ;
  assign n21990 = ~n21772 & ~n21857 ;
  assign n21991 = ~n21989 & n21990 ;
  assign n21993 = ~n21758 & n21991 ;
  assign n21994 = ~n21992 & n21993 ;
  assign n21995 = ~n21988 & ~n21994 ;
  assign n21983 = n21765 & ~n21795 ;
  assign n21984 = ~n21870 & n21983 ;
  assign n21996 = ~n21737 & ~n21984 ;
  assign n21997 = ~n21995 & n21996 ;
  assign n22001 = n21987 & n21991 ;
  assign n22002 = ~n21749 & ~n21797 ;
  assign n22003 = n21782 & ~n22002 ;
  assign n22004 = n21772 & ~n21795 ;
  assign n22005 = ~n22003 & n22004 ;
  assign n22006 = ~n22001 & ~n22005 ;
  assign n21998 = ~n21751 & ~n21772 ;
  assign n21999 = n21757 & ~n21765 ;
  assign n22000 = ~n21998 & n21999 ;
  assign n22007 = n21737 & ~n21859 ;
  assign n22008 = ~n22000 & n22007 ;
  assign n22009 = ~n22006 & n22008 ;
  assign n22010 = ~n21997 & ~n22009 ;
  assign n22011 = ~\u2_L3_reg[28]/NET0131  & n22010 ;
  assign n22012 = \u2_L3_reg[28]/NET0131  & ~n22010 ;
  assign n22013 = ~n22011 & ~n22012 ;
  assign n22029 = n20884 & n20930 ;
  assign n22030 = ~n20887 & ~n20923 ;
  assign n22031 = ~n20883 & ~n22030 ;
  assign n22032 = ~n20864 & n20899 ;
  assign n22033 = n20858 & ~n22032 ;
  assign n22034 = ~n22031 & n22033 ;
  assign n22035 = ~n20890 & ~n20925 ;
  assign n22036 = n20896 & n22035 ;
  assign n22037 = ~n20858 & ~n21365 ;
  assign n22038 = ~n21367 & n22037 ;
  assign n22039 = ~n22036 & n22038 ;
  assign n22040 = ~n22034 & ~n22039 ;
  assign n22041 = ~n22029 & ~n22040 ;
  assign n22042 = n20908 & ~n22041 ;
  assign n22018 = n20887 & n20899 ;
  assign n22020 = n20920 & n21378 ;
  assign n22021 = ~n22018 & ~n22020 ;
  assign n22022 = n20915 & n22021 ;
  assign n22014 = ~n20870 & n20925 ;
  assign n22015 = n20877 & n20920 ;
  assign n22016 = ~n22014 & ~n22015 ;
  assign n22017 = n20858 & ~n22016 ;
  assign n22019 = n21364 & ~n22015 ;
  assign n22023 = ~n22017 & ~n22019 ;
  assign n22024 = n22022 & n22023 ;
  assign n22025 = ~n20908 & ~n22024 ;
  assign n22026 = n20858 & n20913 ;
  assign n22027 = ~n20884 & n20910 ;
  assign n22028 = n20888 & n22027 ;
  assign n22043 = ~n22026 & ~n22028 ;
  assign n22044 = ~n22025 & n22043 ;
  assign n22045 = ~n22042 & n22044 ;
  assign n22046 = \u2_L3_reg[32]/NET0131  & n22045 ;
  assign n22047 = ~\u2_L3_reg[32]/NET0131  & ~n22045 ;
  assign n22048 = ~n22046 & ~n22047 ;
  assign n22082 = decrypt_pad & ~\u2_uk_K_r3_reg[18]/NET0131  ;
  assign n22083 = ~decrypt_pad & ~\u2_uk_K_r3_reg[41]/NET0131  ;
  assign n22084 = ~n22082 & ~n22083 ;
  assign n22085 = \u2_R3_reg[12]/NET0131  & ~n22084 ;
  assign n22086 = ~\u2_R3_reg[12]/NET0131  & n22084 ;
  assign n22087 = ~n22085 & ~n22086 ;
  assign n22049 = decrypt_pad & ~\u2_uk_K_r3_reg[6]/NET0131  ;
  assign n22050 = ~decrypt_pad & ~\u2_uk_K_r3_reg[54]/NET0131  ;
  assign n22051 = ~n22049 & ~n22050 ;
  assign n22052 = \u2_R3_reg[13]/NET0131  & ~n22051 ;
  assign n22053 = ~\u2_R3_reg[13]/NET0131  & n22051 ;
  assign n22054 = ~n22052 & ~n22053 ;
  assign n22062 = decrypt_pad & ~\u2_uk_K_r3_reg[54]/NET0131  ;
  assign n22063 = ~decrypt_pad & ~\u2_uk_K_r3_reg[20]/NET0131  ;
  assign n22064 = ~n22062 & ~n22063 ;
  assign n22065 = \u2_R3_reg[8]/NET0131  & ~n22064 ;
  assign n22066 = ~\u2_R3_reg[8]/NET0131  & n22064 ;
  assign n22067 = ~n22065 & ~n22066 ;
  assign n22069 = ~n22054 & ~n22067 ;
  assign n22070 = n22054 & n22067 ;
  assign n22071 = ~n22069 & ~n22070 ;
  assign n22055 = decrypt_pad & ~\u2_uk_K_r3_reg[26]/NET0131  ;
  assign n22056 = ~decrypt_pad & ~\u2_uk_K_r3_reg[17]/NET0131  ;
  assign n22057 = ~n22055 & ~n22056 ;
  assign n22058 = \u2_R3_reg[9]/NET0131  & ~n22057 ;
  assign n22059 = ~\u2_R3_reg[9]/NET0131  & n22057 ;
  assign n22060 = ~n22058 & ~n22059 ;
  assign n22072 = decrypt_pad & ~\u2_uk_K_r3_reg[34]/NET0131  ;
  assign n22073 = ~decrypt_pad & ~\u2_uk_K_r3_reg[25]/NET0131  ;
  assign n22074 = ~n22072 & ~n22073 ;
  assign n22075 = \u2_R3_reg[10]/NET0131  & ~n22074 ;
  assign n22076 = ~\u2_R3_reg[10]/NET0131  & n22074 ;
  assign n22077 = ~n22075 & ~n22076 ;
  assign n22123 = ~n22060 & n22077 ;
  assign n22124 = ~n22071 & n22123 ;
  assign n22112 = n22054 & ~n22067 ;
  assign n22113 = n22060 & n22112 ;
  assign n22094 = decrypt_pad & ~\u2_uk_K_r3_reg[3]/NET0131  ;
  assign n22095 = ~decrypt_pad & ~\u2_uk_K_r3_reg[26]/NET0131  ;
  assign n22096 = ~n22094 & ~n22095 ;
  assign n22097 = \u2_R3_reg[11]/P0001  & ~n22096 ;
  assign n22098 = ~\u2_R3_reg[11]/P0001  & n22096 ;
  assign n22099 = ~n22097 & ~n22098 ;
  assign n22114 = n22077 & ~n22099 ;
  assign n22115 = n22113 & n22114 ;
  assign n22120 = ~n22054 & n22060 ;
  assign n22121 = n22077 & n22120 ;
  assign n22122 = n22067 & n22121 ;
  assign n22125 = ~n22115 & ~n22122 ;
  assign n22126 = ~n22124 & n22125 ;
  assign n22105 = n22060 & ~n22077 ;
  assign n22116 = n22054 & n22099 ;
  assign n22117 = n22071 & ~n22116 ;
  assign n22118 = n22105 & ~n22117 ;
  assign n22089 = ~n22060 & ~n22077 ;
  assign n22119 = n22089 & n22117 ;
  assign n22127 = ~n22118 & ~n22119 ;
  assign n22128 = n22126 & n22127 ;
  assign n22129 = ~n22087 & ~n22128 ;
  assign n22061 = n22054 & ~n22060 ;
  assign n22068 = ~n22060 & n22067 ;
  assign n22078 = ~n22067 & ~n22077 ;
  assign n22079 = ~n22068 & ~n22078 ;
  assign n22080 = n22071 & n22079 ;
  assign n22081 = ~n22061 & ~n22080 ;
  assign n22088 = ~n22081 & n22087 ;
  assign n22090 = n22069 & n22089 ;
  assign n22091 = n22061 & n22077 ;
  assign n22092 = ~n22090 & ~n22091 ;
  assign n22093 = ~n22088 & n22092 ;
  assign n22100 = ~n22093 & n22099 ;
  assign n22101 = n22077 & n22087 ;
  assign n22102 = n22060 & n22069 ;
  assign n22103 = n22101 & n22102 ;
  assign n22104 = n22087 & ~n22099 ;
  assign n22106 = n22054 & n22105 ;
  assign n22107 = ~n22054 & n22068 ;
  assign n22108 = n22060 & n22070 ;
  assign n22109 = ~n22107 & ~n22108 ;
  assign n22110 = ~n22106 & n22109 ;
  assign n22111 = n22104 & ~n22110 ;
  assign n22130 = ~n22103 & ~n22111 ;
  assign n22131 = ~n22100 & n22130 ;
  assign n22132 = ~n22129 & n22131 ;
  assign n22133 = ~\u2_L3_reg[6]/NET0131  & ~n22132 ;
  assign n22134 = \u2_L3_reg[6]/NET0131  & n22132 ;
  assign n22135 = ~n22133 & ~n22134 ;
  assign n22137 = ~n20930 & n22035 ;
  assign n22136 = n20858 & ~n20908 ;
  assign n22138 = ~n20891 & n22136 ;
  assign n22139 = ~n22018 & n22138 ;
  assign n22140 = ~n22137 & n22139 ;
  assign n22142 = ~n20864 & ~n20916 ;
  assign n22143 = ~n22035 & ~n22142 ;
  assign n22144 = ~n22137 & ~n22143 ;
  assign n22141 = ~n20858 & n20908 ;
  assign n22145 = ~n22136 & ~n22141 ;
  assign n22146 = ~n21365 & n22145 ;
  assign n22147 = ~n22144 & n22146 ;
  assign n22148 = ~n22140 & ~n22147 ;
  assign n22149 = ~n20892 & ~n22148 ;
  assign n22152 = n20870 & n22035 ;
  assign n22151 = ~n20877 & ~n20931 ;
  assign n22150 = n20887 & ~n20899 ;
  assign n22153 = n22141 & ~n22150 ;
  assign n22154 = ~n22151 & n22153 ;
  assign n22155 = ~n22152 & n22154 ;
  assign n22156 = ~n22149 & ~n22155 ;
  assign n22157 = ~\u2_L3_reg[7]/NET0131  & n22156 ;
  assign n22158 = \u2_L3_reg[7]/NET0131  & ~n22156 ;
  assign n22159 = ~n22157 & ~n22158 ;
  assign n22171 = ~n21435 & ~n21694 ;
  assign n22172 = n21396 & ~n22171 ;
  assign n22173 = n21432 & ~n21457 ;
  assign n22174 = ~n21700 & ~n22173 ;
  assign n22175 = ~n21396 & ~n22174 ;
  assign n22176 = ~n21416 & n21719 ;
  assign n22177 = ~n22175 & n22176 ;
  assign n22178 = ~n22172 & n22177 ;
  assign n22179 = ~n21455 & ~n22178 ;
  assign n22164 = ~n21402 & n21465 ;
  assign n22165 = ~n21700 & ~n22164 ;
  assign n22166 = n21396 & ~n22165 ;
  assign n22167 = ~n21402 & n21723 ;
  assign n22168 = n21482 & ~n22167 ;
  assign n22169 = ~n22166 & n22168 ;
  assign n22170 = n21455 & ~n22169 ;
  assign n22160 = n21432 & ~n21458 ;
  assign n22161 = ~n21431 & ~n22160 ;
  assign n22162 = n21396 & ~n22161 ;
  assign n22163 = n21402 & n21708 ;
  assign n22180 = ~n22162 & ~n22163 ;
  assign n22181 = ~n22170 & n22180 ;
  assign n22182 = ~n22179 & n22181 ;
  assign n22183 = ~\u2_L3_reg[8]/NET0131  & ~n22182 ;
  assign n22184 = \u2_L3_reg[8]/NET0131  & n22182 ;
  assign n22185 = ~n22183 & ~n22184 ;
  assign n22186 = n22077 & ~n22113 ;
  assign n22188 = n22099 & n22102 ;
  assign n22187 = n22061 & ~n22067 ;
  assign n22189 = ~n22077 & ~n22187 ;
  assign n22190 = n22109 & n22189 ;
  assign n22191 = ~n22188 & n22190 ;
  assign n22192 = ~n22186 & ~n22191 ;
  assign n22193 = n22069 & n22077 ;
  assign n22194 = ~n22060 & n22193 ;
  assign n22195 = n22099 & ~n22122 ;
  assign n22196 = ~n22194 & n22195 ;
  assign n22197 = n22067 & n22077 ;
  assign n22198 = ~n22054 & ~n22078 ;
  assign n22199 = ~n22197 & n22198 ;
  assign n22200 = ~n22196 & n22199 ;
  assign n22201 = ~n22192 & ~n22200 ;
  assign n22202 = n22087 & ~n22201 ;
  assign n22203 = ~n22060 & n22197 ;
  assign n22204 = ~n22099 & ~n22203 ;
  assign n22205 = ~n22196 & ~n22204 ;
  assign n22210 = n22069 & ~n22077 ;
  assign n22211 = ~n22108 & ~n22187 ;
  assign n22212 = ~n22210 & n22211 ;
  assign n22213 = ~n22099 & ~n22212 ;
  assign n22207 = ~n22069 & n22099 ;
  assign n22206 = ~n22060 & ~n22070 ;
  assign n22208 = ~n22108 & ~n22206 ;
  assign n22209 = n22207 & n22208 ;
  assign n22214 = ~n22090 & ~n22209 ;
  assign n22215 = ~n22213 & n22214 ;
  assign n22216 = ~n22087 & ~n22215 ;
  assign n22217 = ~n22205 & ~n22216 ;
  assign n22218 = ~n22202 & n22217 ;
  assign n22219 = ~\u2_L3_reg[16]/NET0131  & ~n22218 ;
  assign n22220 = \u2_L3_reg[16]/NET0131  & n22218 ;
  assign n22221 = ~n22219 & ~n22220 ;
  assign n22231 = ~n22077 & n22099 ;
  assign n22242 = ~n22060 & ~n22112 ;
  assign n22243 = n22231 & n22242 ;
  assign n22238 = ~n22089 & ~n22099 ;
  assign n22239 = ~n22071 & n22238 ;
  assign n22240 = ~n22068 & n22077 ;
  assign n22241 = n22207 & n22240 ;
  assign n22244 = ~n22239 & ~n22241 ;
  assign n22245 = ~n22243 & n22244 ;
  assign n22246 = ~n22119 & n22245 ;
  assign n22247 = n22087 & ~n22246 ;
  assign n22222 = n22054 & n22078 ;
  assign n22223 = ~n22193 & ~n22222 ;
  assign n22224 = ~n22102 & ~n22203 ;
  assign n22225 = n22223 & n22224 ;
  assign n22226 = n22099 & ~n22225 ;
  assign n22227 = ~n22054 & n22203 ;
  assign n22228 = ~n22226 & ~n22227 ;
  assign n22229 = ~n22087 & ~n22228 ;
  assign n22234 = ~n22071 & n22089 ;
  assign n22235 = ~n22080 & ~n22234 ;
  assign n22236 = ~n22087 & ~n22099 ;
  assign n22237 = ~n22235 & n22236 ;
  assign n22230 = n22108 & n22114 ;
  assign n22232 = ~n22107 & ~n22113 ;
  assign n22233 = n22231 & ~n22232 ;
  assign n22248 = ~n22230 & ~n22233 ;
  assign n22249 = ~n22237 & n22248 ;
  assign n22250 = ~n22229 & n22249 ;
  assign n22251 = ~n22247 & n22250 ;
  assign n22252 = ~\u2_L3_reg[24]/NET0131  & ~n22251 ;
  assign n22253 = \u2_L3_reg[24]/NET0131  & n22251 ;
  assign n22254 = ~n22252 & ~n22253 ;
  assign n22256 = ~n22077 & n22107 ;
  assign n22257 = n22223 & ~n22256 ;
  assign n22258 = n22087 & ~n22257 ;
  assign n22259 = ~n22120 & ~n22197 ;
  assign n22260 = ~n22087 & ~n22121 ;
  assign n22261 = ~n22259 & n22260 ;
  assign n22262 = ~n22258 & ~n22261 ;
  assign n22263 = n22099 & ~n22262 ;
  assign n22267 = n22077 & n22187 ;
  assign n22264 = ~n22060 & ~n22067 ;
  assign n22265 = ~n22099 & ~n22264 ;
  assign n22266 = n22259 & n22265 ;
  assign n22268 = ~n22234 & ~n22266 ;
  assign n22269 = ~n22267 & n22268 ;
  assign n22270 = ~n22087 & ~n22269 ;
  assign n22271 = ~n22102 & ~n22197 ;
  assign n22272 = n22104 & ~n22271 ;
  assign n22274 = n22060 & ~n22070 ;
  assign n22275 = n22101 & n22274 ;
  assign n22255 = n22114 & n22120 ;
  assign n22273 = n22116 & n22203 ;
  assign n22276 = ~n22255 & ~n22273 ;
  assign n22277 = ~n22275 & n22276 ;
  assign n22278 = ~n22272 & n22277 ;
  assign n22279 = ~n22270 & n22278 ;
  assign n22280 = ~n22263 & n22279 ;
  assign n22281 = \u2_L3_reg[30]/NET0131  & ~n22280 ;
  assign n22282 = ~\u2_L3_reg[30]/NET0131  & n22280 ;
  assign n22283 = ~n22281 & ~n22282 ;
  assign n22287 = ~n21402 & n21432 ;
  assign n22288 = ~n21461 & ~n22287 ;
  assign n22289 = n21396 & ~n22288 ;
  assign n22284 = n21396 & ~n21457 ;
  assign n22285 = ~n21443 & ~n21700 ;
  assign n22286 = ~n22284 & ~n22285 ;
  assign n22290 = ~n21455 & ~n22286 ;
  assign n22291 = ~n22289 & n22290 ;
  assign n22294 = n21415 & ~n21442 ;
  assign n22293 = ~n21415 & ~n21426 ;
  assign n22295 = n21396 & ~n22293 ;
  assign n22296 = ~n22294 & n22295 ;
  assign n22297 = ~n21396 & n21464 ;
  assign n22292 = n21402 & n21434 ;
  assign n22298 = ~n21437 & n21455 ;
  assign n22299 = ~n22292 & n22298 ;
  assign n22300 = ~n22297 & n22299 ;
  assign n22301 = ~n22296 & n22300 ;
  assign n22302 = ~n22291 & ~n22301 ;
  assign n22303 = n21436 & n21457 ;
  assign n22304 = ~n21396 & ~n22303 ;
  assign n22305 = ~n21477 & n22304 ;
  assign n22306 = ~n22164 & n22305 ;
  assign n22307 = n21396 & ~n21435 ;
  assign n22308 = ~n21480 & n22307 ;
  assign n22309 = ~n22306 & ~n22308 ;
  assign n22310 = ~n22302 & ~n22309 ;
  assign n22311 = ~\u2_L3_reg[3]/NET0131  & ~n22310 ;
  assign n22312 = \u2_L3_reg[3]/NET0131  & n22310 ;
  assign n22313 = ~n22311 & ~n22312 ;
  assign n22328 = n21494 & n21931 ;
  assign n22329 = n20956 & ~n22328 ;
  assign n22319 = ~n20985 & ~n21940 ;
  assign n22330 = n21001 & ~n22319 ;
  assign n22331 = ~n21505 & ~n22330 ;
  assign n22332 = ~n22329 & n22331 ;
  assign n22333 = n20950 & ~n22332 ;
  assign n22314 = ~n20956 & n21493 ;
  assign n22315 = n20956 & n21940 ;
  assign n22316 = ~n22314 & ~n22315 ;
  assign n22317 = ~n20983 & ~n22316 ;
  assign n22320 = ~n20983 & n22319 ;
  assign n22321 = n20983 & ~n20988 ;
  assign n22322 = ~n20970 & n22321 ;
  assign n22323 = ~n21919 & n22322 ;
  assign n22324 = ~n22320 & ~n22323 ;
  assign n22318 = n21014 & ~n21498 ;
  assign n22325 = ~n22314 & ~n22318 ;
  assign n22326 = ~n22324 & n22325 ;
  assign n22327 = ~n20950 & ~n22326 ;
  assign n22334 = ~n22317 & ~n22327 ;
  assign n22335 = ~n22333 & n22334 ;
  assign n22336 = ~\u2_L3_reg[9]/NET0131  & ~n22335 ;
  assign n22337 = \u2_L3_reg[9]/NET0131  & n22335 ;
  assign n22338 = ~n22336 & ~n22337 ;
  assign n22342 = ~n21795 & ~n21800 ;
  assign n22343 = ~n21772 & ~n22342 ;
  assign n22340 = n21773 & n21806 ;
  assign n22341 = ~n21759 & n21772 ;
  assign n22344 = ~n22340 & ~n22341 ;
  assign n22345 = ~n22343 & n22344 ;
  assign n22346 = n21737 & ~n22345 ;
  assign n22348 = ~n21784 & ~n21798 ;
  assign n22349 = n21805 & n22348 ;
  assign n22350 = ~n21775 & ~n21857 ;
  assign n22347 = n21774 & n21798 ;
  assign n22351 = ~n21877 & ~n22347 ;
  assign n22352 = n22350 & n22351 ;
  assign n22353 = ~n22349 & n22352 ;
  assign n22354 = ~n21737 & ~n22353 ;
  assign n22339 = ~n21772 & n21985 ;
  assign n22355 = n21749 & n21777 ;
  assign n22356 = ~n21883 & ~n22355 ;
  assign n22357 = n21772 & ~n22356 ;
  assign n22358 = ~n22339 & ~n22357 ;
  assign n22359 = ~n22354 & n22358 ;
  assign n22360 = ~n22346 & n22359 ;
  assign n22361 = ~\u2_L3_reg[18]/P0001  & ~n22360 ;
  assign n22362 = \u2_L3_reg[18]/P0001  & n22360 ;
  assign n22363 = ~n22361 & ~n22362 ;
  assign n22364 = decrypt_pad & ~\u2_uk_K_r2_reg[26]/NET0131  ;
  assign n22365 = ~decrypt_pad & ~\u2_uk_K_r2_reg[46]/NET0131  ;
  assign n22366 = ~n22364 & ~n22365 ;
  assign n22367 = \u2_R2_reg[1]/NET0131  & ~n22366 ;
  assign n22368 = ~\u2_R2_reg[1]/NET0131  & n22366 ;
  assign n22369 = ~n22367 & ~n22368 ;
  assign n22370 = decrypt_pad & ~\u2_uk_K_r2_reg[24]/NET0131  ;
  assign n22371 = ~decrypt_pad & ~\u2_uk_K_r2_reg[19]/NET0131  ;
  assign n22372 = ~n22370 & ~n22371 ;
  assign n22373 = \u2_R2_reg[5]/NET0131  & ~n22372 ;
  assign n22374 = ~\u2_R2_reg[5]/NET0131  & n22372 ;
  assign n22375 = ~n22373 & ~n22374 ;
  assign n22376 = ~n22369 & n22375 ;
  assign n22377 = decrypt_pad & ~\u2_uk_K_r2_reg[41]/NET0131  ;
  assign n22378 = ~decrypt_pad & ~\u2_uk_K_r2_reg[4]/NET0131  ;
  assign n22379 = ~n22377 & ~n22378 ;
  assign n22380 = \u2_R2_reg[2]/NET0131  & ~n22379 ;
  assign n22381 = ~\u2_R2_reg[2]/NET0131  & n22379 ;
  assign n22382 = ~n22380 & ~n22381 ;
  assign n22383 = ~n22375 & n22382 ;
  assign n22384 = n22375 & ~n22382 ;
  assign n22385 = ~n22383 & ~n22384 ;
  assign n22386 = decrypt_pad & ~\u2_uk_K_r2_reg[5]/NET0131  ;
  assign n22387 = ~decrypt_pad & ~\u2_uk_K_r2_reg[25]/NET0131  ;
  assign n22388 = ~n22386 & ~n22387 ;
  assign n22389 = \u2_R2_reg[32]/NET0131  & ~n22388 ;
  assign n22390 = ~\u2_R2_reg[32]/NET0131  & n22388 ;
  assign n22391 = ~n22389 & ~n22390 ;
  assign n22392 = ~n22385 & ~n22391 ;
  assign n22393 = ~n22376 & ~n22392 ;
  assign n22394 = decrypt_pad & ~\u2_uk_K_r2_reg[18]/NET0131  ;
  assign n22395 = ~decrypt_pad & ~\u2_uk_K_r2_reg[13]/NET0131  ;
  assign n22396 = ~n22394 & ~n22395 ;
  assign n22397 = \u2_R2_reg[3]/NET0131  & ~n22396 ;
  assign n22398 = ~\u2_R2_reg[3]/NET0131  & n22396 ;
  assign n22399 = ~n22397 & ~n22398 ;
  assign n22400 = ~n22393 & n22399 ;
  assign n22406 = ~n22369 & n22391 ;
  assign n22407 = ~n22369 & n22382 ;
  assign n22408 = n22391 & ~n22399 ;
  assign n22409 = ~n22407 & ~n22408 ;
  assign n22410 = ~n22406 & ~n22409 ;
  assign n22401 = ~n22375 & ~n22391 ;
  assign n22402 = n22375 & n22391 ;
  assign n22403 = ~n22401 & ~n22402 ;
  assign n22404 = ~n22369 & ~n22383 ;
  assign n22405 = n22403 & n22404 ;
  assign n22411 = decrypt_pad & ~\u2_uk_K_r2_reg[53]/P0001  ;
  assign n22412 = ~decrypt_pad & ~\u2_uk_K_r2_reg[48]/NET0131  ;
  assign n22413 = ~n22411 & ~n22412 ;
  assign n22414 = \u2_R2_reg[4]/NET0131  & ~n22413 ;
  assign n22415 = ~\u2_R2_reg[4]/NET0131  & n22413 ;
  assign n22416 = ~n22414 & ~n22415 ;
  assign n22417 = ~n22405 & n22416 ;
  assign n22418 = ~n22410 & n22417 ;
  assign n22419 = ~n22400 & n22418 ;
  assign n22427 = n22382 & n22399 ;
  assign n22428 = ~n22391 & n22427 ;
  assign n22429 = n22375 & n22428 ;
  assign n22424 = ~n22382 & n22401 ;
  assign n22425 = n22383 & n22391 ;
  assign n22426 = n22399 & n22425 ;
  assign n22430 = ~n22424 & ~n22426 ;
  assign n22431 = ~n22429 & n22430 ;
  assign n22432 = n22369 & ~n22431 ;
  assign n22420 = ~n22382 & n22399 ;
  assign n22421 = ~n22369 & ~n22382 ;
  assign n22422 = ~n22420 & ~n22421 ;
  assign n22423 = n22402 & ~n22422 ;
  assign n22433 = ~n22416 & ~n22423 ;
  assign n22434 = ~n22432 & n22433 ;
  assign n22435 = ~n22419 & ~n22434 ;
  assign n22441 = ~n22382 & ~n22391 ;
  assign n22442 = ~n22376 & n22441 ;
  assign n22443 = n22383 & n22406 ;
  assign n22444 = ~n22442 & ~n22443 ;
  assign n22445 = ~n22416 & ~n22444 ;
  assign n22439 = n22375 & ~n22391 ;
  assign n22440 = n22407 & n22439 ;
  assign n22446 = n22369 & ~n22439 ;
  assign n22447 = n22385 & n22446 ;
  assign n22448 = ~n22440 & ~n22447 ;
  assign n22449 = ~n22445 & n22448 ;
  assign n22450 = ~n22399 & ~n22449 ;
  assign n22436 = ~n22369 & ~n22375 ;
  assign n22437 = n22428 & n22436 ;
  assign n22438 = n22406 & n22420 ;
  assign n22451 = ~n22437 & ~n22438 ;
  assign n22452 = ~n22450 & n22451 ;
  assign n22453 = ~n22435 & n22452 ;
  assign n22454 = ~\u2_L2_reg[31]/NET0131  & ~n22453 ;
  assign n22455 = \u2_L2_reg[31]/NET0131  & n22453 ;
  assign n22456 = ~n22454 & ~n22455 ;
  assign n22508 = decrypt_pad & ~\u2_uk_K_r2_reg[52]/NET0131  ;
  assign n22509 = ~decrypt_pad & ~\u2_uk_K_r2_reg[15]/NET0131  ;
  assign n22510 = ~n22508 & ~n22509 ;
  assign n22511 = \u2_R2_reg[24]/NET0131  & ~n22510 ;
  assign n22512 = ~\u2_R2_reg[24]/NET0131  & n22510 ;
  assign n22513 = ~n22511 & ~n22512 ;
  assign n22463 = decrypt_pad & ~\u2_uk_K_r2_reg[31]/NET0131  ;
  assign n22464 = ~decrypt_pad & ~\u2_uk_K_r2_reg[49]/NET0131  ;
  assign n22465 = ~n22463 & ~n22464 ;
  assign n22466 = \u2_R2_reg[20]/NET0131  & ~n22465 ;
  assign n22467 = ~\u2_R2_reg[20]/NET0131  & n22465 ;
  assign n22468 = ~n22466 & ~n22467 ;
  assign n22476 = decrypt_pad & ~\u2_uk_K_r2_reg[9]/NET0131  ;
  assign n22477 = ~decrypt_pad & ~\u2_uk_K_r2_reg[0]/NET0131  ;
  assign n22478 = ~n22476 & ~n22477 ;
  assign n22479 = \u2_R2_reg[22]/NET0131  & ~n22478 ;
  assign n22480 = ~\u2_R2_reg[22]/NET0131  & n22478 ;
  assign n22481 = ~n22479 & ~n22480 ;
  assign n22482 = decrypt_pad & ~\u2_uk_K_r2_reg[42]/NET0131  ;
  assign n22483 = ~decrypt_pad & ~\u2_uk_K_r2_reg[9]/NET0131  ;
  assign n22484 = ~n22482 & ~n22483 ;
  assign n22485 = \u2_R2_reg[21]/NET0131  & ~n22484 ;
  assign n22486 = ~\u2_R2_reg[21]/NET0131  & n22484 ;
  assign n22487 = ~n22485 & ~n22486 ;
  assign n22517 = ~n22481 & n22487 ;
  assign n22533 = n22468 & n22517 ;
  assign n22457 = decrypt_pad & ~\u2_uk_K_r2_reg[22]/NET0131  ;
  assign n22458 = ~decrypt_pad & ~\u2_uk_K_r2_reg[44]/NET0131  ;
  assign n22459 = ~n22457 & ~n22458 ;
  assign n22460 = \u2_R2_reg[23]/NET0131  & ~n22459 ;
  assign n22461 = ~\u2_R2_reg[23]/NET0131  & n22459 ;
  assign n22462 = ~n22460 & ~n22461 ;
  assign n22490 = ~n22468 & n22487 ;
  assign n22491 = n22481 & n22490 ;
  assign n22534 = ~n22462 & ~n22491 ;
  assign n22535 = ~n22533 & n22534 ;
  assign n22469 = decrypt_pad & ~\u2_uk_K_r2_reg[43]/NET0131  ;
  assign n22470 = ~decrypt_pad & ~\u2_uk_K_r2_reg[38]/NET0131  ;
  assign n22471 = ~n22469 & ~n22470 ;
  assign n22472 = \u2_R2_reg[25]/NET0131  & ~n22471 ;
  assign n22473 = ~\u2_R2_reg[25]/NET0131  & n22471 ;
  assign n22474 = ~n22472 & ~n22473 ;
  assign n22525 = n22474 & ~n22487 ;
  assign n22526 = ~n22468 & n22525 ;
  assign n22527 = n22462 & ~n22526 ;
  assign n22536 = n22481 & ~n22487 ;
  assign n22537 = n22468 & n22536 ;
  assign n22538 = ~n22468 & ~n22481 ;
  assign n22539 = ~n22537 & ~n22538 ;
  assign n22540 = n22527 & n22539 ;
  assign n22541 = ~n22535 & ~n22540 ;
  assign n22492 = n22468 & n22474 ;
  assign n22503 = ~n22487 & n22492 ;
  assign n22530 = n22481 & n22503 ;
  assign n22475 = n22468 & ~n22474 ;
  assign n22497 = ~n22462 & ~n22481 ;
  assign n22531 = ~n22497 & ~n22517 ;
  assign n22532 = n22475 & ~n22531 ;
  assign n22542 = ~n22530 & ~n22532 ;
  assign n22543 = ~n22541 & n22542 ;
  assign n22544 = ~n22513 & ~n22543 ;
  assign n22493 = n22487 & n22492 ;
  assign n22488 = ~n22481 & ~n22487 ;
  assign n22489 = n22475 & n22488 ;
  assign n22494 = ~n22489 & ~n22491 ;
  assign n22495 = ~n22493 & n22494 ;
  assign n22496 = n22462 & ~n22495 ;
  assign n22498 = ~n22490 & ~n22492 ;
  assign n22499 = ~n22462 & n22498 ;
  assign n22500 = ~n22497 & ~n22499 ;
  assign n22501 = n22474 & n22487 ;
  assign n22502 = ~n22468 & n22501 ;
  assign n22504 = ~n22481 & ~n22502 ;
  assign n22505 = ~n22503 & n22504 ;
  assign n22506 = ~n22500 & ~n22505 ;
  assign n22507 = ~n22496 & ~n22506 ;
  assign n22514 = ~n22507 & n22513 ;
  assign n22523 = n22475 & n22487 ;
  assign n22524 = ~n22462 & ~n22523 ;
  assign n22528 = ~n22481 & ~n22524 ;
  assign n22529 = ~n22527 & n22528 ;
  assign n22518 = ~n22492 & ~n22517 ;
  assign n22515 = ~n22468 & ~n22474 ;
  assign n22516 = ~n22481 & ~n22515 ;
  assign n22519 = n22462 & ~n22516 ;
  assign n22520 = ~n22518 & n22519 ;
  assign n22521 = ~n22487 & n22515 ;
  assign n22522 = n22497 & n22521 ;
  assign n22545 = ~n22520 & ~n22522 ;
  assign n22546 = ~n22529 & n22545 ;
  assign n22547 = ~n22514 & n22546 ;
  assign n22548 = ~n22544 & n22547 ;
  assign n22549 = ~\u2_L2_reg[11]/NET0131  & n22548 ;
  assign n22550 = \u2_L2_reg[11]/NET0131  & ~n22548 ;
  assign n22551 = ~n22549 & ~n22550 ;
  assign n22581 = decrypt_pad & ~\u2_uk_K_r2_reg[0]/NET0131  ;
  assign n22582 = ~decrypt_pad & ~\u2_uk_K_r2_reg[22]/NET0131  ;
  assign n22583 = ~n22581 & ~n22582 ;
  assign n22584 = \u2_R2_reg[28]/NET0131  & ~n22583 ;
  assign n22585 = ~\u2_R2_reg[28]/NET0131  & n22583 ;
  assign n22586 = ~n22584 & ~n22585 ;
  assign n22552 = decrypt_pad & ~\u2_uk_K_r2_reg[50]/NET0131  ;
  assign n22553 = ~decrypt_pad & ~\u2_uk_K_r2_reg[45]/NET0131  ;
  assign n22554 = ~n22552 & ~n22553 ;
  assign n22555 = \u2_R2_reg[25]/NET0131  & ~n22554 ;
  assign n22556 = ~\u2_R2_reg[25]/NET0131  & n22554 ;
  assign n22557 = ~n22555 & ~n22556 ;
  assign n22565 = decrypt_pad & ~\u2_uk_K_r2_reg[15]/NET0131  ;
  assign n22566 = ~decrypt_pad & ~\u2_uk_K_r2_reg[37]/NET0131  ;
  assign n22567 = ~n22565 & ~n22566 ;
  assign n22568 = \u2_R2_reg[24]/NET0131  & ~n22567 ;
  assign n22569 = ~\u2_R2_reg[24]/NET0131  & n22567 ;
  assign n22570 = ~n22568 & ~n22569 ;
  assign n22587 = decrypt_pad & ~\u2_uk_K_r2_reg[23]/NET0131  ;
  assign n22588 = ~decrypt_pad & ~\u2_uk_K_r2_reg[14]/NET0131  ;
  assign n22589 = ~n22587 & ~n22588 ;
  assign n22590 = \u2_R2_reg[29]/NET0131  & ~n22589 ;
  assign n22591 = ~\u2_R2_reg[29]/NET0131  & n22589 ;
  assign n22592 = ~n22590 & ~n22591 ;
  assign n22593 = ~n22570 & n22592 ;
  assign n22604 = n22557 & n22593 ;
  assign n22606 = ~n22557 & n22570 ;
  assign n22607 = n22592 & n22606 ;
  assign n22608 = ~n22604 & ~n22607 ;
  assign n22558 = decrypt_pad & ~\u2_uk_K_r2_reg[44]/NET0131  ;
  assign n22559 = ~decrypt_pad & ~\u2_uk_K_r2_reg[35]/NET0131  ;
  assign n22560 = ~n22558 & ~n22559 ;
  assign n22561 = \u2_R2_reg[27]/NET0131  & ~n22560 ;
  assign n22562 = ~\u2_R2_reg[27]/NET0131  & n22560 ;
  assign n22563 = ~n22561 & ~n22562 ;
  assign n22571 = decrypt_pad & ~\u2_uk_K_r2_reg[35]/NET0131  ;
  assign n22572 = ~decrypt_pad & ~\u2_uk_K_r2_reg[2]/NET0131  ;
  assign n22573 = ~n22571 & ~n22572 ;
  assign n22574 = \u2_R2_reg[26]/NET0131  & ~n22573 ;
  assign n22575 = ~\u2_R2_reg[26]/NET0131  & n22573 ;
  assign n22576 = ~n22574 & ~n22575 ;
  assign n22605 = n22576 & ~n22604 ;
  assign n22609 = ~n22563 & ~n22605 ;
  assign n22610 = ~n22608 & n22609 ;
  assign n22594 = ~n22557 & n22576 ;
  assign n22599 = n22557 & n22592 ;
  assign n22600 = ~n22576 & n22599 ;
  assign n22601 = ~n22594 & ~n22600 ;
  assign n22602 = n22563 & n22570 ;
  assign n22603 = ~n22601 & n22602 ;
  assign n22595 = n22593 & n22594 ;
  assign n22596 = ~n22557 & ~n22576 ;
  assign n22597 = ~n22570 & ~n22592 ;
  assign n22598 = n22596 & n22597 ;
  assign n22611 = ~n22595 & ~n22598 ;
  assign n22612 = ~n22603 & n22611 ;
  assign n22613 = ~n22610 & n22612 ;
  assign n22614 = n22586 & ~n22613 ;
  assign n22564 = n22557 & ~n22563 ;
  assign n22619 = ~n22564 & ~n22596 ;
  assign n22617 = ~n22563 & ~n22576 ;
  assign n22618 = n22592 & n22617 ;
  assign n22620 = n22570 & ~n22618 ;
  assign n22621 = ~n22619 & n22620 ;
  assign n22615 = n22594 & n22597 ;
  assign n22616 = ~n22563 & n22615 ;
  assign n22577 = ~n22570 & n22576 ;
  assign n22578 = n22570 & ~n22576 ;
  assign n22579 = ~n22577 & ~n22578 ;
  assign n22622 = ~n22557 & n22563 ;
  assign n22623 = n22592 & ~n22622 ;
  assign n22624 = n22579 & n22623 ;
  assign n22625 = ~n22616 & ~n22624 ;
  assign n22626 = ~n22621 & n22625 ;
  assign n22627 = ~n22586 & ~n22626 ;
  assign n22580 = n22564 & n22579 ;
  assign n22628 = n22557 & n22576 ;
  assign n22629 = n22597 & n22628 ;
  assign n22630 = ~n22595 & ~n22629 ;
  assign n22631 = ~n22557 & ~n22592 ;
  assign n22632 = ~n22577 & n22631 ;
  assign n22633 = n22630 & ~n22632 ;
  assign n22634 = n22563 & ~n22633 ;
  assign n22635 = ~n22580 & ~n22634 ;
  assign n22636 = ~n22627 & n22635 ;
  assign n22637 = ~n22614 & n22636 ;
  assign n22638 = ~\u2_L2_reg[22]/NET0131  & ~n22637 ;
  assign n22639 = \u2_L2_reg[22]/NET0131  & n22637 ;
  assign n22640 = ~n22638 & ~n22639 ;
  assign n22659 = ~n22391 & ~n22421 ;
  assign n22660 = n22384 & n22406 ;
  assign n22661 = ~n22659 & ~n22660 ;
  assign n22662 = n22399 & ~n22661 ;
  assign n22656 = ~n22382 & n22391 ;
  assign n22663 = ~n22399 & ~n22656 ;
  assign n22664 = ~n22659 & n22663 ;
  assign n22642 = n22369 & n22375 ;
  assign n22655 = n22382 & n22642 ;
  assign n22657 = ~n22375 & n22656 ;
  assign n22658 = n22369 & n22657 ;
  assign n22665 = ~n22655 & ~n22658 ;
  assign n22666 = ~n22664 & n22665 ;
  assign n22667 = ~n22662 & n22666 ;
  assign n22668 = n22416 & ~n22667 ;
  assign n22641 = n22369 & n22392 ;
  assign n22643 = ~n22436 & ~n22642 ;
  assign n22644 = n22391 & ~n22643 ;
  assign n22645 = ~n22416 & n22644 ;
  assign n22646 = ~n22641 & ~n22645 ;
  assign n22647 = n22399 & ~n22646 ;
  assign n22649 = n22369 & ~n22424 ;
  assign n22650 = ~n22399 & ~n22403 ;
  assign n22651 = ~n22649 & n22650 ;
  assign n22648 = n22369 & n22425 ;
  assign n22652 = ~n22440 & ~n22648 ;
  assign n22653 = ~n22651 & n22652 ;
  assign n22654 = ~n22416 & ~n22653 ;
  assign n22669 = ~n22647 & ~n22654 ;
  assign n22670 = ~n22668 & n22669 ;
  assign n22671 = ~\u2_L2_reg[17]/NET0131  & ~n22670 ;
  assign n22672 = \u2_L2_reg[17]/NET0131  & n22670 ;
  assign n22673 = ~n22671 & ~n22672 ;
  assign n22674 = decrypt_pad & ~\u2_uk_K_r2_reg[47]/NET0131  ;
  assign n22675 = ~decrypt_pad & ~\u2_uk_K_r2_reg[10]/NET0131  ;
  assign n22676 = ~n22674 & ~n22675 ;
  assign n22677 = \u2_R2_reg[15]/NET0131  & ~n22676 ;
  assign n22678 = ~\u2_R2_reg[15]/NET0131  & n22676 ;
  assign n22679 = ~n22677 & ~n22678 ;
  assign n22693 = decrypt_pad & ~\u2_uk_K_r2_reg[13]/NET0131  ;
  assign n22694 = ~decrypt_pad & ~\u2_uk_K_r2_reg[33]/NET0131  ;
  assign n22695 = ~n22693 & ~n22694 ;
  assign n22696 = \u2_R2_reg[13]/NET0131  & ~n22695 ;
  assign n22697 = ~\u2_R2_reg[13]/NET0131  & n22695 ;
  assign n22698 = ~n22696 & ~n22697 ;
  assign n22680 = decrypt_pad & ~\u2_uk_K_r2_reg[3]/NET0131  ;
  assign n22681 = ~decrypt_pad & ~\u2_uk_K_r2_reg[55]/NET0131  ;
  assign n22682 = ~n22680 & ~n22681 ;
  assign n22683 = \u2_R2_reg[17]/NET0131  & ~n22682 ;
  assign n22684 = ~\u2_R2_reg[17]/NET0131  & n22682 ;
  assign n22685 = ~n22683 & ~n22684 ;
  assign n22687 = decrypt_pad & ~\u2_uk_K_r2_reg[19]/NET0131  ;
  assign n22688 = ~decrypt_pad & ~\u2_uk_K_r2_reg[39]/NET0131  ;
  assign n22689 = ~n22687 & ~n22688 ;
  assign n22690 = \u2_R2_reg[12]/NET0131  & ~n22689 ;
  assign n22691 = ~\u2_R2_reg[12]/NET0131  & n22689 ;
  assign n22692 = ~n22690 & ~n22691 ;
  assign n22720 = n22685 & n22692 ;
  assign n22721 = n22698 & n22720 ;
  assign n22722 = n22679 & n22721 ;
  assign n22686 = n22679 & ~n22685 ;
  assign n22699 = ~n22692 & ~n22698 ;
  assign n22700 = n22686 & n22699 ;
  assign n22725 = decrypt_pad & ~\u2_uk_K_r2_reg[55]/NET0131  ;
  assign n22726 = ~decrypt_pad & ~\u2_uk_K_r2_reg[18]/NET0131  ;
  assign n22727 = ~n22725 & ~n22726 ;
  assign n22728 = \u2_R2_reg[16]/NET0131  & ~n22727 ;
  assign n22729 = ~\u2_R2_reg[16]/NET0131  & n22727 ;
  assign n22730 = ~n22728 & ~n22729 ;
  assign n22731 = ~n22700 & ~n22730 ;
  assign n22712 = ~n22692 & n22698 ;
  assign n22703 = decrypt_pad & ~\u2_uk_K_r2_reg[39]/NET0131  ;
  assign n22704 = ~decrypt_pad & ~\u2_uk_K_r2_reg[34]/NET0131  ;
  assign n22705 = ~n22703 & ~n22704 ;
  assign n22706 = \u2_R2_reg[14]/NET0131  & ~n22705 ;
  assign n22707 = ~\u2_R2_reg[14]/NET0131  & n22705 ;
  assign n22708 = ~n22706 & ~n22707 ;
  assign n22718 = n22679 & n22708 ;
  assign n22719 = n22712 & n22718 ;
  assign n22701 = n22685 & ~n22698 ;
  assign n22723 = n22692 & ~n22708 ;
  assign n22724 = n22701 & n22723 ;
  assign n22732 = ~n22719 & ~n22724 ;
  assign n22733 = n22731 & n22732 ;
  assign n22734 = ~n22722 & n22733 ;
  assign n22702 = ~n22685 & n22692 ;
  assign n22709 = n22702 & n22708 ;
  assign n22710 = ~n22701 & ~n22709 ;
  assign n22711 = ~n22679 & ~n22710 ;
  assign n22713 = ~n22685 & n22712 ;
  assign n22714 = n22708 & n22713 ;
  assign n22715 = ~n22685 & ~n22708 ;
  assign n22716 = n22699 & n22715 ;
  assign n22717 = ~n22714 & ~n22716 ;
  assign n22735 = ~n22711 & n22717 ;
  assign n22736 = n22734 & n22735 ;
  assign n22745 = ~n22679 & ~n22685 ;
  assign n22746 = n22699 & n22745 ;
  assign n22747 = ~n22721 & ~n22746 ;
  assign n22748 = n22708 & ~n22747 ;
  assign n22737 = n22685 & ~n22692 ;
  assign n22738 = n22679 & n22737 ;
  assign n22739 = ~n22698 & n22738 ;
  assign n22752 = n22730 & ~n22739 ;
  assign n22740 = n22692 & n22698 ;
  assign n22741 = n22686 & n22740 ;
  assign n22742 = n22698 & ~n22708 ;
  assign n22743 = n22737 & n22742 ;
  assign n22744 = ~n22741 & ~n22743 ;
  assign n22749 = ~n22679 & ~n22708 ;
  assign n22750 = ~n22699 & ~n22740 ;
  assign n22751 = n22749 & n22750 ;
  assign n22753 = n22744 & ~n22751 ;
  assign n22754 = n22752 & n22753 ;
  assign n22755 = ~n22748 & n22754 ;
  assign n22756 = ~n22736 & ~n22755 ;
  assign n22757 = ~n22679 & ~n22743 ;
  assign n22758 = ~n22698 & n22708 ;
  assign n22759 = n22702 & n22758 ;
  assign n22760 = n22679 & ~n22759 ;
  assign n22761 = ~n22716 & n22760 ;
  assign n22762 = ~n22757 & ~n22761 ;
  assign n22763 = ~n22708 & n22740 ;
  assign n22764 = n22686 & n22763 ;
  assign n22765 = ~n22762 & ~n22764 ;
  assign n22766 = ~n22756 & n22765 ;
  assign n22767 = ~\u2_L2_reg[20]/NET0131  & ~n22766 ;
  assign n22768 = \u2_L2_reg[20]/NET0131  & n22766 ;
  assign n22769 = ~n22767 & ~n22768 ;
  assign n22786 = n22475 & ~n22487 ;
  assign n22787 = ~n22493 & ~n22786 ;
  assign n22788 = ~n22488 & ~n22491 ;
  assign n22789 = ~n22474 & ~n22788 ;
  assign n22790 = n22787 & ~n22789 ;
  assign n22791 = n22462 & ~n22790 ;
  assign n22770 = n22481 & n22523 ;
  assign n22777 = ~n22481 & ~n22498 ;
  assign n22792 = ~n22770 & ~n22777 ;
  assign n22793 = ~n22462 & ~n22792 ;
  assign n22794 = n22481 & n22526 ;
  assign n22795 = ~n22793 & ~n22794 ;
  assign n22796 = ~n22791 & n22795 ;
  assign n22797 = ~n22513 & ~n22796 ;
  assign n22771 = n22487 & n22538 ;
  assign n22772 = ~n22502 & ~n22771 ;
  assign n22773 = ~n22770 & n22772 ;
  assign n22774 = n22462 & ~n22773 ;
  assign n22778 = n22462 & ~n22525 ;
  assign n22779 = ~n22536 & n22778 ;
  assign n22775 = n22481 & ~n22492 ;
  assign n22776 = ~n22515 & n22775 ;
  assign n22780 = ~n22776 & ~n22777 ;
  assign n22781 = ~n22779 & n22780 ;
  assign n22782 = ~n22774 & ~n22781 ;
  assign n22783 = n22513 & ~n22782 ;
  assign n22784 = n22462 & n22474 ;
  assign n22785 = n22517 & n22784 ;
  assign n22798 = ~n22489 & ~n22785 ;
  assign n22799 = ~n22783 & n22798 ;
  assign n22800 = ~n22797 & n22799 ;
  assign n22801 = \u2_L2_reg[29]/NET0131  & ~n22800 ;
  assign n22802 = ~\u2_L2_reg[29]/NET0131  & n22800 ;
  assign n22803 = ~n22801 & ~n22802 ;
  assign n22804 = decrypt_pad & ~\u2_uk_K_r2_reg[54]/NET0131  ;
  assign n22805 = ~decrypt_pad & ~\u2_uk_K_r2_reg[17]/NET0131  ;
  assign n22806 = ~n22804 & ~n22805 ;
  assign n22807 = \u2_R2_reg[8]/NET0131  & ~n22806 ;
  assign n22808 = ~\u2_R2_reg[8]/NET0131  & n22806 ;
  assign n22809 = ~n22807 & ~n22808 ;
  assign n22810 = decrypt_pad & ~\u2_uk_K_r2_reg[46]/NET0131  ;
  assign n22811 = ~decrypt_pad & ~\u2_uk_K_r2_reg[41]/NET0131  ;
  assign n22812 = ~n22810 & ~n22811 ;
  assign n22813 = \u2_R2_reg[5]/NET0131  & ~n22812 ;
  assign n22814 = ~\u2_R2_reg[5]/NET0131  & n22812 ;
  assign n22815 = ~n22813 & ~n22814 ;
  assign n22816 = decrypt_pad & ~\u2_uk_K_r2_reg[34]/NET0131  ;
  assign n22817 = ~decrypt_pad & ~\u2_uk_K_r2_reg[54]/NET0131  ;
  assign n22818 = ~n22816 & ~n22817 ;
  assign n22819 = \u2_R2_reg[9]/NET0131  & ~n22818 ;
  assign n22820 = ~\u2_R2_reg[9]/NET0131  & n22818 ;
  assign n22821 = ~n22819 & ~n22820 ;
  assign n22822 = n22815 & ~n22821 ;
  assign n22823 = ~n22815 & n22821 ;
  assign n22824 = decrypt_pad & ~\u2_uk_K_r2_reg[10]/NET0131  ;
  assign n22825 = ~decrypt_pad & ~\u2_uk_K_r2_reg[5]/NET0131  ;
  assign n22826 = ~n22824 & ~n22825 ;
  assign n22827 = \u2_R2_reg[4]/NET0131  & ~n22826 ;
  assign n22828 = ~\u2_R2_reg[4]/NET0131  & n22826 ;
  assign n22829 = ~n22827 & ~n22828 ;
  assign n22830 = n22823 & ~n22829 ;
  assign n22831 = ~n22822 & ~n22830 ;
  assign n22832 = decrypt_pad & ~\u2_uk_K_r2_reg[12]/NET0131  ;
  assign n22833 = ~decrypt_pad & ~\u2_uk_K_r2_reg[32]/NET0131  ;
  assign n22834 = ~n22832 & ~n22833 ;
  assign n22835 = \u2_R2_reg[6]/NET0131  & ~n22834 ;
  assign n22836 = ~\u2_R2_reg[6]/NET0131  & n22834 ;
  assign n22837 = ~n22835 & ~n22836 ;
  assign n22838 = ~n22831 & ~n22837 ;
  assign n22839 = decrypt_pad & ~\u2_uk_K_r2_reg[6]/NET0131  ;
  assign n22840 = ~decrypt_pad & ~\u2_uk_K_r2_reg[26]/NET0131  ;
  assign n22841 = ~n22839 & ~n22840 ;
  assign n22842 = \u2_R2_reg[7]/NET0131  & ~n22841 ;
  assign n22843 = ~\u2_R2_reg[7]/NET0131  & n22841 ;
  assign n22844 = ~n22842 & ~n22843 ;
  assign n22845 = ~n22815 & n22837 ;
  assign n22846 = n22821 & n22829 ;
  assign n22847 = n22845 & n22846 ;
  assign n22848 = n22844 & n22847 ;
  assign n22862 = ~n22838 & ~n22848 ;
  assign n22849 = n22829 & n22837 ;
  assign n22850 = ~n22823 & n22849 ;
  assign n22851 = ~n22830 & ~n22850 ;
  assign n22852 = ~n22844 & ~n22851 ;
  assign n22856 = n22815 & ~n22837 ;
  assign n22857 = ~n22837 & n22844 ;
  assign n22858 = ~n22856 & ~n22857 ;
  assign n22853 = n22821 & ~n22829 ;
  assign n22854 = n22815 & ~n22853 ;
  assign n22855 = ~n22821 & ~n22837 ;
  assign n22859 = ~n22845 & ~n22855 ;
  assign n22860 = ~n22854 & n22859 ;
  assign n22861 = n22858 & n22860 ;
  assign n22863 = ~n22852 & ~n22861 ;
  assign n22864 = n22862 & n22863 ;
  assign n22865 = ~n22809 & ~n22864 ;
  assign n22878 = ~n22821 & ~n22829 ;
  assign n22882 = ~n22847 & ~n22878 ;
  assign n22883 = n22809 & ~n22882 ;
  assign n22884 = ~n22845 & n22853 ;
  assign n22885 = ~n22883 & ~n22884 ;
  assign n22886 = ~n22844 & ~n22856 ;
  assign n22887 = ~n22885 & n22886 ;
  assign n22872 = ~n22837 & n22846 ;
  assign n22873 = n22815 & n22872 ;
  assign n22866 = ~n22821 & n22829 ;
  assign n22867 = ~n22815 & n22866 ;
  assign n22868 = ~n22837 & n22867 ;
  assign n22869 = ~n22829 & n22837 ;
  assign n22870 = n22815 & n22844 ;
  assign n22871 = ~n22869 & n22870 ;
  assign n22874 = ~n22868 & ~n22871 ;
  assign n22875 = ~n22873 & n22874 ;
  assign n22876 = n22809 & ~n22875 ;
  assign n22879 = ~n22856 & ~n22878 ;
  assign n22877 = ~n22829 & ~n22845 ;
  assign n22880 = n22844 & ~n22877 ;
  assign n22881 = ~n22879 & n22880 ;
  assign n22888 = ~n22876 & ~n22881 ;
  assign n22889 = ~n22887 & n22888 ;
  assign n22890 = ~n22865 & n22889 ;
  assign n22891 = \u2_L2_reg[2]/NET0131  & n22890 ;
  assign n22892 = ~\u2_L2_reg[2]/NET0131  & ~n22890 ;
  assign n22893 = ~n22891 & ~n22892 ;
  assign n22903 = n22720 & n22749 ;
  assign n22909 = ~n22746 & ~n22763 ;
  assign n22910 = ~n22903 & n22909 ;
  assign n22904 = ~n22685 & ~n22698 ;
  assign n22905 = ~n22758 & ~n22904 ;
  assign n22906 = n22679 & n22692 ;
  assign n22907 = ~n22905 & n22906 ;
  assign n22908 = ~n22708 & n22738 ;
  assign n22911 = ~n22907 & ~n22908 ;
  assign n22912 = n22910 & n22911 ;
  assign n22913 = n22717 & n22912 ;
  assign n22914 = ~n22730 & ~n22913 ;
  assign n22894 = n22679 & ~n22724 ;
  assign n22895 = ~n22713 & n22894 ;
  assign n22896 = n22702 & ~n22742 ;
  assign n22897 = n22757 & ~n22896 ;
  assign n22898 = ~n22895 & ~n22897 ;
  assign n22899 = n22708 & ~n22750 ;
  assign n22900 = n22685 & n22899 ;
  assign n22901 = ~n22898 & ~n22900 ;
  assign n22902 = n22730 & ~n22901 ;
  assign n22915 = ~n22716 & ~n22900 ;
  assign n22916 = ~n22679 & ~n22915 ;
  assign n22917 = ~n22719 & ~n22764 ;
  assign n22918 = ~n22916 & n22917 ;
  assign n22919 = ~n22902 & n22918 ;
  assign n22920 = ~n22914 & n22919 ;
  assign n22921 = ~\u2_L2_reg[10]/NET0131  & ~n22920 ;
  assign n22922 = \u2_L2_reg[10]/NET0131  & n22920 ;
  assign n22923 = ~n22921 & ~n22922 ;
  assign n22928 = n22570 & n22576 ;
  assign n22930 = n22592 & n22928 ;
  assign n22931 = n22578 & ~n22592 ;
  assign n22932 = ~n22930 & ~n22931 ;
  assign n22933 = ~n22557 & ~n22932 ;
  assign n22924 = ~n22596 & ~n22628 ;
  assign n22925 = n22597 & n22924 ;
  assign n22929 = ~n22563 & n22928 ;
  assign n22936 = ~n22586 & ~n22929 ;
  assign n22937 = ~n22925 & n22936 ;
  assign n22926 = ~n22599 & ~n22631 ;
  assign n22927 = ~n22563 & ~n22926 ;
  assign n22934 = ~n22622 & ~n22628 ;
  assign n22935 = n22593 & ~n22934 ;
  assign n22938 = ~n22927 & ~n22935 ;
  assign n22939 = n22937 & n22938 ;
  assign n22940 = ~n22933 & n22939 ;
  assign n22947 = ~n22592 & n22596 ;
  assign n22948 = ~n22570 & ~n22947 ;
  assign n22949 = n22563 & ~n22606 ;
  assign n22950 = ~n22948 & n22949 ;
  assign n22941 = ~n22576 & ~n22608 ;
  assign n22942 = n22570 & ~n22592 ;
  assign n22943 = ~n22593 & ~n22942 ;
  assign n22944 = n22563 & ~n22570 ;
  assign n22945 = n22594 & ~n22944 ;
  assign n22946 = ~n22943 & n22945 ;
  assign n22951 = n22586 & ~n22629 ;
  assign n22952 = ~n22946 & n22951 ;
  assign n22953 = ~n22941 & n22952 ;
  assign n22954 = ~n22950 & n22953 ;
  assign n22955 = ~n22940 & ~n22954 ;
  assign n22956 = \u2_L2_reg[12]/NET0131  & n22955 ;
  assign n22957 = ~\u2_L2_reg[12]/NET0131  & ~n22955 ;
  assign n22958 = ~n22956 & ~n22957 ;
  assign n22959 = n22822 & n22849 ;
  assign n22960 = ~n22873 & ~n22959 ;
  assign n22961 = n22830 & n22837 ;
  assign n22962 = n22822 & ~n22829 ;
  assign n22963 = ~n22868 & ~n22962 ;
  assign n22964 = ~n22961 & n22963 ;
  assign n22965 = ~n22809 & ~n22964 ;
  assign n22966 = n22960 & ~n22965 ;
  assign n22967 = ~n22844 & ~n22966 ;
  assign n22971 = ~n22815 & ~n22853 ;
  assign n22972 = ~n22866 & ~n22971 ;
  assign n22973 = ~n22856 & n22866 ;
  assign n22974 = n22844 & ~n22973 ;
  assign n22975 = ~n22972 & n22974 ;
  assign n22969 = ~n22822 & n22844 ;
  assign n22970 = n22849 & n22969 ;
  assign n22968 = n22853 & ~n22858 ;
  assign n22976 = ~n22809 & ~n22968 ;
  assign n22977 = ~n22970 & n22976 ;
  assign n22978 = ~n22975 & n22977 ;
  assign n22985 = ~n22837 & n22962 ;
  assign n22986 = n22809 & ~n22985 ;
  assign n22987 = ~n22861 & n22986 ;
  assign n22983 = ~n22855 & n22971 ;
  assign n22984 = ~n22844 & n22983 ;
  assign n22979 = ~n22815 & n22855 ;
  assign n22980 = n22837 & n22853 ;
  assign n22981 = ~n22979 & ~n22980 ;
  assign n22982 = n22844 & ~n22981 ;
  assign n22988 = n22960 & ~n22982 ;
  assign n22989 = ~n22984 & n22988 ;
  assign n22990 = n22987 & n22989 ;
  assign n22991 = ~n22978 & ~n22990 ;
  assign n22992 = ~n22967 & ~n22991 ;
  assign n22993 = ~\u2_L2_reg[13]/NET0131  & n22992 ;
  assign n22994 = \u2_L2_reg[13]/NET0131  & ~n22992 ;
  assign n22995 = ~n22993 & ~n22994 ;
  assign n23055 = decrypt_pad & ~\u2_uk_K_r2_reg[36]/NET0131  ;
  assign n23056 = ~decrypt_pad & ~\u2_uk_K_r2_reg[31]/NET0131  ;
  assign n23057 = ~n23055 & ~n23056 ;
  assign n23058 = \u2_R2_reg[20]/NET0131  & ~n23057 ;
  assign n23059 = ~\u2_R2_reg[20]/NET0131  & n23057 ;
  assign n23060 = ~n23058 & ~n23059 ;
  assign n22996 = decrypt_pad & ~\u2_uk_K_r2_reg[21]/NET0131  ;
  assign n22997 = ~decrypt_pad & ~\u2_uk_K_r2_reg[43]/NET0131  ;
  assign n22998 = ~n22996 & ~n22997 ;
  assign n22999 = \u2_R2_reg[19]/NET0131  & ~n22998 ;
  assign n23000 = ~\u2_R2_reg[19]/NET0131  & n22998 ;
  assign n23001 = ~n22999 & ~n23000 ;
  assign n23022 = decrypt_pad & ~\u2_uk_K_r2_reg[49]/NET0131  ;
  assign n23023 = ~decrypt_pad & ~\u2_uk_K_r2_reg[16]/NET0131  ;
  assign n23024 = ~n23022 & ~n23023 ;
  assign n23025 = \u2_R2_reg[16]/NET0131  & ~n23024 ;
  assign n23026 = ~\u2_R2_reg[16]/NET0131  & n23024 ;
  assign n23027 = ~n23025 & ~n23026 ;
  assign n23002 = decrypt_pad & ~\u2_uk_K_r2_reg[16]/NET0131  ;
  assign n23003 = ~decrypt_pad & ~\u2_uk_K_r2_reg[7]/NET0131  ;
  assign n23004 = ~n23002 & ~n23003 ;
  assign n23005 = \u2_R2_reg[17]/NET0131  & ~n23004 ;
  assign n23006 = ~\u2_R2_reg[17]/NET0131  & n23004 ;
  assign n23007 = ~n23005 & ~n23006 ;
  assign n23008 = decrypt_pad & ~\u2_uk_K_r2_reg[38]/NET0131  ;
  assign n23009 = ~decrypt_pad & ~\u2_uk_K_r2_reg[1]/NET0131  ;
  assign n23010 = ~n23008 & ~n23009 ;
  assign n23011 = \u2_R2_reg[18]/NET0131  & ~n23010 ;
  assign n23012 = ~\u2_R2_reg[18]/NET0131  & n23010 ;
  assign n23013 = ~n23011 & ~n23012 ;
  assign n23043 = n23007 & ~n23013 ;
  assign n23044 = ~n23027 & n23043 ;
  assign n23015 = decrypt_pad & ~\u2_uk_K_r2_reg[37]/NET0131  ;
  assign n23016 = ~decrypt_pad & ~\u2_uk_K_r2_reg[28]/NET0131  ;
  assign n23017 = ~n23015 & ~n23016 ;
  assign n23018 = \u2_R2_reg[21]/NET0131  & ~n23017 ;
  assign n23019 = ~\u2_R2_reg[21]/NET0131  & n23017 ;
  assign n23020 = ~n23018 & ~n23019 ;
  assign n23046 = n23013 & n23027 ;
  assign n23047 = n23020 & ~n23046 ;
  assign n23048 = ~n23044 & n23047 ;
  assign n23028 = ~n23020 & n23027 ;
  assign n23062 = n23007 & n23028 ;
  assign n23063 = ~n23048 & ~n23062 ;
  assign n23064 = n23001 & ~n23063 ;
  assign n23067 = ~n23001 & ~n23013 ;
  assign n23031 = n23007 & n23020 ;
  assign n23068 = ~n23027 & n23031 ;
  assign n23069 = ~n23020 & ~n23027 ;
  assign n23070 = ~n23007 & n23069 ;
  assign n23071 = ~n23068 & ~n23070 ;
  assign n23072 = n23067 & ~n23071 ;
  assign n23075 = ~n23007 & n23013 ;
  assign n23076 = ~n23043 & ~n23075 ;
  assign n23077 = n23028 & ~n23076 ;
  assign n23040 = ~n23007 & n23027 ;
  assign n23065 = ~n23013 & n23020 ;
  assign n23066 = n23040 & n23065 ;
  assign n23032 = n23027 & n23031 ;
  assign n23073 = ~n23001 & n23013 ;
  assign n23074 = n23032 & n23073 ;
  assign n23078 = ~n23066 & ~n23074 ;
  assign n23079 = ~n23077 & n23078 ;
  assign n23080 = ~n23072 & n23079 ;
  assign n23081 = ~n23064 & n23080 ;
  assign n23082 = n23060 & ~n23081 ;
  assign n23033 = ~n23013 & n23032 ;
  assign n23029 = ~n23007 & n23028 ;
  assign n23030 = ~n23013 & n23029 ;
  assign n23014 = n23007 & n23013 ;
  assign n23021 = n23014 & ~n23020 ;
  assign n23034 = ~n23007 & ~n23027 ;
  assign n23035 = n23020 & n23034 ;
  assign n23036 = ~n23021 & ~n23035 ;
  assign n23037 = ~n23030 & n23036 ;
  assign n23038 = ~n23033 & n23037 ;
  assign n23039 = ~n23001 & ~n23038 ;
  assign n23049 = n23001 & ~n23028 ;
  assign n23050 = ~n23021 & n23049 ;
  assign n23051 = ~n23048 & n23050 ;
  assign n23041 = n23020 & n23040 ;
  assign n23042 = n23013 & n23041 ;
  assign n23045 = ~n23020 & n23044 ;
  assign n23052 = ~n23042 & ~n23045 ;
  assign n23053 = ~n23051 & n23052 ;
  assign n23054 = ~n23039 & n23053 ;
  assign n23061 = ~n23054 & ~n23060 ;
  assign n23083 = ~n23013 & n23062 ;
  assign n23084 = n23013 & n23070 ;
  assign n23085 = ~n23083 & ~n23084 ;
  assign n23086 = n23001 & ~n23085 ;
  assign n23087 = n23013 & n23035 ;
  assign n23088 = n23014 & n23069 ;
  assign n23089 = ~n23087 & ~n23088 ;
  assign n23090 = ~n23001 & ~n23089 ;
  assign n23091 = ~n23086 & ~n23090 ;
  assign n23092 = ~n23061 & n23091 ;
  assign n23093 = ~n23082 & n23092 ;
  assign n23094 = ~\u2_L2_reg[14]/NET0131  & ~n23093 ;
  assign n23095 = \u2_L2_reg[14]/NET0131  & n23093 ;
  assign n23096 = ~n23094 & ~n23095 ;
  assign n23097 = decrypt_pad & ~\u2_uk_K_r2_reg[29]/NET0131  ;
  assign n23098 = ~decrypt_pad & ~\u2_uk_K_r2_reg[51]/NET0131  ;
  assign n23099 = ~n23097 & ~n23098 ;
  assign n23100 = \u2_R2_reg[28]/NET0131  & ~n23099 ;
  assign n23101 = ~\u2_R2_reg[28]/NET0131  & n23099 ;
  assign n23102 = ~n23100 & ~n23101 ;
  assign n23103 = decrypt_pad & ~\u2_uk_K_r2_reg[2]/NET0131  ;
  assign n23104 = ~decrypt_pad & ~\u2_uk_K_r2_reg[52]/NET0131  ;
  assign n23105 = ~n23103 & ~n23104 ;
  assign n23106 = \u2_R2_reg[30]/NET0131  & ~n23105 ;
  assign n23107 = ~\u2_R2_reg[30]/NET0131  & n23105 ;
  assign n23108 = ~n23106 & ~n23107 ;
  assign n23109 = ~n23102 & n23108 ;
  assign n23110 = n23102 & ~n23108 ;
  assign n23111 = ~n23109 & ~n23110 ;
  assign n23112 = decrypt_pad & ~\u2_uk_K_r2_reg[45]/NET0131  ;
  assign n23113 = ~decrypt_pad & ~\u2_uk_K_r2_reg[8]/NET0131  ;
  assign n23114 = ~n23112 & ~n23113 ;
  assign n23115 = \u2_R2_reg[1]/NET0131  & ~n23114 ;
  assign n23116 = ~\u2_R2_reg[1]/NET0131  & n23114 ;
  assign n23117 = ~n23115 & ~n23116 ;
  assign n23118 = ~n23102 & n23117 ;
  assign n23119 = decrypt_pad & ~\u2_uk_K_r2_reg[1]/NET0131  ;
  assign n23120 = ~decrypt_pad & ~\u2_uk_K_r2_reg[23]/NET0131  ;
  assign n23121 = ~n23119 & ~n23120 ;
  assign n23122 = \u2_R2_reg[29]/NET0131  & ~n23121 ;
  assign n23123 = ~\u2_R2_reg[29]/NET0131  & n23121 ;
  assign n23124 = ~n23122 & ~n23123 ;
  assign n23125 = ~n23118 & n23124 ;
  assign n23126 = ~n23111 & n23125 ;
  assign n23136 = decrypt_pad & ~\u2_uk_K_r2_reg[51]/NET0131  ;
  assign n23137 = ~decrypt_pad & ~\u2_uk_K_r2_reg[42]/NET0131  ;
  assign n23138 = ~n23136 & ~n23137 ;
  assign n23139 = \u2_R2_reg[32]/NET0131  & ~n23138 ;
  assign n23140 = ~\u2_R2_reg[32]/NET0131  & n23138 ;
  assign n23141 = ~n23139 & ~n23140 ;
  assign n23147 = ~n23126 & n23141 ;
  assign n23127 = ~n23117 & ~n23124 ;
  assign n23128 = ~n23102 & n23127 ;
  assign n23129 = decrypt_pad & ~\u2_uk_K_r2_reg[14]/NET0131  ;
  assign n23130 = ~decrypt_pad & ~\u2_uk_K_r2_reg[36]/NET0131  ;
  assign n23131 = ~n23129 & ~n23130 ;
  assign n23132 = \u2_R2_reg[31]/P0001  & ~n23131 ;
  assign n23133 = ~\u2_R2_reg[31]/P0001  & n23131 ;
  assign n23134 = ~n23132 & ~n23133 ;
  assign n23135 = n23128 & n23134 ;
  assign n23142 = n23117 & ~n23124 ;
  assign n23143 = n23102 & n23108 ;
  assign n23144 = n23108 & ~n23134 ;
  assign n23145 = ~n23143 & ~n23144 ;
  assign n23146 = n23142 & ~n23145 ;
  assign n23148 = ~n23135 & ~n23146 ;
  assign n23149 = n23147 & n23148 ;
  assign n23155 = ~n23124 & ~n23134 ;
  assign n23156 = ~n23108 & n23127 ;
  assign n23157 = ~n23155 & ~n23156 ;
  assign n23158 = n23102 & ~n23157 ;
  assign n23151 = n23118 & ~n23124 ;
  assign n23152 = ~n23125 & ~n23151 ;
  assign n23150 = n23109 & n23124 ;
  assign n23153 = n23134 & ~n23150 ;
  assign n23154 = ~n23152 & n23153 ;
  assign n23159 = ~n23141 & ~n23154 ;
  assign n23160 = ~n23158 & n23159 ;
  assign n23161 = ~n23149 & ~n23160 ;
  assign n23163 = n23111 & n23152 ;
  assign n23162 = ~n23117 & n23150 ;
  assign n23164 = ~n23134 & ~n23162 ;
  assign n23165 = ~n23163 & n23164 ;
  assign n23167 = ~n23108 & n23151 ;
  assign n23166 = n23117 & n23150 ;
  assign n23168 = n23134 & ~n23166 ;
  assign n23169 = ~n23167 & n23168 ;
  assign n23170 = ~n23165 & ~n23169 ;
  assign n23171 = ~n23161 & ~n23170 ;
  assign n23172 = ~\u2_L2_reg[15]/NET0131  & ~n23171 ;
  assign n23173 = \u2_L2_reg[15]/NET0131  & n23171 ;
  assign n23174 = ~n23172 & ~n23173 ;
  assign n23182 = ~n22692 & n22715 ;
  assign n23183 = n22760 & ~n23182 ;
  assign n23184 = ~n22701 & ~n22715 ;
  assign n23185 = n22692 & ~n23184 ;
  assign n23186 = ~n22679 & ~n23185 ;
  assign n23187 = ~n23183 & ~n23186 ;
  assign n23188 = n22708 & n22721 ;
  assign n23189 = ~n22702 & ~n22737 ;
  assign n23190 = n22742 & ~n23189 ;
  assign n23191 = ~n23188 & ~n23190 ;
  assign n23192 = ~n23187 & n23191 ;
  assign n23193 = ~n22730 & ~n23192 ;
  assign n23176 = ~n22698 & n22723 ;
  assign n23177 = ~n22701 & ~n23176 ;
  assign n23178 = n22730 & ~n23177 ;
  assign n23179 = ~n22714 & ~n22900 ;
  assign n23180 = ~n23178 & n23179 ;
  assign n23181 = n22679 & ~n23180 ;
  assign n23175 = n22745 & n22899 ;
  assign n23195 = ~n22702 & n22742 ;
  assign n23196 = n22698 & n22737 ;
  assign n23197 = ~n23195 & ~n23196 ;
  assign n23198 = ~n22679 & ~n23197 ;
  assign n23194 = n22698 & n22709 ;
  assign n23199 = ~n22692 & n22758 ;
  assign n23200 = ~n23194 & ~n23199 ;
  assign n23201 = ~n23198 & n23200 ;
  assign n23202 = n22730 & ~n23201 ;
  assign n23203 = ~n23175 & ~n23202 ;
  assign n23204 = ~n23181 & n23203 ;
  assign n23205 = ~n23193 & n23204 ;
  assign n23206 = ~\u2_L2_reg[1]/NET0131  & ~n23205 ;
  assign n23207 = \u2_L2_reg[1]/NET0131  & n23205 ;
  assign n23208 = ~n23206 & ~n23207 ;
  assign n23212 = ~n23111 & ~n23134 ;
  assign n23213 = ~n23127 & ~n23212 ;
  assign n23214 = ~n23111 & ~n23117 ;
  assign n23215 = ~n23213 & ~n23214 ;
  assign n23220 = ~n23108 & ~n23124 ;
  assign n23219 = n23117 & n23124 ;
  assign n23221 = n23102 & n23134 ;
  assign n23222 = ~n23219 & n23221 ;
  assign n23223 = ~n23220 & n23222 ;
  assign n23224 = ~n23141 & ~n23150 ;
  assign n23209 = ~n23117 & n23124 ;
  assign n23210 = ~n23102 & ~n23134 ;
  assign n23211 = n23209 & n23210 ;
  assign n23216 = ~n23108 & n23124 ;
  assign n23217 = n23102 & n23117 ;
  assign n23218 = n23216 & n23217 ;
  assign n23225 = ~n23211 & ~n23218 ;
  assign n23226 = n23224 & n23225 ;
  assign n23227 = ~n23223 & n23226 ;
  assign n23228 = ~n23215 & n23227 ;
  assign n23230 = n23102 & ~n23117 ;
  assign n23231 = ~n23108 & n23230 ;
  assign n23229 = n23142 & n23143 ;
  assign n23232 = ~n23134 & ~n23229 ;
  assign n23233 = ~n23231 & n23232 ;
  assign n23234 = ~n23118 & ~n23143 ;
  assign n23235 = n23124 & ~n23234 ;
  assign n23236 = n23117 & n23220 ;
  assign n23237 = n23134 & ~n23236 ;
  assign n23238 = ~n23235 & n23237 ;
  assign n23239 = ~n23233 & ~n23238 ;
  assign n23240 = n23124 & n23230 ;
  assign n23241 = ~n23128 & ~n23240 ;
  assign n23242 = n23108 & ~n23241 ;
  assign n23243 = n23141 & ~n23167 ;
  assign n23244 = ~n23242 & n23243 ;
  assign n23245 = ~n23239 & n23244 ;
  assign n23246 = ~n23228 & ~n23245 ;
  assign n23247 = ~n23102 & n23220 ;
  assign n23248 = n23134 & n23247 ;
  assign n23249 = ~n23134 & n23218 ;
  assign n23250 = ~n23248 & ~n23249 ;
  assign n23251 = ~n23246 & n23250 ;
  assign n23252 = ~\u2_L2_reg[21]/NET0131  & ~n23251 ;
  assign n23253 = \u2_L2_reg[21]/NET0131  & n23251 ;
  assign n23254 = ~n23252 & ~n23253 ;
  assign n23255 = ~n22391 & n22643 ;
  assign n23256 = ~n22443 & ~n23255 ;
  assign n23257 = n22416 & ~n23256 ;
  assign n23258 = n22421 & n22439 ;
  assign n23259 = ~n22658 & ~n23258 ;
  assign n23260 = ~n23257 & n23259 ;
  assign n23261 = ~n22399 & ~n23260 ;
  assign n23262 = n22391 & n22655 ;
  assign n23263 = n22369 & n22401 ;
  assign n23264 = ~n22406 & ~n23263 ;
  assign n23265 = n22399 & ~n23264 ;
  assign n23266 = ~n23262 & ~n23265 ;
  assign n23267 = ~n23261 & n23266 ;
  assign n23268 = ~n22427 & ~n23267 ;
  assign n23269 = n22369 & n22399 ;
  assign n23270 = ~n22656 & n23269 ;
  assign n23271 = n22403 & n23270 ;
  assign n23272 = n22416 & ~n22660 ;
  assign n23273 = ~n22437 & n23272 ;
  assign n23274 = ~n23271 & n23273 ;
  assign n23278 = n22401 & n23269 ;
  assign n23279 = ~n22416 & ~n23278 ;
  assign n23280 = ~n22429 & n23279 ;
  assign n23275 = n22408 & ~n22421 ;
  assign n23276 = ~n22436 & n23275 ;
  assign n23277 = n22385 & ~n22643 ;
  assign n23281 = ~n23276 & ~n23277 ;
  assign n23282 = n23280 & n23281 ;
  assign n23283 = ~n23274 & ~n23282 ;
  assign n23284 = ~n23268 & ~n23283 ;
  assign n23285 = \u2_L2_reg[23]/NET0131  & ~n23284 ;
  assign n23286 = ~\u2_L2_reg[23]/NET0131  & n23284 ;
  assign n23287 = ~n23285 & ~n23286 ;
  assign n23289 = ~n23020 & ~n23043 ;
  assign n23290 = ~n23046 & n23289 ;
  assign n23291 = ~n23032 & ~n23034 ;
  assign n23292 = ~n23290 & n23291 ;
  assign n23293 = n23001 & ~n23292 ;
  assign n23294 = ~n23041 & ~n23044 ;
  assign n23295 = ~n23001 & ~n23294 ;
  assign n23288 = n23007 & n23065 ;
  assign n23296 = n23021 & n23027 ;
  assign n23297 = ~n23288 & ~n23296 ;
  assign n23298 = ~n23295 & n23297 ;
  assign n23299 = ~n23293 & n23298 ;
  assign n23300 = n23060 & ~n23299 ;
  assign n23310 = ~n23084 & ~n23296 ;
  assign n23311 = n23034 & n23065 ;
  assign n23312 = n23310 & ~n23311 ;
  assign n23313 = n23001 & ~n23312 ;
  assign n23302 = n23001 & ~n23043 ;
  assign n23301 = ~n23001 & ~n23040 ;
  assign n23303 = ~n23020 & ~n23301 ;
  assign n23304 = ~n23302 & n23303 ;
  assign n23305 = n23001 & ~n23031 ;
  assign n23306 = ~n23027 & n23076 ;
  assign n23307 = ~n23305 & n23306 ;
  assign n23308 = ~n23304 & ~n23307 ;
  assign n23309 = ~n23060 & ~n23308 ;
  assign n23314 = n23040 & n23073 ;
  assign n23315 = ~n23033 & ~n23314 ;
  assign n23316 = ~n23309 & n23315 ;
  assign n23317 = ~n23313 & n23316 ;
  assign n23318 = ~n23300 & n23317 ;
  assign n23319 = ~\u2_L2_reg[25]/NET0131  & ~n23318 ;
  assign n23320 = \u2_L2_reg[25]/NET0131  & n23318 ;
  assign n23321 = ~n23319 & ~n23320 ;
  assign n23322 = ~n22743 & n22894 ;
  assign n23323 = ~n22685 & n22750 ;
  assign n23324 = ~n22721 & ~n23323 ;
  assign n23325 = ~n22708 & ~n23324 ;
  assign n23326 = ~n22904 & ~n23199 ;
  assign n23327 = ~n22730 & ~n23326 ;
  assign n23328 = ~n22679 & ~n23327 ;
  assign n23329 = ~n23325 & n23328 ;
  assign n23330 = ~n23322 & ~n23329 ;
  assign n23331 = n22712 & n22715 ;
  assign n23338 = ~n22700 & n22730 ;
  assign n23339 = ~n23331 & n23338 ;
  assign n23340 = ~n23194 & n23339 ;
  assign n23332 = ~n22738 & ~n23196 ;
  assign n23333 = n22708 & ~n23332 ;
  assign n23334 = n22701 & ~n22708 ;
  assign n23335 = ~n22720 & ~n23334 ;
  assign n23336 = ~n22679 & ~n22723 ;
  assign n23337 = ~n23335 & n23336 ;
  assign n23341 = ~n23333 & ~n23337 ;
  assign n23342 = n23340 & n23341 ;
  assign n23343 = n22698 & n22718 ;
  assign n23344 = ~n22737 & n23343 ;
  assign n23345 = ~n22730 & ~n23176 ;
  assign n23346 = n22744 & n23345 ;
  assign n23347 = ~n23344 & n23346 ;
  assign n23348 = ~n23342 & ~n23347 ;
  assign n23349 = ~n23330 & ~n23348 ;
  assign n23350 = ~\u2_L2_reg[26]/NET0131  & ~n23349 ;
  assign n23351 = \u2_L2_reg[26]/NET0131  & n23349 ;
  assign n23352 = ~n23350 & ~n23351 ;
  assign n23355 = n22815 & n22853 ;
  assign n23356 = ~n22837 & n22878 ;
  assign n23357 = ~n23355 & ~n23356 ;
  assign n23358 = n22844 & n23357 ;
  assign n23362 = n22829 & ~n22983 ;
  assign n23359 = ~n22829 & n22845 ;
  assign n23360 = ~n22844 & ~n22959 ;
  assign n23361 = ~n23359 & n23360 ;
  assign n23363 = ~n22830 & n23361 ;
  assign n23364 = ~n23362 & n23363 ;
  assign n23365 = ~n23358 & ~n23364 ;
  assign n23353 = n22837 & ~n22867 ;
  assign n23354 = ~n22972 & n23353 ;
  assign n23366 = ~n22809 & ~n23354 ;
  assign n23367 = ~n23365 & n23366 ;
  assign n23371 = n23357 & n23361 ;
  assign n23372 = ~n22821 & ~n22869 ;
  assign n23373 = n22854 & ~n23372 ;
  assign n23374 = n22844 & ~n22867 ;
  assign n23375 = ~n23373 & n23374 ;
  assign n23376 = ~n23371 & ~n23375 ;
  assign n23368 = ~n22823 & ~n22844 ;
  assign n23369 = n22829 & ~n22837 ;
  assign n23370 = ~n23368 & n23369 ;
  assign n23377 = n22809 & ~n22961 ;
  assign n23378 = ~n23370 & n23377 ;
  assign n23379 = ~n23376 & n23378 ;
  assign n23380 = ~n23367 & ~n23379 ;
  assign n23381 = ~\u2_L2_reg[28]/NET0131  & n23380 ;
  assign n23382 = \u2_L2_reg[28]/NET0131  & ~n23380 ;
  assign n23383 = ~n23381 & ~n23382 ;
  assign n23387 = n22474 & n22538 ;
  assign n23388 = ~n22523 & ~n23387 ;
  assign n23389 = ~n22530 & n23388 ;
  assign n23390 = n22462 & ~n23389 ;
  assign n23384 = n22487 & n22515 ;
  assign n23385 = ~n22794 & ~n23384 ;
  assign n23386 = ~n22462 & ~n23385 ;
  assign n23391 = n22492 & n22497 ;
  assign n23392 = ~n22489 & ~n23391 ;
  assign n23393 = ~n23386 & n23392 ;
  assign n23394 = ~n23390 & n23393 ;
  assign n23395 = ~n22513 & ~n23394 ;
  assign n23399 = n22462 & n22492 ;
  assign n23400 = ~n23384 & ~n23399 ;
  assign n23401 = ~n22481 & ~n23400 ;
  assign n23396 = ~n22474 & n22517 ;
  assign n23397 = ~n22538 & ~n23396 ;
  assign n23398 = ~n22462 & ~n23397 ;
  assign n23402 = n22481 & n22501 ;
  assign n23403 = ~n23398 & ~n23402 ;
  assign n23404 = ~n23401 & n23403 ;
  assign n23405 = n22513 & ~n23404 ;
  assign n23406 = n22481 & n22787 ;
  assign n23407 = ~n22462 & ~n22516 ;
  assign n23408 = ~n23406 & n23407 ;
  assign n23409 = ~n22502 & ~n22521 ;
  assign n23410 = ~n22523 & n23409 ;
  assign n23411 = n22462 & n22481 ;
  assign n23412 = ~n23410 & n23411 ;
  assign n23413 = ~n23408 & ~n23412 ;
  assign n23414 = ~n23405 & n23413 ;
  assign n23415 = ~n23395 & n23414 ;
  assign n23416 = ~\u2_L2_reg[4]/NET0131  & ~n23415 ;
  assign n23417 = \u2_L2_reg[4]/NET0131  & n23415 ;
  assign n23418 = ~n23416 & ~n23417 ;
  assign n23419 = ~n22462 & n22468 ;
  assign n23420 = ~n23387 & ~n23419 ;
  assign n23421 = ~n22487 & ~n23420 ;
  assign n23425 = n22513 & ~n23396 ;
  assign n23426 = ~n23421 & n23425 ;
  assign n23422 = n22481 & ~n23409 ;
  assign n23423 = ~n22526 & ~n22533 ;
  assign n23424 = n22462 & ~n23423 ;
  assign n23427 = ~n23422 & ~n23424 ;
  assign n23428 = n23426 & n23427 ;
  assign n23431 = n22468 & ~n22517 ;
  assign n23432 = ~n23384 & ~n23431 ;
  assign n23433 = n22462 & ~n23432 ;
  assign n23430 = ~n22462 & ~n23409 ;
  assign n23429 = n22481 & n22493 ;
  assign n23434 = ~n22513 & ~n23429 ;
  assign n23435 = ~n23430 & n23434 ;
  assign n23436 = ~n23433 & n23435 ;
  assign n23437 = ~n23428 & ~n23436 ;
  assign n23438 = ~n22487 & n23391 ;
  assign n23439 = ~n22529 & ~n23438 ;
  assign n23440 = ~n23437 & n23439 ;
  assign n23441 = ~\u2_L2_reg[19]/NET0131  & ~n23440 ;
  assign n23442 = \u2_L2_reg[19]/NET0131  & n23440 ;
  assign n23443 = ~n23441 & ~n23442 ;
  assign n23444 = ~n23118 & ~n23230 ;
  assign n23445 = n23124 & ~n23444 ;
  assign n23446 = ~n23247 & ~n23445 ;
  assign n23447 = ~n23134 & ~n23446 ;
  assign n23453 = ~n23166 & ~n23236 ;
  assign n23448 = n23108 & n23127 ;
  assign n23449 = n23102 & n23448 ;
  assign n23450 = n23124 & n23134 ;
  assign n23451 = ~n23109 & n23450 ;
  assign n23452 = n23444 & n23451 ;
  assign n23454 = ~n23449 & ~n23452 ;
  assign n23455 = n23453 & n23454 ;
  assign n23456 = ~n23447 & n23455 ;
  assign n23457 = n23141 & ~n23456 ;
  assign n23460 = ~n23143 & n23209 ;
  assign n23459 = n23117 & ~n23216 ;
  assign n23461 = n23134 & ~n23459 ;
  assign n23462 = ~n23460 & n23461 ;
  assign n23464 = n23108 & n23151 ;
  assign n23463 = n23144 & n23217 ;
  assign n23465 = ~n23211 & ~n23463 ;
  assign n23466 = ~n23464 & n23465 ;
  assign n23467 = ~n23462 & n23466 ;
  assign n23468 = ~n23141 & ~n23467 ;
  assign n23473 = n23124 & n23231 ;
  assign n23474 = ~n23134 & n23473 ;
  assign n23458 = n23134 & n23448 ;
  assign n23469 = ~n23110 & ~n23209 ;
  assign n23470 = ~n23216 & ~n23230 ;
  assign n23471 = ~n23469 & n23470 ;
  assign n23472 = ~n23134 & n23471 ;
  assign n23475 = ~n23458 & ~n23472 ;
  assign n23476 = ~n23474 & n23475 ;
  assign n23477 = ~n23468 & n23476 ;
  assign n23478 = ~n23457 & n23477 ;
  assign n23479 = ~\u2_L2_reg[27]/NET0131  & ~n23478 ;
  assign n23480 = \u2_L2_reg[27]/NET0131  & n23478 ;
  assign n23481 = ~n23479 & ~n23480 ;
  assign n23486 = ~n22596 & n22926 ;
  assign n23487 = n22943 & n23486 ;
  assign n23485 = n22596 & ~n22943 ;
  assign n23488 = ~n22563 & ~n23485 ;
  assign n23489 = ~n23487 & n23488 ;
  assign n23492 = n22563 & ~n22600 ;
  assign n23490 = ~n22570 & n22631 ;
  assign n23491 = n22576 & n22942 ;
  assign n23493 = ~n23490 & ~n23491 ;
  assign n23494 = n23492 & n23493 ;
  assign n23495 = ~n23489 & ~n23494 ;
  assign n23496 = n22628 & n22942 ;
  assign n23497 = n22586 & ~n23496 ;
  assign n23498 = ~n23495 & n23497 ;
  assign n23499 = n22557 & ~n22932 ;
  assign n23503 = ~n22586 & n22630 ;
  assign n23504 = ~n23499 & n23503 ;
  assign n23500 = n22927 & ~n22931 ;
  assign n23501 = ~n22607 & ~n22931 ;
  assign n23502 = n22563 & ~n23501 ;
  assign n23505 = ~n23500 & ~n23502 ;
  assign n23506 = n23504 & n23505 ;
  assign n23507 = ~n23498 & ~n23506 ;
  assign n23482 = n22564 & ~n22942 ;
  assign n23483 = ~n22579 & n23482 ;
  assign n23484 = n22563 & n22595 ;
  assign n23508 = ~n23483 & ~n23484 ;
  assign n23509 = ~n23507 & n23508 ;
  assign n23510 = \u2_L2_reg[32]/NET0131  & n23509 ;
  assign n23511 = ~\u2_L2_reg[32]/NET0131  & ~n23509 ;
  assign n23512 = ~n23510 & ~n23511 ;
  assign n23513 = decrypt_pad & ~\u2_uk_K_r2_reg[20]/NET0131  ;
  assign n23514 = ~decrypt_pad & ~\u2_uk_K_r2_reg[40]/NET0131  ;
  assign n23515 = ~n23513 & ~n23514 ;
  assign n23516 = \u2_R2_reg[13]/NET0131  & ~n23515 ;
  assign n23517 = ~\u2_R2_reg[13]/NET0131  & n23515 ;
  assign n23518 = ~n23516 & ~n23517 ;
  assign n23526 = decrypt_pad & ~\u2_uk_K_r2_reg[40]/NET0131  ;
  assign n23527 = ~decrypt_pad & ~\u2_uk_K_r2_reg[3]/NET0131  ;
  assign n23528 = ~n23526 & ~n23527 ;
  assign n23529 = \u2_R2_reg[9]/NET0131  & ~n23528 ;
  assign n23530 = ~\u2_R2_reg[9]/NET0131  & n23528 ;
  assign n23531 = ~n23529 & ~n23530 ;
  assign n23540 = ~n23518 & n23531 ;
  assign n23541 = decrypt_pad & ~\u2_uk_K_r2_reg[17]/NET0131  ;
  assign n23542 = ~decrypt_pad & ~\u2_uk_K_r2_reg[12]/NET0131  ;
  assign n23543 = ~n23541 & ~n23542 ;
  assign n23544 = \u2_R2_reg[11]/NET0131  & ~n23543 ;
  assign n23545 = ~\u2_R2_reg[11]/NET0131  & n23543 ;
  assign n23546 = ~n23544 & ~n23545 ;
  assign n23547 = ~n23540 & ~n23546 ;
  assign n23532 = decrypt_pad & ~\u2_uk_K_r2_reg[48]/NET0131  ;
  assign n23533 = ~decrypt_pad & ~\u2_uk_K_r2_reg[11]/NET0131  ;
  assign n23534 = ~n23532 & ~n23533 ;
  assign n23535 = \u2_R2_reg[10]/NET0131  & ~n23534 ;
  assign n23536 = ~\u2_R2_reg[10]/NET0131  & n23534 ;
  assign n23537 = ~n23535 & ~n23536 ;
  assign n23548 = n23531 & ~n23537 ;
  assign n23519 = decrypt_pad & ~\u2_uk_K_r2_reg[11]/NET0131  ;
  assign n23520 = ~decrypt_pad & ~\u2_uk_K_r2_reg[6]/NET0131  ;
  assign n23521 = ~n23519 & ~n23520 ;
  assign n23522 = \u2_R2_reg[8]/NET0131  & ~n23521 ;
  assign n23523 = ~\u2_R2_reg[8]/NET0131  & n23521 ;
  assign n23524 = ~n23522 & ~n23523 ;
  assign n23549 = n23518 & ~n23531 ;
  assign n23550 = n23524 & ~n23549 ;
  assign n23551 = ~n23548 & ~n23550 ;
  assign n23552 = n23547 & ~n23551 ;
  assign n23525 = ~n23518 & ~n23524 ;
  assign n23538 = n23531 & n23537 ;
  assign n23539 = n23525 & n23538 ;
  assign n23553 = decrypt_pad & ~\u2_uk_K_r2_reg[32]/NET0131  ;
  assign n23554 = ~decrypt_pad & ~\u2_uk_K_r2_reg[27]/NET0131  ;
  assign n23555 = ~n23553 & ~n23554 ;
  assign n23556 = \u2_R2_reg[12]/NET0131  & ~n23555 ;
  assign n23557 = ~\u2_R2_reg[12]/NET0131  & n23555 ;
  assign n23558 = ~n23556 & ~n23557 ;
  assign n23559 = ~n23539 & n23558 ;
  assign n23560 = ~n23552 & n23559 ;
  assign n23565 = n23518 & n23524 ;
  assign n23566 = ~n23525 & ~n23565 ;
  assign n23567 = ~n23531 & ~n23537 ;
  assign n23570 = ~n23566 & ~n23567 ;
  assign n23571 = ~n23538 & n23570 ;
  assign n23573 = n23524 & n23537 ;
  assign n23574 = n23540 & n23573 ;
  assign n23564 = ~n23524 & n23546 ;
  assign n23572 = n23548 & n23564 ;
  assign n23575 = ~n23558 & ~n23572 ;
  assign n23576 = ~n23574 & n23575 ;
  assign n23561 = n23518 & ~n23524 ;
  assign n23562 = n23538 & n23561 ;
  assign n23563 = ~n23546 & n23562 ;
  assign n23568 = ~n23564 & n23567 ;
  assign n23569 = n23566 & n23568 ;
  assign n23577 = ~n23563 & ~n23569 ;
  assign n23578 = n23576 & n23577 ;
  assign n23579 = ~n23571 & n23578 ;
  assign n23580 = ~n23560 & ~n23579 ;
  assign n23582 = ~n23524 & ~n23537 ;
  assign n23583 = n23524 & ~n23531 ;
  assign n23584 = ~n23582 & ~n23583 ;
  assign n23585 = n23566 & n23584 ;
  assign n23586 = ~n23549 & ~n23585 ;
  assign n23587 = n23558 & ~n23586 ;
  assign n23581 = n23537 & n23549 ;
  assign n23588 = n23525 & ~n23537 ;
  assign n23589 = ~n23531 & n23588 ;
  assign n23590 = ~n23581 & ~n23589 ;
  assign n23591 = ~n23587 & n23590 ;
  assign n23592 = n23546 & ~n23591 ;
  assign n23593 = ~n23580 & ~n23592 ;
  assign n23594 = ~\u2_L2_reg[6]/NET0131  & ~n23593 ;
  assign n23595 = \u2_L2_reg[6]/NET0131  & n23593 ;
  assign n23596 = ~n23594 & ~n23595 ;
  assign n23611 = n23001 & ~n23030 ;
  assign n23612 = ~n23032 & n23611 ;
  assign n23599 = n23020 & ~n23027 ;
  assign n23613 = ~n23075 & n23599 ;
  assign n23614 = ~n23001 & ~n23041 ;
  assign n23615 = ~n23613 & n23614 ;
  assign n23616 = ~n23612 & ~n23615 ;
  assign n23617 = ~n23044 & n23310 ;
  assign n23618 = ~n23616 & n23617 ;
  assign n23619 = ~n23060 & ~n23618 ;
  assign n23597 = n23013 & n23029 ;
  assign n23598 = ~n23001 & ~n23597 ;
  assign n23600 = n23001 & ~n23599 ;
  assign n23601 = ~n23076 & ~n23600 ;
  assign n23602 = ~n23021 & ~n23601 ;
  assign n23603 = ~n23598 & ~n23602 ;
  assign n23604 = ~n23013 & n23070 ;
  assign n23605 = ~n23041 & ~n23604 ;
  assign n23606 = n23001 & ~n23605 ;
  assign n23607 = n23027 & n23067 ;
  assign n23608 = n23089 & ~n23607 ;
  assign n23609 = ~n23606 & n23608 ;
  assign n23610 = n23060 & ~n23609 ;
  assign n23620 = ~n23603 & ~n23610 ;
  assign n23621 = ~n23619 & n23620 ;
  assign n23622 = ~\u2_L2_reg[8]/NET0131  & ~n23621 ;
  assign n23623 = \u2_L2_reg[8]/NET0131  & n23621 ;
  assign n23624 = ~n23622 & ~n23623 ;
  assign n23625 = n22557 & ~n22943 ;
  assign n23626 = ~n22607 & ~n23625 ;
  assign n23627 = n22576 & ~n23626 ;
  assign n23628 = ~n22576 & ~n22631 ;
  assign n23629 = n22943 & n23628 ;
  assign n23630 = n22563 & ~n23629 ;
  assign n23631 = ~n22570 & ~n22924 ;
  assign n23632 = ~n22563 & ~n23491 ;
  assign n23633 = ~n23625 & n23632 ;
  assign n23634 = ~n23631 & n23633 ;
  assign n23635 = ~n23630 & ~n23634 ;
  assign n23636 = ~n23627 & ~n23635 ;
  assign n23637 = n22586 & ~n23636 ;
  assign n23641 = n22628 & ~n22943 ;
  assign n23639 = n22576 & ~n22606 ;
  assign n23640 = n22943 & ~n23639 ;
  assign n23642 = ~n22586 & ~n23640 ;
  assign n23643 = ~n23641 & n23642 ;
  assign n23644 = ~n22615 & ~n23643 ;
  assign n23645 = n22563 & ~n23644 ;
  assign n23638 = ~n22563 & n23627 ;
  assign n23646 = ~n22563 & n23629 ;
  assign n23647 = ~n22615 & ~n23646 ;
  assign n23648 = ~n22586 & ~n23647 ;
  assign n23649 = ~n23638 & ~n23648 ;
  assign n23650 = ~n23645 & n23649 ;
  assign n23651 = ~n23637 & n23650 ;
  assign n23652 = ~\u2_L2_reg[7]/NET0131  & ~n23651 ;
  assign n23653 = \u2_L2_reg[7]/NET0131  & n23651 ;
  assign n23654 = ~n23652 & ~n23653 ;
  assign n23668 = ~n22644 & ~n23255 ;
  assign n23669 = n22382 & ~n23668 ;
  assign n23657 = ~n22402 & ~n22643 ;
  assign n23670 = n22420 & n23657 ;
  assign n23671 = ~n22658 & ~n23670 ;
  assign n23672 = ~n23669 & n23671 ;
  assign n23673 = n22416 & ~n23672 ;
  assign n23658 = ~n22399 & n23657 ;
  assign n23655 = n22399 & n22643 ;
  assign n23656 = ~n22657 & n23655 ;
  assign n23659 = ~n22403 & n22407 ;
  assign n23660 = n22642 & n22656 ;
  assign n23661 = ~n23659 & ~n23660 ;
  assign n23662 = ~n23656 & n23661 ;
  assign n23663 = ~n23658 & n23662 ;
  assign n23664 = ~n22416 & ~n23663 ;
  assign n23665 = ~n22391 & n22655 ;
  assign n23666 = ~n23660 & ~n23665 ;
  assign n23667 = ~n22399 & ~n23666 ;
  assign n23674 = ~n23664 & ~n23667 ;
  assign n23675 = ~n23673 & n23674 ;
  assign n23676 = ~\u2_L2_reg[9]/NET0131  & ~n23675 ;
  assign n23677 = \u2_L2_reg[9]/NET0131  & n23675 ;
  assign n23678 = ~n23676 & ~n23677 ;
  assign n23681 = n23531 & ~n23565 ;
  assign n23682 = ~n23531 & n23565 ;
  assign n23683 = ~n23681 & ~n23682 ;
  assign n23684 = ~n23525 & n23683 ;
  assign n23685 = n23540 & n23564 ;
  assign n23686 = ~n23684 & ~n23685 ;
  assign n23687 = ~n23537 & ~n23686 ;
  assign n23688 = ~n23546 & ~n23573 ;
  assign n23689 = ~n23518 & ~n23582 ;
  assign n23690 = n23688 & n23689 ;
  assign n23691 = ~n23562 & ~n23690 ;
  assign n23692 = ~n23687 & n23691 ;
  assign n23693 = n23558 & ~n23692 ;
  assign n23694 = ~n23525 & n23546 ;
  assign n23695 = ~n23683 & n23694 ;
  assign n23696 = n23546 & ~n23589 ;
  assign n23697 = ~n23531 & ~n23561 ;
  assign n23698 = ~n23681 & ~n23697 ;
  assign n23699 = ~n23588 & ~n23698 ;
  assign n23700 = ~n23696 & ~n23699 ;
  assign n23701 = ~n23695 & ~n23700 ;
  assign n23702 = ~n23558 & ~n23701 ;
  assign n23679 = ~n23546 & n23573 ;
  assign n23680 = ~n23531 & n23679 ;
  assign n23703 = n23525 & n23537 ;
  assign n23704 = ~n23531 & n23703 ;
  assign n23705 = ~n23574 & ~n23704 ;
  assign n23706 = n23546 & ~n23705 ;
  assign n23707 = ~n23680 & ~n23706 ;
  assign n23708 = ~n23702 & n23707 ;
  assign n23709 = ~n23693 & n23708 ;
  assign n23710 = ~\u2_L2_reg[16]/NET0131  & ~n23709 ;
  assign n23711 = \u2_L2_reg[16]/NET0131  & n23709 ;
  assign n23712 = ~n23710 & ~n23711 ;
  assign n23716 = ~n22867 & ~n22872 ;
  assign n23717 = ~n22844 & ~n23716 ;
  assign n23714 = n22845 & n22878 ;
  assign n23715 = ~n22831 & n22844 ;
  assign n23718 = ~n23714 & ~n23715 ;
  assign n23719 = ~n23717 & n23718 ;
  assign n23720 = n22809 & ~n23719 ;
  assign n23722 = ~n22856 & ~n22870 ;
  assign n23723 = n22877 & n23722 ;
  assign n23724 = ~n22847 & ~n22959 ;
  assign n23721 = n22846 & n22870 ;
  assign n23725 = ~n22979 & ~n23721 ;
  assign n23726 = n23724 & n23725 ;
  assign n23727 = ~n23723 & n23726 ;
  assign n23728 = ~n22809 & ~n23727 ;
  assign n23713 = ~n22844 & n23355 ;
  assign n23729 = n22821 & n22849 ;
  assign n23730 = ~n22985 & ~n23729 ;
  assign n23731 = n22844 & ~n23730 ;
  assign n23732 = ~n23713 & ~n23731 ;
  assign n23733 = ~n23728 & n23732 ;
  assign n23734 = ~n23720 & n23733 ;
  assign n23735 = ~\u2_L2_reg[18]/P0001  & ~n23734 ;
  assign n23736 = \u2_L2_reg[18]/P0001  & n23734 ;
  assign n23737 = ~n23735 & ~n23736 ;
  assign n23745 = ~n23537 & n23561 ;
  assign n23746 = ~n23703 & ~n23745 ;
  assign n23747 = n23537 & n23583 ;
  assign n23744 = n23525 & n23531 ;
  assign n23748 = n23546 & ~n23744 ;
  assign n23749 = ~n23747 & n23748 ;
  assign n23750 = n23746 & n23749 ;
  assign n23753 = ~n23566 & n23567 ;
  assign n23751 = ~n23537 & ~n23540 ;
  assign n23752 = n23566 & ~n23751 ;
  assign n23754 = ~n23546 & ~n23752 ;
  assign n23755 = ~n23753 & n23754 ;
  assign n23756 = ~n23750 & ~n23755 ;
  assign n23757 = ~n23558 & ~n23756 ;
  assign n23758 = ~n23546 & n23570 ;
  assign n23762 = n23558 & ~n23569 ;
  assign n23759 = n23537 & ~n23583 ;
  assign n23760 = n23694 & n23759 ;
  assign n23740 = ~n23537 & n23546 ;
  assign n23761 = n23697 & n23740 ;
  assign n23763 = ~n23760 & ~n23761 ;
  assign n23764 = n23762 & n23763 ;
  assign n23765 = ~n23758 & n23764 ;
  assign n23766 = ~n23757 & ~n23765 ;
  assign n23738 = n23518 & n23531 ;
  assign n23739 = ~n23583 & ~n23738 ;
  assign n23741 = ~n23565 & n23740 ;
  assign n23742 = ~n23739 & n23741 ;
  assign n23743 = n23679 & n23738 ;
  assign n23767 = ~n23742 & ~n23743 ;
  assign n23768 = ~n23766 & n23767 ;
  assign n23769 = ~\u2_L2_reg[24]/NET0131  & ~n23768 ;
  assign n23770 = \u2_L2_reg[24]/NET0131  & n23768 ;
  assign n23771 = ~n23769 & ~n23770 ;
  assign n23788 = ~n23540 & n23573 ;
  assign n23783 = ~n23518 & ~n23537 ;
  assign n23787 = n23531 & n23783 ;
  assign n23789 = ~n23558 & ~n23787 ;
  assign n23790 = ~n23788 & n23789 ;
  assign n23784 = n23583 & n23783 ;
  assign n23785 = n23558 & ~n23784 ;
  assign n23786 = n23746 & n23785 ;
  assign n23791 = n23546 & ~n23786 ;
  assign n23792 = ~n23790 & n23791 ;
  assign n23773 = ~n23573 & ~n23744 ;
  assign n23774 = ~n23546 & ~n23773 ;
  assign n23772 = n23537 & n23681 ;
  assign n23775 = n23558 & ~n23772 ;
  assign n23776 = ~n23774 & n23775 ;
  assign n23779 = ~n23558 & ~n23753 ;
  assign n23777 = ~n23524 & n23581 ;
  assign n23778 = n23688 & ~n23739 ;
  assign n23780 = ~n23777 & ~n23778 ;
  assign n23781 = n23779 & n23780 ;
  assign n23782 = ~n23776 & ~n23781 ;
  assign n23793 = n23546 & ~n23682 ;
  assign n23794 = n23537 & ~n23547 ;
  assign n23795 = ~n23793 & n23794 ;
  assign n23796 = ~n23782 & ~n23795 ;
  assign n23797 = ~n23792 & n23796 ;
  assign n23798 = \u2_L2_reg[30]/NET0131  & ~n23797 ;
  assign n23799 = ~\u2_L2_reg[30]/NET0131  & n23797 ;
  assign n23800 = ~n23798 & ~n23799 ;
  assign n23804 = n23001 & ~n23075 ;
  assign n23805 = ~n23028 & ~n23065 ;
  assign n23806 = ~n23041 & ~n23805 ;
  assign n23807 = ~n23804 & ~n23806 ;
  assign n23801 = ~n23027 & n23065 ;
  assign n23802 = ~n23062 & ~n23801 ;
  assign n23803 = n23001 & ~n23802 ;
  assign n23808 = ~n23060 & ~n23803 ;
  assign n23809 = ~n23807 & n23808 ;
  assign n23810 = n23027 & ~n23065 ;
  assign n23811 = ~n23034 & n23600 ;
  assign n23812 = ~n23810 & n23811 ;
  assign n23814 = ~n23033 & n23060 ;
  assign n23813 = ~n23001 & n23068 ;
  assign n23815 = ~n23597 & ~n23813 ;
  assign n23816 = n23814 & n23815 ;
  assign n23817 = ~n23812 & n23816 ;
  assign n23818 = ~n23809 & ~n23817 ;
  assign n23819 = ~n23087 & n23611 ;
  assign n23820 = ~n23001 & ~n23042 ;
  assign n23821 = ~n23083 & ~n23604 ;
  assign n23822 = n23820 & n23821 ;
  assign n23823 = ~n23819 & ~n23822 ;
  assign n23824 = ~n23818 & ~n23823 ;
  assign n23825 = ~\u2_L2_reg[3]/NET0131  & ~n23824 ;
  assign n23826 = \u2_L2_reg[3]/NET0131  & n23824 ;
  assign n23827 = ~n23825 & ~n23826 ;
  assign n23828 = decrypt_pad & ~\u2_uk_K_r1_reg[49]/NET0131  ;
  assign n23829 = ~decrypt_pad & ~\u2_uk_K_r1_reg[43]/NET0131  ;
  assign n23830 = ~n23828 & ~n23829 ;
  assign n23831 = \u2_R1_reg[26]/NET0131  & ~n23830 ;
  assign n23832 = ~\u2_R1_reg[26]/NET0131  & n23830 ;
  assign n23833 = ~n23831 & ~n23832 ;
  assign n23834 = decrypt_pad & ~\u2_uk_K_r1_reg[9]/NET0131  ;
  assign n23835 = ~decrypt_pad & ~\u2_uk_K_r1_reg[31]/NET0131  ;
  assign n23836 = ~n23834 & ~n23835 ;
  assign n23837 = \u2_R1_reg[25]/NET0131  & ~n23836 ;
  assign n23838 = ~\u2_R1_reg[25]/NET0131  & n23836 ;
  assign n23839 = ~n23837 & ~n23838 ;
  assign n23840 = n23833 & ~n23839 ;
  assign n23841 = decrypt_pad & ~\u2_uk_K_r1_reg[29]/NET0131  ;
  assign n23842 = ~decrypt_pad & ~\u2_uk_K_r1_reg[23]/NET0131  ;
  assign n23843 = ~n23841 & ~n23842 ;
  assign n23844 = \u2_R1_reg[24]/NET0131  & ~n23843 ;
  assign n23845 = ~\u2_R1_reg[24]/NET0131  & n23843 ;
  assign n23846 = ~n23844 & ~n23845 ;
  assign n23847 = decrypt_pad & ~\u2_uk_K_r1_reg[37]/NET0131  ;
  assign n23848 = ~decrypt_pad & ~\u2_uk_K_r1_reg[0]/NET0131  ;
  assign n23849 = ~n23847 & ~n23848 ;
  assign n23850 = \u2_R1_reg[29]/NET0131  & ~n23849 ;
  assign n23851 = ~\u2_R1_reg[29]/NET0131  & n23849 ;
  assign n23852 = ~n23850 & ~n23851 ;
  assign n23853 = ~n23846 & n23852 ;
  assign n23854 = n23840 & n23853 ;
  assign n23855 = ~n23846 & ~n23852 ;
  assign n23856 = n23833 & n23855 ;
  assign n23857 = n23839 & n23856 ;
  assign n23858 = ~n23854 & ~n23857 ;
  assign n23859 = ~n23839 & ~n23852 ;
  assign n23860 = n23839 & n23852 ;
  assign n23861 = ~n23833 & n23860 ;
  assign n23862 = ~n23840 & ~n23861 ;
  assign n23863 = decrypt_pad & ~\u2_uk_K_r1_reg[14]/NET0131  ;
  assign n23864 = ~decrypt_pad & ~\u2_uk_K_r1_reg[8]/NET0131  ;
  assign n23865 = ~n23863 & ~n23864 ;
  assign n23866 = \u2_R1_reg[28]/NET0131  & ~n23865 ;
  assign n23867 = ~\u2_R1_reg[28]/NET0131  & n23865 ;
  assign n23868 = ~n23866 & ~n23867 ;
  assign n23869 = ~n23862 & n23868 ;
  assign n23870 = ~n23859 & ~n23869 ;
  assign n23871 = n23846 & ~n23870 ;
  assign n23872 = n23858 & ~n23871 ;
  assign n23873 = decrypt_pad & ~\u2_uk_K_r1_reg[31]/NET0131  ;
  assign n23874 = ~decrypt_pad & ~\u2_uk_K_r1_reg[21]/NET0131  ;
  assign n23875 = ~n23873 & ~n23874 ;
  assign n23876 = \u2_R1_reg[27]/NET0131  & ~n23875 ;
  assign n23877 = ~\u2_R1_reg[27]/NET0131  & n23875 ;
  assign n23878 = ~n23876 & ~n23877 ;
  assign n23879 = ~n23872 & n23878 ;
  assign n23880 = ~n23839 & n23878 ;
  assign n23881 = ~n23833 & n23880 ;
  assign n23882 = ~n23852 & ~n23878 ;
  assign n23883 = ~n23840 & n23882 ;
  assign n23884 = ~n23881 & ~n23883 ;
  assign n23885 = n23846 & ~n23884 ;
  assign n23886 = ~n23833 & ~n23846 ;
  assign n23887 = n23833 & n23846 ;
  assign n23888 = ~n23886 & ~n23887 ;
  assign n23889 = n23852 & ~n23888 ;
  assign n23890 = ~n23839 & n23856 ;
  assign n23891 = ~n23889 & ~n23890 ;
  assign n23892 = ~n23880 & ~n23891 ;
  assign n23893 = ~n23885 & ~n23892 ;
  assign n23894 = ~n23868 & ~n23893 ;
  assign n23898 = n23846 & n23852 ;
  assign n23899 = ~n23833 & ~n23839 ;
  assign n23900 = n23898 & n23899 ;
  assign n23901 = ~n23846 & n23860 ;
  assign n23902 = ~n23900 & ~n23901 ;
  assign n23903 = ~n23878 & ~n23902 ;
  assign n23904 = n23855 & n23899 ;
  assign n23905 = ~n23854 & ~n23904 ;
  assign n23906 = ~n23903 & n23905 ;
  assign n23907 = n23868 & ~n23906 ;
  assign n23895 = ~n23852 & n23881 ;
  assign n23896 = n23839 & ~n23878 ;
  assign n23897 = ~n23888 & n23896 ;
  assign n23908 = ~n23895 & ~n23897 ;
  assign n23909 = ~n23907 & n23908 ;
  assign n23910 = ~n23894 & n23909 ;
  assign n23911 = ~n23879 & n23910 ;
  assign n23912 = ~\u2_L1_reg[22]/NET0131  & ~n23911 ;
  assign n23913 = \u2_L1_reg[22]/NET0131  & n23911 ;
  assign n23914 = ~n23912 & ~n23913 ;
  assign n23915 = decrypt_pad & ~\u2_uk_K_r1_reg[10]/P0001  ;
  assign n23916 = ~decrypt_pad & ~\u2_uk_K_r1_reg[34]/NET0131  ;
  assign n23917 = ~n23915 & ~n23916 ;
  assign n23918 = \u2_R1_reg[4]/NET0131  & ~n23917 ;
  assign n23919 = ~\u2_R1_reg[4]/NET0131  & n23917 ;
  assign n23920 = ~n23918 & ~n23919 ;
  assign n23948 = decrypt_pad & ~\u2_uk_K_r1_reg[32]/NET0131  ;
  assign n23949 = ~decrypt_pad & ~\u2_uk_K_r1_reg[24]/NET0131  ;
  assign n23950 = ~n23948 & ~n23949 ;
  assign n23951 = \u2_R1_reg[3]/NET0131  & ~n23950 ;
  assign n23952 = ~\u2_R1_reg[3]/NET0131  & n23950 ;
  assign n23953 = ~n23951 & ~n23952 ;
  assign n23921 = decrypt_pad & ~\u2_uk_K_r1_reg[55]/NET0131  ;
  assign n23922 = ~decrypt_pad & ~\u2_uk_K_r1_reg[47]/NET0131  ;
  assign n23923 = ~n23921 & ~n23922 ;
  assign n23924 = \u2_R1_reg[2]/NET0131  & ~n23923 ;
  assign n23925 = ~\u2_R1_reg[2]/NET0131  & n23923 ;
  assign n23926 = ~n23924 & ~n23925 ;
  assign n23941 = decrypt_pad & ~\u2_uk_K_r1_reg[19]/NET0131  ;
  assign n23942 = ~decrypt_pad & ~\u2_uk_K_r1_reg[11]/NET0131  ;
  assign n23943 = ~n23941 & ~n23942 ;
  assign n23944 = \u2_R1_reg[32]/NET0131  & ~n23943 ;
  assign n23945 = ~\u2_R1_reg[32]/NET0131  & n23943 ;
  assign n23946 = ~n23944 & ~n23945 ;
  assign n23927 = decrypt_pad & ~\u2_uk_K_r1_reg[40]/NET0131  ;
  assign n23928 = ~decrypt_pad & ~\u2_uk_K_r1_reg[32]/NET0131  ;
  assign n23929 = ~n23927 & ~n23928 ;
  assign n23930 = \u2_R1_reg[1]/NET0131  & ~n23929 ;
  assign n23931 = ~\u2_R1_reg[1]/NET0131  & n23929 ;
  assign n23932 = ~n23930 & ~n23931 ;
  assign n23934 = decrypt_pad & ~\u2_uk_K_r1_reg[13]/NET0131  ;
  assign n23935 = ~decrypt_pad & ~\u2_uk_K_r1_reg[5]/NET0131  ;
  assign n23936 = ~n23934 & ~n23935 ;
  assign n23937 = \u2_R1_reg[5]/NET0131  & ~n23936 ;
  assign n23938 = ~\u2_R1_reg[5]/NET0131  & n23936 ;
  assign n23939 = ~n23937 & ~n23938 ;
  assign n23955 = ~n23932 & ~n23939 ;
  assign n23956 = n23946 & n23955 ;
  assign n23957 = n23926 & n23956 ;
  assign n23958 = ~n23932 & n23939 ;
  assign n23959 = ~n23926 & ~n23946 ;
  assign n23960 = ~n23958 & n23959 ;
  assign n23961 = ~n23957 & ~n23960 ;
  assign n23962 = ~n23953 & ~n23961 ;
  assign n23963 = n23939 & ~n23946 ;
  assign n23964 = n23926 & n23953 ;
  assign n23965 = n23963 & n23964 ;
  assign n23966 = ~n23939 & n23959 ;
  assign n23967 = ~n23965 & ~n23966 ;
  assign n23968 = n23932 & ~n23967 ;
  assign n23933 = n23926 & n23932 ;
  assign n23940 = n23933 & ~n23939 ;
  assign n23947 = n23940 & n23946 ;
  assign n23954 = n23947 & n23953 ;
  assign n23969 = n23939 & n23946 ;
  assign n23970 = ~n23926 & n23953 ;
  assign n23971 = ~n23926 & ~n23932 ;
  assign n23972 = ~n23970 & ~n23971 ;
  assign n23973 = n23969 & ~n23972 ;
  assign n23974 = ~n23954 & ~n23973 ;
  assign n23975 = ~n23968 & n23974 ;
  assign n23976 = ~n23962 & n23975 ;
  assign n23977 = ~n23920 & ~n23976 ;
  assign n23988 = ~n23939 & ~n23946 ;
  assign n23989 = n23926 & n23988 ;
  assign n23992 = ~n23958 & ~n23989 ;
  assign n23993 = n23953 & ~n23992 ;
  assign n24002 = ~n23926 & n23956 ;
  assign n23994 = ~n23932 & ~n23946 ;
  assign n23995 = n23932 & n23946 ;
  assign n23996 = ~n23994 & ~n23995 ;
  assign n23997 = n23932 & n23953 ;
  assign n23998 = ~n23971 & ~n23997 ;
  assign n23999 = ~n23996 & n23998 ;
  assign n24000 = n23932 & ~n23970 ;
  assign n24001 = n23963 & ~n24000 ;
  assign n24003 = ~n23999 & ~n24001 ;
  assign n24004 = ~n24002 & n24003 ;
  assign n24005 = ~n23993 & n24004 ;
  assign n24006 = n23920 & ~n24005 ;
  assign n23978 = ~n23932 & n23963 ;
  assign n23979 = n23926 & n23978 ;
  assign n23980 = ~n23926 & ~n23939 ;
  assign n23981 = n23926 & n23969 ;
  assign n23982 = ~n23980 & ~n23981 ;
  assign n23983 = n23932 & ~n23982 ;
  assign n23984 = ~n23979 & ~n23983 ;
  assign n23985 = ~n23953 & ~n23984 ;
  assign n23986 = ~n23932 & n23953 ;
  assign n23987 = ~n23926 & n23946 ;
  assign n23990 = ~n23987 & ~n23989 ;
  assign n23991 = n23986 & ~n23990 ;
  assign n24007 = ~n23985 & ~n23991 ;
  assign n24008 = ~n24006 & n24007 ;
  assign n24009 = ~n23977 & n24008 ;
  assign n24010 = ~\u2_L1_reg[31]/NET0131  & ~n24009 ;
  assign n24011 = \u2_L1_reg[31]/NET0131  & n24009 ;
  assign n24012 = ~n24010 & ~n24011 ;
  assign n24064 = decrypt_pad & ~\u2_uk_K_r1_reg[7]/P0001  ;
  assign n24065 = ~decrypt_pad & ~\u2_uk_K_r1_reg[1]/NET0131  ;
  assign n24066 = ~n24064 & ~n24065 ;
  assign n24067 = \u2_R1_reg[24]/NET0131  & ~n24066 ;
  assign n24068 = ~\u2_R1_reg[24]/NET0131  & n24066 ;
  assign n24069 = ~n24067 & ~n24068 ;
  assign n24013 = decrypt_pad & ~\u2_uk_K_r1_reg[36]/NET0131  ;
  assign n24014 = ~decrypt_pad & ~\u2_uk_K_r1_reg[30]/NET0131  ;
  assign n24015 = ~n24013 & ~n24014 ;
  assign n24016 = \u2_R1_reg[23]/NET0131  & ~n24015 ;
  assign n24017 = ~\u2_R1_reg[23]/NET0131  & n24015 ;
  assign n24018 = ~n24016 & ~n24017 ;
  assign n24039 = decrypt_pad & ~\u2_uk_K_r1_reg[23]/NET0131  ;
  assign n24040 = ~decrypt_pad & ~\u2_uk_K_r1_reg[45]/NET0131  ;
  assign n24041 = ~n24039 & ~n24040 ;
  assign n24042 = \u2_R1_reg[22]/NET0131  & ~n24041 ;
  assign n24043 = ~\u2_R1_reg[22]/NET0131  & n24041 ;
  assign n24044 = ~n24042 & ~n24043 ;
  assign n24019 = decrypt_pad & ~\u2_uk_K_r1_reg[45]/NET0131  ;
  assign n24020 = ~decrypt_pad & ~\u2_uk_K_r1_reg[35]/NET0131  ;
  assign n24021 = ~n24019 & ~n24020 ;
  assign n24022 = \u2_R1_reg[20]/NET0131  & ~n24021 ;
  assign n24023 = ~\u2_R1_reg[20]/NET0131  & n24021 ;
  assign n24024 = ~n24022 & ~n24023 ;
  assign n24032 = decrypt_pad & ~\u2_uk_K_r1_reg[1]/NET0131  ;
  assign n24033 = ~decrypt_pad & ~\u2_uk_K_r1_reg[50]/NET0131  ;
  assign n24034 = ~n24032 & ~n24033 ;
  assign n24035 = \u2_R1_reg[21]/NET0131  & ~n24034 ;
  assign n24036 = ~\u2_R1_reg[21]/NET0131  & n24034 ;
  assign n24037 = ~n24035 & ~n24036 ;
  assign n24056 = n24024 & ~n24037 ;
  assign n24092 = n24044 & n24056 ;
  assign n24071 = ~n24024 & ~n24044 ;
  assign n24025 = decrypt_pad & ~\u2_uk_K_r1_reg[2]/NET0131  ;
  assign n24026 = ~decrypt_pad & ~\u2_uk_K_r1_reg[51]/NET0131  ;
  assign n24027 = ~n24025 & ~n24026 ;
  assign n24028 = \u2_R1_reg[25]/NET0131  & ~n24027 ;
  assign n24029 = ~\u2_R1_reg[25]/NET0131  & n24027 ;
  assign n24030 = ~n24028 & ~n24029 ;
  assign n24082 = ~n24024 & ~n24037 ;
  assign n24091 = n24030 & n24082 ;
  assign n24093 = ~n24071 & ~n24091 ;
  assign n24094 = ~n24092 & n24093 ;
  assign n24095 = n24018 & ~n24094 ;
  assign n24045 = n24037 & n24044 ;
  assign n24046 = ~n24024 & n24045 ;
  assign n24076 = n24037 & ~n24044 ;
  assign n24086 = n24024 & n24076 ;
  assign n24087 = ~n24046 & ~n24086 ;
  assign n24088 = ~n24018 & ~n24087 ;
  assign n24047 = n24024 & ~n24030 ;
  assign n24080 = ~n24018 & ~n24044 ;
  assign n24089 = ~n24076 & ~n24080 ;
  assign n24090 = n24047 & ~n24089 ;
  assign n24096 = n24030 & n24092 ;
  assign n24097 = ~n24090 & ~n24096 ;
  assign n24098 = ~n24088 & n24097 ;
  assign n24099 = ~n24095 & n24098 ;
  assign n24100 = ~n24069 & ~n24099 ;
  assign n24048 = ~n24037 & n24047 ;
  assign n24049 = ~n24044 & n24048 ;
  assign n24031 = n24024 & n24030 ;
  assign n24038 = n24031 & n24037 ;
  assign n24050 = ~n24038 & ~n24046 ;
  assign n24051 = ~n24049 & n24050 ;
  assign n24052 = n24018 & ~n24051 ;
  assign n24057 = n24030 & n24056 ;
  assign n24054 = n24030 & n24037 ;
  assign n24055 = ~n24024 & n24054 ;
  assign n24058 = ~n24044 & ~n24055 ;
  assign n24059 = ~n24057 & n24058 ;
  assign n24053 = n24031 & n24044 ;
  assign n24060 = ~n24018 & ~n24046 ;
  assign n24061 = ~n24053 & n24060 ;
  assign n24062 = ~n24059 & n24061 ;
  assign n24063 = ~n24052 & ~n24062 ;
  assign n24070 = ~n24063 & n24069 ;
  assign n24081 = n24037 & n24047 ;
  assign n24083 = ~n24030 & n24082 ;
  assign n24084 = ~n24081 & ~n24083 ;
  assign n24085 = n24080 & ~n24084 ;
  assign n24072 = n24030 & n24071 ;
  assign n24073 = ~n24037 & n24072 ;
  assign n24074 = n24018 & n24073 ;
  assign n24075 = ~n24024 & ~n24030 ;
  assign n24077 = n24075 & n24076 ;
  assign n24078 = ~n24053 & ~n24077 ;
  assign n24079 = n24018 & ~n24078 ;
  assign n24101 = ~n24074 & ~n24079 ;
  assign n24102 = ~n24085 & n24101 ;
  assign n24103 = ~n24070 & n24102 ;
  assign n24104 = ~n24100 & n24103 ;
  assign n24105 = ~\u2_L1_reg[11]/NET0131  & n24104 ;
  assign n24106 = \u2_L1_reg[11]/NET0131  & ~n24104 ;
  assign n24107 = ~n24105 & ~n24106 ;
  assign n24108 = decrypt_pad & ~\u2_uk_K_r1_reg[38]/NET0131  ;
  assign n24109 = ~decrypt_pad & ~\u2_uk_K_r1_reg[28]/NET0131  ;
  assign n24110 = ~n24108 & ~n24109 ;
  assign n24111 = \u2_R1_reg[32]/NET0131  & ~n24110 ;
  assign n24112 = ~\u2_R1_reg[32]/NET0131  & n24110 ;
  assign n24113 = ~n24111 & ~n24112 ;
  assign n24152 = decrypt_pad & ~\u2_uk_K_r1_reg[28]/NET0131  ;
  assign n24153 = ~decrypt_pad & ~\u2_uk_K_r1_reg[22]/NET0131  ;
  assign n24154 = ~n24152 & ~n24153 ;
  assign n24155 = \u2_R1_reg[31]/P0001  & ~n24154 ;
  assign n24156 = ~\u2_R1_reg[31]/P0001  & n24154 ;
  assign n24157 = ~n24155 & ~n24156 ;
  assign n24127 = decrypt_pad & ~\u2_uk_K_r1_reg[43]/NET0131  ;
  assign n24128 = ~decrypt_pad & ~\u2_uk_K_r1_reg[37]/NET0131  ;
  assign n24129 = ~n24127 & ~n24128 ;
  assign n24130 = \u2_R1_reg[28]/NET0131  & ~n24129 ;
  assign n24131 = ~\u2_R1_reg[28]/NET0131  & n24129 ;
  assign n24132 = ~n24130 & ~n24131 ;
  assign n24114 = decrypt_pad & ~\u2_uk_K_r1_reg[15]/NET0131  ;
  assign n24115 = ~decrypt_pad & ~\u2_uk_K_r1_reg[9]/NET0131  ;
  assign n24116 = ~n24114 & ~n24115 ;
  assign n24117 = \u2_R1_reg[29]/NET0131  & ~n24116 ;
  assign n24118 = ~\u2_R1_reg[29]/NET0131  & n24116 ;
  assign n24119 = ~n24117 & ~n24118 ;
  assign n24120 = decrypt_pad & ~\u2_uk_K_r1_reg[0]/NET0131  ;
  assign n24121 = ~decrypt_pad & ~\u2_uk_K_r1_reg[49]/NET0131  ;
  assign n24122 = ~n24120 & ~n24121 ;
  assign n24123 = \u2_R1_reg[1]/NET0131  & ~n24122 ;
  assign n24124 = ~\u2_R1_reg[1]/NET0131  & n24122 ;
  assign n24125 = ~n24123 & ~n24124 ;
  assign n24160 = ~n24119 & n24125 ;
  assign n24161 = ~n24132 & n24160 ;
  assign n24133 = decrypt_pad & ~\u2_uk_K_r1_reg[16]/NET0131  ;
  assign n24134 = ~decrypt_pad & ~\u2_uk_K_r1_reg[38]/NET0131  ;
  assign n24135 = ~n24133 & ~n24134 ;
  assign n24136 = \u2_R1_reg[30]/NET0131  & ~n24135 ;
  assign n24137 = ~\u2_R1_reg[30]/NET0131  & n24135 ;
  assign n24138 = ~n24136 & ~n24137 ;
  assign n24181 = ~n24119 & ~n24125 ;
  assign n24182 = n24138 & n24181 ;
  assign n24183 = n24132 & n24182 ;
  assign n24184 = ~n24161 & ~n24183 ;
  assign n24185 = n24157 & ~n24184 ;
  assign n24126 = n24119 & n24125 ;
  assign n24167 = n24132 & ~n24138 ;
  assign n24139 = ~n24132 & n24138 ;
  assign n24175 = ~n24125 & n24139 ;
  assign n24176 = ~n24167 & ~n24175 ;
  assign n24177 = ~n24126 & n24176 ;
  assign n24178 = ~n24157 & ~n24177 ;
  assign n24148 = n24119 & n24132 ;
  assign n24149 = ~n24138 & n24148 ;
  assign n24150 = ~n24125 & n24149 ;
  assign n24179 = n24138 & n24148 ;
  assign n24180 = n24125 & n24179 ;
  assign n24186 = ~n24150 & ~n24180 ;
  assign n24187 = ~n24178 & n24186 ;
  assign n24188 = ~n24185 & n24187 ;
  assign n24189 = ~n24113 & ~n24188 ;
  assign n24163 = n24119 & ~n24138 ;
  assign n24164 = ~n24125 & n24132 ;
  assign n24165 = ~n24163 & ~n24164 ;
  assign n24166 = ~n24113 & ~n24165 ;
  assign n24168 = n24119 & ~n24125 ;
  assign n24169 = ~n24167 & ~n24168 ;
  assign n24170 = ~n24150 & ~n24169 ;
  assign n24171 = ~n24166 & n24170 ;
  assign n24144 = ~n24132 & ~n24138 ;
  assign n24145 = ~n24119 & n24144 ;
  assign n24159 = ~n24125 & n24145 ;
  assign n24162 = n24138 & n24161 ;
  assign n24172 = ~n24159 & ~n24162 ;
  assign n24173 = ~n24171 & n24172 ;
  assign n24174 = n24157 & ~n24173 ;
  assign n24140 = n24126 & n24139 ;
  assign n24141 = n24113 & n24140 ;
  assign n24142 = ~n24119 & n24132 ;
  assign n24143 = n24138 & n24142 ;
  assign n24146 = ~n24143 & ~n24145 ;
  assign n24147 = n24113 & ~n24146 ;
  assign n24151 = ~n24147 & ~n24150 ;
  assign n24158 = ~n24151 & ~n24157 ;
  assign n24190 = ~n24141 & ~n24158 ;
  assign n24191 = ~n24174 & n24190 ;
  assign n24192 = ~n24189 & n24191 ;
  assign n24193 = \u2_L1_reg[5]/NET0131  & ~n24192 ;
  assign n24194 = ~\u2_L1_reg[5]/NET0131  & n24192 ;
  assign n24195 = ~n24193 & ~n24194 ;
  assign n24198 = n23833 & n23839 ;
  assign n24206 = ~n23899 & ~n24198 ;
  assign n24196 = n23846 & ~n23852 ;
  assign n24204 = ~n23853 & ~n24196 ;
  assign n24205 = n23839 & n23846 ;
  assign n24207 = n24204 & ~n24205 ;
  assign n24208 = n24206 & n24207 ;
  assign n24201 = ~n23860 & ~n23887 ;
  assign n24202 = ~n23859 & n24201 ;
  assign n24203 = ~n23878 & ~n24202 ;
  assign n24199 = ~n23880 & ~n24198 ;
  assign n24200 = n23853 & ~n24199 ;
  assign n24197 = n23899 & n24196 ;
  assign n24209 = ~n23868 & ~n24197 ;
  assign n24210 = ~n24200 & n24209 ;
  assign n24211 = ~n24203 & n24210 ;
  assign n24212 = ~n24208 & n24211 ;
  assign n24216 = ~n23904 & ~n24205 ;
  assign n24217 = n23878 & ~n24216 ;
  assign n24218 = n23868 & ~n23900 ;
  assign n24219 = ~n23857 & n24218 ;
  assign n24213 = n23854 & ~n23878 ;
  assign n24214 = ~n23898 & ~n24198 ;
  assign n24215 = ~n24201 & n24214 ;
  assign n24220 = ~n24213 & ~n24215 ;
  assign n24221 = n24219 & n24220 ;
  assign n24222 = ~n24217 & n24221 ;
  assign n24223 = ~n24212 & ~n24222 ;
  assign n24224 = \u2_L1_reg[12]/NET0131  & n24223 ;
  assign n24225 = ~\u2_L1_reg[12]/NET0131  & ~n24223 ;
  assign n24226 = ~n24224 & ~n24225 ;
  assign n24245 = ~n23969 & ~n23988 ;
  assign n24246 = ~n23932 & ~n24245 ;
  assign n24247 = ~n23966 & ~n24246 ;
  assign n24248 = ~n23953 & ~n24247 ;
  assign n24242 = n23939 & n23995 ;
  assign n24243 = ~n23956 & ~n24242 ;
  assign n24244 = n23953 & ~n24243 ;
  assign n24249 = ~n23947 & ~n23979 ;
  assign n24250 = ~n24244 & n24249 ;
  assign n24251 = ~n24248 & n24250 ;
  assign n24252 = ~n23920 & ~n24251 ;
  assign n24227 = ~n23926 & n23963 ;
  assign n24228 = ~n23989 & ~n24227 ;
  assign n24229 = n23997 & ~n24228 ;
  assign n24232 = ~n23946 & ~n23971 ;
  assign n24233 = n23969 & n23971 ;
  assign n24234 = ~n24232 & ~n24233 ;
  assign n24235 = n23953 & ~n24234 ;
  assign n24236 = ~n23953 & ~n23987 ;
  assign n24237 = ~n24232 & n24236 ;
  assign n24230 = n23933 & n23939 ;
  assign n24231 = n23980 & n23995 ;
  assign n24238 = ~n24230 & ~n24231 ;
  assign n24239 = ~n24237 & n24238 ;
  assign n24240 = ~n24235 & n24239 ;
  assign n24241 = n23920 & ~n24240 ;
  assign n24253 = ~n24229 & ~n24241 ;
  assign n24254 = ~n24252 & n24253 ;
  assign n24255 = ~\u2_L1_reg[17]/NET0131  & ~n24254 ;
  assign n24256 = \u2_L1_reg[17]/NET0131  & n24254 ;
  assign n24257 = ~n24255 & ~n24256 ;
  assign n24258 = decrypt_pad & ~\u2_uk_K_r1_reg[17]/NET0131  ;
  assign n24259 = ~decrypt_pad & ~\u2_uk_K_r1_reg[41]/NET0131  ;
  assign n24260 = ~n24258 & ~n24259 ;
  assign n24261 = \u2_R1_reg[17]/NET0131  & ~n24260 ;
  assign n24262 = ~\u2_R1_reg[17]/NET0131  & n24260 ;
  assign n24263 = ~n24261 & ~n24262 ;
  assign n24264 = decrypt_pad & ~\u2_uk_K_r1_reg[33]/NET0131  ;
  assign n24265 = ~decrypt_pad & ~\u2_uk_K_r1_reg[25]/NET0131  ;
  assign n24266 = ~n24264 & ~n24265 ;
  assign n24267 = \u2_R1_reg[12]/NET0131  & ~n24266 ;
  assign n24268 = ~\u2_R1_reg[12]/NET0131  & n24266 ;
  assign n24269 = ~n24267 & ~n24268 ;
  assign n24270 = ~n24263 & ~n24269 ;
  assign n24271 = decrypt_pad & ~\u2_uk_K_r1_reg[27]/NET0131  ;
  assign n24272 = ~decrypt_pad & ~\u2_uk_K_r1_reg[19]/NET0131  ;
  assign n24273 = ~n24271 & ~n24272 ;
  assign n24274 = \u2_R1_reg[13]/NET0131  & ~n24273 ;
  assign n24275 = ~\u2_R1_reg[13]/NET0131  & n24273 ;
  assign n24276 = ~n24274 & ~n24275 ;
  assign n24303 = n24270 & ~n24276 ;
  assign n24295 = n24263 & n24269 ;
  assign n24296 = n24276 & n24295 ;
  assign n24297 = decrypt_pad & ~\u2_uk_K_r1_reg[4]/NET0131  ;
  assign n24298 = ~decrypt_pad & ~\u2_uk_K_r1_reg[53]/NET0131  ;
  assign n24299 = ~n24297 & ~n24298 ;
  assign n24300 = \u2_R1_reg[15]/NET0131  & ~n24299 ;
  assign n24301 = ~\u2_R1_reg[15]/NET0131  & n24299 ;
  assign n24302 = ~n24300 & ~n24301 ;
  assign n24304 = ~n24296 & n24302 ;
  assign n24305 = ~n24303 & n24304 ;
  assign n24278 = decrypt_pad & ~\u2_uk_K_r1_reg[53]/NET0131  ;
  assign n24279 = ~decrypt_pad & ~\u2_uk_K_r1_reg[20]/NET0131  ;
  assign n24280 = ~n24278 & ~n24279 ;
  assign n24281 = \u2_R1_reg[14]/NET0131  & ~n24280 ;
  assign n24282 = ~\u2_R1_reg[14]/NET0131  & n24280 ;
  assign n24283 = ~n24281 & ~n24282 ;
  assign n24306 = ~n24263 & n24269 ;
  assign n24307 = n24283 & n24306 ;
  assign n24308 = n24263 & ~n24276 ;
  assign n24309 = ~n24302 & ~n24308 ;
  assign n24310 = ~n24307 & n24309 ;
  assign n24311 = ~n24305 & ~n24310 ;
  assign n24277 = n24270 & n24276 ;
  assign n24284 = n24277 & n24283 ;
  assign n24285 = ~n24263 & ~n24283 ;
  assign n24286 = ~n24269 & n24285 ;
  assign n24287 = ~n24276 & n24286 ;
  assign n24288 = ~n24284 & ~n24287 ;
  assign n24315 = ~n24283 & n24308 ;
  assign n24316 = n24269 & n24315 ;
  assign n24289 = decrypt_pad & ~\u2_uk_K_r1_reg[12]/NET0131  ;
  assign n24290 = ~decrypt_pad & ~\u2_uk_K_r1_reg[4]/NET0131  ;
  assign n24291 = ~n24289 & ~n24290 ;
  assign n24292 = \u2_R1_reg[16]/NET0131  & ~n24291 ;
  assign n24293 = ~\u2_R1_reg[16]/NET0131  & n24291 ;
  assign n24294 = ~n24292 & ~n24293 ;
  assign n24312 = n24276 & n24302 ;
  assign n24313 = n24283 & n24312 ;
  assign n24314 = ~n24269 & n24313 ;
  assign n24317 = ~n24294 & ~n24314 ;
  assign n24318 = ~n24316 & n24317 ;
  assign n24319 = n24288 & n24318 ;
  assign n24320 = ~n24311 & n24319 ;
  assign n24331 = n24283 & n24296 ;
  assign n24324 = ~n24276 & ~n24302 ;
  assign n24325 = n24270 & n24324 ;
  assign n24326 = n24283 & n24325 ;
  assign n24321 = ~n24276 & n24302 ;
  assign n24322 = n24263 & ~n24269 ;
  assign n24323 = n24321 & n24322 ;
  assign n24338 = n24294 & ~n24323 ;
  assign n24339 = ~n24326 & n24338 ;
  assign n24340 = ~n24331 & n24339 ;
  assign n24327 = n24306 & n24312 ;
  assign n24328 = ~n24283 & n24322 ;
  assign n24329 = n24276 & n24328 ;
  assign n24330 = ~n24327 & ~n24329 ;
  assign n24332 = n24276 & ~n24283 ;
  assign n24333 = ~n24269 & n24332 ;
  assign n24334 = n24269 & ~n24283 ;
  assign n24335 = ~n24276 & n24334 ;
  assign n24336 = ~n24333 & ~n24335 ;
  assign n24337 = ~n24302 & ~n24336 ;
  assign n24341 = n24330 & ~n24337 ;
  assign n24342 = n24340 & n24341 ;
  assign n24343 = ~n24320 & ~n24342 ;
  assign n24346 = ~n24302 & n24329 ;
  assign n24344 = ~n24286 & ~n24307 ;
  assign n24345 = n24321 & ~n24344 ;
  assign n24347 = ~n24283 & n24327 ;
  assign n24348 = ~n24345 & ~n24347 ;
  assign n24349 = ~n24346 & n24348 ;
  assign n24350 = ~n24343 & n24349 ;
  assign n24351 = ~\u2_L1_reg[20]/NET0131  & ~n24350 ;
  assign n24352 = \u2_L1_reg[20]/NET0131  & n24350 ;
  assign n24353 = ~n24351 & ~n24352 ;
  assign n24391 = decrypt_pad & ~\u2_uk_K_r1_reg[11]/NET0131  ;
  assign n24392 = ~decrypt_pad & ~\u2_uk_K_r1_reg[3]/NET0131  ;
  assign n24393 = ~n24391 & ~n24392 ;
  assign n24394 = \u2_R1_reg[8]/NET0131  & ~n24393 ;
  assign n24395 = ~\u2_R1_reg[8]/NET0131  & n24393 ;
  assign n24396 = ~n24394 & ~n24395 ;
  assign n24384 = decrypt_pad & ~\u2_uk_K_r1_reg[20]/NET0131  ;
  assign n24385 = ~decrypt_pad & ~\u2_uk_K_r1_reg[12]/NET0131  ;
  assign n24386 = ~n24384 & ~n24385 ;
  assign n24387 = \u2_R1_reg[7]/NET0131  & ~n24386 ;
  assign n24388 = ~\u2_R1_reg[7]/NET0131  & n24386 ;
  assign n24389 = ~n24387 & ~n24388 ;
  assign n24354 = decrypt_pad & ~\u2_uk_K_r1_reg[3]/NET0131  ;
  assign n24355 = ~decrypt_pad & ~\u2_uk_K_r1_reg[27]/NET0131  ;
  assign n24356 = ~n24354 & ~n24355 ;
  assign n24357 = \u2_R1_reg[5]/NET0131  & ~n24356 ;
  assign n24358 = ~\u2_R1_reg[5]/NET0131  & n24356 ;
  assign n24359 = ~n24357 & ~n24358 ;
  assign n24360 = decrypt_pad & ~\u2_uk_K_r1_reg[26]/NET0131  ;
  assign n24361 = ~decrypt_pad & ~\u2_uk_K_r1_reg[18]/NET0131  ;
  assign n24362 = ~n24360 & ~n24361 ;
  assign n24363 = \u2_R1_reg[6]/NET0131  & ~n24362 ;
  assign n24364 = ~\u2_R1_reg[6]/NET0131  & n24362 ;
  assign n24365 = ~n24363 & ~n24364 ;
  assign n24381 = n24359 & n24365 ;
  assign n24367 = decrypt_pad & ~\u2_uk_K_r1_reg[24]/NET0131  ;
  assign n24368 = ~decrypt_pad & ~\u2_uk_K_r1_reg[48]/NET0131  ;
  assign n24369 = ~n24367 & ~n24368 ;
  assign n24370 = \u2_R1_reg[4]/NET0131  & ~n24369 ;
  assign n24371 = ~\u2_R1_reg[4]/NET0131  & n24369 ;
  assign n24372 = ~n24370 & ~n24371 ;
  assign n24374 = decrypt_pad & ~\u2_uk_K_r1_reg[48]/NET0131  ;
  assign n24375 = ~decrypt_pad & ~\u2_uk_K_r1_reg[40]/NET0131  ;
  assign n24376 = ~n24374 & ~n24375 ;
  assign n24377 = \u2_R1_reg[9]/NET0131  & ~n24376 ;
  assign n24378 = ~\u2_R1_reg[9]/NET0131  & n24376 ;
  assign n24379 = ~n24377 & ~n24378 ;
  assign n24397 = ~n24372 & ~n24379 ;
  assign n24423 = n24381 & n24397 ;
  assign n24411 = n24372 & n24379 ;
  assign n24421 = n24359 & n24411 ;
  assign n24380 = n24372 & ~n24379 ;
  assign n24422 = ~n24359 & n24380 ;
  assign n24424 = ~n24421 & ~n24422 ;
  assign n24425 = ~n24423 & n24424 ;
  assign n24426 = n24389 & ~n24425 ;
  assign n24398 = ~n24365 & n24397 ;
  assign n24399 = ~n24372 & n24379 ;
  assign n24400 = n24359 & n24399 ;
  assign n24401 = ~n24398 & ~n24400 ;
  assign n24420 = ~n24389 & ~n24401 ;
  assign n24404 = ~n24365 & n24372 ;
  assign n24417 = ~n24359 & n24411 ;
  assign n24418 = ~n24389 & ~n24417 ;
  assign n24419 = n24404 & ~n24418 ;
  assign n24406 = ~n24359 & n24399 ;
  assign n24427 = n24365 & n24406 ;
  assign n24428 = ~n24419 & ~n24427 ;
  assign n24429 = ~n24420 & n24428 ;
  assign n24430 = ~n24426 & n24429 ;
  assign n24431 = n24396 & ~n24430 ;
  assign n24366 = ~n24359 & n24365 ;
  assign n24373 = n24366 & ~n24372 ;
  assign n24382 = n24380 & n24381 ;
  assign n24383 = ~n24373 & ~n24382 ;
  assign n24390 = ~n24383 & ~n24389 ;
  assign n24402 = n24389 & n24401 ;
  assign n24405 = ~n24379 & n24404 ;
  assign n24403 = n24359 & n24372 ;
  assign n24407 = ~n24389 & ~n24403 ;
  assign n24408 = ~n24405 & n24407 ;
  assign n24409 = ~n24406 & n24408 ;
  assign n24410 = ~n24402 & ~n24409 ;
  assign n24412 = ~n24397 & ~n24411 ;
  assign n24413 = n24366 & ~n24412 ;
  assign n24414 = ~n24382 & ~n24413 ;
  assign n24415 = ~n24410 & n24414 ;
  assign n24416 = ~n24396 & ~n24415 ;
  assign n24432 = ~n24390 & ~n24416 ;
  assign n24433 = ~n24431 & n24432 ;
  assign n24434 = ~\u2_L1_reg[28]/NET0131  & ~n24433 ;
  assign n24435 = \u2_L1_reg[28]/NET0131  & n24433 ;
  assign n24436 = ~n24434 & ~n24435 ;
  assign n24442 = ~n24038 & ~n24048 ;
  assign n24443 = ~n24030 & ~n24044 ;
  assign n24444 = n24037 & n24075 ;
  assign n24445 = ~n24443 & ~n24444 ;
  assign n24446 = ~n24076 & ~n24445 ;
  assign n24447 = n24442 & ~n24446 ;
  assign n24448 = n24018 & ~n24447 ;
  assign n24437 = n24044 & n24081 ;
  assign n24438 = ~n24044 & ~n24047 ;
  assign n24439 = ~n24082 & n24438 ;
  assign n24440 = ~n24437 & ~n24439 ;
  assign n24441 = ~n24018 & ~n24440 ;
  assign n24449 = n24044 & n24091 ;
  assign n24450 = ~n24441 & ~n24449 ;
  assign n24451 = ~n24448 & n24450 ;
  assign n24452 = ~n24069 & ~n24451 ;
  assign n24453 = n24037 & n24071 ;
  assign n24454 = ~n24055 & ~n24453 ;
  assign n24455 = ~n24437 & n24454 ;
  assign n24456 = n24018 & ~n24455 ;
  assign n24459 = ~n24031 & n24044 ;
  assign n24460 = ~n24075 & n24459 ;
  assign n24457 = ~n24037 & ~n24443 ;
  assign n24458 = n24018 & ~n24457 ;
  assign n24461 = ~n24439 & ~n24458 ;
  assign n24462 = ~n24460 & n24461 ;
  assign n24463 = ~n24456 & ~n24462 ;
  assign n24464 = n24069 & ~n24463 ;
  assign n24465 = n24018 & ~n24044 ;
  assign n24466 = n24054 & n24465 ;
  assign n24467 = ~n24049 & ~n24466 ;
  assign n24468 = ~n24464 & n24467 ;
  assign n24469 = ~n24452 & n24468 ;
  assign n24470 = \u2_L1_reg[29]/NET0131  & ~n24469 ;
  assign n24471 = ~\u2_L1_reg[29]/NET0131  & n24469 ;
  assign n24472 = ~n24470 & ~n24471 ;
  assign n24475 = ~n24380 & ~n24403 ;
  assign n24476 = n24365 & ~n24475 ;
  assign n24477 = ~n24406 & ~n24476 ;
  assign n24478 = ~n24389 & ~n24477 ;
  assign n24482 = ~n24359 & ~n24389 ;
  assign n24483 = ~n24365 & n24379 ;
  assign n24484 = n24482 & n24483 ;
  assign n24485 = n24365 & n24400 ;
  assign n24486 = ~n24484 & ~n24485 ;
  assign n24473 = n24365 & n24417 ;
  assign n24474 = n24389 & n24473 ;
  assign n24479 = n24359 & ~n24379 ;
  assign n24480 = ~n24406 & ~n24479 ;
  assign n24481 = ~n24365 & ~n24480 ;
  assign n24487 = ~n24474 & ~n24481 ;
  assign n24488 = n24486 & n24487 ;
  assign n24489 = ~n24478 & n24488 ;
  assign n24490 = ~n24396 & ~n24489 ;
  assign n24496 = ~n24397 & ~n24405 ;
  assign n24497 = ~n24359 & ~n24496 ;
  assign n24494 = n24365 & ~n24403 ;
  assign n24495 = ~n24412 & n24494 ;
  assign n24498 = ~n24365 & n24421 ;
  assign n24499 = ~n24495 & ~n24498 ;
  assign n24500 = ~n24497 & n24499 ;
  assign n24501 = n24396 & ~n24500 ;
  assign n24491 = ~n24359 & ~n24365 ;
  assign n24492 = ~n24381 & ~n24491 ;
  assign n24493 = n24399 & ~n24492 ;
  assign n24502 = ~n24389 & ~n24493 ;
  assign n24503 = ~n24501 & n24502 ;
  assign n24505 = ~n24359 & ~n24380 ;
  assign n24506 = n24396 & ~n24494 ;
  assign n24507 = ~n24505 & n24506 ;
  assign n24508 = n24366 & ~n24379 ;
  assign n24509 = ~n24372 & n24508 ;
  assign n24504 = n24359 & n24404 ;
  assign n24510 = n24389 & ~n24504 ;
  assign n24511 = ~n24509 & n24510 ;
  assign n24512 = ~n24507 & n24511 ;
  assign n24513 = ~n24503 & ~n24512 ;
  assign n24514 = ~n24490 & ~n24513 ;
  assign n24515 = \u2_L1_reg[2]/NET0131  & n24514 ;
  assign n24516 = ~\u2_L1_reg[2]/NET0131  & ~n24514 ;
  assign n24517 = ~n24515 & ~n24516 ;
  assign n24532 = ~n24072 & ~n24081 ;
  assign n24533 = ~n24096 & n24532 ;
  assign n24534 = n24018 & ~n24533 ;
  assign n24535 = n24031 & n24080 ;
  assign n24536 = ~n24049 & ~n24535 ;
  assign n24537 = ~n24534 & n24536 ;
  assign n24538 = ~n24069 & ~n24537 ;
  assign n24519 = ~n24444 & ~n24449 ;
  assign n24520 = ~n24069 & ~n24519 ;
  assign n24518 = ~n24030 & n24071 ;
  assign n24521 = ~n24030 & n24076 ;
  assign n24522 = ~n24071 & ~n24521 ;
  assign n24523 = n24069 & ~n24522 ;
  assign n24524 = ~n24518 & ~n24523 ;
  assign n24525 = ~n24520 & n24524 ;
  assign n24526 = ~n24018 & ~n24525 ;
  assign n24527 = n24024 & n24465 ;
  assign n24528 = ~n24045 & ~n24527 ;
  assign n24529 = n24030 & ~n24528 ;
  assign n24530 = ~n24077 & ~n24529 ;
  assign n24531 = n24069 & ~n24530 ;
  assign n24540 = ~n24055 & ~n24083 ;
  assign n24541 = n24018 & ~n24081 ;
  assign n24542 = n24540 & n24541 ;
  assign n24539 = ~n24018 & n24442 ;
  assign n24543 = n24044 & ~n24539 ;
  assign n24544 = ~n24542 & n24543 ;
  assign n24545 = ~n24531 & ~n24544 ;
  assign n24546 = ~n24526 & n24545 ;
  assign n24547 = ~n24538 & n24546 ;
  assign n24548 = ~\u2_L1_reg[4]/NET0131  & ~n24547 ;
  assign n24549 = \u2_L1_reg[4]/NET0131  & n24547 ;
  assign n24550 = ~n24548 & ~n24549 ;
  assign n24569 = n24306 & ~n24332 ;
  assign n24570 = ~n24329 & ~n24569 ;
  assign n24571 = ~n24302 & ~n24570 ;
  assign n24552 = ~n24276 & n24283 ;
  assign n24565 = n24322 & n24552 ;
  assign n24566 = ~n24331 & ~n24565 ;
  assign n24567 = ~n24277 & ~n24316 ;
  assign n24568 = n24302 & ~n24567 ;
  assign n24572 = n24566 & ~n24568 ;
  assign n24573 = ~n24571 & n24572 ;
  assign n24574 = n24294 & ~n24573 ;
  assign n24551 = ~n24263 & ~n24276 ;
  assign n24553 = ~n24551 & ~n24552 ;
  assign n24554 = n24269 & ~n24553 ;
  assign n24555 = ~n24328 & ~n24554 ;
  assign n24556 = n24302 & ~n24555 ;
  assign n24559 = n24269 & n24332 ;
  assign n24557 = ~n24283 & ~n24302 ;
  assign n24558 = n24295 & n24557 ;
  assign n24560 = ~n24325 & ~n24558 ;
  assign n24561 = ~n24559 & n24560 ;
  assign n24562 = n24288 & n24561 ;
  assign n24563 = ~n24556 & n24562 ;
  assign n24564 = ~n24294 & ~n24563 ;
  assign n24575 = ~n24287 & n24566 ;
  assign n24576 = ~n24302 & ~n24575 ;
  assign n24577 = ~n24314 & ~n24347 ;
  assign n24578 = ~n24576 & n24577 ;
  assign n24579 = ~n24564 & n24578 ;
  assign n24580 = ~n24574 & n24579 ;
  assign n24581 = ~\u2_L1_reg[10]/NET0131  & ~n24580 ;
  assign n24582 = \u2_L1_reg[10]/NET0131  & n24580 ;
  assign n24583 = ~n24581 & ~n24582 ;
  assign n24584 = ~n24382 & ~n24498 ;
  assign n24585 = ~n24372 & n24479 ;
  assign n24586 = n24380 & n24491 ;
  assign n24587 = ~n24585 & ~n24586 ;
  assign n24588 = ~n24427 & n24587 ;
  assign n24589 = ~n24396 & ~n24588 ;
  assign n24590 = n24584 & ~n24589 ;
  assign n24591 = ~n24389 & ~n24590 ;
  assign n24598 = ~n24359 & n24412 ;
  assign n24597 = n24359 & ~n24405 ;
  assign n24599 = n24389 & ~n24597 ;
  assign n24600 = ~n24598 & n24599 ;
  assign n24594 = n24365 & n24389 ;
  assign n24595 = n24372 & ~n24479 ;
  assign n24596 = n24594 & n24595 ;
  assign n24592 = ~n24365 & n24399 ;
  assign n24593 = ~n24482 & n24592 ;
  assign n24601 = ~n24396 & ~n24593 ;
  assign n24602 = ~n24596 & n24601 ;
  assign n24603 = ~n24600 & n24602 ;
  assign n24605 = n24418 & ~n24508 ;
  assign n24607 = ~n24379 & n24491 ;
  assign n24606 = n24365 & n24399 ;
  assign n24608 = n24389 & ~n24606 ;
  assign n24609 = ~n24607 & n24608 ;
  assign n24610 = ~n24605 & ~n24609 ;
  assign n24604 = n24359 & n24398 ;
  assign n24611 = n24396 & ~n24604 ;
  assign n24612 = n24486 & n24611 ;
  assign n24613 = n24584 & n24612 ;
  assign n24614 = ~n24610 & n24613 ;
  assign n24615 = ~n24603 & ~n24614 ;
  assign n24616 = ~n24591 & ~n24615 ;
  assign n24617 = ~\u2_L1_reg[13]/NET0131  & n24616 ;
  assign n24618 = \u2_L1_reg[13]/NET0131  & ~n24616 ;
  assign n24619 = ~n24617 & ~n24618 ;
  assign n24621 = n24119 & ~n24176 ;
  assign n24622 = ~n24132 & n24181 ;
  assign n24623 = n24157 & n24622 ;
  assign n24620 = n24125 & n24143 ;
  assign n24624 = n24138 & ~n24157 ;
  assign n24625 = n24160 & n24624 ;
  assign n24626 = n24113 & ~n24625 ;
  assign n24627 = ~n24620 & n24626 ;
  assign n24628 = ~n24623 & n24627 ;
  assign n24629 = ~n24621 & n24628 ;
  assign n24631 = ~n24138 & n24168 ;
  assign n24632 = ~n24148 & ~n24631 ;
  assign n24633 = ~n24161 & n24632 ;
  assign n24634 = n24157 & ~n24633 ;
  assign n24630 = n24167 & n24181 ;
  assign n24635 = ~n24113 & ~n24630 ;
  assign n24636 = ~n24634 & n24635 ;
  assign n24637 = ~n24629 & ~n24636 ;
  assign n24639 = n24144 & ~n24160 ;
  assign n24640 = ~n24168 & n24639 ;
  assign n24641 = n24113 & ~n24138 ;
  assign n24642 = n24142 & ~n24641 ;
  assign n24638 = n24139 & n24168 ;
  assign n24643 = ~n24157 & ~n24638 ;
  assign n24644 = ~n24642 & n24643 ;
  assign n24645 = ~n24640 & n24644 ;
  assign n24646 = ~n24138 & n24160 ;
  assign n24647 = ~n24132 & n24646 ;
  assign n24648 = ~n24140 & n24157 ;
  assign n24649 = ~n24647 & n24648 ;
  assign n24650 = ~n24645 & ~n24649 ;
  assign n24651 = ~n24637 & ~n24650 ;
  assign n24652 = ~\u2_L1_reg[15]/NET0131  & ~n24651 ;
  assign n24653 = \u2_L1_reg[15]/NET0131  & n24651 ;
  assign n24654 = ~n24652 & ~n24653 ;
  assign n24712 = decrypt_pad & ~\u2_uk_K_r1_reg[50]/NET0131  ;
  assign n24713 = ~decrypt_pad & ~\u2_uk_K_r1_reg[44]/P0001  ;
  assign n24714 = ~n24712 & ~n24713 ;
  assign n24715 = \u2_R1_reg[20]/NET0131  & ~n24714 ;
  assign n24716 = ~\u2_R1_reg[20]/NET0131  & n24714 ;
  assign n24717 = ~n24715 & ~n24716 ;
  assign n24687 = decrypt_pad & ~\u2_uk_K_r1_reg[35]/NET0131  ;
  assign n24688 = ~decrypt_pad & ~\u2_uk_K_r1_reg[29]/NET0131  ;
  assign n24689 = ~n24687 & ~n24688 ;
  assign n24690 = \u2_R1_reg[19]/NET0131  & ~n24689 ;
  assign n24691 = ~\u2_R1_reg[19]/NET0131  & n24689 ;
  assign n24692 = ~n24690 & ~n24691 ;
  assign n24675 = decrypt_pad & ~\u2_uk_K_r1_reg[52]/NET0131  ;
  assign n24676 = ~decrypt_pad & ~\u2_uk_K_r1_reg[42]/NET0131  ;
  assign n24677 = ~n24675 & ~n24676 ;
  assign n24678 = \u2_R1_reg[18]/NET0131  & ~n24677 ;
  assign n24679 = ~\u2_R1_reg[18]/NET0131  & n24677 ;
  assign n24680 = ~n24678 & ~n24679 ;
  assign n24668 = decrypt_pad & ~\u2_uk_K_r1_reg[30]/NET0131  ;
  assign n24669 = ~decrypt_pad & ~\u2_uk_K_r1_reg[52]/NET0131  ;
  assign n24670 = ~n24668 & ~n24669 ;
  assign n24671 = \u2_R1_reg[17]/NET0131  & ~n24670 ;
  assign n24672 = ~\u2_R1_reg[17]/NET0131  & n24670 ;
  assign n24673 = ~n24671 & ~n24672 ;
  assign n24655 = decrypt_pad & ~\u2_uk_K_r1_reg[51]/NET0131  ;
  assign n24656 = ~decrypt_pad & ~\u2_uk_K_r1_reg[14]/NET0131  ;
  assign n24657 = ~n24655 & ~n24656 ;
  assign n24658 = \u2_R1_reg[21]/NET0131  & ~n24657 ;
  assign n24659 = ~\u2_R1_reg[21]/NET0131  & n24657 ;
  assign n24660 = ~n24658 & ~n24659 ;
  assign n24661 = decrypt_pad & ~\u2_uk_K_r1_reg[8]/NET0131  ;
  assign n24662 = ~decrypt_pad & ~\u2_uk_K_r1_reg[2]/NET0131  ;
  assign n24663 = ~n24661 & ~n24662 ;
  assign n24664 = \u2_R1_reg[16]/NET0131  & ~n24663 ;
  assign n24665 = ~\u2_R1_reg[16]/NET0131  & n24663 ;
  assign n24666 = ~n24664 & ~n24665 ;
  assign n24694 = n24660 & n24666 ;
  assign n24726 = n24673 & n24694 ;
  assign n24727 = ~n24680 & n24726 ;
  assign n24704 = ~n24666 & ~n24673 ;
  assign n24730 = n24660 & n24704 ;
  assign n24719 = n24673 & n24680 ;
  assign n24720 = ~n24660 & n24719 ;
  assign n24667 = ~n24660 & n24666 ;
  assign n24728 = ~n24673 & ~n24680 ;
  assign n24729 = n24667 & n24728 ;
  assign n24731 = ~n24720 & ~n24729 ;
  assign n24732 = ~n24730 & n24731 ;
  assign n24733 = ~n24727 & n24732 ;
  assign n24734 = ~n24692 & ~n24733 ;
  assign n24681 = n24673 & ~n24680 ;
  assign n24682 = ~n24666 & n24681 ;
  assign n24683 = n24666 & n24680 ;
  assign n24684 = n24660 & ~n24683 ;
  assign n24685 = ~n24682 & n24684 ;
  assign n24721 = ~n24667 & n24692 ;
  assign n24722 = ~n24720 & n24721 ;
  assign n24723 = ~n24685 & n24722 ;
  assign n24699 = ~n24673 & n24680 ;
  assign n24724 = n24694 & n24699 ;
  assign n24725 = ~n24660 & n24682 ;
  assign n24735 = ~n24724 & ~n24725 ;
  assign n24736 = ~n24723 & n24735 ;
  assign n24737 = ~n24734 & n24736 ;
  assign n24738 = ~n24717 & ~n24737 ;
  assign n24674 = n24667 & n24673 ;
  assign n24686 = ~n24674 & ~n24685 ;
  assign n24693 = ~n24686 & n24692 ;
  assign n24695 = n24673 & ~n24692 ;
  assign n24702 = n24660 & ~n24666 ;
  assign n24703 = n24695 & n24702 ;
  assign n24705 = ~n24660 & ~n24692 ;
  assign n24706 = n24704 & n24705 ;
  assign n24707 = ~n24703 & ~n24706 ;
  assign n24708 = ~n24680 & ~n24707 ;
  assign n24696 = n24680 & ~n24695 ;
  assign n24697 = ~n24681 & n24694 ;
  assign n24698 = ~n24696 & n24697 ;
  assign n24700 = ~n24681 & ~n24699 ;
  assign n24701 = n24667 & ~n24700 ;
  assign n24709 = ~n24698 & ~n24701 ;
  assign n24710 = ~n24708 & n24709 ;
  assign n24711 = ~n24693 & n24710 ;
  assign n24718 = ~n24711 & n24717 ;
  assign n24739 = ~n24660 & ~n24666 ;
  assign n24740 = n24699 & n24739 ;
  assign n24741 = n24674 & ~n24680 ;
  assign n24742 = ~n24740 & ~n24741 ;
  assign n24743 = n24692 & ~n24742 ;
  assign n24744 = n24660 & n24680 ;
  assign n24745 = n24704 & n24744 ;
  assign n24746 = n24719 & n24739 ;
  assign n24747 = ~n24745 & ~n24746 ;
  assign n24748 = ~n24692 & ~n24747 ;
  assign n24749 = ~n24743 & ~n24748 ;
  assign n24750 = ~n24718 & n24749 ;
  assign n24751 = ~n24738 & n24750 ;
  assign n24752 = ~\u2_L1_reg[14]/NET0131  & ~n24751 ;
  assign n24753 = \u2_L1_reg[14]/NET0131  & n24751 ;
  assign n24754 = ~n24752 & ~n24753 ;
  assign n24755 = ~n24018 & n24056 ;
  assign n24759 = n24069 & ~n24521 ;
  assign n24760 = ~n24755 & n24759 ;
  assign n24761 = ~n24073 & n24760 ;
  assign n24756 = ~n24086 & ~n24091 ;
  assign n24757 = n24018 & ~n24756 ;
  assign n24758 = n24044 & ~n24540 ;
  assign n24762 = ~n24757 & ~n24758 ;
  assign n24763 = n24761 & n24762 ;
  assign n24766 = n24024 & ~n24076 ;
  assign n24767 = ~n24444 & ~n24766 ;
  assign n24768 = n24018 & ~n24767 ;
  assign n24765 = ~n24018 & ~n24540 ;
  assign n24764 = n24037 & n24053 ;
  assign n24769 = ~n24069 & ~n24764 ;
  assign n24770 = ~n24765 & n24769 ;
  assign n24771 = ~n24768 & n24770 ;
  assign n24772 = ~n24763 & ~n24771 ;
  assign n24773 = ~n24057 & ~n24081 ;
  assign n24774 = n24080 & ~n24773 ;
  assign n24775 = ~n24074 & ~n24774 ;
  assign n24776 = ~n24772 & n24775 ;
  assign n24777 = ~\u2_L1_reg[19]/NET0131  & ~n24776 ;
  assign n24778 = \u2_L1_reg[19]/NET0131  & n24776 ;
  assign n24779 = ~n24777 & ~n24778 ;
  assign n24783 = ~n24125 & n24167 ;
  assign n24784 = ~n24157 & ~n24783 ;
  assign n24785 = ~n24620 & n24784 ;
  assign n24787 = n24157 & ~n24179 ;
  assign n24786 = n24126 & ~n24132 ;
  assign n24788 = ~n24646 & ~n24786 ;
  assign n24789 = n24787 & n24788 ;
  assign n24790 = ~n24785 & ~n24789 ;
  assign n24791 = ~n24125 & n24148 ;
  assign n24792 = ~n24622 & ~n24791 ;
  assign n24793 = n24138 & ~n24792 ;
  assign n24794 = n24113 & ~n24647 ;
  assign n24795 = ~n24793 & n24794 ;
  assign n24796 = ~n24790 & n24795 ;
  assign n24781 = n24125 & ~n24157 ;
  assign n24801 = ~n24126 & ~n24781 ;
  assign n24802 = n24167 & ~n24801 ;
  assign n24797 = ~n24119 & ~n24781 ;
  assign n24798 = n24139 & ~n24797 ;
  assign n24807 = ~n24183 & ~n24798 ;
  assign n24808 = ~n24802 & n24807 ;
  assign n24799 = ~n24143 & ~n24791 ;
  assign n24800 = n24157 & ~n24799 ;
  assign n24803 = ~n24132 & ~n24157 ;
  assign n24804 = n24168 & n24803 ;
  assign n24805 = ~n24113 & ~n24804 ;
  assign n24806 = ~n24159 & n24805 ;
  assign n24809 = ~n24800 & n24806 ;
  assign n24810 = n24808 & n24809 ;
  assign n24811 = ~n24796 & ~n24810 ;
  assign n24780 = n24145 & n24157 ;
  assign n24782 = n24149 & n24781 ;
  assign n24812 = ~n24780 & ~n24782 ;
  assign n24813 = ~n24811 & n24812 ;
  assign n24814 = ~\u2_L1_reg[21]/NET0131  & ~n24813 ;
  assign n24815 = \u2_L1_reg[21]/NET0131  & n24813 ;
  assign n24816 = ~n24814 & ~n24815 ;
  assign n24832 = ~n24263 & ~n24333 ;
  assign n24831 = n24269 & n24283 ;
  assign n24833 = n24276 & ~n24302 ;
  assign n24834 = ~n24831 & n24833 ;
  assign n24835 = ~n24832 & n24834 ;
  assign n24836 = ~n24263 & ~n24334 ;
  assign n24837 = n24321 & ~n24836 ;
  assign n24817 = n24276 & n24307 ;
  assign n24838 = ~n24269 & n24552 ;
  assign n24839 = ~n24817 & ~n24838 ;
  assign n24840 = ~n24837 & n24839 ;
  assign n24841 = ~n24835 & n24840 ;
  assign n24842 = n24294 & ~n24841 ;
  assign n24819 = ~n24285 & ~n24308 ;
  assign n24820 = n24269 & ~n24819 ;
  assign n24821 = ~n24302 & ~n24820 ;
  assign n24822 = n24306 & n24552 ;
  assign n24823 = ~n24286 & n24302 ;
  assign n24824 = ~n24822 & n24823 ;
  assign n24825 = ~n24821 & ~n24824 ;
  assign n24826 = ~n24270 & ~n24295 ;
  assign n24827 = n24332 & n24826 ;
  assign n24828 = ~n24331 & ~n24827 ;
  assign n24829 = ~n24825 & n24828 ;
  assign n24830 = ~n24294 & ~n24829 ;
  assign n24843 = ~n24284 & n24566 ;
  assign n24844 = n24302 & ~n24843 ;
  assign n24818 = ~n24302 & n24817 ;
  assign n24845 = ~n24326 & ~n24818 ;
  assign n24846 = ~n24844 & n24845 ;
  assign n24847 = ~n24830 & n24846 ;
  assign n24848 = ~n24842 & n24847 ;
  assign n24849 = ~\u2_L1_reg[1]/NET0131  & ~n24848 ;
  assign n24850 = \u2_L1_reg[1]/NET0131  & n24848 ;
  assign n24851 = ~n24849 & ~n24850 ;
  assign n24856 = ~n23957 & ~n24231 ;
  assign n24852 = n23932 & n23988 ;
  assign n24853 = ~n23978 & ~n24852 ;
  assign n24854 = n23958 & n23959 ;
  assign n24855 = ~n23953 & ~n24854 ;
  assign n24857 = n24853 & n24855 ;
  assign n24858 = n24856 & n24857 ;
  assign n24859 = n23932 & n23963 ;
  assign n24860 = n23953 & ~n24859 ;
  assign n24861 = ~n23947 & n24860 ;
  assign n24862 = ~n24858 & ~n24861 ;
  assign n24863 = n23986 & n23989 ;
  assign n24864 = n23920 & ~n24233 ;
  assign n24865 = ~n24863 & n24864 ;
  assign n24866 = ~n24862 & n24865 ;
  assign n24868 = n23953 & ~n24852 ;
  assign n24869 = ~n23981 & ~n23995 ;
  assign n24870 = n24855 & n24869 ;
  assign n24871 = ~n24868 & ~n24870 ;
  assign n24872 = ~n23920 & ~n23965 ;
  assign n24867 = ~n23932 & n23980 ;
  assign n24873 = ~n24230 & ~n24867 ;
  assign n24874 = n24872 & n24873 ;
  assign n24875 = ~n24871 & n24874 ;
  assign n24876 = ~n24866 & ~n24875 ;
  assign n24877 = ~n23963 & n23970 ;
  assign n24878 = n23996 & n24877 ;
  assign n24879 = n23933 & ~n23953 ;
  assign n24880 = n23969 & n24879 ;
  assign n24881 = ~n24878 & ~n24880 ;
  assign n24882 = ~n24876 & n24881 ;
  assign n24883 = \u2_L1_reg[23]/NET0131  & ~n24882 ;
  assign n24884 = ~\u2_L1_reg[23]/NET0131  & n24882 ;
  assign n24885 = ~n24883 & ~n24884 ;
  assign n24888 = ~n24660 & ~n24681 ;
  assign n24889 = ~n24683 & n24888 ;
  assign n24890 = ~n24704 & ~n24726 ;
  assign n24891 = ~n24889 & n24890 ;
  assign n24892 = n24692 & ~n24891 ;
  assign n24893 = ~n24673 & n24694 ;
  assign n24894 = ~n24682 & ~n24893 ;
  assign n24895 = ~n24692 & ~n24894 ;
  assign n24886 = n24660 & ~n24680 ;
  assign n24887 = n24673 & n24886 ;
  assign n24896 = n24674 & n24680 ;
  assign n24897 = ~n24887 & ~n24896 ;
  assign n24898 = ~n24895 & n24897 ;
  assign n24899 = ~n24892 & n24898 ;
  assign n24900 = n24717 & ~n24899 ;
  assign n24910 = ~n24740 & ~n24896 ;
  assign n24911 = ~n24680 & n24702 ;
  assign n24912 = ~n24673 & n24911 ;
  assign n24913 = n24910 & ~n24912 ;
  assign n24914 = n24692 & ~n24913 ;
  assign n24901 = n24666 & ~n24692 ;
  assign n24902 = ~n24681 & ~n24901 ;
  assign n24903 = ~n24660 & ~n24695 ;
  assign n24904 = ~n24902 & n24903 ;
  assign n24905 = n24692 & ~n24744 ;
  assign n24906 = ~n24666 & n24700 ;
  assign n24907 = ~n24905 & n24906 ;
  assign n24908 = ~n24904 & ~n24907 ;
  assign n24909 = ~n24717 & ~n24908 ;
  assign n24915 = n24699 & n24901 ;
  assign n24916 = ~n24727 & ~n24915 ;
  assign n24917 = ~n24909 & n24916 ;
  assign n24918 = ~n24914 & n24917 ;
  assign n24919 = ~n24900 & n24918 ;
  assign n24920 = ~\u2_L1_reg[25]/NET0131  & ~n24919 ;
  assign n24921 = \u2_L1_reg[25]/NET0131  & n24919 ;
  assign n24922 = ~n24920 & ~n24921 ;
  assign n24924 = n24276 & ~n24344 ;
  assign n24923 = n24283 & n24322 ;
  assign n24925 = ~n24303 & ~n24923 ;
  assign n24926 = ~n24924 & n24925 ;
  assign n24927 = ~n24324 & ~n24926 ;
  assign n24928 = ~n24295 & ~n24315 ;
  assign n24929 = ~n24302 & ~n24334 ;
  assign n24930 = ~n24928 & n24929 ;
  assign n24931 = n24294 & ~n24930 ;
  assign n24932 = ~n24927 & n24931 ;
  assign n24933 = ~n24551 & ~n24838 ;
  assign n24934 = ~n24302 & ~n24933 ;
  assign n24935 = n24313 & ~n24322 ;
  assign n24936 = ~n24294 & ~n24335 ;
  assign n24937 = ~n24935 & n24936 ;
  assign n24938 = n24330 & n24937 ;
  assign n24939 = ~n24934 & n24938 ;
  assign n24940 = ~n24932 & ~n24939 ;
  assign n24941 = ~n24276 & n24306 ;
  assign n24942 = ~n24277 & ~n24296 ;
  assign n24943 = ~n24941 & n24942 ;
  assign n24944 = n24557 & ~n24943 ;
  assign n24945 = n24263 & n24302 ;
  assign n24946 = ~n24336 & n24945 ;
  assign n24947 = ~n24944 & ~n24946 ;
  assign n24948 = ~n24940 & n24947 ;
  assign n24949 = ~\u2_L1_reg[26]/NET0131  & ~n24948 ;
  assign n24950 = \u2_L1_reg[26]/NET0131  & n24948 ;
  assign n24951 = ~n24949 & ~n24950 ;
  assign n24952 = ~n24145 & ~n24786 ;
  assign n24953 = ~n24791 & n24952 ;
  assign n24954 = ~n24157 & ~n24953 ;
  assign n24955 = n24157 & ~n24164 ;
  assign n24956 = ~n24632 & n24955 ;
  assign n24957 = ~n24140 & ~n24646 ;
  assign n24958 = ~n24183 & n24957 ;
  assign n24959 = ~n24956 & n24958 ;
  assign n24960 = ~n24954 & n24959 ;
  assign n24961 = n24113 & ~n24960 ;
  assign n24968 = n24165 & ~n24181 ;
  assign n24969 = n24157 & ~n24631 ;
  assign n24970 = ~n24968 & n24969 ;
  assign n24966 = n24125 & n24132 ;
  assign n24967 = n24624 & n24966 ;
  assign n24971 = ~n24804 & ~n24967 ;
  assign n24972 = ~n24162 & n24971 ;
  assign n24973 = ~n24970 & n24972 ;
  assign n24974 = ~n24113 & ~n24973 ;
  assign n24962 = n24157 & n24182 ;
  assign n24963 = n24165 & ~n24169 ;
  assign n24964 = ~n24150 & ~n24963 ;
  assign n24965 = ~n24157 & ~n24964 ;
  assign n24975 = ~n24962 & ~n24965 ;
  assign n24976 = ~n24974 & n24975 ;
  assign n24977 = ~n24961 & n24976 ;
  assign n24978 = ~\u2_L1_reg[27]/NET0131  & ~n24977 ;
  assign n24979 = \u2_L1_reg[27]/NET0131  & n24977 ;
  assign n24980 = ~n24978 & ~n24979 ;
  assign n24998 = ~n23855 & ~n23899 ;
  assign n24999 = ~n23839 & n24204 ;
  assign n25000 = ~n24998 & ~n24999 ;
  assign n24985 = ~n23839 & n23898 ;
  assign n25001 = n23833 & n24985 ;
  assign n25002 = ~n25000 & ~n25001 ;
  assign n25003 = ~n23878 & ~n25002 ;
  assign n25004 = n23833 & n24196 ;
  assign n25005 = ~n23839 & ~n23878 ;
  assign n25006 = n25004 & ~n25005 ;
  assign n25007 = ~n23839 & n23855 ;
  assign n25008 = ~n23861 & ~n25007 ;
  assign n25009 = n23878 & ~n25008 ;
  assign n25010 = ~n25006 & ~n25009 ;
  assign n25011 = ~n25003 & n25010 ;
  assign n25012 = n23868 & ~n25011 ;
  assign n24981 = ~n23833 & n24196 ;
  assign n24982 = ~n23859 & ~n23860 ;
  assign n24983 = ~n24981 & ~n24982 ;
  assign n24984 = ~n23878 & ~n24983 ;
  assign n24986 = n23878 & ~n24981 ;
  assign n24987 = ~n24985 & n24986 ;
  assign n24988 = ~n24984 & ~n24987 ;
  assign n24989 = n23839 & n24981 ;
  assign n24990 = n23860 & n23887 ;
  assign n24991 = ~n24989 & ~n24990 ;
  assign n24992 = n23858 & n24991 ;
  assign n24993 = ~n24988 & n24992 ;
  assign n24994 = ~n23868 & ~n24993 ;
  assign n24995 = n23854 & n23878 ;
  assign n24996 = n23896 & ~n24196 ;
  assign n24997 = n23888 & n24996 ;
  assign n25013 = ~n24995 & ~n24997 ;
  assign n25014 = ~n24994 & n25013 ;
  assign n25015 = ~n25012 & n25014 ;
  assign n25016 = \u2_L1_reg[32]/NET0131  & n25015 ;
  assign n25017 = ~\u2_L1_reg[32]/NET0131  & ~n25015 ;
  assign n25018 = ~n25016 & ~n25017 ;
  assign n25052 = decrypt_pad & ~\u2_uk_K_r1_reg[46]/NET0131  ;
  assign n25053 = ~decrypt_pad & ~\u2_uk_K_r1_reg[13]/NET0131  ;
  assign n25054 = ~n25052 & ~n25053 ;
  assign n25055 = \u2_R1_reg[12]/NET0131  & ~n25054 ;
  assign n25056 = ~\u2_R1_reg[12]/NET0131  & n25054 ;
  assign n25057 = ~n25055 & ~n25056 ;
  assign n25019 = decrypt_pad & ~\u2_uk_K_r1_reg[34]/NET0131  ;
  assign n25020 = ~decrypt_pad & ~\u2_uk_K_r1_reg[26]/NET0131  ;
  assign n25021 = ~n25019 & ~n25020 ;
  assign n25022 = \u2_R1_reg[13]/NET0131  & ~n25021 ;
  assign n25023 = ~\u2_R1_reg[13]/NET0131  & n25021 ;
  assign n25024 = ~n25022 & ~n25023 ;
  assign n25032 = decrypt_pad & ~\u2_uk_K_r1_reg[25]/NET0131  ;
  assign n25033 = ~decrypt_pad & ~\u2_uk_K_r1_reg[17]/NET0131  ;
  assign n25034 = ~n25032 & ~n25033 ;
  assign n25035 = \u2_R1_reg[8]/NET0131  & ~n25034 ;
  assign n25036 = ~\u2_R1_reg[8]/NET0131  & n25034 ;
  assign n25037 = ~n25035 & ~n25036 ;
  assign n25039 = ~n25024 & ~n25037 ;
  assign n25040 = n25024 & n25037 ;
  assign n25041 = ~n25039 & ~n25040 ;
  assign n25025 = decrypt_pad & ~\u2_uk_K_r1_reg[54]/NET0131  ;
  assign n25026 = ~decrypt_pad & ~\u2_uk_K_r1_reg[46]/NET0131  ;
  assign n25027 = ~n25025 & ~n25026 ;
  assign n25028 = \u2_R1_reg[9]/NET0131  & ~n25027 ;
  assign n25029 = ~\u2_R1_reg[9]/NET0131  & n25027 ;
  assign n25030 = ~n25028 & ~n25029 ;
  assign n25042 = decrypt_pad & ~\u2_uk_K_r1_reg[5]/NET0131  ;
  assign n25043 = ~decrypt_pad & ~\u2_uk_K_r1_reg[54]/NET0131  ;
  assign n25044 = ~n25042 & ~n25043 ;
  assign n25045 = \u2_R1_reg[10]/NET0131  & ~n25044 ;
  assign n25046 = ~\u2_R1_reg[10]/NET0131  & n25044 ;
  assign n25047 = ~n25045 & ~n25046 ;
  assign n25093 = ~n25030 & n25047 ;
  assign n25094 = ~n25041 & n25093 ;
  assign n25082 = n25024 & ~n25037 ;
  assign n25083 = n25030 & n25082 ;
  assign n25064 = decrypt_pad & ~\u2_uk_K_r1_reg[6]/NET0131  ;
  assign n25065 = ~decrypt_pad & ~\u2_uk_K_r1_reg[55]/NET0131  ;
  assign n25066 = ~n25064 & ~n25065 ;
  assign n25067 = \u2_R1_reg[11]/P0001  & ~n25066 ;
  assign n25068 = ~\u2_R1_reg[11]/P0001  & n25066 ;
  assign n25069 = ~n25067 & ~n25068 ;
  assign n25084 = n25047 & ~n25069 ;
  assign n25085 = n25083 & n25084 ;
  assign n25090 = ~n25024 & n25030 ;
  assign n25091 = n25047 & n25090 ;
  assign n25092 = n25037 & n25091 ;
  assign n25095 = ~n25085 & ~n25092 ;
  assign n25096 = ~n25094 & n25095 ;
  assign n25075 = n25030 & ~n25047 ;
  assign n25086 = n25024 & n25069 ;
  assign n25087 = n25041 & ~n25086 ;
  assign n25088 = n25075 & ~n25087 ;
  assign n25059 = ~n25030 & ~n25047 ;
  assign n25089 = n25059 & n25087 ;
  assign n25097 = ~n25088 & ~n25089 ;
  assign n25098 = n25096 & n25097 ;
  assign n25099 = ~n25057 & ~n25098 ;
  assign n25031 = n25024 & ~n25030 ;
  assign n25038 = ~n25030 & n25037 ;
  assign n25048 = ~n25037 & ~n25047 ;
  assign n25049 = ~n25038 & ~n25048 ;
  assign n25050 = n25041 & n25049 ;
  assign n25051 = ~n25031 & ~n25050 ;
  assign n25058 = ~n25051 & n25057 ;
  assign n25060 = n25039 & n25059 ;
  assign n25061 = n25031 & n25047 ;
  assign n25062 = ~n25060 & ~n25061 ;
  assign n25063 = ~n25058 & n25062 ;
  assign n25070 = ~n25063 & n25069 ;
  assign n25071 = n25047 & n25057 ;
  assign n25072 = n25030 & n25039 ;
  assign n25073 = n25071 & n25072 ;
  assign n25074 = n25057 & ~n25069 ;
  assign n25076 = n25024 & n25075 ;
  assign n25077 = ~n25024 & n25038 ;
  assign n25078 = n25030 & n25040 ;
  assign n25079 = ~n25077 & ~n25078 ;
  assign n25080 = ~n25076 & n25079 ;
  assign n25081 = n25074 & ~n25080 ;
  assign n25100 = ~n25073 & ~n25081 ;
  assign n25101 = ~n25070 & n25100 ;
  assign n25102 = ~n25099 & n25101 ;
  assign n25103 = ~\u2_L1_reg[6]/NET0131  & ~n25102 ;
  assign n25104 = \u2_L1_reg[6]/NET0131  & n25102 ;
  assign n25105 = ~n25103 & ~n25104 ;
  assign n25106 = n23839 & ~n24204 ;
  assign n25107 = ~n24985 & ~n25106 ;
  assign n25108 = n23833 & ~n25107 ;
  assign n25109 = ~n23833 & ~n23859 ;
  assign n25110 = n24204 & n25109 ;
  assign n25111 = n23878 & ~n25110 ;
  assign n25112 = ~n23846 & ~n24206 ;
  assign n25113 = ~n23878 & ~n25004 ;
  assign n25114 = ~n25106 & n25113 ;
  assign n25115 = ~n25112 & n25114 ;
  assign n25116 = ~n25111 & ~n25115 ;
  assign n25117 = ~n25108 & ~n25116 ;
  assign n25118 = n23868 & ~n25117 ;
  assign n25126 = ~n23878 & n25110 ;
  assign n25127 = ~n23890 & ~n25126 ;
  assign n25128 = ~n23868 & ~n25127 ;
  assign n25120 = ~n24198 & ~n24204 ;
  assign n25121 = ~n23856 & ~n24990 ;
  assign n25122 = ~n25120 & n25121 ;
  assign n25119 = n23868 & ~n23890 ;
  assign n25123 = n23878 & ~n25119 ;
  assign n25124 = ~n25122 & n25123 ;
  assign n25125 = ~n23878 & n25108 ;
  assign n25129 = ~n25124 & ~n25125 ;
  assign n25130 = ~n25128 & n25129 ;
  assign n25131 = ~n25118 & n25130 ;
  assign n25132 = ~\u2_L1_reg[7]/NET0131  & ~n25131 ;
  assign n25133 = \u2_L1_reg[7]/NET0131  & n25131 ;
  assign n25134 = ~n25132 & ~n25133 ;
  assign n25139 = n24692 & ~n24729 ;
  assign n25140 = ~n24726 & n25139 ;
  assign n25141 = ~n24699 & n24702 ;
  assign n25142 = ~n24692 & ~n24893 ;
  assign n25143 = ~n25141 & n25142 ;
  assign n25144 = ~n25140 & ~n25143 ;
  assign n25145 = ~n24682 & n24910 ;
  assign n25146 = ~n25144 & n25145 ;
  assign n25147 = ~n24717 & ~n25146 ;
  assign n25148 = n24728 & n24739 ;
  assign n25149 = ~n24893 & ~n25148 ;
  assign n25150 = n24692 & ~n25149 ;
  assign n25151 = ~n24680 & n24901 ;
  assign n25152 = n24747 & ~n25151 ;
  assign n25153 = ~n25150 & n25152 ;
  assign n25154 = n24717 & ~n25153 ;
  assign n25135 = ~n24700 & n24702 ;
  assign n25136 = ~n24720 & ~n25135 ;
  assign n25137 = n24692 & ~n25136 ;
  assign n25138 = ~n24660 & n24915 ;
  assign n25155 = ~n25137 & ~n25138 ;
  assign n25156 = ~n25154 & n25155 ;
  assign n25157 = ~n25147 & n25156 ;
  assign n25158 = ~\u2_L1_reg[8]/NET0131  & ~n25157 ;
  assign n25159 = \u2_L1_reg[8]/NET0131  & n25157 ;
  assign n25160 = ~n25158 & ~n25159 ;
  assign n25161 = n25047 & ~n25083 ;
  assign n25163 = n25069 & n25072 ;
  assign n25162 = n25031 & ~n25037 ;
  assign n25164 = ~n25047 & ~n25162 ;
  assign n25165 = n25079 & n25164 ;
  assign n25166 = ~n25163 & n25165 ;
  assign n25167 = ~n25161 & ~n25166 ;
  assign n25168 = n25039 & n25047 ;
  assign n25169 = ~n25030 & n25168 ;
  assign n25170 = n25069 & ~n25092 ;
  assign n25171 = ~n25169 & n25170 ;
  assign n25172 = n25037 & n25047 ;
  assign n25173 = ~n25024 & ~n25048 ;
  assign n25174 = ~n25172 & n25173 ;
  assign n25175 = ~n25171 & n25174 ;
  assign n25176 = ~n25167 & ~n25175 ;
  assign n25177 = n25057 & ~n25176 ;
  assign n25178 = ~n25030 & n25172 ;
  assign n25179 = ~n25069 & ~n25178 ;
  assign n25180 = ~n25171 & ~n25179 ;
  assign n25185 = n25039 & ~n25047 ;
  assign n25186 = ~n25078 & ~n25162 ;
  assign n25187 = ~n25185 & n25186 ;
  assign n25188 = ~n25069 & ~n25187 ;
  assign n25182 = ~n25039 & n25069 ;
  assign n25181 = ~n25030 & ~n25040 ;
  assign n25183 = ~n25078 & ~n25181 ;
  assign n25184 = n25182 & n25183 ;
  assign n25189 = ~n25060 & ~n25184 ;
  assign n25190 = ~n25188 & n25189 ;
  assign n25191 = ~n25057 & ~n25190 ;
  assign n25192 = ~n25180 & ~n25191 ;
  assign n25193 = ~n25177 & n25192 ;
  assign n25194 = ~\u2_L1_reg[16]/NET0131  & ~n25193 ;
  assign n25195 = \u2_L1_reg[16]/NET0131  & n25193 ;
  assign n25196 = ~n25194 & ~n25195 ;
  assign n25206 = ~n25047 & n25069 ;
  assign n25217 = ~n25030 & ~n25082 ;
  assign n25218 = n25206 & n25217 ;
  assign n25213 = ~n25059 & ~n25069 ;
  assign n25214 = ~n25041 & n25213 ;
  assign n25215 = ~n25038 & n25047 ;
  assign n25216 = n25182 & n25215 ;
  assign n25219 = ~n25214 & ~n25216 ;
  assign n25220 = ~n25218 & n25219 ;
  assign n25221 = ~n25089 & n25220 ;
  assign n25222 = n25057 & ~n25221 ;
  assign n25197 = n25024 & n25048 ;
  assign n25198 = ~n25168 & ~n25197 ;
  assign n25199 = ~n25072 & ~n25178 ;
  assign n25200 = n25198 & n25199 ;
  assign n25201 = n25069 & ~n25200 ;
  assign n25202 = ~n25024 & n25178 ;
  assign n25203 = ~n25201 & ~n25202 ;
  assign n25204 = ~n25057 & ~n25203 ;
  assign n25209 = ~n25041 & n25059 ;
  assign n25210 = ~n25050 & ~n25209 ;
  assign n25211 = ~n25057 & ~n25069 ;
  assign n25212 = ~n25210 & n25211 ;
  assign n25205 = n25078 & n25084 ;
  assign n25207 = ~n25077 & ~n25083 ;
  assign n25208 = n25206 & ~n25207 ;
  assign n25223 = ~n25205 & ~n25208 ;
  assign n25224 = ~n25212 & n25223 ;
  assign n25225 = ~n25204 & n25224 ;
  assign n25226 = ~n25222 & n25225 ;
  assign n25227 = ~\u2_L1_reg[24]/NET0131  & ~n25226 ;
  assign n25228 = \u2_L1_reg[24]/NET0131  & n25226 ;
  assign n25229 = ~n25227 & ~n25228 ;
  assign n25231 = ~n25047 & n25077 ;
  assign n25232 = n25198 & ~n25231 ;
  assign n25233 = n25057 & ~n25232 ;
  assign n25234 = ~n25090 & ~n25172 ;
  assign n25235 = ~n25057 & ~n25091 ;
  assign n25236 = ~n25234 & n25235 ;
  assign n25237 = ~n25233 & ~n25236 ;
  assign n25238 = n25069 & ~n25237 ;
  assign n25242 = n25047 & n25162 ;
  assign n25239 = ~n25030 & ~n25037 ;
  assign n25240 = ~n25069 & ~n25239 ;
  assign n25241 = n25234 & n25240 ;
  assign n25243 = ~n25209 & ~n25241 ;
  assign n25244 = ~n25242 & n25243 ;
  assign n25245 = ~n25057 & ~n25244 ;
  assign n25246 = ~n25072 & ~n25172 ;
  assign n25247 = n25074 & ~n25246 ;
  assign n25249 = n25030 & ~n25040 ;
  assign n25250 = n25071 & n25249 ;
  assign n25230 = n25084 & n25090 ;
  assign n25248 = n25086 & n25178 ;
  assign n25251 = ~n25230 & ~n25248 ;
  assign n25252 = ~n25250 & n25251 ;
  assign n25253 = ~n25247 & n25252 ;
  assign n25254 = ~n25245 & n25253 ;
  assign n25255 = ~n25238 & n25254 ;
  assign n25256 = \u2_L1_reg[30]/NET0131  & ~n25255 ;
  assign n25257 = ~\u2_L1_reg[30]/NET0131  & n25255 ;
  assign n25258 = ~n25256 & ~n25257 ;
  assign n25260 = n24666 & ~n24886 ;
  assign n25261 = n24692 & ~n24702 ;
  assign n25262 = ~n24704 & n25261 ;
  assign n25263 = ~n25260 & n25262 ;
  assign n25259 = n24667 & n24699 ;
  assign n25264 = ~n24703 & n24717 ;
  assign n25265 = ~n25259 & n25264 ;
  assign n25266 = ~n24727 & n25265 ;
  assign n25267 = ~n25263 & n25266 ;
  assign n25272 = ~n24674 & ~n24911 ;
  assign n25273 = n24692 & ~n25272 ;
  assign n25268 = n24692 & ~n24699 ;
  assign n25269 = ~n24739 & ~n24744 ;
  assign n25270 = ~n24893 & n25269 ;
  assign n25271 = ~n25268 & ~n25270 ;
  assign n25274 = ~n24717 & ~n25271 ;
  assign n25275 = ~n25273 & n25274 ;
  assign n25276 = ~n25267 & ~n25275 ;
  assign n25277 = ~n24745 & n25139 ;
  assign n25278 = ~n24692 & ~n24724 ;
  assign n25279 = ~n25148 & n25278 ;
  assign n25280 = ~n24741 & n25279 ;
  assign n25281 = ~n25277 & ~n25280 ;
  assign n25282 = ~n25276 & ~n25281 ;
  assign n25283 = ~\u2_L1_reg[3]/NET0131  & ~n25282 ;
  assign n25284 = \u2_L1_reg[3]/NET0131  & n25282 ;
  assign n25285 = ~n25283 & ~n25284 ;
  assign n25286 = ~n23926 & n24242 ;
  assign n25287 = ~n23955 & ~n24859 ;
  assign n25288 = ~n23953 & n25287 ;
  assign n25289 = ~n23940 & ~n23958 ;
  assign n25290 = n24868 & n25289 ;
  assign n25291 = ~n25288 & ~n25290 ;
  assign n25292 = ~n25286 & ~n25291 ;
  assign n25293 = ~n23920 & ~n25292 ;
  assign n25301 = n23920 & n24243 ;
  assign n25302 = n24853 & n25301 ;
  assign n25300 = ~n23920 & ~n24246 ;
  assign n25303 = n23926 & ~n25300 ;
  assign n25304 = ~n25302 & n25303 ;
  assign n25294 = n23970 & ~n25287 ;
  assign n25295 = ~n24231 & ~n25294 ;
  assign n25296 = n23920 & ~n25295 ;
  assign n25297 = n23926 & n24859 ;
  assign n25298 = ~n25286 & ~n25297 ;
  assign n25299 = ~n23953 & ~n25298 ;
  assign n25305 = ~n25296 & ~n25299 ;
  assign n25306 = ~n25304 & n25305 ;
  assign n25307 = ~n25293 & n25306 ;
  assign n25308 = ~\u2_L1_reg[9]/NET0131  & ~n25307 ;
  assign n25309 = \u2_L1_reg[9]/NET0131  & n25307 ;
  assign n25310 = ~n25308 & ~n25309 ;
  assign n25314 = n24389 & ~n24480 ;
  assign n25311 = n24379 & n24404 ;
  assign n25312 = ~n24422 & ~n25311 ;
  assign n25313 = ~n24389 & ~n25312 ;
  assign n25315 = ~n24509 & ~n25313 ;
  assign n25316 = ~n25314 & n25315 ;
  assign n25317 = n24396 & ~n25316 ;
  assign n25321 = ~n24382 & ~n24607 ;
  assign n25322 = ~n24473 & n25321 ;
  assign n25318 = n24389 & n24421 ;
  assign n25319 = ~n24372 & ~n24594 ;
  assign n25320 = ~n24492 & n25319 ;
  assign n25323 = ~n25318 & ~n25320 ;
  assign n25324 = n25322 & n25323 ;
  assign n25325 = ~n24396 & ~n25324 ;
  assign n25326 = ~n24389 & n24400 ;
  assign n25327 = n24365 & n24411 ;
  assign n25328 = ~n24604 & ~n25327 ;
  assign n25329 = n24389 & ~n25328 ;
  assign n25330 = ~n25326 & ~n25329 ;
  assign n25331 = ~n25325 & n25330 ;
  assign n25332 = ~n25317 & n25331 ;
  assign n25333 = ~\u2_L1_reg[18]/P0001  & ~n25332 ;
  assign n25334 = \u2_L1_reg[18]/P0001  & n25332 ;
  assign n25335 = ~n25333 & ~n25334 ;
  assign n25342 = decrypt_pad & ~\u2_uk_K_r0_reg[50]/NET0131  ;
  assign n25343 = ~decrypt_pad & ~\u2_uk_K_r0_reg[16]/NET0131  ;
  assign n25344 = ~n25342 & ~n25343 ;
  assign n25345 = \u2_R0_reg[23]/NET0131  & ~n25344 ;
  assign n25346 = ~\u2_R0_reg[23]/NET0131  & n25344 ;
  assign n25347 = ~n25345 & ~n25346 ;
  assign n25348 = decrypt_pad & ~\u2_uk_K_r0_reg[37]/NET0131  ;
  assign n25349 = ~decrypt_pad & ~\u2_uk_K_r0_reg[31]/NET0131  ;
  assign n25350 = ~n25348 & ~n25349 ;
  assign n25351 = \u2_R0_reg[22]/NET0131  & ~n25350 ;
  assign n25352 = ~\u2_R0_reg[22]/NET0131  & n25350 ;
  assign n25353 = ~n25351 & ~n25352 ;
  assign n25355 = decrypt_pad & ~\u2_uk_K_r0_reg[0]/NET0131  ;
  assign n25356 = ~decrypt_pad & ~\u2_uk_K_r0_reg[21]/NET0131  ;
  assign n25357 = ~n25355 & ~n25356 ;
  assign n25358 = \u2_R0_reg[20]/NET0131  & ~n25357 ;
  assign n25359 = ~\u2_R0_reg[20]/NET0131  & n25357 ;
  assign n25360 = ~n25358 & ~n25359 ;
  assign n25377 = decrypt_pad & ~\u2_uk_K_r0_reg[16]/NET0131  ;
  assign n25378 = ~decrypt_pad & ~\u2_uk_K_r0_reg[37]/NET0131  ;
  assign n25379 = ~n25377 & ~n25378 ;
  assign n25380 = \u2_R0_reg[25]/NET0131  & ~n25379 ;
  assign n25381 = ~\u2_R0_reg[25]/NET0131  & n25379 ;
  assign n25382 = ~n25380 & ~n25381 ;
  assign n25383 = n25360 & ~n25382 ;
  assign n25362 = decrypt_pad & ~\u2_uk_K_r0_reg[15]/NET0131  ;
  assign n25363 = ~decrypt_pad & ~\u2_uk_K_r0_reg[36]/NET0131  ;
  assign n25364 = ~n25362 & ~n25363 ;
  assign n25365 = \u2_R0_reg[21]/NET0131  & ~n25364 ;
  assign n25366 = ~\u2_R0_reg[21]/NET0131  & n25364 ;
  assign n25367 = ~n25365 & ~n25366 ;
  assign n25389 = ~n25360 & ~n25367 ;
  assign n25417 = ~n25383 & ~n25389 ;
  assign n25418 = n25353 & n25417 ;
  assign n25419 = n25367 & n25382 ;
  assign n25420 = ~n25360 & n25419 ;
  assign n25386 = n25360 & n25382 ;
  assign n25387 = ~n25367 & n25386 ;
  assign n25421 = ~n25353 & ~n25387 ;
  assign n25422 = ~n25420 & n25421 ;
  assign n25423 = ~n25418 & ~n25422 ;
  assign n25424 = ~n25347 & ~n25423 ;
  assign n25336 = decrypt_pad & ~\u2_uk_K_r0_reg[21]/NET0131  ;
  assign n25337 = ~decrypt_pad & ~\u2_uk_K_r0_reg[42]/NET0131  ;
  assign n25338 = ~n25336 & ~n25337 ;
  assign n25339 = \u2_R0_reg[24]/NET0131  & ~n25338 ;
  assign n25340 = ~\u2_R0_reg[24]/NET0131  & n25338 ;
  assign n25341 = ~n25339 & ~n25340 ;
  assign n25368 = n25353 & ~n25360 ;
  assign n25369 = n25367 & n25368 ;
  assign n25414 = n25347 & ~n25369 ;
  assign n25411 = ~n25353 & ~n25367 ;
  assign n25412 = n25383 & n25411 ;
  assign n25413 = n25367 & n25386 ;
  assign n25415 = ~n25412 & ~n25413 ;
  assign n25416 = n25414 & n25415 ;
  assign n25425 = n25341 & ~n25416 ;
  assign n25426 = ~n25424 & n25425 ;
  assign n25370 = ~n25353 & n25367 ;
  assign n25392 = n25370 & ~n25382 ;
  assign n25393 = n25360 & n25392 ;
  assign n25388 = n25353 & n25387 ;
  assign n25390 = n25382 & n25389 ;
  assign n25391 = n25347 & n25390 ;
  assign n25396 = ~n25388 & ~n25391 ;
  assign n25397 = ~n25393 & n25396 ;
  assign n25371 = n25360 & n25370 ;
  assign n25372 = ~n25369 & ~n25371 ;
  assign n25373 = ~n25347 & ~n25372 ;
  assign n25384 = ~n25347 & ~n25353 ;
  assign n25385 = n25383 & n25384 ;
  assign n25354 = n25347 & ~n25353 ;
  assign n25361 = n25354 & ~n25360 ;
  assign n25374 = n25360 & ~n25367 ;
  assign n25375 = n25347 & n25353 ;
  assign n25376 = n25374 & n25375 ;
  assign n25394 = ~n25361 & ~n25376 ;
  assign n25395 = ~n25385 & n25394 ;
  assign n25398 = ~n25373 & n25395 ;
  assign n25399 = n25397 & n25398 ;
  assign n25400 = ~n25341 & ~n25399 ;
  assign n25405 = n25367 & n25383 ;
  assign n25406 = ~n25347 & n25405 ;
  assign n25407 = ~n25391 & ~n25406 ;
  assign n25408 = ~n25353 & ~n25407 ;
  assign n25401 = n25353 & n25386 ;
  assign n25402 = ~n25360 & n25392 ;
  assign n25403 = ~n25401 & ~n25402 ;
  assign n25404 = n25347 & ~n25403 ;
  assign n25409 = ~n25382 & n25389 ;
  assign n25410 = n25384 & n25409 ;
  assign n25427 = ~n25404 & ~n25410 ;
  assign n25428 = ~n25408 & n25427 ;
  assign n25429 = ~n25400 & n25428 ;
  assign n25430 = ~n25426 & n25429 ;
  assign n25431 = ~\u2_L0_reg[11]/NET0131  & n25430 ;
  assign n25432 = \u2_L0_reg[11]/NET0131  & ~n25430 ;
  assign n25433 = ~n25431 & ~n25432 ;
  assign n25434 = decrypt_pad & ~\u2_uk_K_r0_reg[8]/NET0131  ;
  assign n25435 = ~decrypt_pad & ~\u2_uk_K_r0_reg[29]/NET0131  ;
  assign n25436 = ~n25434 & ~n25435 ;
  assign n25437 = \u2_R0_reg[26]/NET0131  & ~n25436 ;
  assign n25438 = ~\u2_R0_reg[26]/NET0131  & n25436 ;
  assign n25439 = ~n25437 & ~n25438 ;
  assign n25440 = decrypt_pad & ~\u2_uk_K_r0_reg[23]/NET0131  ;
  assign n25441 = ~decrypt_pad & ~\u2_uk_K_r0_reg[44]/NET0131  ;
  assign n25442 = ~n25440 & ~n25441 ;
  assign n25443 = \u2_R0_reg[25]/NET0131  & ~n25442 ;
  assign n25444 = ~\u2_R0_reg[25]/NET0131  & n25442 ;
  assign n25445 = ~n25443 & ~n25444 ;
  assign n25446 = n25439 & ~n25445 ;
  assign n25447 = decrypt_pad & ~\u2_uk_K_r0_reg[43]/NET0131  ;
  assign n25448 = ~decrypt_pad & ~\u2_uk_K_r0_reg[9]/NET0131  ;
  assign n25449 = ~n25447 & ~n25448 ;
  assign n25450 = \u2_R0_reg[24]/NET0131  & ~n25449 ;
  assign n25451 = ~\u2_R0_reg[24]/NET0131  & n25449 ;
  assign n25452 = ~n25450 & ~n25451 ;
  assign n25453 = decrypt_pad & ~\u2_uk_K_r0_reg[51]/NET0131  ;
  assign n25454 = ~decrypt_pad & ~\u2_uk_K_r0_reg[45]/NET0131  ;
  assign n25455 = ~n25453 & ~n25454 ;
  assign n25456 = \u2_R0_reg[29]/NET0131  & ~n25455 ;
  assign n25457 = ~\u2_R0_reg[29]/NET0131  & n25455 ;
  assign n25458 = ~n25456 & ~n25457 ;
  assign n25459 = ~n25452 & n25458 ;
  assign n25460 = n25446 & n25459 ;
  assign n25461 = ~n25452 & ~n25458 ;
  assign n25462 = n25439 & n25461 ;
  assign n25463 = n25445 & n25462 ;
  assign n25464 = ~n25460 & ~n25463 ;
  assign n25465 = ~n25445 & ~n25458 ;
  assign n25466 = n25445 & n25458 ;
  assign n25467 = ~n25439 & n25466 ;
  assign n25468 = ~n25446 & ~n25467 ;
  assign n25469 = decrypt_pad & ~\u2_uk_K_r0_reg[28]/NET0131  ;
  assign n25470 = ~decrypt_pad & ~\u2_uk_K_r0_reg[49]/NET0131  ;
  assign n25471 = ~n25469 & ~n25470 ;
  assign n25472 = \u2_R0_reg[28]/NET0131  & ~n25471 ;
  assign n25473 = ~\u2_R0_reg[28]/NET0131  & n25471 ;
  assign n25474 = ~n25472 & ~n25473 ;
  assign n25475 = ~n25468 & n25474 ;
  assign n25476 = ~n25465 & ~n25475 ;
  assign n25477 = n25452 & ~n25476 ;
  assign n25478 = n25464 & ~n25477 ;
  assign n25479 = decrypt_pad & ~\u2_uk_K_r0_reg[45]/NET0131  ;
  assign n25480 = ~decrypt_pad & ~\u2_uk_K_r0_reg[7]/NET0131  ;
  assign n25481 = ~n25479 & ~n25480 ;
  assign n25482 = \u2_R0_reg[27]/NET0131  & ~n25481 ;
  assign n25483 = ~\u2_R0_reg[27]/NET0131  & n25481 ;
  assign n25484 = ~n25482 & ~n25483 ;
  assign n25485 = ~n25478 & n25484 ;
  assign n25486 = ~n25445 & n25484 ;
  assign n25487 = ~n25439 & n25486 ;
  assign n25488 = ~n25458 & ~n25484 ;
  assign n25489 = ~n25446 & n25488 ;
  assign n25490 = ~n25487 & ~n25489 ;
  assign n25491 = n25452 & ~n25490 ;
  assign n25492 = ~n25439 & ~n25452 ;
  assign n25493 = n25439 & n25452 ;
  assign n25494 = ~n25492 & ~n25493 ;
  assign n25495 = n25458 & ~n25494 ;
  assign n25496 = ~n25445 & n25462 ;
  assign n25497 = ~n25495 & ~n25496 ;
  assign n25498 = ~n25486 & ~n25497 ;
  assign n25499 = ~n25491 & ~n25498 ;
  assign n25500 = ~n25474 & ~n25499 ;
  assign n25504 = n25452 & n25458 ;
  assign n25505 = ~n25439 & ~n25445 ;
  assign n25506 = n25504 & n25505 ;
  assign n25507 = ~n25452 & n25466 ;
  assign n25508 = ~n25506 & ~n25507 ;
  assign n25509 = ~n25484 & ~n25508 ;
  assign n25510 = n25461 & n25505 ;
  assign n25511 = ~n25460 & ~n25510 ;
  assign n25512 = ~n25509 & n25511 ;
  assign n25513 = n25474 & ~n25512 ;
  assign n25501 = ~n25458 & n25487 ;
  assign n25502 = n25445 & ~n25484 ;
  assign n25503 = ~n25494 & n25502 ;
  assign n25514 = ~n25501 & ~n25503 ;
  assign n25515 = ~n25513 & n25514 ;
  assign n25516 = ~n25500 & n25515 ;
  assign n25517 = ~n25485 & n25516 ;
  assign n25518 = ~\u2_L0_reg[22]/NET0131  & ~n25517 ;
  assign n25519 = \u2_L0_reg[22]/NET0131  & n25517 ;
  assign n25520 = ~n25518 & ~n25519 ;
  assign n25521 = decrypt_pad & ~\u2_uk_K_r0_reg[24]/P0001  ;
  assign n25522 = ~decrypt_pad & ~\u2_uk_K_r0_reg[20]/NET0131  ;
  assign n25523 = ~n25521 & ~n25522 ;
  assign n25524 = \u2_R0_reg[4]/NET0131  & ~n25523 ;
  assign n25525 = ~\u2_R0_reg[4]/NET0131  & n25523 ;
  assign n25526 = ~n25524 & ~n25525 ;
  assign n25554 = decrypt_pad & ~\u2_uk_K_r0_reg[46]/NET0131  ;
  assign n25555 = ~decrypt_pad & ~\u2_uk_K_r0_reg[10]/NET0131  ;
  assign n25556 = ~n25554 & ~n25555 ;
  assign n25557 = \u2_R0_reg[3]/NET0131  & ~n25556 ;
  assign n25558 = ~\u2_R0_reg[3]/NET0131  & n25556 ;
  assign n25559 = ~n25557 & ~n25558 ;
  assign n25527 = decrypt_pad & ~\u2_uk_K_r0_reg[12]/NET0131  ;
  assign n25528 = ~decrypt_pad & ~\u2_uk_K_r0_reg[33]/NET0131  ;
  assign n25529 = ~n25527 & ~n25528 ;
  assign n25530 = \u2_R0_reg[2]/NET0131  & ~n25529 ;
  assign n25531 = ~\u2_R0_reg[2]/NET0131  & n25529 ;
  assign n25532 = ~n25530 & ~n25531 ;
  assign n25547 = decrypt_pad & ~\u2_uk_K_r0_reg[33]/NET0131  ;
  assign n25548 = ~decrypt_pad & ~\u2_uk_K_r0_reg[54]/NET0131  ;
  assign n25549 = ~n25547 & ~n25548 ;
  assign n25550 = \u2_R0_reg[32]/NET0131  & ~n25549 ;
  assign n25551 = ~\u2_R0_reg[32]/NET0131  & n25549 ;
  assign n25552 = ~n25550 & ~n25551 ;
  assign n25533 = decrypt_pad & ~\u2_uk_K_r0_reg[54]/NET0131  ;
  assign n25534 = ~decrypt_pad & ~\u2_uk_K_r0_reg[18]/NET0131  ;
  assign n25535 = ~n25533 & ~n25534 ;
  assign n25536 = \u2_R0_reg[1]/NET0131  & ~n25535 ;
  assign n25537 = ~\u2_R0_reg[1]/NET0131  & n25535 ;
  assign n25538 = ~n25536 & ~n25537 ;
  assign n25540 = decrypt_pad & ~\u2_uk_K_r0_reg[27]/NET0131  ;
  assign n25541 = ~decrypt_pad & ~\u2_uk_K_r0_reg[48]/NET0131  ;
  assign n25542 = ~n25540 & ~n25541 ;
  assign n25543 = \u2_R0_reg[5]/NET0131  & ~n25542 ;
  assign n25544 = ~\u2_R0_reg[5]/NET0131  & n25542 ;
  assign n25545 = ~n25543 & ~n25544 ;
  assign n25561 = ~n25538 & ~n25545 ;
  assign n25562 = n25552 & n25561 ;
  assign n25563 = n25532 & n25562 ;
  assign n25564 = ~n25538 & n25545 ;
  assign n25565 = ~n25532 & ~n25552 ;
  assign n25566 = ~n25564 & n25565 ;
  assign n25567 = ~n25563 & ~n25566 ;
  assign n25568 = ~n25559 & ~n25567 ;
  assign n25569 = n25545 & ~n25552 ;
  assign n25570 = n25532 & n25559 ;
  assign n25571 = n25569 & n25570 ;
  assign n25572 = ~n25545 & ~n25552 ;
  assign n25573 = ~n25532 & n25572 ;
  assign n25574 = ~n25571 & ~n25573 ;
  assign n25575 = n25538 & ~n25574 ;
  assign n25539 = n25532 & n25538 ;
  assign n25546 = n25539 & ~n25545 ;
  assign n25553 = n25546 & n25552 ;
  assign n25560 = n25553 & n25559 ;
  assign n25576 = n25545 & n25552 ;
  assign n25577 = ~n25532 & n25559 ;
  assign n25578 = ~n25532 & ~n25538 ;
  assign n25579 = ~n25577 & ~n25578 ;
  assign n25580 = n25576 & ~n25579 ;
  assign n25581 = ~n25560 & ~n25580 ;
  assign n25582 = ~n25575 & n25581 ;
  assign n25583 = ~n25568 & n25582 ;
  assign n25584 = ~n25526 & ~n25583 ;
  assign n25586 = n25532 & n25572 ;
  assign n25587 = ~n25564 & ~n25586 ;
  assign n25588 = n25559 & ~n25587 ;
  assign n25594 = n25538 & ~n25577 ;
  assign n25595 = n25569 & ~n25594 ;
  assign n25585 = ~n25532 & n25562 ;
  assign n25589 = ~n25538 & n25552 ;
  assign n25590 = n25532 & ~n25538 ;
  assign n25591 = n25552 & ~n25559 ;
  assign n25592 = ~n25590 & ~n25591 ;
  assign n25593 = ~n25589 & ~n25592 ;
  assign n25596 = ~n25585 & ~n25593 ;
  assign n25597 = ~n25595 & n25596 ;
  assign n25598 = ~n25588 & n25597 ;
  assign n25599 = n25526 & ~n25598 ;
  assign n25600 = ~n25538 & n25559 ;
  assign n25601 = ~n25532 & n25552 ;
  assign n25602 = ~n25586 & ~n25601 ;
  assign n25603 = n25600 & ~n25602 ;
  assign n25608 = ~n25538 & n25569 ;
  assign n25609 = n25532 & n25608 ;
  assign n25604 = n25539 & n25545 ;
  assign n25605 = n25552 & n25604 ;
  assign n25606 = ~n25532 & n25538 ;
  assign n25607 = ~n25545 & n25606 ;
  assign n25610 = ~n25605 & ~n25607 ;
  assign n25611 = ~n25609 & n25610 ;
  assign n25612 = ~n25559 & ~n25611 ;
  assign n25613 = ~n25603 & ~n25612 ;
  assign n25614 = ~n25599 & n25613 ;
  assign n25615 = ~n25584 & n25614 ;
  assign n25616 = ~\u2_L0_reg[31]/NET0131  & ~n25615 ;
  assign n25617 = \u2_L0_reg[31]/NET0131  & n25615 ;
  assign n25618 = ~n25616 & ~n25617 ;
  assign n25619 = decrypt_pad & ~\u2_uk_K_r0_reg[41]/NET0131  ;
  assign n25620 = ~decrypt_pad & ~\u2_uk_K_r0_reg[5]/NET0131  ;
  assign n25621 = ~n25619 & ~n25620 ;
  assign n25622 = \u2_R0_reg[13]/NET0131  & ~n25621 ;
  assign n25623 = ~\u2_R0_reg[13]/NET0131  & n25621 ;
  assign n25624 = ~n25622 & ~n25623 ;
  assign n25632 = decrypt_pad & ~\u2_uk_K_r0_reg[47]/NET0131  ;
  assign n25633 = ~decrypt_pad & ~\u2_uk_K_r0_reg[11]/NET0131  ;
  assign n25634 = ~n25632 & ~n25633 ;
  assign n25635 = \u2_R0_reg[12]/NET0131  & ~n25634 ;
  assign n25636 = ~\u2_R0_reg[12]/NET0131  & n25634 ;
  assign n25637 = ~n25635 & ~n25636 ;
  assign n25665 = n25624 & ~n25637 ;
  assign n25666 = ~n25624 & n25637 ;
  assign n25667 = ~n25665 & ~n25666 ;
  assign n25639 = decrypt_pad & ~\u2_uk_K_r0_reg[18]/NET0131  ;
  assign n25640 = ~decrypt_pad & ~\u2_uk_K_r0_reg[39]/NET0131  ;
  assign n25641 = ~n25639 & ~n25640 ;
  assign n25642 = \u2_R0_reg[15]/NET0131  & ~n25641 ;
  assign n25643 = ~\u2_R0_reg[15]/NET0131  & n25641 ;
  assign n25644 = ~n25642 & ~n25643 ;
  assign n25646 = decrypt_pad & ~\u2_uk_K_r0_reg[10]/NET0131  ;
  assign n25647 = ~decrypt_pad & ~\u2_uk_K_r0_reg[6]/NET0131  ;
  assign n25648 = ~n25646 & ~n25647 ;
  assign n25649 = \u2_R0_reg[14]/NET0131  & ~n25648 ;
  assign n25650 = ~\u2_R0_reg[14]/NET0131  & n25648 ;
  assign n25651 = ~n25649 & ~n25650 ;
  assign n25668 = ~n25644 & ~n25651 ;
  assign n25669 = ~n25667 & n25668 ;
  assign n25656 = ~n25624 & n25644 ;
  assign n25625 = decrypt_pad & ~\u2_uk_K_r0_reg[6]/NET0131  ;
  assign n25626 = ~decrypt_pad & ~\u2_uk_K_r0_reg[27]/NET0131  ;
  assign n25627 = ~n25625 & ~n25626 ;
  assign n25628 = \u2_R0_reg[17]/NET0131  & ~n25627 ;
  assign n25629 = ~\u2_R0_reg[17]/NET0131  & n25627 ;
  assign n25630 = ~n25628 & ~n25629 ;
  assign n25657 = n25630 & ~n25637 ;
  assign n25658 = n25656 & n25657 ;
  assign n25653 = ~n25630 & n25637 ;
  assign n25654 = n25624 & n25644 ;
  assign n25655 = n25653 & n25654 ;
  assign n25670 = decrypt_pad & ~\u2_uk_K_r0_reg[26]/NET0131  ;
  assign n25671 = ~decrypt_pad & ~\u2_uk_K_r0_reg[47]/NET0131  ;
  assign n25672 = ~n25670 & ~n25671 ;
  assign n25673 = \u2_R0_reg[16]/NET0131  & ~n25672 ;
  assign n25674 = ~\u2_R0_reg[16]/NET0131  & n25672 ;
  assign n25675 = ~n25673 & ~n25674 ;
  assign n25676 = ~n25655 & n25675 ;
  assign n25677 = ~n25658 & n25676 ;
  assign n25678 = ~n25669 & n25677 ;
  assign n25631 = ~n25624 & ~n25630 ;
  assign n25638 = n25631 & ~n25637 ;
  assign n25645 = n25638 & ~n25644 ;
  assign n25652 = n25645 & n25651 ;
  assign n25659 = n25624 & ~n25651 ;
  assign n25660 = n25657 & n25659 ;
  assign n25661 = n25630 & n25637 ;
  assign n25662 = n25651 & n25661 ;
  assign n25663 = n25624 & n25662 ;
  assign n25664 = ~n25660 & ~n25663 ;
  assign n25679 = ~n25652 & n25664 ;
  assign n25680 = n25678 & n25679 ;
  assign n25688 = n25624 & n25661 ;
  assign n25689 = ~n25638 & n25644 ;
  assign n25690 = ~n25688 & n25689 ;
  assign n25692 = n25651 & n25653 ;
  assign n25691 = ~n25624 & n25630 ;
  assign n25693 = ~n25644 & ~n25691 ;
  assign n25694 = ~n25692 & n25693 ;
  assign n25695 = ~n25690 & ~n25694 ;
  assign n25681 = ~n25630 & n25665 ;
  assign n25682 = n25651 & n25681 ;
  assign n25683 = ~n25637 & ~n25651 ;
  assign n25684 = n25631 & n25683 ;
  assign n25685 = ~n25682 & ~n25684 ;
  assign n25696 = n25630 & ~n25651 ;
  assign n25697 = n25666 & n25696 ;
  assign n25686 = ~n25637 & n25651 ;
  assign n25687 = n25654 & n25686 ;
  assign n25698 = ~n25675 & ~n25687 ;
  assign n25699 = ~n25697 & n25698 ;
  assign n25700 = n25685 & n25699 ;
  assign n25701 = ~n25695 & n25700 ;
  assign n25702 = ~n25680 & ~n25701 ;
  assign n25703 = ~n25630 & n25683 ;
  assign n25704 = ~n25692 & ~n25703 ;
  assign n25705 = n25656 & ~n25704 ;
  assign n25706 = ~n25651 & n25653 ;
  assign n25707 = n25654 & n25706 ;
  assign n25708 = ~n25644 & n25696 ;
  assign n25709 = n25665 & n25708 ;
  assign n25710 = ~n25707 & ~n25709 ;
  assign n25711 = ~n25705 & n25710 ;
  assign n25712 = ~n25702 & n25711 ;
  assign n25713 = ~\u2_L0_reg[20]/NET0131  & ~n25712 ;
  assign n25714 = \u2_L0_reg[20]/NET0131  & n25712 ;
  assign n25715 = ~n25713 & ~n25714 ;
  assign n25739 = ~n25367 & n25383 ;
  assign n25740 = ~n25413 & ~n25739 ;
  assign n25741 = ~n25369 & ~n25411 ;
  assign n25742 = ~n25382 & ~n25741 ;
  assign n25743 = n25740 & ~n25742 ;
  assign n25744 = n25347 & ~n25743 ;
  assign n25716 = n25353 & n25405 ;
  assign n25736 = ~n25353 & n25417 ;
  assign n25737 = ~n25716 & ~n25736 ;
  assign n25738 = ~n25347 & ~n25737 ;
  assign n25745 = n25353 & n25390 ;
  assign n25746 = ~n25738 & ~n25745 ;
  assign n25747 = ~n25744 & n25746 ;
  assign n25748 = ~n25341 & ~n25747 ;
  assign n25717 = ~n25353 & ~n25360 ;
  assign n25718 = n25367 & n25717 ;
  assign n25719 = ~n25420 & ~n25718 ;
  assign n25720 = ~n25716 & n25719 ;
  assign n25721 = n25347 & ~n25720 ;
  assign n25722 = ~n25360 & ~n25382 ;
  assign n25726 = n25353 & n25722 ;
  assign n25727 = n25382 & n25717 ;
  assign n25728 = ~n25726 & ~n25727 ;
  assign n25729 = ~n25367 & ~n25728 ;
  assign n25723 = ~n25370 & n25722 ;
  assign n25724 = ~n25401 & ~n25723 ;
  assign n25725 = ~n25347 & ~n25724 ;
  assign n25730 = ~n25385 & ~n25388 ;
  assign n25731 = ~n25725 & n25730 ;
  assign n25732 = ~n25729 & n25731 ;
  assign n25733 = ~n25721 & n25732 ;
  assign n25734 = n25341 & ~n25733 ;
  assign n25735 = n25354 & n25419 ;
  assign n25749 = ~n25412 & ~n25735 ;
  assign n25750 = ~n25734 & n25749 ;
  assign n25751 = ~n25748 & n25750 ;
  assign n25752 = \u2_L0_reg[29]/NET0131  & ~n25751 ;
  assign n25753 = ~\u2_L0_reg[29]/NET0131  & n25751 ;
  assign n25754 = ~n25752 & ~n25753 ;
  assign n25759 = ~n25405 & ~n25727 ;
  assign n25760 = ~n25388 & n25759 ;
  assign n25761 = n25347 & ~n25760 ;
  assign n25755 = n25367 & n25722 ;
  assign n25756 = ~n25745 & ~n25755 ;
  assign n25757 = ~n25347 & ~n25756 ;
  assign n25758 = n25384 & n25386 ;
  assign n25762 = ~n25412 & ~n25758 ;
  assign n25763 = ~n25757 & n25762 ;
  assign n25764 = ~n25761 & n25763 ;
  assign n25765 = ~n25341 & ~n25764 ;
  assign n25773 = ~n25392 & ~n25717 ;
  assign n25774 = ~n25347 & ~n25773 ;
  assign n25775 = n25353 & n25419 ;
  assign n25776 = n25354 & n25386 ;
  assign n25777 = ~n25775 & ~n25776 ;
  assign n25778 = ~n25402 & n25777 ;
  assign n25779 = ~n25774 & n25778 ;
  assign n25780 = n25341 & ~n25779 ;
  assign n25766 = ~n25409 & ~n25420 ;
  assign n25767 = ~n25405 & n25766 ;
  assign n25768 = n25375 & ~n25767 ;
  assign n25769 = n25353 & n25740 ;
  assign n25770 = ~n25353 & ~n25722 ;
  assign n25771 = ~n25347 & ~n25770 ;
  assign n25772 = ~n25769 & n25771 ;
  assign n25781 = ~n25768 & ~n25772 ;
  assign n25782 = ~n25780 & n25781 ;
  assign n25783 = ~n25765 & n25782 ;
  assign n25784 = ~\u2_L0_reg[4]/NET0131  & ~n25783 ;
  assign n25785 = \u2_L0_reg[4]/NET0131  & n25783 ;
  assign n25786 = ~n25784 & ~n25785 ;
  assign n25787 = decrypt_pad & ~\u2_uk_K_r0_reg[52]/P0001  ;
  assign n25788 = ~decrypt_pad & ~\u2_uk_K_r0_reg[14]/NET0131  ;
  assign n25789 = ~n25787 & ~n25788 ;
  assign n25790 = \u2_R0_reg[32]/NET0131  & ~n25789 ;
  assign n25791 = ~\u2_R0_reg[32]/NET0131  & n25789 ;
  assign n25792 = ~n25790 & ~n25791 ;
  assign n25831 = decrypt_pad & ~\u2_uk_K_r0_reg[42]/NET0131  ;
  assign n25832 = ~decrypt_pad & ~\u2_uk_K_r0_reg[8]/NET0131  ;
  assign n25833 = ~n25831 & ~n25832 ;
  assign n25834 = \u2_R0_reg[31]/P0001  & ~n25833 ;
  assign n25835 = ~\u2_R0_reg[31]/P0001  & n25833 ;
  assign n25836 = ~n25834 & ~n25835 ;
  assign n25806 = decrypt_pad & ~\u2_uk_K_r0_reg[2]/NET0131  ;
  assign n25807 = ~decrypt_pad & ~\u2_uk_K_r0_reg[23]/NET0131  ;
  assign n25808 = ~n25806 & ~n25807 ;
  assign n25809 = \u2_R0_reg[28]/NET0131  & ~n25808 ;
  assign n25810 = ~\u2_R0_reg[28]/NET0131  & n25808 ;
  assign n25811 = ~n25809 & ~n25810 ;
  assign n25793 = decrypt_pad & ~\u2_uk_K_r0_reg[29]/NET0131  ;
  assign n25794 = ~decrypt_pad & ~\u2_uk_K_r0_reg[50]/NET0131  ;
  assign n25795 = ~n25793 & ~n25794 ;
  assign n25796 = \u2_R0_reg[29]/NET0131  & ~n25795 ;
  assign n25797 = ~\u2_R0_reg[29]/NET0131  & n25795 ;
  assign n25798 = ~n25796 & ~n25797 ;
  assign n25799 = decrypt_pad & ~\u2_uk_K_r0_reg[14]/NET0131  ;
  assign n25800 = ~decrypt_pad & ~\u2_uk_K_r0_reg[35]/NET0131  ;
  assign n25801 = ~n25799 & ~n25800 ;
  assign n25802 = \u2_R0_reg[1]/NET0131  & ~n25801 ;
  assign n25803 = ~\u2_R0_reg[1]/NET0131  & n25801 ;
  assign n25804 = ~n25802 & ~n25803 ;
  assign n25839 = ~n25798 & n25804 ;
  assign n25840 = ~n25811 & n25839 ;
  assign n25812 = decrypt_pad & ~\u2_uk_K_r0_reg[30]/NET0131  ;
  assign n25813 = ~decrypt_pad & ~\u2_uk_K_r0_reg[51]/NET0131  ;
  assign n25814 = ~n25812 & ~n25813 ;
  assign n25815 = \u2_R0_reg[30]/NET0131  & ~n25814 ;
  assign n25816 = ~\u2_R0_reg[30]/NET0131  & n25814 ;
  assign n25817 = ~n25815 & ~n25816 ;
  assign n25860 = ~n25798 & ~n25804 ;
  assign n25861 = n25817 & n25860 ;
  assign n25862 = n25811 & n25861 ;
  assign n25863 = ~n25840 & ~n25862 ;
  assign n25864 = n25836 & ~n25863 ;
  assign n25805 = n25798 & n25804 ;
  assign n25846 = n25811 & ~n25817 ;
  assign n25818 = ~n25811 & n25817 ;
  assign n25854 = ~n25804 & n25818 ;
  assign n25855 = ~n25846 & ~n25854 ;
  assign n25856 = ~n25805 & n25855 ;
  assign n25857 = ~n25836 & ~n25856 ;
  assign n25827 = n25798 & n25811 ;
  assign n25828 = ~n25817 & n25827 ;
  assign n25829 = ~n25804 & n25828 ;
  assign n25858 = n25817 & n25827 ;
  assign n25859 = n25804 & n25858 ;
  assign n25865 = ~n25829 & ~n25859 ;
  assign n25866 = ~n25857 & n25865 ;
  assign n25867 = ~n25864 & n25866 ;
  assign n25868 = ~n25792 & ~n25867 ;
  assign n25842 = n25798 & ~n25817 ;
  assign n25843 = ~n25804 & n25811 ;
  assign n25844 = ~n25842 & ~n25843 ;
  assign n25845 = ~n25792 & ~n25844 ;
  assign n25847 = n25798 & ~n25804 ;
  assign n25848 = ~n25846 & ~n25847 ;
  assign n25849 = ~n25829 & ~n25848 ;
  assign n25850 = ~n25845 & n25849 ;
  assign n25823 = ~n25811 & ~n25817 ;
  assign n25824 = ~n25798 & n25823 ;
  assign n25838 = ~n25804 & n25824 ;
  assign n25841 = n25817 & n25840 ;
  assign n25851 = ~n25838 & ~n25841 ;
  assign n25852 = ~n25850 & n25851 ;
  assign n25853 = n25836 & ~n25852 ;
  assign n25819 = n25805 & n25818 ;
  assign n25820 = n25792 & n25819 ;
  assign n25821 = ~n25798 & n25811 ;
  assign n25822 = n25817 & n25821 ;
  assign n25825 = ~n25822 & ~n25824 ;
  assign n25826 = n25792 & ~n25825 ;
  assign n25830 = ~n25826 & ~n25829 ;
  assign n25837 = ~n25830 & ~n25836 ;
  assign n25869 = ~n25820 & ~n25837 ;
  assign n25870 = ~n25853 & n25869 ;
  assign n25871 = ~n25868 & n25870 ;
  assign n25872 = \u2_L0_reg[5]/NET0131  & ~n25871 ;
  assign n25873 = ~\u2_L0_reg[5]/NET0131  & n25871 ;
  assign n25874 = ~n25872 & ~n25873 ;
  assign n25886 = n25656 & ~n25696 ;
  assign n25887 = ~n25659 & ~n25708 ;
  assign n25888 = ~n25886 & n25887 ;
  assign n25889 = n25637 & ~n25888 ;
  assign n25890 = ~n25637 & n25696 ;
  assign n25891 = n25644 & n25890 ;
  assign n25892 = ~n25645 & ~n25891 ;
  assign n25893 = n25685 & n25892 ;
  assign n25894 = ~n25889 & n25893 ;
  assign n25895 = ~n25675 & ~n25894 ;
  assign n25880 = n25653 & ~n25659 ;
  assign n25881 = ~n25660 & ~n25880 ;
  assign n25882 = ~n25644 & ~n25881 ;
  assign n25875 = ~n25624 & n25651 ;
  assign n25876 = n25657 & n25875 ;
  assign n25877 = ~n25663 & ~n25876 ;
  assign n25878 = ~n25681 & ~n25697 ;
  assign n25879 = n25644 & ~n25878 ;
  assign n25883 = n25877 & ~n25879 ;
  assign n25884 = ~n25882 & n25883 ;
  assign n25885 = n25675 & ~n25884 ;
  assign n25896 = ~n25684 & n25877 ;
  assign n25897 = ~n25644 & ~n25896 ;
  assign n25898 = ~n25687 & ~n25707 ;
  assign n25899 = ~n25897 & n25898 ;
  assign n25900 = ~n25885 & n25899 ;
  assign n25901 = ~n25895 & n25900 ;
  assign n25902 = ~\u2_L0_reg[10]/NET0131  & ~n25901 ;
  assign n25903 = \u2_L0_reg[10]/NET0131  & n25901 ;
  assign n25904 = ~n25902 & ~n25903 ;
  assign n25911 = n25445 & n25452 ;
  assign n25912 = ~n25510 & ~n25911 ;
  assign n25913 = n25484 & ~n25912 ;
  assign n25905 = n25466 & n25492 ;
  assign n25914 = n25474 & ~n25506 ;
  assign n25915 = ~n25905 & n25914 ;
  assign n25907 = n25452 & ~n25458 ;
  assign n25908 = ~n25459 & ~n25907 ;
  assign n25906 = ~n25452 & n25484 ;
  assign n25909 = n25446 & ~n25906 ;
  assign n25910 = ~n25908 & n25909 ;
  assign n25916 = ~n25463 & ~n25910 ;
  assign n25917 = n25915 & n25916 ;
  assign n25918 = ~n25913 & n25917 ;
  assign n25921 = n25439 & n25445 ;
  assign n25922 = ~n25486 & ~n25921 ;
  assign n25923 = n25459 & ~n25922 ;
  assign n25919 = ~n25439 & n25907 ;
  assign n25920 = ~n25445 & n25919 ;
  assign n25930 = ~n25474 & ~n25920 ;
  assign n25931 = ~n25923 & n25930 ;
  assign n25924 = ~n25465 & ~n25466 ;
  assign n25925 = ~n25493 & n25924 ;
  assign n25926 = ~n25484 & ~n25925 ;
  assign n25927 = ~n25505 & ~n25921 ;
  assign n25928 = ~n25466 & n25908 ;
  assign n25929 = n25927 & n25928 ;
  assign n25932 = ~n25926 & ~n25929 ;
  assign n25933 = n25931 & n25932 ;
  assign n25934 = ~n25918 & ~n25933 ;
  assign n25935 = \u2_L0_reg[12]/NET0131  & n25934 ;
  assign n25936 = ~\u2_L0_reg[12]/NET0131  & ~n25934 ;
  assign n25937 = ~n25935 & ~n25936 ;
  assign n25938 = decrypt_pad & ~\u2_uk_K_r0_reg[9]/NET0131  ;
  assign n25939 = ~decrypt_pad & ~\u2_uk_K_r0_reg[30]/NET0131  ;
  assign n25940 = ~n25938 & ~n25939 ;
  assign n25941 = \u2_R0_reg[20]/NET0131  & ~n25940 ;
  assign n25942 = ~\u2_R0_reg[20]/NET0131  & n25940 ;
  assign n25943 = ~n25941 & ~n25942 ;
  assign n25944 = decrypt_pad & ~\u2_uk_K_r0_reg[22]/NET0131  ;
  assign n25945 = ~decrypt_pad & ~\u2_uk_K_r0_reg[43]/NET0131  ;
  assign n25946 = ~n25944 & ~n25945 ;
  assign n25947 = \u2_R0_reg[16]/NET0131  & ~n25946 ;
  assign n25948 = ~\u2_R0_reg[16]/NET0131  & n25946 ;
  assign n25949 = ~n25947 & ~n25948 ;
  assign n25950 = decrypt_pad & ~\u2_uk_K_r0_reg[44]/NET0131  ;
  assign n25951 = ~decrypt_pad & ~\u2_uk_K_r0_reg[38]/NET0131  ;
  assign n25952 = ~n25950 & ~n25951 ;
  assign n25953 = \u2_R0_reg[17]/NET0131  & ~n25952 ;
  assign n25954 = ~\u2_R0_reg[17]/NET0131  & n25952 ;
  assign n25955 = ~n25953 & ~n25954 ;
  assign n25956 = n25949 & ~n25955 ;
  assign n25963 = decrypt_pad & ~\u2_uk_K_r0_reg[7]/NET0131  ;
  assign n25964 = ~decrypt_pad & ~\u2_uk_K_r0_reg[28]/NET0131  ;
  assign n25965 = ~n25963 & ~n25964 ;
  assign n25966 = \u2_R0_reg[18]/NET0131  & ~n25965 ;
  assign n25967 = ~\u2_R0_reg[18]/NET0131  & n25965 ;
  assign n25968 = ~n25966 & ~n25967 ;
  assign n25981 = n25955 & ~n25968 ;
  assign n26004 = ~n25956 & ~n25981 ;
  assign n25957 = decrypt_pad & ~\u2_uk_K_r0_reg[38]/NET0131  ;
  assign n25958 = ~decrypt_pad & ~\u2_uk_K_r0_reg[0]/NET0131  ;
  assign n25959 = ~n25957 & ~n25958 ;
  assign n25960 = \u2_R0_reg[21]/NET0131  & ~n25959 ;
  assign n25961 = ~\u2_R0_reg[21]/NET0131  & n25959 ;
  assign n25962 = ~n25960 & ~n25961 ;
  assign n25969 = n25962 & n25968 ;
  assign n25991 = ~n25949 & ~n25962 ;
  assign n26005 = ~n25969 & ~n25991 ;
  assign n26006 = ~n26004 & ~n26005 ;
  assign n26007 = ~n25949 & ~n25955 ;
  assign n25970 = ~n25962 & ~n25968 ;
  assign n26008 = ~n25955 & n25970 ;
  assign n26009 = ~n26007 & ~n26008 ;
  assign n26010 = ~n25991 & ~n26009 ;
  assign n25984 = n25949 & n25962 ;
  assign n25985 = ~n25968 & n25984 ;
  assign n26013 = n25955 & n25985 ;
  assign n25973 = decrypt_pad & ~\u2_uk_K_r0_reg[49]/NET0131  ;
  assign n25974 = ~decrypt_pad & ~\u2_uk_K_r0_reg[15]/NET0131  ;
  assign n25975 = ~n25973 & ~n25974 ;
  assign n25976 = \u2_R0_reg[19]/NET0131  & ~n25975 ;
  assign n25977 = ~\u2_R0_reg[19]/NET0131  & n25975 ;
  assign n25978 = ~n25976 & ~n25977 ;
  assign n26011 = n25955 & ~n25962 ;
  assign n26012 = n25968 & n26011 ;
  assign n26014 = ~n25978 & ~n26012 ;
  assign n26015 = ~n26013 & n26014 ;
  assign n26016 = ~n26010 & n26015 ;
  assign n25992 = ~n25955 & n25991 ;
  assign n26019 = n25978 & ~n25992 ;
  assign n26017 = n25949 & n25969 ;
  assign n26018 = ~n25949 & n25981 ;
  assign n26020 = ~n26017 & ~n26018 ;
  assign n26021 = n26019 & n26020 ;
  assign n26022 = ~n26016 & ~n26021 ;
  assign n26023 = ~n26006 & ~n26022 ;
  assign n26024 = ~n25943 & ~n26023 ;
  assign n25979 = n25949 & ~n25962 ;
  assign n25980 = n25955 & n25979 ;
  assign n25982 = ~n25949 & n25962 ;
  assign n25983 = ~n25981 & n25982 ;
  assign n25986 = ~n25980 & ~n25983 ;
  assign n25987 = ~n25985 & n25986 ;
  assign n25988 = n25978 & ~n25987 ;
  assign n25989 = ~n25968 & ~n25978 ;
  assign n25990 = n25955 & n25982 ;
  assign n25993 = ~n25990 & ~n25992 ;
  assign n25994 = n25989 & ~n25993 ;
  assign n25995 = n25955 & n25984 ;
  assign n25996 = n25968 & ~n25978 ;
  assign n25997 = n25995 & n25996 ;
  assign n25971 = ~n25969 & ~n25970 ;
  assign n25972 = n25956 & n25971 ;
  assign n25998 = n25979 & n25981 ;
  assign n25999 = ~n25972 & ~n25998 ;
  assign n26000 = ~n25997 & n25999 ;
  assign n26001 = ~n25994 & n26000 ;
  assign n26002 = ~n25988 & n26001 ;
  assign n26003 = n25943 & ~n26002 ;
  assign n26025 = n25968 & n25992 ;
  assign n26026 = ~n25998 & ~n26025 ;
  assign n26027 = n25978 & ~n26026 ;
  assign n26028 = ~n25955 & n25968 ;
  assign n26029 = n25982 & n26028 ;
  assign n26030 = ~n25949 & n25968 ;
  assign n26031 = n26011 & n26030 ;
  assign n26032 = ~n26029 & ~n26031 ;
  assign n26033 = ~n25978 & ~n26032 ;
  assign n26034 = ~n26027 & ~n26033 ;
  assign n26035 = ~n26003 & n26034 ;
  assign n26036 = ~n26024 & n26035 ;
  assign n26037 = ~\u2_L0_reg[14]/NET0131  & ~n26036 ;
  assign n26038 = \u2_L0_reg[14]/NET0131  & n26036 ;
  assign n26039 = ~n26037 & ~n26038 ;
  assign n26056 = ~n25552 & ~n25578 ;
  assign n26057 = n25576 & n25578 ;
  assign n26058 = ~n26056 & ~n26057 ;
  assign n26059 = n25559 & ~n26058 ;
  assign n26060 = ~n25559 & ~n25601 ;
  assign n26061 = ~n26056 & n26060 ;
  assign n26055 = n25552 & n25607 ;
  assign n26062 = ~n25604 & ~n26055 ;
  assign n26063 = ~n26061 & n26062 ;
  assign n26064 = ~n26059 & n26063 ;
  assign n26065 = n25526 & ~n26064 ;
  assign n26040 = ~n25532 & n25569 ;
  assign n26041 = ~n25586 & ~n26040 ;
  assign n26042 = n25538 & ~n26041 ;
  assign n26043 = n25538 & n25576 ;
  assign n26044 = ~n25562 & ~n26043 ;
  assign n26045 = ~n25526 & ~n26044 ;
  assign n26046 = ~n26042 & ~n26045 ;
  assign n26047 = n25559 & ~n26046 ;
  assign n26049 = n25538 & ~n25573 ;
  assign n26048 = ~n25572 & ~n25576 ;
  assign n26050 = ~n25559 & ~n26048 ;
  assign n26051 = ~n26049 & n26050 ;
  assign n26052 = ~n25553 & ~n25609 ;
  assign n26053 = ~n26051 & n26052 ;
  assign n26054 = ~n25526 & ~n26053 ;
  assign n26066 = ~n26047 & ~n26054 ;
  assign n26067 = ~n26065 & n26066 ;
  assign n26068 = ~\u2_L0_reg[17]/NET0131  & ~n26067 ;
  assign n26069 = \u2_L0_reg[17]/NET0131  & n26067 ;
  assign n26070 = ~n26068 & ~n26069 ;
  assign n26073 = n25360 & ~n25370 ;
  assign n26074 = ~n25755 & ~n26073 ;
  assign n26075 = n25347 & ~n26074 ;
  assign n26072 = ~n25347 & ~n25766 ;
  assign n26071 = n25353 & n25413 ;
  assign n26076 = ~n25341 & ~n26071 ;
  assign n26077 = ~n26072 & n26076 ;
  assign n26078 = ~n26075 & n26077 ;
  assign n26081 = n25353 & n25420 ;
  assign n26082 = ~n25347 & n25374 ;
  assign n26083 = n25341 & ~n25392 ;
  assign n26084 = ~n26082 & n26083 ;
  assign n26085 = ~n26081 & n26084 ;
  assign n26079 = ~n25371 & ~n25390 ;
  assign n26080 = n25347 & ~n26079 ;
  assign n26086 = ~n25729 & ~n26080 ;
  assign n26087 = n26085 & n26086 ;
  assign n26088 = ~n26078 & ~n26087 ;
  assign n26089 = n25384 & n25387 ;
  assign n26090 = ~n25408 & ~n26089 ;
  assign n26091 = ~n26088 & n26090 ;
  assign n26092 = ~\u2_L0_reg[19]/NET0131  & ~n26091 ;
  assign n26093 = \u2_L0_reg[19]/NET0131  & n26091 ;
  assign n26094 = ~n26092 & ~n26093 ;
  assign n26111 = n25637 & n25691 ;
  assign n26112 = ~n25644 & ~n25706 ;
  assign n26113 = ~n26111 & n26112 ;
  assign n26114 = n25653 & n25875 ;
  assign n26115 = n25644 & ~n25703 ;
  assign n26116 = ~n26114 & n26115 ;
  assign n26117 = ~n26113 & ~n26116 ;
  assign n26118 = n25624 & n25706 ;
  assign n26119 = n25664 & ~n26118 ;
  assign n26120 = ~n26117 & n26119 ;
  assign n26121 = ~n25675 & ~n26120 ;
  assign n26104 = n25651 & ~n25657 ;
  assign n26105 = n25624 & ~n25644 ;
  assign n26106 = ~n25653 & n26105 ;
  assign n26107 = ~n26104 & n26106 ;
  assign n26097 = n25624 & n25692 ;
  assign n26103 = ~n25637 & n25875 ;
  assign n26108 = ~n26097 & ~n26103 ;
  assign n26109 = ~n26107 & n26108 ;
  assign n26110 = n25675 & ~n26109 ;
  assign n26095 = ~n25682 & n25877 ;
  assign n26096 = n25644 & ~n26095 ;
  assign n26099 = ~n25651 & n25666 ;
  assign n26100 = ~n25691 & ~n26099 ;
  assign n26101 = n25644 & n25675 ;
  assign n26102 = ~n26100 & n26101 ;
  assign n26098 = ~n25644 & n26097 ;
  assign n26122 = ~n25652 & ~n26098 ;
  assign n26123 = ~n26102 & n26122 ;
  assign n26124 = ~n26096 & n26123 ;
  assign n26125 = ~n26110 & n26124 ;
  assign n26126 = ~n26121 & n26125 ;
  assign n26127 = ~\u2_L0_reg[1]/NET0131  & ~n26126 ;
  assign n26128 = \u2_L0_reg[1]/NET0131  & n26126 ;
  assign n26129 = ~n26127 & ~n26128 ;
  assign n26131 = n25798 & ~n25855 ;
  assign n26132 = ~n25811 & n25860 ;
  assign n26133 = n25836 & n26132 ;
  assign n26130 = n25804 & n25822 ;
  assign n26134 = n25817 & ~n25836 ;
  assign n26135 = n25839 & n26134 ;
  assign n26136 = n25792 & ~n26135 ;
  assign n26137 = ~n26130 & n26136 ;
  assign n26138 = ~n26133 & n26137 ;
  assign n26139 = ~n26131 & n26138 ;
  assign n26141 = ~n25817 & n25847 ;
  assign n26142 = ~n25827 & ~n26141 ;
  assign n26143 = ~n25840 & n26142 ;
  assign n26144 = n25836 & ~n26143 ;
  assign n26140 = n25846 & n25860 ;
  assign n26145 = ~n25792 & ~n26140 ;
  assign n26146 = ~n26144 & n26145 ;
  assign n26147 = ~n26139 & ~n26146 ;
  assign n26149 = n25823 & ~n25839 ;
  assign n26150 = ~n25847 & n26149 ;
  assign n26151 = n25792 & ~n25817 ;
  assign n26152 = n25821 & ~n26151 ;
  assign n26148 = n25818 & n25847 ;
  assign n26153 = ~n25836 & ~n26148 ;
  assign n26154 = ~n26152 & n26153 ;
  assign n26155 = ~n26150 & n26154 ;
  assign n26156 = ~n25817 & n25839 ;
  assign n26157 = ~n25811 & n26156 ;
  assign n26158 = ~n25819 & n25836 ;
  assign n26159 = ~n26157 & n26158 ;
  assign n26160 = ~n26155 & ~n26159 ;
  assign n26161 = ~n26147 & ~n26160 ;
  assign n26162 = ~\u2_L0_reg[15]/NET0131  & ~n26161 ;
  assign n26163 = \u2_L0_reg[15]/NET0131  & n26161 ;
  assign n26164 = ~n26162 & ~n26163 ;
  assign n26168 = ~n25804 & n25846 ;
  assign n26169 = ~n25836 & ~n26168 ;
  assign n26170 = ~n26130 & n26169 ;
  assign n26172 = n25836 & ~n25858 ;
  assign n26171 = n25805 & ~n25811 ;
  assign n26173 = ~n26156 & ~n26171 ;
  assign n26174 = n26172 & n26173 ;
  assign n26175 = ~n26170 & ~n26174 ;
  assign n26176 = ~n25804 & n25827 ;
  assign n26177 = ~n26132 & ~n26176 ;
  assign n26178 = n25817 & ~n26177 ;
  assign n26179 = n25792 & ~n26157 ;
  assign n26180 = ~n26178 & n26179 ;
  assign n26181 = ~n26175 & n26180 ;
  assign n26166 = n25804 & ~n25836 ;
  assign n26186 = ~n25805 & ~n26166 ;
  assign n26187 = n25846 & ~n26186 ;
  assign n26182 = ~n25798 & ~n26166 ;
  assign n26183 = n25818 & ~n26182 ;
  assign n26192 = ~n25862 & ~n26183 ;
  assign n26193 = ~n26187 & n26192 ;
  assign n26184 = ~n25822 & ~n26176 ;
  assign n26185 = n25836 & ~n26184 ;
  assign n26188 = ~n25811 & ~n25836 ;
  assign n26189 = n25847 & n26188 ;
  assign n26190 = ~n25792 & ~n26189 ;
  assign n26191 = ~n25838 & n26190 ;
  assign n26194 = ~n26185 & n26191 ;
  assign n26195 = n26193 & n26194 ;
  assign n26196 = ~n26181 & ~n26195 ;
  assign n26165 = n25824 & n25836 ;
  assign n26167 = n25828 & n26166 ;
  assign n26197 = ~n26165 & ~n26167 ;
  assign n26198 = ~n26196 & n26197 ;
  assign n26199 = ~\u2_L0_reg[21]/NET0131  & ~n26198 ;
  assign n26200 = \u2_L0_reg[21]/NET0131  & n26198 ;
  assign n26201 = ~n26199 & ~n26200 ;
  assign n26202 = n25955 & ~n26030 ;
  assign n26203 = n25971 & n26202 ;
  assign n26204 = ~n25955 & n25984 ;
  assign n26205 = ~n25978 & ~n26204 ;
  assign n26206 = ~n26018 & n26205 ;
  assign n26207 = n25978 & ~n25995 ;
  assign n26208 = ~n25962 & n26030 ;
  assign n26209 = n26009 & ~n26208 ;
  assign n26210 = n26207 & n26209 ;
  assign n26211 = ~n26206 & ~n26210 ;
  assign n26212 = ~n26203 & ~n26211 ;
  assign n26213 = n25943 & ~n26212 ;
  assign n26219 = ~n25978 & ~n26007 ;
  assign n26218 = n25978 & ~n26011 ;
  assign n26220 = ~n25968 & ~n26218 ;
  assign n26221 = ~n26219 & n26220 ;
  assign n26214 = n25968 & n25990 ;
  assign n26215 = ~n25955 & ~n25979 ;
  assign n26216 = ~n25978 & ~n26202 ;
  assign n26217 = ~n26215 & n26216 ;
  assign n26222 = ~n26214 & ~n26217 ;
  assign n26223 = ~n26221 & n26222 ;
  assign n26224 = ~n25943 & ~n26223 ;
  assign n26225 = n25971 & n26007 ;
  assign n26226 = n25968 & n25980 ;
  assign n26227 = ~n26225 & ~n26226 ;
  assign n26228 = n25978 & ~n26227 ;
  assign n26229 = n25956 & n25996 ;
  assign n26230 = ~n26013 & ~n26229 ;
  assign n26231 = ~n26228 & n26230 ;
  assign n26232 = ~n26224 & n26231 ;
  assign n26233 = ~n26213 & n26232 ;
  assign n26234 = ~\u2_L0_reg[25]/NET0131  & ~n26233 ;
  assign n26235 = \u2_L0_reg[25]/NET0131  & n26233 ;
  assign n26236 = ~n26234 & ~n26235 ;
  assign n26237 = ~n25630 & ~n25667 ;
  assign n26238 = ~n25688 & ~n26237 ;
  assign n26239 = ~n25651 & ~n26238 ;
  assign n26240 = ~n25631 & ~n26103 ;
  assign n26241 = ~n25675 & ~n26240 ;
  assign n26242 = ~n25644 & ~n26241 ;
  assign n26243 = ~n26239 & n26242 ;
  assign n26244 = n25644 & ~n25660 ;
  assign n26245 = ~n25697 & n26244 ;
  assign n26246 = ~n26243 & ~n26245 ;
  assign n26248 = ~n25624 & n25890 ;
  assign n26249 = ~n25644 & ~n25662 ;
  assign n26250 = ~n26248 & n26249 ;
  assign n26251 = ~n25689 & ~n26250 ;
  assign n26247 = n25624 & ~n25704 ;
  assign n26252 = ~n25624 & ~n25644 ;
  assign n26253 = n25651 & n25657 ;
  assign n26254 = ~n26252 & n26253 ;
  assign n26255 = n25675 & ~n26254 ;
  assign n26256 = ~n26247 & n26255 ;
  assign n26257 = ~n26251 & n26256 ;
  assign n26258 = n25654 & n26104 ;
  assign n26259 = ~n25655 & ~n25675 ;
  assign n26260 = ~n25660 & ~n26099 ;
  assign n26261 = n26259 & n26260 ;
  assign n26262 = ~n26258 & n26261 ;
  assign n26263 = ~n26257 & ~n26262 ;
  assign n26264 = ~n26246 & ~n26263 ;
  assign n26265 = ~\u2_L0_reg[26]/NET0131  & ~n26264 ;
  assign n26266 = \u2_L0_reg[26]/NET0131  & n26264 ;
  assign n26267 = ~n26265 & ~n26266 ;
  assign n26305 = decrypt_pad & ~\u2_uk_K_r0_reg[25]/P0001  ;
  assign n26306 = ~decrypt_pad & ~\u2_uk_K_r0_reg[46]/NET0131  ;
  assign n26307 = ~n26305 & ~n26306 ;
  assign n26308 = \u2_R0_reg[8]/NET0131  & ~n26307 ;
  assign n26309 = ~\u2_R0_reg[8]/NET0131  & n26307 ;
  assign n26310 = ~n26308 & ~n26309 ;
  assign n26298 = decrypt_pad & ~\u2_uk_K_r0_reg[34]/NET0131  ;
  assign n26299 = ~decrypt_pad & ~\u2_uk_K_r0_reg[55]/NET0131  ;
  assign n26300 = ~n26298 & ~n26299 ;
  assign n26301 = \u2_R0_reg[7]/NET0131  & ~n26300 ;
  assign n26302 = ~\u2_R0_reg[7]/NET0131  & n26300 ;
  assign n26303 = ~n26301 & ~n26302 ;
  assign n26274 = decrypt_pad & ~\u2_uk_K_r0_reg[40]/NET0131  ;
  assign n26275 = ~decrypt_pad & ~\u2_uk_K_r0_reg[4]/NET0131  ;
  assign n26276 = ~n26274 & ~n26275 ;
  assign n26277 = \u2_R0_reg[6]/NET0131  & ~n26276 ;
  assign n26278 = ~\u2_R0_reg[6]/NET0131  & n26276 ;
  assign n26279 = ~n26277 & ~n26278 ;
  assign n26281 = decrypt_pad & ~\u2_uk_K_r0_reg[13]/NET0131  ;
  assign n26282 = ~decrypt_pad & ~\u2_uk_K_r0_reg[34]/NET0131  ;
  assign n26283 = ~n26281 & ~n26282 ;
  assign n26284 = \u2_R0_reg[4]/NET0131  & ~n26283 ;
  assign n26285 = ~\u2_R0_reg[4]/NET0131  & n26283 ;
  assign n26286 = ~n26284 & ~n26285 ;
  assign n26288 = decrypt_pad & ~\u2_uk_K_r0_reg[5]/NET0131  ;
  assign n26289 = ~decrypt_pad & ~\u2_uk_K_r0_reg[26]/NET0131  ;
  assign n26290 = ~n26288 & ~n26289 ;
  assign n26291 = \u2_R0_reg[9]/NET0131  & ~n26290 ;
  assign n26292 = ~\u2_R0_reg[9]/NET0131  & n26290 ;
  assign n26293 = ~n26291 & ~n26292 ;
  assign n26315 = n26286 & ~n26293 ;
  assign n26340 = ~n26279 & n26315 ;
  assign n26268 = decrypt_pad & ~\u2_uk_K_r0_reg[17]/NET0131  ;
  assign n26269 = ~decrypt_pad & ~\u2_uk_K_r0_reg[13]/NET0131  ;
  assign n26270 = ~n26268 & ~n26269 ;
  assign n26271 = \u2_R0_reg[5]/NET0131  & ~n26270 ;
  assign n26272 = ~\u2_R0_reg[5]/NET0131  & n26270 ;
  assign n26273 = ~n26271 & ~n26272 ;
  assign n26338 = n26273 & n26286 ;
  assign n26311 = ~n26286 & n26293 ;
  assign n26339 = ~n26273 & n26311 ;
  assign n26341 = ~n26338 & ~n26339 ;
  assign n26342 = ~n26340 & n26341 ;
  assign n26343 = ~n26303 & ~n26342 ;
  assign n26322 = ~n26286 & ~n26293 ;
  assign n26323 = ~n26279 & n26322 ;
  assign n26324 = n26273 & n26311 ;
  assign n26325 = ~n26323 & ~n26324 ;
  assign n26344 = n26303 & ~n26325 ;
  assign n26294 = n26273 & ~n26293 ;
  assign n26295 = n26286 & n26294 ;
  assign n26296 = n26279 & n26295 ;
  assign n26335 = ~n26273 & ~n26315 ;
  assign n26336 = n26279 & ~n26311 ;
  assign n26337 = n26335 & n26336 ;
  assign n26345 = ~n26296 & ~n26337 ;
  assign n26346 = ~n26344 & n26345 ;
  assign n26347 = ~n26343 & n26346 ;
  assign n26348 = ~n26310 & ~n26347 ;
  assign n26280 = ~n26273 & n26279 ;
  assign n26287 = n26280 & ~n26286 ;
  assign n26297 = ~n26287 & ~n26296 ;
  assign n26304 = ~n26297 & ~n26303 ;
  assign n26313 = ~n26286 & n26294 ;
  assign n26314 = n26279 & n26313 ;
  assign n26316 = ~n26273 & n26315 ;
  assign n26317 = n26286 & n26293 ;
  assign n26318 = n26273 & n26317 ;
  assign n26319 = ~n26316 & ~n26318 ;
  assign n26320 = ~n26314 & n26319 ;
  assign n26321 = n26303 & ~n26320 ;
  assign n26326 = ~n26303 & ~n26325 ;
  assign n26312 = n26280 & n26311 ;
  assign n26327 = ~n26273 & n26293 ;
  assign n26328 = ~n26303 & ~n26327 ;
  assign n26329 = ~n26279 & n26286 ;
  assign n26330 = ~n26328 & n26329 ;
  assign n26331 = ~n26312 & ~n26330 ;
  assign n26332 = ~n26326 & n26331 ;
  assign n26333 = ~n26321 & n26332 ;
  assign n26334 = n26310 & ~n26333 ;
  assign n26349 = ~n26304 & ~n26334 ;
  assign n26350 = ~n26348 & n26349 ;
  assign n26351 = ~\u2_L0_reg[28]/NET0131  & ~n26350 ;
  assign n26352 = \u2_L0_reg[28]/NET0131  & n26350 ;
  assign n26353 = ~n26351 & ~n26352 ;
  assign n26386 = ~n26294 & ~n26339 ;
  assign n26387 = ~n26279 & ~n26386 ;
  assign n26377 = n26279 & n26324 ;
  assign n26378 = ~n26273 & ~n26279 ;
  assign n26379 = n26293 & ~n26303 ;
  assign n26380 = n26378 & n26379 ;
  assign n26381 = ~n26377 & ~n26380 ;
  assign n26361 = n26279 & n26286 ;
  assign n26382 = ~n26327 & ~n26361 ;
  assign n26383 = ~n26273 & n26317 ;
  assign n26384 = ~n26303 & ~n26383 ;
  assign n26385 = ~n26382 & n26384 ;
  assign n26388 = n26381 & ~n26385 ;
  assign n26389 = ~n26387 & n26388 ;
  assign n26390 = ~n26310 & ~n26389 ;
  assign n26354 = ~n26279 & ~n26319 ;
  assign n26355 = n26273 & ~n26279 ;
  assign n26356 = ~n26338 & ~n26355 ;
  assign n26357 = n26303 & ~n26356 ;
  assign n26358 = ~n26354 & ~n26357 ;
  assign n26359 = n26310 & ~n26358 ;
  assign n26364 = n26280 & ~n26293 ;
  assign n26365 = ~n26286 & n26364 ;
  assign n26362 = n26327 & n26361 ;
  assign n26363 = ~n26310 & n26362 ;
  assign n26360 = ~n26279 & n26338 ;
  assign n26366 = n26303 & ~n26360 ;
  assign n26367 = ~n26363 & n26366 ;
  assign n26368 = ~n26365 & n26367 ;
  assign n26369 = n26322 & ~n26355 ;
  assign n26370 = ~n26362 & ~n26369 ;
  assign n26371 = n26310 & ~n26370 ;
  assign n26372 = ~n26280 & ~n26355 ;
  assign n26373 = n26311 & n26372 ;
  assign n26374 = ~n26303 & ~n26373 ;
  assign n26375 = ~n26371 & n26374 ;
  assign n26376 = ~n26368 & ~n26375 ;
  assign n26391 = ~n26359 & ~n26376 ;
  assign n26392 = ~n26390 & n26391 ;
  assign n26393 = \u2_L0_reg[2]/NET0131  & n26392 ;
  assign n26394 = ~\u2_L0_reg[2]/NET0131  & ~n26392 ;
  assign n26395 = ~n26393 & ~n26394 ;
  assign n26403 = n25949 & n26008 ;
  assign n26404 = n26207 & ~n26403 ;
  assign n26405 = n25982 & ~n26028 ;
  assign n26406 = n26205 & ~n26405 ;
  assign n26407 = ~n26404 & ~n26406 ;
  assign n26408 = ~n26018 & ~n26025 ;
  assign n26409 = ~n26226 & n26408 ;
  assign n26410 = ~n26407 & n26409 ;
  assign n26411 = ~n25943 & ~n26410 ;
  assign n26396 = n25979 & n26028 ;
  assign n26397 = ~n25978 & ~n26396 ;
  assign n26398 = n25978 & ~n26029 ;
  assign n26399 = n25981 & n25982 ;
  assign n26400 = ~n26012 & ~n26399 ;
  assign n26401 = n26398 & n26400 ;
  assign n26402 = ~n26397 & ~n26401 ;
  assign n26412 = n25970 & n26007 ;
  assign n26413 = ~n26204 & ~n26412 ;
  assign n26414 = n25978 & ~n26413 ;
  assign n26415 = n25949 & n25989 ;
  assign n26416 = n26032 & ~n26415 ;
  assign n26417 = ~n26414 & n26416 ;
  assign n26418 = n25943 & ~n26417 ;
  assign n26419 = ~n26402 & ~n26418 ;
  assign n26420 = ~n26411 & n26419 ;
  assign n26421 = ~\u2_L0_reg[8]/NET0131  & ~n26420 ;
  assign n26422 = \u2_L0_reg[8]/NET0131  & n26420 ;
  assign n26423 = ~n26421 & ~n26422 ;
  assign n26425 = ~n26364 & n26384 ;
  assign n26427 = ~n26293 & n26378 ;
  assign n26426 = n26279 & n26311 ;
  assign n26428 = n26303 & ~n26426 ;
  assign n26429 = ~n26427 & n26428 ;
  assign n26430 = ~n26425 & ~n26429 ;
  assign n26424 = n26273 & n26323 ;
  assign n26431 = n26310 & ~n26424 ;
  assign n26432 = n26381 & n26431 ;
  assign n26433 = ~n26430 & n26432 ;
  assign n26435 = n26311 & ~n26372 ;
  assign n26434 = n26315 & n26378 ;
  assign n26436 = ~n26303 & ~n26310 ;
  assign n26437 = ~n26313 & n26436 ;
  assign n26438 = ~n26434 & n26437 ;
  assign n26439 = ~n26435 & n26438 ;
  assign n26440 = ~n26433 & ~n26439 ;
  assign n26441 = ~n26279 & n26317 ;
  assign n26442 = n26273 & n26441 ;
  assign n26443 = ~n26296 & ~n26442 ;
  assign n26444 = ~n26440 & n26443 ;
  assign n26445 = ~n26295 & ~n26311 ;
  assign n26446 = ~n26335 & n26445 ;
  assign n26447 = ~n26279 & ~n26446 ;
  assign n26448 = ~n26294 & n26336 ;
  assign n26449 = n26303 & ~n26310 ;
  assign n26450 = ~n26448 & n26449 ;
  assign n26451 = ~n26447 & n26450 ;
  assign n26452 = ~n26444 & ~n26451 ;
  assign n26453 = ~\u2_L0_reg[13]/NET0131  & ~n26452 ;
  assign n26454 = \u2_L0_reg[13]/NET0131  & n26452 ;
  assign n26455 = ~n26453 & ~n26454 ;
  assign n26477 = n25538 & n25569 ;
  assign n26478 = ~n25553 & ~n26477 ;
  assign n26479 = n25559 & ~n26478 ;
  assign n26476 = n25586 & n25600 ;
  assign n26480 = ~n26057 & ~n26476 ;
  assign n26481 = ~n26479 & n26480 ;
  assign n26482 = n25526 & ~n26481 ;
  assign n26472 = ~n25538 & n26040 ;
  assign n26473 = ~n25605 & ~n26055 ;
  assign n26474 = ~n26472 & n26473 ;
  assign n26475 = ~n25559 & ~n26474 ;
  assign n26458 = ~n25545 & n25578 ;
  assign n26461 = ~n25571 & ~n25604 ;
  assign n26462 = ~n26458 & n26461 ;
  assign n26456 = n25538 & n25572 ;
  assign n26457 = n25559 & n26456 ;
  assign n26459 = ~n25561 & ~n25578 ;
  assign n26460 = n25591 & n26459 ;
  assign n26463 = ~n26457 & ~n26460 ;
  assign n26464 = n26462 & n26463 ;
  assign n26465 = ~n25526 & ~n26464 ;
  assign n26466 = ~n25589 & ~n26456 ;
  assign n26467 = n25577 & ~n26466 ;
  assign n26468 = ~n25608 & ~n26456 ;
  assign n26469 = ~n25563 & n26468 ;
  assign n26470 = n25526 & ~n25559 ;
  assign n26471 = ~n26469 & n26470 ;
  assign n26483 = ~n26467 & ~n26471 ;
  assign n26484 = ~n26465 & n26483 ;
  assign n26485 = ~n26475 & n26484 ;
  assign n26486 = ~n26482 & n26485 ;
  assign n26487 = \u2_L0_reg[23]/NET0131  & ~n26486 ;
  assign n26488 = ~\u2_L0_reg[23]/NET0131  & n26486 ;
  assign n26489 = ~n26487 & ~n26488 ;
  assign n26490 = ~n25824 & ~n26171 ;
  assign n26491 = ~n26176 & n26490 ;
  assign n26492 = ~n25836 & ~n26491 ;
  assign n26493 = n25836 & ~n25843 ;
  assign n26494 = ~n26142 & n26493 ;
  assign n26495 = ~n25819 & ~n26156 ;
  assign n26496 = ~n25862 & n26495 ;
  assign n26497 = ~n26494 & n26496 ;
  assign n26498 = ~n26492 & n26497 ;
  assign n26499 = n25792 & ~n26498 ;
  assign n26506 = n25844 & ~n25860 ;
  assign n26507 = n25836 & ~n26141 ;
  assign n26508 = ~n26506 & n26507 ;
  assign n26504 = n25804 & n25811 ;
  assign n26505 = n26134 & n26504 ;
  assign n26509 = ~n26189 & ~n26505 ;
  assign n26510 = ~n25841 & n26509 ;
  assign n26511 = ~n26508 & n26510 ;
  assign n26512 = ~n25792 & ~n26511 ;
  assign n26500 = n25836 & n25861 ;
  assign n26501 = n25844 & ~n25848 ;
  assign n26502 = ~n25829 & ~n26501 ;
  assign n26503 = ~n25836 & ~n26502 ;
  assign n26513 = ~n26500 & ~n26503 ;
  assign n26514 = ~n26512 & n26513 ;
  assign n26515 = ~n26499 & n26514 ;
  assign n26516 = ~\u2_L0_reg[27]/NET0131  & ~n26515 ;
  assign n26517 = \u2_L0_reg[27]/NET0131  & n26515 ;
  assign n26518 = ~n26516 & ~n26517 ;
  assign n26534 = ~n25461 & ~n25505 ;
  assign n26535 = ~n25445 & n25908 ;
  assign n26536 = ~n26534 & ~n26535 ;
  assign n26521 = ~n25445 & n25504 ;
  assign n26537 = n25439 & n26521 ;
  assign n26538 = ~n26536 & ~n26537 ;
  assign n26539 = ~n25484 & ~n26538 ;
  assign n26540 = n25439 & n25907 ;
  assign n26541 = ~n25445 & ~n25484 ;
  assign n26542 = n26540 & ~n26541 ;
  assign n26543 = ~n25445 & n25461 ;
  assign n26544 = ~n25467 & ~n26543 ;
  assign n26545 = n25484 & ~n26544 ;
  assign n26546 = ~n26542 & ~n26545 ;
  assign n26547 = ~n26539 & n26546 ;
  assign n26548 = n25474 & ~n26547 ;
  assign n26519 = ~n25919 & ~n25924 ;
  assign n26520 = ~n25484 & ~n26519 ;
  assign n26522 = n25484 & ~n25919 ;
  assign n26523 = ~n26521 & n26522 ;
  assign n26524 = ~n26520 & ~n26523 ;
  assign n26525 = n25445 & n25919 ;
  assign n26526 = n25466 & n25493 ;
  assign n26527 = ~n26525 & ~n26526 ;
  assign n26528 = n25464 & n26527 ;
  assign n26529 = ~n26524 & n26528 ;
  assign n26530 = ~n25474 & ~n26529 ;
  assign n26531 = n25460 & n25484 ;
  assign n26532 = n25502 & ~n25907 ;
  assign n26533 = n25494 & n26532 ;
  assign n26549 = ~n26531 & ~n26533 ;
  assign n26550 = ~n26530 & n26549 ;
  assign n26551 = ~n26548 & n26550 ;
  assign n26552 = \u2_L0_reg[32]/NET0131  & n26551 ;
  assign n26553 = ~\u2_L0_reg[32]/NET0131  & ~n26551 ;
  assign n26554 = ~n26552 & ~n26553 ;
  assign n26556 = n26005 & n26205 ;
  assign n26557 = ~n25968 & n25982 ;
  assign n26558 = n25978 & ~n25980 ;
  assign n26559 = ~n26557 & n26558 ;
  assign n26560 = ~n26556 & ~n26559 ;
  assign n26555 = ~n25979 & n26028 ;
  assign n26561 = ~n25943 & ~n26555 ;
  assign n26562 = ~n26560 & n26561 ;
  assign n26563 = ~n25949 & n26011 ;
  assign n26564 = ~n25985 & ~n26563 ;
  assign n26565 = n25978 & ~n26564 ;
  assign n26566 = ~n25978 & n25990 ;
  assign n26567 = n25943 & ~n26396 ;
  assign n26568 = ~n26013 & n26567 ;
  assign n26569 = ~n26566 & n26568 ;
  assign n26570 = ~n26565 & n26569 ;
  assign n26571 = ~n26562 & ~n26570 ;
  assign n26572 = n26398 & ~n26403 ;
  assign n26573 = ~n25989 & ~n26205 ;
  assign n26574 = ~n25998 & ~n26412 ;
  assign n26575 = ~n26573 & n26574 ;
  assign n26576 = ~n26572 & ~n26575 ;
  assign n26577 = ~n26571 & ~n26576 ;
  assign n26578 = ~\u2_L0_reg[3]/NET0131  & ~n26577 ;
  assign n26579 = \u2_L0_reg[3]/NET0131  & n26577 ;
  assign n26580 = ~n26578 & ~n26579 ;
  assign n26615 = decrypt_pad & ~\u2_uk_K_r0_reg[20]/NET0131  ;
  assign n26616 = ~decrypt_pad & ~\u2_uk_K_r0_reg[41]/NET0131  ;
  assign n26617 = ~n26615 & ~n26616 ;
  assign n26618 = \u2_R0_reg[11]/P0001  & ~n26617 ;
  assign n26619 = ~\u2_R0_reg[11]/P0001  & n26617 ;
  assign n26620 = ~n26618 & ~n26619 ;
  assign n26581 = decrypt_pad & ~\u2_uk_K_r0_reg[3]/NET0131  ;
  assign n26582 = ~decrypt_pad & ~\u2_uk_K_r0_reg[24]/P0001  ;
  assign n26583 = ~n26581 & ~n26582 ;
  assign n26584 = \u2_R0_reg[12]/NET0131  & ~n26583 ;
  assign n26585 = ~\u2_R0_reg[12]/NET0131  & n26583 ;
  assign n26586 = ~n26584 & ~n26585 ;
  assign n26594 = decrypt_pad & ~\u2_uk_K_r0_reg[48]/NET0131  ;
  assign n26595 = ~decrypt_pad & ~\u2_uk_K_r0_reg[12]/NET0131  ;
  assign n26596 = ~n26594 & ~n26595 ;
  assign n26597 = \u2_R0_reg[13]/NET0131  & ~n26596 ;
  assign n26598 = ~\u2_R0_reg[13]/NET0131  & n26596 ;
  assign n26599 = ~n26597 & ~n26598 ;
  assign n26607 = decrypt_pad & ~\u2_uk_K_r0_reg[11]/NET0131  ;
  assign n26608 = ~decrypt_pad & ~\u2_uk_K_r0_reg[32]/NET0131  ;
  assign n26609 = ~n26607 & ~n26608 ;
  assign n26610 = \u2_R0_reg[9]/NET0131  & ~n26609 ;
  assign n26611 = ~\u2_R0_reg[9]/NET0131  & n26609 ;
  assign n26612 = ~n26610 & ~n26611 ;
  assign n26652 = n26599 & ~n26612 ;
  assign n26600 = decrypt_pad & ~\u2_uk_K_r0_reg[39]/NET0131  ;
  assign n26601 = ~decrypt_pad & ~\u2_uk_K_r0_reg[3]/NET0131  ;
  assign n26602 = ~n26600 & ~n26601 ;
  assign n26603 = \u2_R0_reg[8]/NET0131  & ~n26602 ;
  assign n26604 = ~\u2_R0_reg[8]/NET0131  & n26602 ;
  assign n26605 = ~n26603 & ~n26604 ;
  assign n26606 = ~n26599 & ~n26605 ;
  assign n26622 = n26599 & n26605 ;
  assign n26631 = ~n26606 & ~n26622 ;
  assign n26626 = n26605 & ~n26612 ;
  assign n26587 = decrypt_pad & ~\u2_uk_K_r0_reg[19]/NET0131  ;
  assign n26588 = ~decrypt_pad & ~\u2_uk_K_r0_reg[40]/NET0131  ;
  assign n26589 = ~n26587 & ~n26588 ;
  assign n26590 = \u2_R0_reg[10]/NET0131  & ~n26589 ;
  assign n26591 = ~\u2_R0_reg[10]/NET0131  & n26589 ;
  assign n26592 = ~n26590 & ~n26591 ;
  assign n26653 = ~n26592 & ~n26605 ;
  assign n26654 = ~n26626 & ~n26653 ;
  assign n26655 = n26631 & n26654 ;
  assign n26656 = ~n26652 & ~n26655 ;
  assign n26657 = n26586 & ~n26656 ;
  assign n26640 = ~n26592 & ~n26612 ;
  assign n26651 = n26606 & n26640 ;
  assign n26632 = n26592 & ~n26612 ;
  assign n26658 = n26599 & n26632 ;
  assign n26659 = ~n26651 & ~n26658 ;
  assign n26660 = ~n26657 & n26659 ;
  assign n26661 = n26620 & ~n26660 ;
  assign n26642 = n26599 & ~n26605 ;
  assign n26643 = n26612 & n26642 ;
  assign n26644 = n26592 & ~n26620 ;
  assign n26645 = n26643 & n26644 ;
  assign n26633 = ~n26631 & n26632 ;
  assign n26634 = ~n26599 & n26612 ;
  assign n26635 = n26592 & n26605 ;
  assign n26636 = n26634 & n26635 ;
  assign n26646 = ~n26633 & ~n26636 ;
  assign n26647 = ~n26645 & n26646 ;
  assign n26624 = ~n26592 & n26612 ;
  assign n26637 = n26599 & n26620 ;
  assign n26638 = n26631 & ~n26637 ;
  assign n26639 = n26624 & ~n26638 ;
  assign n26641 = n26638 & n26640 ;
  assign n26648 = ~n26639 & ~n26641 ;
  assign n26649 = n26647 & n26648 ;
  assign n26650 = ~n26586 & ~n26649 ;
  assign n26593 = n26586 & n26592 ;
  assign n26613 = n26606 & n26612 ;
  assign n26614 = n26593 & n26613 ;
  assign n26621 = n26586 & ~n26620 ;
  assign n26627 = ~n26599 & n26626 ;
  assign n26623 = n26612 & n26622 ;
  assign n26625 = n26599 & n26624 ;
  assign n26628 = ~n26623 & ~n26625 ;
  assign n26629 = ~n26627 & n26628 ;
  assign n26630 = n26621 & ~n26629 ;
  assign n26662 = ~n26614 & ~n26630 ;
  assign n26663 = ~n26650 & n26662 ;
  assign n26664 = ~n26661 & n26663 ;
  assign n26665 = ~\u2_L0_reg[6]/NET0131  & ~n26664 ;
  assign n26666 = \u2_L0_reg[6]/NET0131  & n26664 ;
  assign n26667 = ~n26665 & ~n26666 ;
  assign n26668 = n25445 & ~n25908 ;
  assign n26669 = ~n26521 & ~n26668 ;
  assign n26670 = n25439 & ~n26669 ;
  assign n26671 = ~n25439 & ~n25465 ;
  assign n26672 = n25908 & n26671 ;
  assign n26673 = n25484 & ~n26672 ;
  assign n26674 = ~n25452 & ~n25927 ;
  assign n26675 = ~n25484 & ~n26540 ;
  assign n26676 = ~n26668 & n26675 ;
  assign n26677 = ~n26674 & n26676 ;
  assign n26678 = ~n26673 & ~n26677 ;
  assign n26679 = ~n26670 & ~n26678 ;
  assign n26680 = n25474 & ~n26679 ;
  assign n26688 = ~n25484 & n26672 ;
  assign n26689 = ~n25496 & ~n26688 ;
  assign n26690 = ~n25474 & ~n26689 ;
  assign n26682 = ~n25908 & ~n25921 ;
  assign n26683 = ~n25462 & ~n26526 ;
  assign n26684 = ~n26682 & n26683 ;
  assign n26681 = n25474 & ~n25496 ;
  assign n26685 = n25484 & ~n26681 ;
  assign n26686 = ~n26684 & n26685 ;
  assign n26687 = ~n25484 & n26670 ;
  assign n26691 = ~n26686 & ~n26687 ;
  assign n26692 = ~n26690 & n26691 ;
  assign n26693 = ~n26680 & n26692 ;
  assign n26694 = ~\u2_L0_reg[7]/NET0131  & ~n26693 ;
  assign n26695 = \u2_L0_reg[7]/NET0131  & n26693 ;
  assign n26696 = ~n26694 & ~n26695 ;
  assign n26699 = n26592 & n26606 ;
  assign n26700 = ~n26612 & n26699 ;
  assign n26701 = n26620 & ~n26636 ;
  assign n26702 = ~n26700 & n26701 ;
  assign n26722 = ~n26599 & ~n26635 ;
  assign n26723 = ~n26653 & n26722 ;
  assign n26724 = ~n26702 & n26723 ;
  assign n26708 = ~n26612 & ~n26642 ;
  assign n26709 = n26612 & ~n26622 ;
  assign n26710 = ~n26708 & ~n26709 ;
  assign n26717 = n26613 & n26620 ;
  assign n26718 = ~n26710 & ~n26717 ;
  assign n26719 = ~n26592 & ~n26718 ;
  assign n26720 = n26592 & n26643 ;
  assign n26721 = ~n26592 & n26627 ;
  assign n26725 = ~n26720 & ~n26721 ;
  assign n26726 = ~n26719 & n26725 ;
  assign n26727 = ~n26724 & n26726 ;
  assign n26728 = n26586 & ~n26727 ;
  assign n26697 = n26592 & n26626 ;
  assign n26698 = ~n26620 & ~n26697 ;
  assign n26703 = ~n26698 & ~n26702 ;
  assign n26711 = ~n26592 & n26606 ;
  assign n26712 = ~n26710 & ~n26711 ;
  assign n26713 = ~n26620 & ~n26712 ;
  assign n26705 = ~n26606 & n26620 ;
  assign n26704 = ~n26612 & ~n26622 ;
  assign n26706 = ~n26623 & ~n26704 ;
  assign n26707 = n26705 & n26706 ;
  assign n26714 = ~n26651 & ~n26707 ;
  assign n26715 = ~n26713 & n26714 ;
  assign n26716 = ~n26586 & ~n26715 ;
  assign n26729 = ~n26703 & ~n26716 ;
  assign n26730 = ~n26728 & n26729 ;
  assign n26731 = ~\u2_L0_reg[16]/NET0131  & ~n26730 ;
  assign n26732 = \u2_L0_reg[16]/NET0131  & n26730 ;
  assign n26733 = ~n26731 & ~n26732 ;
  assign n26750 = n26599 & n26653 ;
  assign n26751 = ~n26699 & ~n26750 ;
  assign n26752 = ~n26613 & ~n26697 ;
  assign n26753 = n26751 & n26752 ;
  assign n26754 = n26620 & ~n26753 ;
  assign n26755 = ~n26599 & n26697 ;
  assign n26756 = ~n26754 & ~n26755 ;
  assign n26757 = ~n26586 & ~n26756 ;
  assign n26735 = ~n26631 & n26640 ;
  assign n26736 = ~n26655 & ~n26735 ;
  assign n26737 = ~n26620 & ~n26736 ;
  assign n26738 = ~n26586 & ~n26737 ;
  assign n26739 = ~n26592 & n26620 ;
  assign n26740 = n26708 & n26739 ;
  assign n26745 = n26586 & ~n26740 ;
  assign n26741 = n26592 & ~n26626 ;
  assign n26742 = n26705 & n26741 ;
  assign n26743 = ~n26620 & ~n26640 ;
  assign n26744 = ~n26631 & n26743 ;
  assign n26746 = ~n26742 & ~n26744 ;
  assign n26747 = n26745 & n26746 ;
  assign n26748 = ~n26641 & n26747 ;
  assign n26749 = ~n26738 & ~n26748 ;
  assign n26734 = n26623 & n26644 ;
  assign n26758 = ~n26627 & ~n26643 ;
  assign n26759 = n26739 & ~n26758 ;
  assign n26760 = ~n26734 & ~n26759 ;
  assign n26761 = ~n26749 & n26760 ;
  assign n26762 = ~n26757 & n26761 ;
  assign n26763 = ~\u2_L0_reg[24]/NET0131  & ~n26762 ;
  assign n26764 = \u2_L0_reg[24]/NET0131  & n26762 ;
  assign n26765 = ~n26763 & ~n26764 ;
  assign n26767 = ~n26721 & n26751 ;
  assign n26768 = n26586 & ~n26767 ;
  assign n26770 = n26592 & n26634 ;
  assign n26769 = ~n26634 & ~n26635 ;
  assign n26771 = ~n26586 & ~n26769 ;
  assign n26772 = ~n26770 & n26771 ;
  assign n26773 = ~n26768 & ~n26772 ;
  assign n26774 = n26620 & ~n26773 ;
  assign n26775 = ~n26605 & ~n26612 ;
  assign n26776 = ~n26620 & ~n26775 ;
  assign n26777 = n26769 & n26776 ;
  assign n26778 = n26632 & n26642 ;
  assign n26779 = ~n26735 & ~n26778 ;
  assign n26780 = ~n26777 & n26779 ;
  assign n26781 = ~n26586 & ~n26780 ;
  assign n26782 = ~n26613 & ~n26635 ;
  assign n26783 = n26621 & ~n26782 ;
  assign n26785 = n26593 & n26709 ;
  assign n26766 = n26634 & n26644 ;
  assign n26784 = n26637 & n26697 ;
  assign n26786 = ~n26766 & ~n26784 ;
  assign n26787 = ~n26785 & n26786 ;
  assign n26788 = ~n26783 & n26787 ;
  assign n26789 = ~n26781 & n26788 ;
  assign n26790 = ~n26774 & n26789 ;
  assign n26791 = \u2_L0_reg[30]/NET0131  & ~n26790 ;
  assign n26792 = ~\u2_L0_reg[30]/NET0131  & n26790 ;
  assign n26793 = ~n26791 & ~n26792 ;
  assign n26808 = n26044 & n26468 ;
  assign n26809 = n25532 & ~n26808 ;
  assign n26799 = ~n25561 & ~n26477 ;
  assign n26810 = n25577 & ~n26799 ;
  assign n26811 = ~n26055 & ~n26810 ;
  assign n26812 = ~n26809 & n26811 ;
  assign n26813 = n25526 & ~n26812 ;
  assign n26794 = ~n25532 & n26043 ;
  assign n26795 = n25532 & n26477 ;
  assign n26796 = ~n26794 & ~n26795 ;
  assign n26797 = ~n25559 & ~n26796 ;
  assign n26800 = ~n25559 & n26799 ;
  assign n26801 = n25559 & ~n25564 ;
  assign n26802 = ~n25546 & n26801 ;
  assign n26803 = ~n26456 & n26802 ;
  assign n26804 = ~n26800 & ~n26803 ;
  assign n26798 = n25590 & ~n26048 ;
  assign n26805 = ~n26794 & ~n26798 ;
  assign n26806 = ~n26804 & n26805 ;
  assign n26807 = ~n25526 & ~n26806 ;
  assign n26814 = ~n26797 & ~n26807 ;
  assign n26815 = ~n26813 & n26814 ;
  assign n26816 = ~\u2_L0_reg[9]/NET0131  & ~n26815 ;
  assign n26817 = \u2_L0_reg[9]/NET0131  & n26815 ;
  assign n26818 = ~n26816 & ~n26817 ;
  assign n26821 = n26303 & ~n26386 ;
  assign n26819 = ~n26316 & ~n26441 ;
  assign n26820 = ~n26303 & ~n26819 ;
  assign n26822 = ~n26365 & ~n26820 ;
  assign n26823 = ~n26821 & n26822 ;
  assign n26824 = n26310 & ~n26823 ;
  assign n26829 = ~n26362 & ~n26427 ;
  assign n26830 = ~n26296 & n26829 ;
  assign n26825 = n26303 & n26318 ;
  assign n26826 = n26279 & n26303 ;
  assign n26827 = ~n26286 & ~n26826 ;
  assign n26828 = n26372 & n26827 ;
  assign n26831 = ~n26825 & ~n26828 ;
  assign n26832 = n26830 & n26831 ;
  assign n26833 = ~n26310 & ~n26832 ;
  assign n26834 = ~n26303 & n26324 ;
  assign n26835 = n26279 & n26317 ;
  assign n26836 = ~n26424 & ~n26835 ;
  assign n26837 = n26303 & ~n26836 ;
  assign n26838 = ~n26834 & ~n26837 ;
  assign n26839 = ~n26833 & n26838 ;
  assign n26840 = ~n26824 & n26839 ;
  assign n26841 = ~\u2_L0_reg[18]/P0001  & ~n26840 ;
  assign n26842 = \u2_L0_reg[18]/P0001  & n26840 ;
  assign n26843 = ~n26841 & ~n26842 ;
  assign n26844 = decrypt_pad & ~\u1_uk_K_r1_reg[44]/P0001  ;
  assign n26845 = ~decrypt_pad & ~\u1_uk_K_r1_reg[50]/NET0131  ;
  assign n26846 = ~n26844 & ~n26845 ;
  assign n26847 = \u1_R1_reg[20]/NET0131  & ~n26846 ;
  assign n26848 = ~\u1_R1_reg[20]/NET0131  & n26846 ;
  assign n26849 = ~n26847 & ~n26848 ;
  assign n26870 = decrypt_pad & ~\u1_uk_K_r1_reg[29]/NET0131  ;
  assign n26871 = ~decrypt_pad & ~\u1_uk_K_r1_reg[35]/NET0131  ;
  assign n26872 = ~n26870 & ~n26871 ;
  assign n26873 = \u1_R1_reg[19]/NET0131  & ~n26872 ;
  assign n26874 = ~\u1_R1_reg[19]/NET0131  & n26872 ;
  assign n26875 = ~n26873 & ~n26874 ;
  assign n26850 = decrypt_pad & ~\u1_uk_K_r1_reg[42]/NET0131  ;
  assign n26851 = ~decrypt_pad & ~\u1_uk_K_r1_reg[52]/NET0131  ;
  assign n26852 = ~n26850 & ~n26851 ;
  assign n26853 = \u1_R1_reg[18]/NET0131  & ~n26852 ;
  assign n26854 = ~\u1_R1_reg[18]/NET0131  & n26852 ;
  assign n26855 = ~n26853 & ~n26854 ;
  assign n26876 = decrypt_pad & ~\u1_uk_K_r1_reg[2]/NET0131  ;
  assign n26877 = ~decrypt_pad & ~\u1_uk_K_r1_reg[8]/NET0131  ;
  assign n26878 = ~n26876 & ~n26877 ;
  assign n26879 = \u1_R1_reg[16]/NET0131  & ~n26878 ;
  assign n26880 = ~\u1_R1_reg[16]/NET0131  & n26878 ;
  assign n26881 = ~n26879 & ~n26880 ;
  assign n26886 = n26855 & n26881 ;
  assign n26856 = decrypt_pad & ~\u1_uk_K_r1_reg[14]/NET0131  ;
  assign n26857 = ~decrypt_pad & ~\u1_uk_K_r1_reg[51]/NET0131  ;
  assign n26858 = ~n26856 & ~n26857 ;
  assign n26859 = \u1_R1_reg[21]/NET0131  & ~n26858 ;
  assign n26860 = ~\u1_R1_reg[21]/NET0131  & n26858 ;
  assign n26861 = ~n26859 & ~n26860 ;
  assign n26863 = decrypt_pad & ~\u1_uk_K_r1_reg[52]/NET0131  ;
  assign n26864 = ~decrypt_pad & ~\u1_uk_K_r1_reg[30]/NET0131  ;
  assign n26865 = ~n26863 & ~n26864 ;
  assign n26866 = \u1_R1_reg[17]/NET0131  & ~n26865 ;
  assign n26867 = ~\u1_R1_reg[17]/NET0131  & n26865 ;
  assign n26868 = ~n26866 & ~n26867 ;
  assign n26885 = ~n26855 & n26868 ;
  assign n26887 = ~n26861 & ~n26885 ;
  assign n26888 = ~n26886 & n26887 ;
  assign n26882 = ~n26868 & ~n26881 ;
  assign n26883 = n26861 & n26881 ;
  assign n26884 = n26868 & n26883 ;
  assign n26889 = ~n26882 & ~n26884 ;
  assign n26890 = ~n26888 & n26889 ;
  assign n26891 = n26875 & ~n26890 ;
  assign n26892 = ~n26881 & n26885 ;
  assign n26893 = ~n26868 & n26883 ;
  assign n26894 = ~n26892 & ~n26893 ;
  assign n26895 = ~n26875 & ~n26894 ;
  assign n26862 = ~n26855 & n26861 ;
  assign n26869 = n26862 & n26868 ;
  assign n26896 = n26855 & n26868 ;
  assign n26897 = ~n26861 & n26881 ;
  assign n26898 = n26896 & n26897 ;
  assign n26899 = ~n26869 & ~n26898 ;
  assign n26900 = ~n26895 & n26899 ;
  assign n26901 = ~n26891 & n26900 ;
  assign n26902 = n26849 & ~n26901 ;
  assign n26918 = ~n26861 & n26882 ;
  assign n26919 = n26855 & n26918 ;
  assign n26920 = ~n26898 & ~n26919 ;
  assign n26921 = n26862 & n26882 ;
  assign n26922 = n26920 & ~n26921 ;
  assign n26923 = n26875 & ~n26922 ;
  assign n26903 = ~n26881 & n26896 ;
  assign n26904 = ~n26868 & n26897 ;
  assign n26905 = ~n26903 & ~n26904 ;
  assign n26906 = ~n26861 & n26875 ;
  assign n26907 = ~n26905 & ~n26906 ;
  assign n26909 = ~n26861 & n26868 ;
  assign n26910 = n26875 & ~n26909 ;
  assign n26908 = ~n26875 & ~n26882 ;
  assign n26911 = ~n26855 & ~n26908 ;
  assign n26912 = ~n26910 & n26911 ;
  assign n26913 = ~n26907 & ~n26912 ;
  assign n26914 = ~n26849 & ~n26913 ;
  assign n26915 = n26855 & ~n26868 ;
  assign n26916 = ~n26875 & n26881 ;
  assign n26917 = n26915 & n26916 ;
  assign n26924 = ~n26855 & n26884 ;
  assign n26925 = ~n26917 & ~n26924 ;
  assign n26926 = ~n26914 & n26925 ;
  assign n26927 = ~n26923 & n26926 ;
  assign n26928 = ~n26902 & n26927 ;
  assign n26929 = \u1_L1_reg[25]/NET0131  & n26928 ;
  assign n26930 = ~\u1_L1_reg[25]/NET0131  & ~n26928 ;
  assign n26931 = ~n26929 & ~n26930 ;
  assign n26973 = decrypt_pad & ~\u2_key_r_reg[35]/P0001  ;
  assign n26974 = ~decrypt_pad & ~\u2_key_r_reg[42]/P0001  ;
  assign n26975 = ~n26973 & ~n26974 ;
  assign n26976 = \u2_desIn_r_reg[25]/NET0131  & ~n26975 ;
  assign n26977 = ~\u2_desIn_r_reg[25]/NET0131  & n26975 ;
  assign n26978 = ~n26976 & ~n26977 ;
  assign n26966 = decrypt_pad & ~\u2_key_r_reg[52]/NET0131  ;
  assign n26967 = ~decrypt_pad & ~\u2_key_r_reg[0]/NET0131  ;
  assign n26968 = ~n26966 & ~n26967 ;
  assign n26969 = \u2_desIn_r_reg[17]/NET0131  & ~n26968 ;
  assign n26970 = ~\u2_desIn_r_reg[17]/NET0131  & n26968 ;
  assign n26971 = ~n26969 & ~n26970 ;
  assign n26945 = decrypt_pad & ~\u2_key_r_reg[15]/NET0131  ;
  assign n26946 = ~decrypt_pad & ~\u2_key_r_reg[22]/NET0131  ;
  assign n26947 = ~n26945 & ~n26946 ;
  assign n26948 = \u2_desIn_r_reg[9]/NET0131  & ~n26947 ;
  assign n26949 = ~\u2_desIn_r_reg[9]/NET0131  & n26947 ;
  assign n26950 = ~n26948 & ~n26949 ;
  assign n26932 = decrypt_pad & ~\u2_key_r_reg[31]/NET0131  ;
  assign n26933 = ~decrypt_pad & ~\u2_key_r_reg[38]/NET0131  ;
  assign n26934 = ~n26932 & ~n26933 ;
  assign n26935 = \u2_desIn_r_reg[33]/NET0131  & ~n26934 ;
  assign n26936 = ~\u2_desIn_r_reg[33]/NET0131  & n26934 ;
  assign n26937 = ~n26935 & ~n26936 ;
  assign n26938 = decrypt_pad & ~\u2_key_r_reg[50]/NET0131  ;
  assign n26939 = ~decrypt_pad & ~\u2_key_r_reg[2]/NET0131  ;
  assign n26940 = ~n26938 & ~n26939 ;
  assign n26941 = \u2_desIn_r_reg[59]/NET0131  & ~n26940 ;
  assign n26942 = ~\u2_desIn_r_reg[59]/NET0131  & n26940 ;
  assign n26943 = ~n26941 & ~n26942 ;
  assign n26951 = decrypt_pad & ~\u2_key_r_reg[30]/NET0131  ;
  assign n26952 = ~decrypt_pad & ~\u2_key_r_reg[37]/NET0131  ;
  assign n26953 = ~n26951 & ~n26952 ;
  assign n26954 = \u2_desIn_r_reg[1]/NET0131  & ~n26953 ;
  assign n26955 = ~\u2_desIn_r_reg[1]/NET0131  & n26953 ;
  assign n26956 = ~n26954 & ~n26955 ;
  assign n26998 = n26943 & ~n26956 ;
  assign n26999 = n26937 & n26998 ;
  assign n27000 = ~n26950 & n26999 ;
  assign n26944 = n26937 & ~n26943 ;
  assign n27001 = n26944 & n26956 ;
  assign n27002 = ~n27000 & ~n27001 ;
  assign n27003 = ~n26971 & ~n27002 ;
  assign n26957 = n26950 & ~n26956 ;
  assign n27004 = n26937 & n26956 ;
  assign n27005 = ~n26950 & n27004 ;
  assign n27006 = ~n26957 & ~n27005 ;
  assign n27007 = n26943 & n26971 ;
  assign n27008 = ~n27006 & n27007 ;
  assign n26958 = n26944 & n26957 ;
  assign n26963 = ~n26937 & ~n26956 ;
  assign n26979 = ~n26943 & n26963 ;
  assign n26997 = ~n26950 & n26979 ;
  assign n27009 = ~n26958 & ~n26997 ;
  assign n27010 = ~n27008 & n27009 ;
  assign n27011 = ~n27003 & n27010 ;
  assign n27012 = n26978 & ~n27011 ;
  assign n26980 = n26950 & n26979 ;
  assign n26981 = ~n26971 & n26980 ;
  assign n26982 = ~n26956 & n26971 ;
  assign n26983 = ~n26937 & ~n26971 ;
  assign n26984 = ~n26982 & ~n26983 ;
  assign n26985 = n26943 & ~n26957 ;
  assign n26986 = ~n26984 & n26985 ;
  assign n26987 = ~n26981 & ~n26986 ;
  assign n26988 = ~n26978 & ~n26987 ;
  assign n26959 = ~n26943 & n26950 ;
  assign n26960 = n26956 & n26959 ;
  assign n26961 = ~n26937 & n26960 ;
  assign n26962 = ~n26958 & ~n26961 ;
  assign n26964 = ~n26959 & n26963 ;
  assign n26965 = n26962 & ~n26964 ;
  assign n26972 = ~n26965 & n26971 ;
  assign n26992 = n26956 & ~n26971 ;
  assign n26993 = n26937 & ~n26978 ;
  assign n26994 = ~n26992 & ~n26993 ;
  assign n26989 = ~n26943 & ~n26950 ;
  assign n26990 = n26943 & n26950 ;
  assign n26991 = ~n26989 & ~n26990 ;
  assign n26995 = ~n26982 & ~n26991 ;
  assign n26996 = ~n26994 & n26995 ;
  assign n27013 = ~n26972 & ~n26996 ;
  assign n27014 = ~n26988 & n27013 ;
  assign n27015 = ~n27012 & n27014 ;
  assign n27016 = ~\u2_desIn_r_reg[42]/NET0131  & ~n27015 ;
  assign n27017 = \u2_desIn_r_reg[42]/NET0131  & n27015 ;
  assign n27018 = ~n27016 & ~n27017 ;
  assign n27032 = decrypt_pad & ~\u2_key_r_reg[53]/NET0131  ;
  assign n27033 = ~decrypt_pad & ~\u2_key_r_reg[3]/NET0131  ;
  assign n27034 = ~n27032 & ~n27033 ;
  assign n27035 = \u2_desIn_r_reg[23]/NET0131  & ~n27034 ;
  assign n27036 = ~\u2_desIn_r_reg[23]/NET0131  & n27034 ;
  assign n27037 = ~n27035 & ~n27036 ;
  assign n27039 = decrypt_pad & ~\u2_key_r_reg[4]/NET0131  ;
  assign n27040 = ~decrypt_pad & ~\u2_key_r_reg[11]/NET0131  ;
  assign n27041 = ~n27039 & ~n27040 ;
  assign n27042 = \u2_desIn_r_reg[7]/NET0131  & ~n27041 ;
  assign n27043 = ~\u2_desIn_r_reg[7]/NET0131  & n27041 ;
  assign n27044 = ~n27042 & ~n27043 ;
  assign n27045 = decrypt_pad & ~\u2_key_r_reg[34]/NET0131  ;
  assign n27046 = ~decrypt_pad & ~\u2_key_r_reg[41]/NET0131  ;
  assign n27047 = ~n27045 & ~n27046 ;
  assign n27048 = \u2_desIn_r_reg[39]/NET0131  & ~n27047 ;
  assign n27049 = ~\u2_desIn_r_reg[39]/NET0131  & n27047 ;
  assign n27050 = ~n27048 & ~n27049 ;
  assign n27056 = ~n27044 & n27050 ;
  assign n27019 = decrypt_pad & ~\u2_key_r_reg[19]/NET0131  ;
  assign n27020 = ~decrypt_pad & ~\u2_key_r_reg[26]/NET0131  ;
  assign n27021 = ~n27019 & ~n27020 ;
  assign n27022 = \u2_desIn_r_reg[15]/NET0131  & ~n27021 ;
  assign n27023 = ~\u2_desIn_r_reg[15]/NET0131  & n27021 ;
  assign n27024 = ~n27022 & ~n27023 ;
  assign n27025 = decrypt_pad & ~\u2_key_r_reg[40]/NET0131  ;
  assign n27026 = ~decrypt_pad & ~\u2_key_r_reg[47]/NET0131  ;
  assign n27027 = ~n27025 & ~n27026 ;
  assign n27028 = \u2_desIn_r_reg[57]/NET0131  & ~n27027 ;
  assign n27029 = ~\u2_desIn_r_reg[57]/NET0131  & n27027 ;
  assign n27030 = ~n27028 & ~n27029 ;
  assign n27031 = n27024 & ~n27030 ;
  assign n27057 = n27031 & ~n27050 ;
  assign n27058 = ~n27056 & ~n27057 ;
  assign n27059 = n27037 & ~n27058 ;
  assign n27072 = ~n27024 & n27030 ;
  assign n27073 = ~n27031 & ~n27072 ;
  assign n27071 = n27030 & n27050 ;
  assign n27074 = ~n27044 & ~n27071 ;
  assign n27075 = ~n27073 & n27074 ;
  assign n27060 = ~n27030 & n27050 ;
  assign n27054 = ~n27024 & n27037 ;
  assign n27061 = n27044 & ~n27054 ;
  assign n27062 = n27060 & ~n27061 ;
  assign n27063 = n27030 & ~n27037 ;
  assign n27064 = n27044 & n27063 ;
  assign n27065 = decrypt_pad & ~\u2_key_r_reg[6]/NET0131  ;
  assign n27066 = ~decrypt_pad & ~\u2_key_r_reg[13]/NET0131  ;
  assign n27067 = ~n27065 & ~n27066 ;
  assign n27068 = \u2_desIn_r_reg[31]/NET0131  & ~n27067 ;
  assign n27069 = ~\u2_desIn_r_reg[31]/NET0131  & n27067 ;
  assign n27070 = ~n27068 & ~n27069 ;
  assign n27076 = ~n27064 & n27070 ;
  assign n27077 = ~n27062 & n27076 ;
  assign n27078 = ~n27075 & n27077 ;
  assign n27079 = ~n27059 & n27078 ;
  assign n27038 = n27031 & n27037 ;
  assign n27080 = n27038 & n27050 ;
  assign n27081 = ~n27030 & ~n27050 ;
  assign n27082 = ~n27024 & n27081 ;
  assign n27083 = ~n27080 & ~n27082 ;
  assign n27084 = n27044 & ~n27083 ;
  assign n27051 = ~n27044 & ~n27050 ;
  assign n27093 = n27030 & n27051 ;
  assign n27094 = n27024 & ~n27093 ;
  assign n27092 = ~n27037 & ~n27072 ;
  assign n27095 = ~n27044 & n27060 ;
  assign n27096 = n27092 & ~n27095 ;
  assign n27097 = ~n27094 & n27096 ;
  assign n27085 = n27044 & ~n27050 ;
  assign n27086 = n27030 & n27085 ;
  assign n27087 = n27024 & n27086 ;
  assign n27088 = n27037 & n27087 ;
  assign n27089 = ~n27024 & ~n27044 ;
  assign n27090 = ~n27054 & ~n27089 ;
  assign n27091 = n27071 & ~n27090 ;
  assign n27098 = ~n27070 & ~n27091 ;
  assign n27099 = ~n27088 & n27098 ;
  assign n27100 = ~n27097 & n27099 ;
  assign n27101 = ~n27084 & n27100 ;
  assign n27102 = ~n27079 & ~n27101 ;
  assign n27103 = n27044 & n27071 ;
  assign n27104 = n27024 & ~n27095 ;
  assign n27105 = ~n27103 & n27104 ;
  assign n27106 = ~n27024 & ~n27085 ;
  assign n27107 = ~n27037 & ~n27106 ;
  assign n27108 = ~n27105 & n27107 ;
  assign n27052 = n27038 & n27051 ;
  assign n27053 = n27030 & ~n27044 ;
  assign n27055 = n27053 & n27054 ;
  assign n27109 = ~n27052 & ~n27055 ;
  assign n27110 = ~n27108 & n27109 ;
  assign n27111 = ~n27102 & n27110 ;
  assign n27112 = ~\u2_desIn_r_reg[48]/NET0131  & ~n27111 ;
  assign n27113 = \u2_desIn_r_reg[48]/NET0131  & n27111 ;
  assign n27114 = ~n27112 & ~n27113 ;
  assign n27115 = decrypt_pad & ~\u2_key_r_reg[28]/NET0131  ;
  assign n27116 = ~decrypt_pad & ~\u2_key_r_reg[35]/P0001  ;
  assign n27117 = ~n27115 & ~n27116 ;
  assign n27118 = \u2_desIn_r_reg[59]/NET0131  & ~n27117 ;
  assign n27119 = ~\u2_desIn_r_reg[59]/NET0131  & n27117 ;
  assign n27120 = ~n27118 & ~n27119 ;
  assign n27121 = decrypt_pad & ~\u2_key_r_reg[2]/NET0131  ;
  assign n27122 = ~decrypt_pad & ~\u2_key_r_reg[9]/NET0131  ;
  assign n27123 = ~n27121 & ~n27122 ;
  assign n27124 = \u2_desIn_r_reg[51]/NET0131  & ~n27123 ;
  assign n27125 = ~\u2_desIn_r_reg[51]/NET0131  & n27123 ;
  assign n27126 = ~n27124 & ~n27125 ;
  assign n27140 = decrypt_pad & ~\u2_key_r_reg[44]/NET0131  ;
  assign n27141 = ~decrypt_pad & ~\u2_key_r_reg[51]/NET0131  ;
  assign n27142 = ~n27140 & ~n27141 ;
  assign n27143 = \u2_desIn_r_reg[43]/NET0131  & ~n27142 ;
  assign n27144 = ~\u2_desIn_r_reg[43]/NET0131  & n27142 ;
  assign n27145 = ~n27143 & ~n27144 ;
  assign n27127 = decrypt_pad & ~\u2_key_r_reg[7]/NET0131  ;
  assign n27128 = ~decrypt_pad & ~\u2_key_r_reg[14]/NET0131  ;
  assign n27129 = ~n27127 & ~n27128 ;
  assign n27130 = \u2_desIn_r_reg[27]/NET0131  & ~n27129 ;
  assign n27131 = ~\u2_desIn_r_reg[27]/NET0131  & n27129 ;
  assign n27132 = ~n27130 & ~n27131 ;
  assign n27133 = decrypt_pad & ~\u2_key_r_reg[22]/NET0131  ;
  assign n27134 = ~decrypt_pad & ~\u2_key_r_reg[29]/NET0131  ;
  assign n27135 = ~n27133 & ~n27134 ;
  assign n27136 = \u2_desIn_r_reg[35]/NET0131  & ~n27135 ;
  assign n27137 = ~\u2_desIn_r_reg[35]/NET0131  & n27135 ;
  assign n27138 = ~n27136 & ~n27137 ;
  assign n27154 = ~n27132 & n27138 ;
  assign n27155 = n27145 & n27154 ;
  assign n27161 = ~n27126 & ~n27155 ;
  assign n27188 = n27138 & ~n27145 ;
  assign n27189 = n27132 & n27188 ;
  assign n27190 = n27161 & ~n27189 ;
  assign n27146 = decrypt_pad & ~\u2_key_r_reg[23]/NET0131  ;
  assign n27147 = ~decrypt_pad & ~\u2_key_r_reg[30]/NET0131  ;
  assign n27148 = ~n27146 & ~n27147 ;
  assign n27149 = \u2_desIn_r_reg[1]/NET0131  & ~n27148 ;
  assign n27150 = ~\u2_desIn_r_reg[1]/NET0131  & n27148 ;
  assign n27151 = ~n27149 & ~n27150 ;
  assign n27180 = ~n27132 & n27151 ;
  assign n27181 = ~n27138 & n27180 ;
  assign n27182 = n27126 & ~n27181 ;
  assign n27191 = ~n27132 & ~n27145 ;
  assign n27139 = n27132 & ~n27138 ;
  assign n27192 = n27139 & n27145 ;
  assign n27193 = ~n27191 & ~n27192 ;
  assign n27194 = n27182 & n27193 ;
  assign n27195 = ~n27190 & ~n27194 ;
  assign n27183 = n27132 & ~n27151 ;
  assign n27177 = ~n27126 & ~n27145 ;
  assign n27196 = ~n27177 & ~n27188 ;
  assign n27197 = n27183 & ~n27196 ;
  assign n27156 = n27132 & n27151 ;
  assign n27162 = n27145 & n27156 ;
  assign n27198 = ~n27138 & n27162 ;
  assign n27199 = ~n27197 & ~n27198 ;
  assign n27200 = ~n27195 & n27199 ;
  assign n27201 = ~n27120 & ~n27200 ;
  assign n27157 = n27138 & n27156 ;
  assign n27152 = ~n27145 & ~n27151 ;
  assign n27153 = n27139 & n27152 ;
  assign n27158 = ~n27153 & ~n27155 ;
  assign n27159 = ~n27157 & n27158 ;
  assign n27160 = n27126 & ~n27159 ;
  assign n27165 = n27139 & n27151 ;
  assign n27163 = n27138 & n27151 ;
  assign n27164 = ~n27132 & n27163 ;
  assign n27166 = ~n27145 & ~n27164 ;
  assign n27167 = ~n27165 & n27166 ;
  assign n27168 = n27161 & ~n27162 ;
  assign n27169 = ~n27167 & n27168 ;
  assign n27170 = ~n27160 & ~n27169 ;
  assign n27171 = n27120 & ~n27170 ;
  assign n27184 = n27138 & n27183 ;
  assign n27185 = ~n27126 & ~n27184 ;
  assign n27186 = ~n27145 & ~n27182 ;
  assign n27187 = ~n27185 & n27186 ;
  assign n27172 = ~n27132 & ~n27151 ;
  assign n27173 = n27138 & n27172 ;
  assign n27174 = ~n27145 & n27173 ;
  assign n27175 = ~n27162 & ~n27174 ;
  assign n27176 = n27126 & ~n27175 ;
  assign n27178 = ~n27138 & n27172 ;
  assign n27179 = n27177 & n27178 ;
  assign n27202 = ~n27176 & ~n27179 ;
  assign n27203 = ~n27187 & n27202 ;
  assign n27204 = ~n27171 & n27203 ;
  assign n27205 = ~n27201 & n27204 ;
  assign n27206 = ~\u2_desIn_r_reg[20]/NET0131  & n27205 ;
  assign n27207 = \u2_desIn_r_reg[20]/NET0131  & ~n27205 ;
  assign n27208 = ~n27206 & ~n27207 ;
  assign n27209 = decrypt_pad & ~\u2_key_r_reg[13]/NET0131  ;
  assign n27210 = ~decrypt_pad & ~\u2_key_r_reg[20]/NET0131  ;
  assign n27211 = ~n27209 & ~n27210 ;
  assign n27212 = \u2_desIn_r_reg[3]/NET0131  & ~n27211 ;
  assign n27213 = ~\u2_desIn_r_reg[3]/NET0131  & n27211 ;
  assign n27214 = ~n27212 & ~n27213 ;
  assign n27215 = decrypt_pad & ~\u2_key_r_reg[54]/NET0131  ;
  assign n27216 = ~decrypt_pad & ~\u2_key_r_reg[4]/NET0131  ;
  assign n27217 = ~n27215 & ~n27216 ;
  assign n27218 = \u2_desIn_r_reg[29]/NET0131  & ~n27217 ;
  assign n27219 = ~\u2_desIn_r_reg[29]/NET0131  & n27217 ;
  assign n27220 = ~n27218 & ~n27219 ;
  assign n27221 = ~n27214 & ~n27220 ;
  assign n27222 = decrypt_pad & ~\u2_key_r_reg[48]/NET0131  ;
  assign n27223 = ~decrypt_pad & ~\u2_key_r_reg[55]/NET0131  ;
  assign n27224 = ~n27222 & ~n27223 ;
  assign n27225 = \u2_desIn_r_reg[37]/NET0131  & ~n27224 ;
  assign n27226 = ~\u2_desIn_r_reg[37]/NET0131  & n27224 ;
  assign n27227 = ~n27225 & ~n27226 ;
  assign n27254 = n27221 & ~n27227 ;
  assign n27246 = n27214 & n27220 ;
  assign n27247 = n27227 & n27246 ;
  assign n27248 = decrypt_pad & ~\u2_key_r_reg[25]/NET0131  ;
  assign n27249 = ~decrypt_pad & ~\u2_key_r_reg[32]/NET0131  ;
  assign n27250 = ~n27248 & ~n27249 ;
  assign n27251 = \u2_desIn_r_reg[53]/NET0131  & ~n27250 ;
  assign n27252 = ~\u2_desIn_r_reg[53]/NET0131  & n27250 ;
  assign n27253 = ~n27251 & ~n27252 ;
  assign n27255 = ~n27247 & n27253 ;
  assign n27256 = ~n27254 & n27255 ;
  assign n27229 = decrypt_pad & ~\u2_key_r_reg[17]/NET0131  ;
  assign n27230 = ~decrypt_pad & ~\u2_key_r_reg[24]/NET0131  ;
  assign n27231 = ~n27229 & ~n27230 ;
  assign n27232 = \u2_desIn_r_reg[45]/NET0131  & ~n27231 ;
  assign n27233 = ~\u2_desIn_r_reg[45]/NET0131  & n27231 ;
  assign n27234 = ~n27232 & ~n27233 ;
  assign n27257 = ~n27214 & n27220 ;
  assign n27258 = n27234 & n27257 ;
  assign n27259 = n27214 & ~n27227 ;
  assign n27260 = ~n27253 & ~n27259 ;
  assign n27261 = ~n27258 & n27260 ;
  assign n27262 = ~n27256 & ~n27261 ;
  assign n27228 = n27221 & n27227 ;
  assign n27235 = n27228 & n27234 ;
  assign n27236 = ~n27214 & ~n27234 ;
  assign n27237 = ~n27220 & n27236 ;
  assign n27238 = ~n27227 & n27237 ;
  assign n27239 = ~n27235 & ~n27238 ;
  assign n27266 = ~n27234 & n27259 ;
  assign n27267 = n27220 & n27266 ;
  assign n27240 = decrypt_pad & ~\u2_key_r_reg[33]/NET0131  ;
  assign n27241 = ~decrypt_pad & ~\u2_key_r_reg[40]/NET0131  ;
  assign n27242 = ~n27240 & ~n27241 ;
  assign n27243 = \u2_desIn_r_reg[61]/NET0131  & ~n27242 ;
  assign n27244 = ~\u2_desIn_r_reg[61]/NET0131  & n27242 ;
  assign n27245 = ~n27243 & ~n27244 ;
  assign n27263 = n27227 & n27253 ;
  assign n27264 = n27234 & n27263 ;
  assign n27265 = ~n27220 & n27264 ;
  assign n27268 = ~n27245 & ~n27265 ;
  assign n27269 = ~n27267 & n27268 ;
  assign n27270 = n27239 & n27269 ;
  assign n27271 = ~n27262 & n27270 ;
  assign n27282 = n27234 & n27247 ;
  assign n27275 = ~n27227 & ~n27253 ;
  assign n27276 = n27221 & n27275 ;
  assign n27277 = n27234 & n27276 ;
  assign n27272 = ~n27227 & n27253 ;
  assign n27273 = n27214 & ~n27220 ;
  assign n27274 = n27272 & n27273 ;
  assign n27289 = n27245 & ~n27274 ;
  assign n27290 = ~n27277 & n27289 ;
  assign n27291 = ~n27282 & n27290 ;
  assign n27278 = n27257 & n27263 ;
  assign n27279 = ~n27234 & n27273 ;
  assign n27280 = n27227 & n27279 ;
  assign n27281 = ~n27278 & ~n27280 ;
  assign n27283 = n27227 & ~n27234 ;
  assign n27284 = ~n27220 & n27283 ;
  assign n27285 = n27220 & ~n27234 ;
  assign n27286 = ~n27227 & n27285 ;
  assign n27287 = ~n27284 & ~n27286 ;
  assign n27288 = ~n27253 & ~n27287 ;
  assign n27292 = n27281 & ~n27288 ;
  assign n27293 = n27291 & n27292 ;
  assign n27294 = ~n27271 & ~n27293 ;
  assign n27297 = ~n27253 & n27280 ;
  assign n27295 = ~n27237 & ~n27258 ;
  assign n27296 = n27272 & ~n27295 ;
  assign n27298 = ~n27234 & n27278 ;
  assign n27299 = ~n27296 & ~n27298 ;
  assign n27300 = ~n27297 & n27299 ;
  assign n27301 = ~n27294 & n27300 ;
  assign n27302 = ~\u2_desIn_r_reg[26]/NET0131  & ~n27301 ;
  assign n27303 = \u2_desIn_r_reg[26]/NET0131  & n27301 ;
  assign n27304 = ~n27302 & ~n27303 ;
  assign n27323 = n27257 & ~n27283 ;
  assign n27324 = ~n27280 & ~n27323 ;
  assign n27325 = ~n27253 & ~n27324 ;
  assign n27306 = ~n27227 & n27234 ;
  assign n27319 = n27273 & n27306 ;
  assign n27320 = ~n27282 & ~n27319 ;
  assign n27321 = ~n27228 & ~n27267 ;
  assign n27322 = n27253 & ~n27321 ;
  assign n27326 = n27320 & ~n27322 ;
  assign n27327 = ~n27325 & n27326 ;
  assign n27328 = n27245 & ~n27327 ;
  assign n27305 = ~n27214 & ~n27227 ;
  assign n27307 = ~n27305 & ~n27306 ;
  assign n27308 = n27220 & ~n27307 ;
  assign n27309 = ~n27279 & ~n27308 ;
  assign n27310 = n27253 & ~n27309 ;
  assign n27313 = n27220 & n27283 ;
  assign n27311 = ~n27234 & ~n27253 ;
  assign n27312 = n27246 & n27311 ;
  assign n27314 = ~n27276 & ~n27312 ;
  assign n27315 = ~n27313 & n27314 ;
  assign n27316 = n27239 & n27315 ;
  assign n27317 = ~n27310 & n27316 ;
  assign n27318 = ~n27245 & ~n27317 ;
  assign n27329 = ~n27238 & n27320 ;
  assign n27330 = ~n27253 & ~n27329 ;
  assign n27331 = ~n27265 & ~n27298 ;
  assign n27332 = ~n27330 & n27331 ;
  assign n27333 = ~n27318 & n27332 ;
  assign n27334 = ~n27328 & n27333 ;
  assign n27335 = ~\u2_desIn_r_reg[12]/NET0131  & ~n27334 ;
  assign n27336 = \u2_desIn_r_reg[12]/NET0131  & n27334 ;
  assign n27337 = ~n27335 & ~n27336 ;
  assign n27344 = n26943 & n26956 ;
  assign n27345 = ~n26997 & ~n27344 ;
  assign n27346 = n26971 & ~n27345 ;
  assign n27343 = n26989 & n27004 ;
  assign n27347 = n26978 & ~n27343 ;
  assign n27348 = ~n26961 & n27347 ;
  assign n27338 = ~n26937 & n26943 ;
  assign n27339 = ~n26944 & ~n27338 ;
  assign n27340 = ~n26943 & n26971 ;
  assign n27341 = n26957 & ~n27340 ;
  assign n27342 = ~n27339 & n27341 ;
  assign n27349 = ~n27000 & ~n27342 ;
  assign n27350 = n27348 & n27349 ;
  assign n27351 = ~n27346 & n27350 ;
  assign n27353 = ~n26950 & ~n26956 ;
  assign n27357 = n27338 & n27353 ;
  assign n27352 = ~n26971 & n26990 ;
  assign n27363 = ~n26978 & ~n27352 ;
  assign n27364 = ~n27357 & n27363 ;
  assign n27354 = ~n26959 & ~n27004 ;
  assign n27355 = ~n27338 & ~n27353 ;
  assign n27356 = n27354 & n27355 ;
  assign n27365 = ~n26980 & ~n27356 ;
  assign n27358 = n26950 & n26956 ;
  assign n27359 = ~n26982 & ~n27358 ;
  assign n27360 = n26944 & ~n27359 ;
  assign n27361 = ~n26963 & ~n27004 ;
  assign n27362 = ~n26971 & ~n27361 ;
  assign n27366 = ~n27360 & ~n27362 ;
  assign n27367 = n27365 & n27366 ;
  assign n27368 = n27364 & n27367 ;
  assign n27369 = ~n27351 & ~n27368 ;
  assign n27370 = \u2_desIn_r_reg[28]/NET0131  & n27369 ;
  assign n27371 = ~\u2_desIn_r_reg[28]/NET0131  & ~n27369 ;
  assign n27372 = ~n27370 & ~n27371 ;
  assign n27431 = decrypt_pad & ~\u2_key_r_reg[16]/NET0131  ;
  assign n27432 = ~decrypt_pad & ~\u2_key_r_reg[23]/NET0131  ;
  assign n27433 = ~n27431 & ~n27432 ;
  assign n27434 = \u2_desIn_r_reg[27]/NET0131  & ~n27433 ;
  assign n27435 = ~\u2_desIn_r_reg[27]/NET0131  & n27433 ;
  assign n27436 = ~n27434 & ~n27435 ;
  assign n27386 = decrypt_pad & ~\u2_key_r_reg[14]/NET0131  ;
  assign n27387 = ~decrypt_pad & ~\u2_key_r_reg[21]/NET0131  ;
  assign n27388 = ~n27386 & ~n27387 ;
  assign n27389 = \u2_desIn_r_reg[11]/NET0131  & ~n27388 ;
  assign n27390 = ~\u2_desIn_r_reg[11]/NET0131  & n27388 ;
  assign n27391 = ~n27389 & ~n27390 ;
  assign n27406 = decrypt_pad & ~\u2_key_r_reg[1]/NET0131  ;
  assign n27407 = ~decrypt_pad & ~\u2_key_r_reg[8]/NET0131  ;
  assign n27408 = ~n27406 & ~n27407 ;
  assign n27409 = \u2_desIn_r_reg[19]/NET0131  & ~n27408 ;
  assign n27410 = ~\u2_desIn_r_reg[19]/NET0131  & n27408 ;
  assign n27411 = ~n27409 & ~n27410 ;
  assign n27373 = decrypt_pad & ~\u2_key_r_reg[45]/NET0131  ;
  assign n27374 = ~decrypt_pad & ~\u2_key_r_reg[52]/NET0131  ;
  assign n27375 = ~n27373 & ~n27374 ;
  assign n27376 = \u2_desIn_r_reg[35]/NET0131  & ~n27375 ;
  assign n27377 = ~\u2_desIn_r_reg[35]/NET0131  & n27375 ;
  assign n27378 = ~n27376 & ~n27377 ;
  assign n27379 = decrypt_pad & ~\u2_key_r_reg[29]/NET0131  ;
  assign n27380 = ~decrypt_pad & ~\u2_key_r_reg[36]/NET0131  ;
  assign n27381 = ~n27379 & ~n27380 ;
  assign n27382 = \u2_desIn_r_reg[61]/NET0131  & ~n27381 ;
  assign n27383 = ~\u2_desIn_r_reg[61]/NET0131  & n27381 ;
  assign n27384 = ~n27382 & ~n27383 ;
  assign n27394 = decrypt_pad & ~\u2_key_r_reg[51]/NET0131  ;
  assign n27395 = ~decrypt_pad & ~\u2_key_r_reg[31]/NET0131  ;
  assign n27396 = ~n27394 & ~n27395 ;
  assign n27397 = \u2_desIn_r_reg[3]/NET0131  & ~n27396 ;
  assign n27398 = ~\u2_desIn_r_reg[3]/NET0131  & n27396 ;
  assign n27399 = ~n27397 & ~n27398 ;
  assign n27413 = ~n27384 & ~n27399 ;
  assign n27414 = ~n27378 & n27413 ;
  assign n27452 = ~n27411 & n27414 ;
  assign n27449 = ~n27384 & n27399 ;
  assign n27450 = n27378 & n27449 ;
  assign n27451 = ~n27411 & n27450 ;
  assign n27422 = ~n27378 & n27399 ;
  assign n27441 = n27384 & n27422 ;
  assign n27400 = n27384 & ~n27399 ;
  assign n27448 = n27378 & n27400 ;
  assign n27453 = ~n27441 & ~n27448 ;
  assign n27454 = ~n27451 & n27453 ;
  assign n27455 = ~n27452 & n27454 ;
  assign n27456 = ~n27391 & ~n27455 ;
  assign n27401 = ~n27391 & n27399 ;
  assign n27412 = ~n27384 & n27401 ;
  assign n27438 = n27384 & n27391 ;
  assign n27439 = n27378 & ~n27438 ;
  assign n27440 = ~n27412 & n27439 ;
  assign n27442 = ~n27440 & ~n27441 ;
  assign n27443 = n27411 & ~n27442 ;
  assign n27404 = n27378 & n27384 ;
  assign n27420 = n27399 & n27404 ;
  assign n27444 = n27391 & ~n27411 ;
  assign n27445 = n27420 & n27444 ;
  assign n27385 = ~n27378 & n27384 ;
  assign n27446 = n27391 & ~n27399 ;
  assign n27447 = n27385 & n27446 ;
  assign n27457 = ~n27445 & ~n27447 ;
  assign n27458 = ~n27443 & n27457 ;
  assign n27459 = ~n27456 & n27458 ;
  assign n27460 = n27436 & ~n27459 ;
  assign n27392 = n27378 & ~n27391 ;
  assign n27393 = ~n27385 & ~n27392 ;
  assign n27402 = ~n27400 & ~n27401 ;
  assign n27403 = n27393 & ~n27402 ;
  assign n27405 = n27391 & n27404 ;
  assign n27415 = ~n27405 & n27411 ;
  assign n27416 = ~n27412 & ~n27414 ;
  assign n27417 = n27415 & n27416 ;
  assign n27424 = n27378 & n27413 ;
  assign n27423 = n27391 & n27422 ;
  assign n27425 = ~n27411 & ~n27423 ;
  assign n27426 = ~n27424 & n27425 ;
  assign n27418 = ~n27378 & n27400 ;
  assign n27419 = ~n27391 & n27418 ;
  assign n27421 = ~n27391 & n27420 ;
  assign n27427 = ~n27419 & ~n27421 ;
  assign n27428 = n27426 & n27427 ;
  assign n27429 = ~n27417 & ~n27428 ;
  assign n27430 = ~n27403 & ~n27429 ;
  assign n27437 = ~n27430 & ~n27436 ;
  assign n27461 = n27391 & n27414 ;
  assign n27462 = n27384 & ~n27391 ;
  assign n27463 = n27422 & n27462 ;
  assign n27464 = ~n27461 & ~n27463 ;
  assign n27465 = n27411 & ~n27464 ;
  assign n27466 = n27391 & n27424 ;
  assign n27467 = ~n27384 & n27423 ;
  assign n27468 = ~n27466 & ~n27467 ;
  assign n27469 = ~n27411 & ~n27468 ;
  assign n27470 = ~n27465 & ~n27469 ;
  assign n27471 = ~n27437 & n27470 ;
  assign n27472 = ~n27460 & n27471 ;
  assign n27473 = ~\u2_desIn_r_reg[44]/NET0131  & ~n27472 ;
  assign n27474 = \u2_desIn_r_reg[44]/NET0131  & n27472 ;
  assign n27475 = ~n27473 & ~n27474 ;
  assign n27482 = decrypt_pad & ~\u2_key_r_reg[21]/NET0131  ;
  assign n27483 = ~decrypt_pad & ~\u2_key_r_reg[28]/NET0131  ;
  assign n27484 = ~n27482 & ~n27483 ;
  assign n27485 = \u2_desIn_r_reg[7]/NET0131  & ~n27484 ;
  assign n27486 = ~\u2_desIn_r_reg[7]/NET0131  & n27484 ;
  assign n27487 = ~n27485 & ~n27486 ;
  assign n27501 = decrypt_pad & ~\u2_key_r_reg[37]/NET0131  ;
  assign n27502 = ~decrypt_pad & ~\u2_key_r_reg[44]/NET0131  ;
  assign n27503 = ~n27501 & ~n27502 ;
  assign n27504 = \u2_desIn_r_reg[41]/NET0131  & ~n27503 ;
  assign n27505 = ~\u2_desIn_r_reg[41]/NET0131  & n27503 ;
  assign n27506 = ~n27504 & ~n27505 ;
  assign n27488 = decrypt_pad & ~\u2_key_r_reg[9]/NET0131  ;
  assign n27489 = ~decrypt_pad & ~\u2_key_r_reg[16]/NET0131  ;
  assign n27490 = ~n27488 & ~n27489 ;
  assign n27491 = \u2_desIn_r_reg[25]/NET0131  & ~n27490 ;
  assign n27492 = ~\u2_desIn_r_reg[25]/NET0131  & n27490 ;
  assign n27493 = ~n27491 & ~n27492 ;
  assign n27495 = decrypt_pad & ~\u2_key_r_reg[36]/NET0131  ;
  assign n27496 = ~decrypt_pad & ~\u2_key_r_reg[43]/NET0131  ;
  assign n27497 = ~n27495 & ~n27496 ;
  assign n27498 = \u2_desIn_r_reg[33]/NET0131  & ~n27497 ;
  assign n27499 = ~\u2_desIn_r_reg[33]/NET0131  & n27497 ;
  assign n27500 = ~n27498 & ~n27499 ;
  assign n27514 = n27493 & ~n27500 ;
  assign n27535 = n27506 & n27514 ;
  assign n27476 = decrypt_pad & ~\u2_key_r_reg[49]/NET0131  ;
  assign n27477 = ~decrypt_pad & ~\u2_key_r_reg[1]/NET0131  ;
  assign n27478 = ~n27476 & ~n27477 ;
  assign n27479 = \u2_desIn_r_reg[49]/NET0131  & ~n27478 ;
  assign n27480 = ~\u2_desIn_r_reg[49]/NET0131  & n27478 ;
  assign n27481 = ~n27479 & ~n27480 ;
  assign n27536 = ~n27481 & n27506 ;
  assign n27537 = ~n27500 & n27536 ;
  assign n27538 = ~n27535 & ~n27537 ;
  assign n27539 = n27487 & ~n27538 ;
  assign n27528 = n27493 & ~n27506 ;
  assign n27529 = ~n27487 & n27506 ;
  assign n27530 = ~n27493 & n27529 ;
  assign n27531 = ~n27528 & ~n27530 ;
  assign n27532 = n27500 & ~n27531 ;
  assign n27515 = decrypt_pad & ~\u2_key_r_reg[0]/NET0131  ;
  assign n27516 = ~decrypt_pad & ~\u2_key_r_reg[7]/NET0131  ;
  assign n27517 = ~n27515 & ~n27516 ;
  assign n27518 = \u2_desIn_r_reg[57]/NET0131  & ~n27517 ;
  assign n27519 = ~\u2_desIn_r_reg[57]/NET0131  & n27517 ;
  assign n27520 = ~n27518 & ~n27519 ;
  assign n27509 = ~n27487 & ~n27493 ;
  assign n27533 = n27481 & ~n27500 ;
  assign n27534 = n27509 & n27533 ;
  assign n27540 = n27520 & ~n27534 ;
  assign n27541 = ~n27532 & n27540 ;
  assign n27542 = ~n27539 & n27541 ;
  assign n27545 = n27493 & n27500 ;
  assign n27507 = n27500 & ~n27506 ;
  assign n27546 = ~n27487 & n27507 ;
  assign n27547 = ~n27545 & ~n27546 ;
  assign n27494 = n27487 & ~n27493 ;
  assign n27548 = n27494 & ~n27500 ;
  assign n27549 = n27547 & ~n27548 ;
  assign n27550 = n27481 & ~n27549 ;
  assign n27510 = ~n27500 & ~n27506 ;
  assign n27543 = ~n27487 & n27493 ;
  assign n27544 = n27510 & n27543 ;
  assign n27551 = ~n27520 & ~n27544 ;
  assign n27552 = ~n27550 & n27551 ;
  assign n27553 = ~n27542 & ~n27552 ;
  assign n27511 = n27500 & n27506 ;
  assign n27512 = ~n27510 & ~n27511 ;
  assign n27513 = n27509 & ~n27512 ;
  assign n27508 = n27494 & n27507 ;
  assign n27521 = ~n27506 & n27520 ;
  assign n27522 = n27514 & ~n27521 ;
  assign n27523 = ~n27508 & ~n27522 ;
  assign n27524 = ~n27513 & n27523 ;
  assign n27525 = ~n27481 & ~n27524 ;
  assign n27526 = n27481 & n27494 ;
  assign n27527 = ~n27512 & n27526 ;
  assign n27554 = ~n27525 & ~n27527 ;
  assign n27555 = ~n27553 & n27554 ;
  assign n27556 = ~\u2_desIn_r_reg[52]/NET0131  & ~n27555 ;
  assign n27557 = \u2_desIn_r_reg[52]/NET0131  & n27555 ;
  assign n27558 = ~n27556 & ~n27557 ;
  assign n27563 = ~n27164 & ~n27178 ;
  assign n27578 = n27145 & ~n27563 ;
  assign n27575 = n27138 & n27152 ;
  assign n27576 = ~n27181 & ~n27189 ;
  assign n27577 = n27126 & ~n27576 ;
  assign n27579 = ~n27575 & ~n27577 ;
  assign n27580 = ~n27578 & n27579 ;
  assign n27581 = n27120 & ~n27580 ;
  assign n27564 = ~n27126 & ~n27563 ;
  assign n27559 = n27145 & n27157 ;
  assign n27560 = n27132 & ~n27188 ;
  assign n27561 = ~n27173 & ~n27560 ;
  assign n27562 = n27126 & ~n27561 ;
  assign n27565 = ~n27559 & ~n27562 ;
  assign n27566 = ~n27564 & n27565 ;
  assign n27567 = ~n27120 & ~n27566 ;
  assign n27570 = ~n27126 & n27132 ;
  assign n27571 = ~n27145 & n27180 ;
  assign n27572 = ~n27570 & ~n27571 ;
  assign n27568 = n27156 & n27177 ;
  assign n27569 = ~n27120 & ~n27568 ;
  assign n27573 = ~n27138 & ~n27569 ;
  assign n27574 = ~n27572 & n27573 ;
  assign n27582 = ~n27187 & ~n27574 ;
  assign n27583 = ~n27567 & n27582 ;
  assign n27584 = ~n27581 & n27583 ;
  assign n27585 = ~\u2_desIn_r_reg[18]/NET0131  & ~n27584 ;
  assign n27586 = \u2_desIn_r_reg[18]/NET0131  & n27584 ;
  assign n27587 = ~n27585 & ~n27586 ;
  assign n27604 = ~n27030 & ~n27089 ;
  assign n27605 = n27071 & n27089 ;
  assign n27606 = ~n27604 & ~n27605 ;
  assign n27607 = n27037 & ~n27606 ;
  assign n27608 = n27092 & ~n27604 ;
  assign n27603 = ~n27024 & n27086 ;
  assign n27609 = n27044 & n27050 ;
  assign n27610 = n27024 & n27609 ;
  assign n27611 = ~n27603 & ~n27610 ;
  assign n27612 = ~n27608 & n27611 ;
  assign n27613 = ~n27607 & n27612 ;
  assign n27614 = n27070 & ~n27613 ;
  assign n27588 = ~n27071 & ~n27081 ;
  assign n27589 = ~n27044 & ~n27588 ;
  assign n27590 = ~n27082 & ~n27589 ;
  assign n27591 = ~n27037 & ~n27590 ;
  assign n27592 = ~n27086 & ~n27095 ;
  assign n27593 = n27024 & ~n27592 ;
  assign n27594 = ~n27591 & ~n27593 ;
  assign n27595 = ~n27070 & ~n27594 ;
  assign n27596 = ~n27024 & n27060 ;
  assign n27597 = ~n27057 & ~n27596 ;
  assign n27598 = n27044 & ~n27597 ;
  assign n27599 = ~n27093 & ~n27103 ;
  assign n27600 = ~n27070 & ~n27599 ;
  assign n27601 = ~n27598 & ~n27600 ;
  assign n27602 = n27037 & ~n27601 ;
  assign n27615 = ~n27595 & ~n27602 ;
  assign n27616 = ~n27614 & n27615 ;
  assign n27617 = ~\u2_desIn_r_reg[2]/NET0131  & ~n27616 ;
  assign n27618 = \u2_desIn_r_reg[2]/NET0131  & n27616 ;
  assign n27619 = ~n27617 & ~n27618 ;
  assign n27635 = ~n27214 & ~n27284 ;
  assign n27634 = n27220 & n27234 ;
  assign n27636 = n27227 & ~n27253 ;
  assign n27637 = ~n27634 & n27636 ;
  assign n27638 = ~n27635 & n27637 ;
  assign n27639 = ~n27214 & ~n27285 ;
  assign n27640 = n27272 & ~n27639 ;
  assign n27620 = n27227 & n27258 ;
  assign n27641 = ~n27220 & n27306 ;
  assign n27642 = ~n27620 & ~n27641 ;
  assign n27643 = ~n27640 & n27642 ;
  assign n27644 = ~n27638 & n27643 ;
  assign n27645 = n27245 & ~n27644 ;
  assign n27622 = ~n27236 & ~n27259 ;
  assign n27623 = n27220 & ~n27622 ;
  assign n27624 = ~n27253 & ~n27623 ;
  assign n27625 = n27257 & n27306 ;
  assign n27626 = ~n27237 & n27253 ;
  assign n27627 = ~n27625 & n27626 ;
  assign n27628 = ~n27624 & ~n27627 ;
  assign n27629 = ~n27221 & ~n27246 ;
  assign n27630 = n27283 & n27629 ;
  assign n27631 = ~n27282 & ~n27630 ;
  assign n27632 = ~n27628 & n27631 ;
  assign n27633 = ~n27245 & ~n27632 ;
  assign n27646 = ~n27235 & n27320 ;
  assign n27647 = n27253 & ~n27646 ;
  assign n27621 = ~n27253 & n27620 ;
  assign n27648 = ~n27277 & ~n27621 ;
  assign n27649 = ~n27647 & n27648 ;
  assign n27650 = ~n27633 & n27649 ;
  assign n27651 = ~n27645 & n27650 ;
  assign n27652 = ~\u2_desIn_r_reg[6]/NET0131  & ~n27651 ;
  assign n27653 = \u2_desIn_r_reg[6]/NET0131  & n27651 ;
  assign n27654 = ~n27652 & ~n27653 ;
  assign n27657 = ~n27481 & n27500 ;
  assign n27662 = n27509 & n27657 ;
  assign n27661 = n27514 & n27529 ;
  assign n27671 = ~n27520 & ~n27661 ;
  assign n27672 = ~n27662 & n27671 ;
  assign n27655 = ~n27493 & n27510 ;
  assign n27663 = ~n27487 & n27655 ;
  assign n27658 = n27487 & n27493 ;
  assign n27659 = ~n27506 & n27658 ;
  assign n27664 = ~n27533 & n27659 ;
  assign n27673 = ~n27663 & ~n27664 ;
  assign n27674 = n27672 & n27673 ;
  assign n27665 = ~n27487 & n27545 ;
  assign n27666 = ~n27535 & ~n27665 ;
  assign n27667 = n27481 & ~n27666 ;
  assign n27668 = n27487 & n27536 ;
  assign n27669 = ~n27511 & ~n27668 ;
  assign n27670 = ~n27493 & ~n27669 ;
  assign n27675 = ~n27667 & ~n27670 ;
  assign n27676 = n27674 & n27675 ;
  assign n27678 = ~n27535 & ~n27543 ;
  assign n27679 = ~n27529 & ~n27678 ;
  assign n27680 = ~n27481 & ~n27679 ;
  assign n27681 = n27487 & n27510 ;
  assign n27685 = n27481 & ~n27681 ;
  assign n27682 = n27487 & n27500 ;
  assign n27683 = ~n27493 & n27682 ;
  assign n27684 = n27493 & n27511 ;
  assign n27686 = ~n27683 & ~n27684 ;
  assign n27687 = n27685 & n27686 ;
  assign n27688 = ~n27680 & ~n27687 ;
  assign n27689 = ~n27487 & ~n27500 ;
  assign n27690 = ~n27543 & ~n27689 ;
  assign n27691 = n27506 & ~n27514 ;
  assign n27692 = ~n27690 & n27691 ;
  assign n27677 = n27487 & n27655 ;
  assign n27693 = n27520 & ~n27677 ;
  assign n27694 = ~n27692 & n27693 ;
  assign n27695 = ~n27688 & n27694 ;
  assign n27696 = ~n27676 & ~n27695 ;
  assign n27656 = n27481 & n27655 ;
  assign n27660 = n27657 & n27659 ;
  assign n27697 = ~n27656 & ~n27660 ;
  assign n27698 = ~n27696 & n27697 ;
  assign n27699 = ~\u2_desIn_r_reg[34]/NET0131  & ~n27698 ;
  assign n27700 = \u2_desIn_r_reg[34]/NET0131  & n27698 ;
  assign n27701 = ~n27699 & ~n27700 ;
  assign n27703 = n27227 & ~n27295 ;
  assign n27702 = n27234 & n27273 ;
  assign n27704 = ~n27254 & ~n27702 ;
  assign n27705 = ~n27703 & n27704 ;
  assign n27706 = ~n27275 & ~n27705 ;
  assign n27707 = ~n27246 & ~n27266 ;
  assign n27708 = ~n27253 & ~n27285 ;
  assign n27709 = ~n27707 & n27708 ;
  assign n27710 = n27245 & ~n27709 ;
  assign n27711 = ~n27706 & n27710 ;
  assign n27712 = ~n27305 & ~n27641 ;
  assign n27713 = ~n27253 & ~n27712 ;
  assign n27714 = n27264 & ~n27273 ;
  assign n27715 = ~n27245 & ~n27286 ;
  assign n27716 = ~n27714 & n27715 ;
  assign n27717 = n27281 & n27716 ;
  assign n27718 = ~n27713 & n27717 ;
  assign n27719 = ~n27711 & ~n27718 ;
  assign n27720 = ~n27227 & n27257 ;
  assign n27721 = ~n27228 & ~n27247 ;
  assign n27722 = ~n27720 & n27721 ;
  assign n27723 = n27311 & ~n27722 ;
  assign n27724 = n27214 & n27253 ;
  assign n27725 = ~n27287 & n27724 ;
  assign n27726 = ~n27723 & ~n27725 ;
  assign n27727 = ~n27719 & n27726 ;
  assign n27728 = ~\u2_desIn_r_reg[8]/NET0131  & ~n27727 ;
  assign n27729 = \u2_desIn_r_reg[8]/NET0131  & n27727 ;
  assign n27730 = ~n27728 & ~n27729 ;
  assign n27768 = decrypt_pad & ~\u2_key_r_reg[32]/NET0131  ;
  assign n27769 = ~decrypt_pad & ~\u2_key_r_reg[39]/P0001  ;
  assign n27770 = ~n27768 & ~n27769 ;
  assign n27771 = \u2_desIn_r_reg[63]/NET0131  & ~n27770 ;
  assign n27772 = ~\u2_desIn_r_reg[63]/NET0131  & n27770 ;
  assign n27773 = ~n27771 & ~n27772 ;
  assign n27761 = decrypt_pad & ~\u2_key_r_reg[41]/NET0131  ;
  assign n27762 = ~decrypt_pad & ~\u2_key_r_reg[48]/NET0131  ;
  assign n27763 = ~n27761 & ~n27762 ;
  assign n27764 = \u2_desIn_r_reg[55]/NET0131  & ~n27763 ;
  assign n27765 = ~\u2_desIn_r_reg[55]/NET0131  & n27763 ;
  assign n27766 = ~n27764 & ~n27765 ;
  assign n27737 = decrypt_pad & ~\u2_key_r_reg[47]/NET0131  ;
  assign n27738 = ~decrypt_pad & ~\u2_key_r_reg[54]/NET0131  ;
  assign n27739 = ~n27737 & ~n27738 ;
  assign n27740 = \u2_desIn_r_reg[47]/NET0131  & ~n27739 ;
  assign n27741 = ~\u2_desIn_r_reg[47]/NET0131  & n27739 ;
  assign n27742 = ~n27740 & ~n27741 ;
  assign n27744 = decrypt_pad & ~\u2_key_r_reg[20]/NET0131  ;
  assign n27745 = ~decrypt_pad & ~\u2_key_r_reg[27]/NET0131  ;
  assign n27746 = ~n27744 & ~n27745 ;
  assign n27747 = \u2_desIn_r_reg[31]/NET0131  & ~n27746 ;
  assign n27748 = ~\u2_desIn_r_reg[31]/NET0131  & n27746 ;
  assign n27749 = ~n27747 & ~n27748 ;
  assign n27751 = decrypt_pad & ~\u2_key_r_reg[12]/NET0131  ;
  assign n27752 = ~decrypt_pad & ~\u2_key_r_reg[19]/NET0131  ;
  assign n27753 = ~n27751 & ~n27752 ;
  assign n27754 = \u2_desIn_r_reg[5]/NET0131  & ~n27753 ;
  assign n27755 = ~\u2_desIn_r_reg[5]/NET0131  & n27753 ;
  assign n27756 = ~n27754 & ~n27755 ;
  assign n27778 = n27749 & ~n27756 ;
  assign n27803 = ~n27742 & n27778 ;
  assign n27731 = decrypt_pad & ~\u2_key_r_reg[24]/NET0131  ;
  assign n27732 = ~decrypt_pad & ~\u2_key_r_reg[6]/NET0131  ;
  assign n27733 = ~n27731 & ~n27732 ;
  assign n27734 = \u2_desIn_r_reg[39]/NET0131  & ~n27733 ;
  assign n27735 = ~\u2_desIn_r_reg[39]/NET0131  & n27733 ;
  assign n27736 = ~n27734 & ~n27735 ;
  assign n27801 = n27736 & n27749 ;
  assign n27774 = ~n27749 & n27756 ;
  assign n27802 = ~n27736 & n27774 ;
  assign n27804 = ~n27801 & ~n27802 ;
  assign n27805 = ~n27803 & n27804 ;
  assign n27806 = ~n27766 & ~n27805 ;
  assign n27785 = ~n27749 & ~n27756 ;
  assign n27786 = ~n27742 & n27785 ;
  assign n27787 = n27736 & n27774 ;
  assign n27788 = ~n27786 & ~n27787 ;
  assign n27807 = n27766 & ~n27788 ;
  assign n27757 = n27736 & ~n27756 ;
  assign n27758 = n27749 & n27757 ;
  assign n27759 = n27742 & n27758 ;
  assign n27798 = ~n27736 & ~n27778 ;
  assign n27799 = n27742 & ~n27774 ;
  assign n27800 = n27798 & n27799 ;
  assign n27808 = ~n27759 & ~n27800 ;
  assign n27809 = ~n27807 & n27808 ;
  assign n27810 = ~n27806 & n27809 ;
  assign n27811 = ~n27773 & ~n27810 ;
  assign n27743 = ~n27736 & n27742 ;
  assign n27750 = n27743 & ~n27749 ;
  assign n27760 = ~n27750 & ~n27759 ;
  assign n27767 = ~n27760 & ~n27766 ;
  assign n27776 = ~n27749 & n27757 ;
  assign n27777 = n27742 & n27776 ;
  assign n27779 = ~n27736 & n27778 ;
  assign n27780 = n27749 & n27756 ;
  assign n27781 = n27736 & n27780 ;
  assign n27782 = ~n27779 & ~n27781 ;
  assign n27783 = ~n27777 & n27782 ;
  assign n27784 = n27766 & ~n27783 ;
  assign n27789 = ~n27766 & ~n27788 ;
  assign n27775 = n27743 & n27774 ;
  assign n27790 = ~n27736 & n27756 ;
  assign n27791 = ~n27766 & ~n27790 ;
  assign n27792 = ~n27742 & n27749 ;
  assign n27793 = ~n27791 & n27792 ;
  assign n27794 = ~n27775 & ~n27793 ;
  assign n27795 = ~n27789 & n27794 ;
  assign n27796 = ~n27784 & n27795 ;
  assign n27797 = n27773 & ~n27796 ;
  assign n27812 = ~n27767 & ~n27797 ;
  assign n27813 = ~n27811 & n27812 ;
  assign n27814 = ~\u2_desIn_r_reg[24]/NET0131  & ~n27813 ;
  assign n27815 = \u2_desIn_r_reg[24]/NET0131  & n27813 ;
  assign n27816 = ~n27814 & ~n27815 ;
  assign n27836 = n27139 & ~n27151 ;
  assign n27837 = ~n27157 & ~n27836 ;
  assign n27838 = n27145 & ~n27154 ;
  assign n27839 = ~n27151 & ~n27188 ;
  assign n27840 = ~n27838 & n27839 ;
  assign n27841 = n27837 & ~n27840 ;
  assign n27842 = n27126 & ~n27841 ;
  assign n27817 = n27145 & n27184 ;
  assign n27822 = ~n27154 & ~n27156 ;
  assign n27823 = ~n27145 & ~n27822 ;
  assign n27834 = ~n27817 & ~n27823 ;
  assign n27835 = ~n27126 & ~n27834 ;
  assign n27843 = n27145 & n27181 ;
  assign n27844 = ~n27835 & ~n27843 ;
  assign n27845 = ~n27842 & n27844 ;
  assign n27846 = ~n27120 & ~n27845 ;
  assign n27818 = n27138 & n27191 ;
  assign n27819 = ~n27164 & ~n27818 ;
  assign n27820 = ~n27817 & n27819 ;
  assign n27821 = n27126 & ~n27820 ;
  assign n27826 = n27145 & ~n27156 ;
  assign n27827 = ~n27172 & n27826 ;
  assign n27824 = ~n27138 & ~n27152 ;
  assign n27825 = n27126 & ~n27824 ;
  assign n27828 = ~n27823 & ~n27825 ;
  assign n27829 = ~n27827 & n27828 ;
  assign n27830 = ~n27821 & ~n27829 ;
  assign n27831 = n27120 & ~n27830 ;
  assign n27832 = n27126 & ~n27145 ;
  assign n27833 = n27163 & n27832 ;
  assign n27847 = ~n27153 & ~n27833 ;
  assign n27848 = ~n27831 & n27847 ;
  assign n27849 = ~n27846 & n27848 ;
  assign n27850 = \u2_desIn_r_reg[32]/NET0131  & ~n27849 ;
  assign n27851 = ~\u2_desIn_r_reg[32]/NET0131  & n27849 ;
  assign n27852 = ~n27850 & ~n27851 ;
  assign n27885 = ~n27757 & ~n27802 ;
  assign n27886 = ~n27742 & ~n27885 ;
  assign n27876 = n27742 & n27787 ;
  assign n27877 = ~n27736 & ~n27742 ;
  assign n27878 = n27756 & ~n27766 ;
  assign n27879 = n27877 & n27878 ;
  assign n27880 = ~n27876 & ~n27879 ;
  assign n27860 = n27742 & n27749 ;
  assign n27881 = ~n27790 & ~n27860 ;
  assign n27882 = ~n27736 & n27780 ;
  assign n27883 = ~n27766 & ~n27882 ;
  assign n27884 = ~n27881 & n27883 ;
  assign n27887 = n27880 & ~n27884 ;
  assign n27888 = ~n27886 & n27887 ;
  assign n27889 = ~n27773 & ~n27888 ;
  assign n27853 = ~n27742 & ~n27782 ;
  assign n27854 = n27736 & ~n27742 ;
  assign n27855 = ~n27801 & ~n27854 ;
  assign n27856 = n27766 & ~n27855 ;
  assign n27857 = ~n27853 & ~n27856 ;
  assign n27858 = n27773 & ~n27857 ;
  assign n27863 = n27743 & ~n27756 ;
  assign n27864 = ~n27749 & n27863 ;
  assign n27861 = n27790 & n27860 ;
  assign n27862 = ~n27773 & n27861 ;
  assign n27859 = ~n27742 & n27801 ;
  assign n27865 = n27766 & ~n27859 ;
  assign n27866 = ~n27862 & n27865 ;
  assign n27867 = ~n27864 & n27866 ;
  assign n27868 = n27785 & ~n27854 ;
  assign n27869 = ~n27861 & ~n27868 ;
  assign n27870 = n27773 & ~n27869 ;
  assign n27871 = ~n27743 & ~n27854 ;
  assign n27872 = n27774 & n27871 ;
  assign n27873 = ~n27766 & ~n27872 ;
  assign n27874 = ~n27870 & n27873 ;
  assign n27875 = ~n27867 & ~n27874 ;
  assign n27890 = ~n27858 & ~n27875 ;
  assign n27891 = ~n27889 & n27890 ;
  assign n27892 = \u2_desIn_r_reg[14]/NET0131  & n27891 ;
  assign n27893 = ~\u2_desIn_r_reg[14]/NET0131  & ~n27891 ;
  assign n27894 = ~n27892 & ~n27893 ;
  assign n27896 = ~n27378 & ~n27401 ;
  assign n27897 = ~n27438 & n27896 ;
  assign n27898 = ~n27413 & ~n27420 ;
  assign n27899 = ~n27897 & n27898 ;
  assign n27900 = n27411 & ~n27899 ;
  assign n27901 = ~n27412 & ~n27448 ;
  assign n27902 = ~n27411 & ~n27901 ;
  assign n27895 = n27392 & n27399 ;
  assign n27903 = n27391 & n27441 ;
  assign n27904 = ~n27895 & ~n27903 ;
  assign n27905 = ~n27902 & n27904 ;
  assign n27906 = ~n27900 & n27905 ;
  assign n27907 = n27436 & ~n27906 ;
  assign n27918 = ~n27461 & ~n27903 ;
  assign n27919 = ~n27384 & n27392 ;
  assign n27920 = ~n27399 & n27919 ;
  assign n27921 = n27918 & ~n27920 ;
  assign n27922 = n27411 & ~n27921 ;
  assign n27908 = n27391 & n27449 ;
  assign n27909 = ~n27418 & ~n27908 ;
  assign n27910 = ~n27378 & n27411 ;
  assign n27911 = ~n27909 & ~n27910 ;
  assign n27913 = n27411 & ~n27422 ;
  assign n27912 = ~n27411 & ~n27413 ;
  assign n27914 = ~n27391 & ~n27912 ;
  assign n27915 = ~n27913 & n27914 ;
  assign n27916 = ~n27911 & ~n27915 ;
  assign n27917 = ~n27436 & ~n27916 ;
  assign n27923 = n27400 & n27444 ;
  assign n27924 = ~n27421 & ~n27923 ;
  assign n27925 = ~n27917 & n27924 ;
  assign n27926 = ~n27922 & n27925 ;
  assign n27927 = ~n27907 & n27926 ;
  assign n27928 = ~\u2_desIn_r_reg[0]/NET0131  & ~n27927 ;
  assign n27929 = \u2_desIn_r_reg[0]/NET0131  & n27927 ;
  assign n27930 = ~n27928 & ~n27929 ;
  assign n27945 = n27145 & n27163 ;
  assign n27944 = n27156 & n27832 ;
  assign n27946 = n27120 & ~n27944 ;
  assign n27947 = ~n27945 & n27946 ;
  assign n27948 = ~n27174 & n27947 ;
  assign n27949 = ~n27184 & ~n27571 ;
  assign n27950 = ~n27198 & n27949 ;
  assign n27951 = n27126 & ~n27950 ;
  assign n27952 = ~n27153 & n27569 ;
  assign n27953 = ~n27951 & n27952 ;
  assign n27954 = ~n27948 & ~n27953 ;
  assign n27932 = ~n27173 & ~n27843 ;
  assign n27933 = ~n27120 & ~n27932 ;
  assign n27931 = ~n27145 & n27172 ;
  assign n27934 = ~n27191 & ~n27575 ;
  assign n27935 = n27120 & ~n27934 ;
  assign n27936 = ~n27931 & ~n27935 ;
  assign n27937 = ~n27933 & n27936 ;
  assign n27938 = ~n27126 & ~n27937 ;
  assign n27941 = ~n27126 & n27837 ;
  assign n27939 = n27126 & ~n27184 ;
  assign n27940 = n27563 & n27939 ;
  assign n27942 = n27145 & ~n27940 ;
  assign n27943 = ~n27941 & n27942 ;
  assign n27955 = ~n27938 & ~n27943 ;
  assign n27956 = ~n27954 & n27955 ;
  assign n27957 = ~\u2_desIn_r_reg[30]/NET0131  & ~n27956 ;
  assign n27958 = \u2_desIn_r_reg[30]/NET0131  & n27956 ;
  assign n27959 = ~n27957 & ~n27958 ;
  assign n27979 = n27481 & ~n27548 ;
  assign n27980 = ~n27661 & n27979 ;
  assign n27981 = ~n27481 & ~n27682 ;
  assign n27982 = n27531 & n27981 ;
  assign n27983 = ~n27980 & ~n27982 ;
  assign n27962 = n27507 & n27543 ;
  assign n27984 = n27511 & n27658 ;
  assign n27985 = ~n27962 & ~n27984 ;
  assign n27986 = ~n27983 & n27985 ;
  assign n27987 = ~n27520 & ~n27986 ;
  assign n27960 = ~n27487 & n27500 ;
  assign n27961 = ~n27528 & ~n27960 ;
  assign n27963 = ~n27961 & ~n27962 ;
  assign n27964 = n27481 & ~n27963 ;
  assign n27965 = ~n27481 & ~n27655 ;
  assign n27966 = ~n27964 & ~n27965 ;
  assign n27967 = n27506 & n27683 ;
  assign n27968 = ~n27966 & ~n27967 ;
  assign n27969 = n27520 & ~n27968 ;
  assign n27975 = n27506 & n27548 ;
  assign n27973 = ~n27507 & ~n27543 ;
  assign n27974 = ~n27961 & n27973 ;
  assign n27976 = ~n27663 & ~n27974 ;
  assign n27977 = ~n27975 & n27976 ;
  assign n27978 = n27481 & ~n27977 ;
  assign n27970 = n27493 & n27520 ;
  assign n27971 = n27537 & n27970 ;
  assign n27972 = ~n27481 & n27962 ;
  assign n27988 = ~n27971 & ~n27972 ;
  assign n27989 = ~n27978 & n27988 ;
  assign n27990 = ~n27969 & n27989 ;
  assign n27991 = ~n27987 & n27990 ;
  assign n27992 = \u2_desIn_r_reg[38]/NET0131  & ~n27991 ;
  assign n27993 = ~\u2_desIn_r_reg[38]/NET0131  & n27991 ;
  assign n27994 = ~n27992 & ~n27993 ;
  assign n27996 = ~n27863 & n27883 ;
  assign n27998 = ~n27756 & n27877 ;
  assign n27997 = n27742 & n27774 ;
  assign n27999 = n27766 & ~n27997 ;
  assign n28000 = ~n27998 & n27999 ;
  assign n28001 = ~n27996 & ~n28000 ;
  assign n27995 = n27736 & n27786 ;
  assign n28002 = n27773 & ~n27995 ;
  assign n28003 = n27880 & n28002 ;
  assign n28004 = ~n28001 & n28003 ;
  assign n28006 = n27774 & ~n27871 ;
  assign n28005 = n27778 & n27877 ;
  assign n28007 = ~n27766 & ~n27773 ;
  assign n28008 = ~n27776 & n28007 ;
  assign n28009 = ~n28005 & n28008 ;
  assign n28010 = ~n28006 & n28009 ;
  assign n28011 = ~n28004 & ~n28010 ;
  assign n28012 = ~n27742 & n27780 ;
  assign n28013 = n27736 & n28012 ;
  assign n28014 = ~n27759 & ~n28013 ;
  assign n28015 = ~n28011 & n28014 ;
  assign n28016 = ~n27758 & ~n27774 ;
  assign n28017 = ~n27798 & n28016 ;
  assign n28018 = ~n27742 & ~n28017 ;
  assign n28019 = ~n27757 & n27799 ;
  assign n28020 = n27766 & ~n27773 ;
  assign n28021 = ~n28019 & n28020 ;
  assign n28022 = ~n28018 & n28021 ;
  assign n28023 = ~n28015 & ~n28022 ;
  assign n28024 = ~\u2_desIn_r_reg[36]/NET0131  & ~n28023 ;
  assign n28025 = \u2_desIn_r_reg[36]/NET0131  & n28023 ;
  assign n28026 = ~n28024 & ~n28025 ;
  assign n28048 = n27044 & n27060 ;
  assign n28049 = ~n27087 & ~n28048 ;
  assign n28050 = n27037 & ~n28049 ;
  assign n28051 = ~n27052 & ~n27605 ;
  assign n28052 = ~n28050 & n28051 ;
  assign n28053 = n27070 & ~n28052 ;
  assign n28031 = ~n27070 & ~n27103 ;
  assign n28032 = n27024 & ~n27599 ;
  assign n28033 = ~n28031 & n28032 ;
  assign n28027 = n27044 & n27081 ;
  assign n28028 = ~n27095 & ~n28027 ;
  assign n28029 = n27070 & ~n28028 ;
  assign n28030 = ~n27024 & ~n27592 ;
  assign n28034 = ~n28029 & ~n28030 ;
  assign n28035 = ~n28033 & n28034 ;
  assign n28036 = ~n27037 & ~n28035 ;
  assign n28037 = ~n27053 & ~n28027 ;
  assign n28038 = n27054 & ~n28037 ;
  assign n28039 = ~n27050 & n27089 ;
  assign n28043 = ~n27610 & ~n28039 ;
  assign n28044 = ~n27080 & n28043 ;
  assign n28040 = n27037 & n28027 ;
  assign n28041 = ~n27051 & n27063 ;
  assign n28042 = ~n27089 & n28041 ;
  assign n28045 = ~n28040 & ~n28042 ;
  assign n28046 = n28044 & n28045 ;
  assign n28047 = ~n27070 & ~n28046 ;
  assign n28054 = ~n28038 & ~n28047 ;
  assign n28055 = ~n28036 & n28054 ;
  assign n28056 = ~n28053 & n28055 ;
  assign n28057 = \u2_desIn_r_reg[50]/NET0131  & ~n28056 ;
  assign n28058 = ~\u2_desIn_r_reg[50]/NET0131  & n28056 ;
  assign n28059 = ~n28057 & ~n28058 ;
  assign n28082 = n26950 & n27338 ;
  assign n28083 = ~n26979 & ~n27005 ;
  assign n28084 = ~n28082 & n28083 ;
  assign n28085 = n26971 & ~n28084 ;
  assign n28076 = n27338 & n27358 ;
  assign n28078 = n27339 & n27361 ;
  assign n28079 = ~n27353 & ~n28078 ;
  assign n28077 = n27339 & n27353 ;
  assign n28080 = ~n26971 & ~n28077 ;
  assign n28081 = ~n28079 & n28080 ;
  assign n28086 = ~n28076 & ~n28081 ;
  assign n28087 = ~n28085 & n28086 ;
  assign n28088 = n26978 & ~n28087 ;
  assign n28060 = ~n26958 & n26971 ;
  assign n28061 = n26943 & n27005 ;
  assign n28062 = ~n26960 & ~n26971 ;
  assign n28063 = ~n28061 & n28062 ;
  assign n28064 = ~n28060 & ~n28063 ;
  assign n28065 = ~n26950 & n27338 ;
  assign n28066 = ~n26999 & ~n28065 ;
  assign n28067 = n26971 & ~n28066 ;
  assign n28072 = n26962 & ~n28067 ;
  assign n28068 = n26937 & n26990 ;
  assign n28069 = ~n28065 & ~n28068 ;
  assign n28070 = n26956 & ~n28069 ;
  assign n28071 = n27362 & ~n28065 ;
  assign n28073 = ~n28070 & ~n28071 ;
  assign n28074 = n28072 & n28073 ;
  assign n28075 = ~n26978 & ~n28074 ;
  assign n28089 = ~n28064 & ~n28075 ;
  assign n28090 = ~n28088 & n28089 ;
  assign n28091 = \u2_desIn_r_reg[56]/NET0131  & n28090 ;
  assign n28092 = ~\u2_desIn_r_reg[56]/NET0131  & ~n28090 ;
  assign n28093 = ~n28091 & ~n28092 ;
  assign n28127 = decrypt_pad & ~\u2_key_r_reg[10]/NET0131  ;
  assign n28128 = ~decrypt_pad & ~\u2_key_r_reg[17]/NET0131  ;
  assign n28129 = ~n28127 & ~n28128 ;
  assign n28130 = \u2_desIn_r_reg[29]/NET0131  & ~n28129 ;
  assign n28131 = ~\u2_desIn_r_reg[29]/NET0131  & n28129 ;
  assign n28132 = ~n28130 & ~n28131 ;
  assign n28094 = decrypt_pad & ~\u2_key_r_reg[55]/NET0131  ;
  assign n28095 = ~decrypt_pad & ~\u2_key_r_reg[5]/NET0131  ;
  assign n28096 = ~n28094 & ~n28095 ;
  assign n28097 = \u2_desIn_r_reg[37]/NET0131  & ~n28096 ;
  assign n28098 = ~\u2_desIn_r_reg[37]/NET0131  & n28096 ;
  assign n28099 = ~n28097 & ~n28098 ;
  assign n28107 = decrypt_pad & ~\u2_key_r_reg[46]/NET0131  ;
  assign n28108 = ~decrypt_pad & ~\u2_key_r_reg[53]/NET0131  ;
  assign n28109 = ~n28107 & ~n28108 ;
  assign n28110 = \u2_desIn_r_reg[63]/NET0131  & ~n28109 ;
  assign n28111 = ~\u2_desIn_r_reg[63]/NET0131  & n28109 ;
  assign n28112 = ~n28110 & ~n28111 ;
  assign n28114 = ~n28099 & ~n28112 ;
  assign n28115 = n28099 & n28112 ;
  assign n28116 = ~n28114 & ~n28115 ;
  assign n28100 = decrypt_pad & ~\u2_key_r_reg[18]/NET0131  ;
  assign n28101 = ~decrypt_pad & ~\u2_key_r_reg[25]/NET0131  ;
  assign n28102 = ~n28100 & ~n28101 ;
  assign n28103 = \u2_desIn_r_reg[5]/NET0131  & ~n28102 ;
  assign n28104 = ~\u2_desIn_r_reg[5]/NET0131  & n28102 ;
  assign n28105 = ~n28103 & ~n28104 ;
  assign n28117 = decrypt_pad & ~\u2_key_r_reg[26]/NET0131  ;
  assign n28118 = ~decrypt_pad & ~\u2_key_r_reg[33]/NET0131  ;
  assign n28119 = ~n28117 & ~n28118 ;
  assign n28120 = \u2_desIn_r_reg[13]/NET0131  & ~n28119 ;
  assign n28121 = ~\u2_desIn_r_reg[13]/NET0131  & n28119 ;
  assign n28122 = ~n28120 & ~n28121 ;
  assign n28168 = ~n28105 & n28122 ;
  assign n28169 = ~n28116 & n28168 ;
  assign n28157 = n28099 & ~n28112 ;
  assign n28158 = n28105 & n28157 ;
  assign n28139 = decrypt_pad & ~\u2_key_r_reg[27]/NET0131  ;
  assign n28140 = ~decrypt_pad & ~\u2_key_r_reg[34]/NET0131  ;
  assign n28141 = ~n28139 & ~n28140 ;
  assign n28142 = \u2_desIn_r_reg[21]/NET0131  & ~n28141 ;
  assign n28143 = ~\u2_desIn_r_reg[21]/NET0131  & n28141 ;
  assign n28144 = ~n28142 & ~n28143 ;
  assign n28159 = n28122 & ~n28144 ;
  assign n28160 = n28158 & n28159 ;
  assign n28165 = ~n28099 & n28105 ;
  assign n28166 = n28122 & n28165 ;
  assign n28167 = n28112 & n28166 ;
  assign n28170 = ~n28160 & ~n28167 ;
  assign n28171 = ~n28169 & n28170 ;
  assign n28150 = n28105 & ~n28122 ;
  assign n28161 = n28099 & n28144 ;
  assign n28162 = n28116 & ~n28161 ;
  assign n28163 = n28150 & ~n28162 ;
  assign n28134 = ~n28105 & ~n28122 ;
  assign n28164 = n28134 & n28162 ;
  assign n28172 = ~n28163 & ~n28164 ;
  assign n28173 = n28171 & n28172 ;
  assign n28174 = ~n28132 & ~n28173 ;
  assign n28106 = n28099 & ~n28105 ;
  assign n28113 = ~n28105 & n28112 ;
  assign n28123 = ~n28112 & ~n28122 ;
  assign n28124 = ~n28113 & ~n28123 ;
  assign n28125 = n28116 & n28124 ;
  assign n28126 = ~n28106 & ~n28125 ;
  assign n28133 = ~n28126 & n28132 ;
  assign n28135 = n28114 & n28134 ;
  assign n28136 = n28106 & n28122 ;
  assign n28137 = ~n28135 & ~n28136 ;
  assign n28138 = ~n28133 & n28137 ;
  assign n28145 = ~n28138 & n28144 ;
  assign n28146 = n28122 & n28132 ;
  assign n28147 = n28105 & n28114 ;
  assign n28148 = n28146 & n28147 ;
  assign n28149 = n28132 & ~n28144 ;
  assign n28151 = n28099 & n28150 ;
  assign n28152 = ~n28099 & n28113 ;
  assign n28153 = n28105 & n28115 ;
  assign n28154 = ~n28152 & ~n28153 ;
  assign n28155 = ~n28151 & n28154 ;
  assign n28156 = n28149 & ~n28155 ;
  assign n28175 = ~n28148 & ~n28156 ;
  assign n28176 = ~n28145 & n28175 ;
  assign n28177 = ~n28174 & n28176 ;
  assign n28178 = ~\u2_desIn_r_reg[46]/NET0131  & ~n28177 ;
  assign n28179 = \u2_desIn_r_reg[46]/NET0131  & n28177 ;
  assign n28180 = ~n28178 & ~n28179 ;
  assign n28181 = n26956 & ~n27339 ;
  assign n28182 = ~n26999 & ~n28181 ;
  assign n28183 = n26950 & ~n28182 ;
  assign n28184 = ~n26950 & ~n26963 ;
  assign n28185 = n27339 & n28184 ;
  assign n28186 = n26971 & ~n28185 ;
  assign n28187 = ~n26956 & n26989 ;
  assign n28188 = ~n28082 & ~n28187 ;
  assign n28189 = n28062 & n28188 ;
  assign n28190 = ~n28181 & n28189 ;
  assign n28191 = ~n28186 & ~n28190 ;
  assign n28192 = ~n28183 & ~n28191 ;
  assign n28193 = n26978 & ~n28192 ;
  assign n28201 = n26978 & ~n26980 ;
  assign n28199 = n26950 & ~n26998 ;
  assign n28200 = n27339 & ~n28199 ;
  assign n28198 = ~n27339 & n27358 ;
  assign n28202 = n26971 & ~n28198 ;
  assign n28203 = ~n28200 & n28202 ;
  assign n28204 = ~n28201 & n28203 ;
  assign n28194 = ~n26971 & n28183 ;
  assign n28195 = ~n26971 & n28185 ;
  assign n28196 = ~n26980 & ~n28195 ;
  assign n28197 = ~n26978 & ~n28196 ;
  assign n28205 = ~n28194 & ~n28197 ;
  assign n28206 = ~n28204 & n28205 ;
  assign n28207 = ~n28193 & n28206 ;
  assign n28208 = ~\u2_desIn_r_reg[54]/NET0131  & ~n28207 ;
  assign n28209 = \u2_desIn_r_reg[54]/NET0131  & n28207 ;
  assign n28210 = ~n28208 & ~n28209 ;
  assign n28226 = ~n27448 & ~n27450 ;
  assign n28227 = ~n27919 & n28226 ;
  assign n28228 = ~n27411 & ~n28227 ;
  assign n28224 = ~n27419 & ~n27420 ;
  assign n28225 = n27411 & ~n28224 ;
  assign n28229 = ~n27412 & n27918 ;
  assign n28230 = ~n28225 & n28229 ;
  assign n28231 = ~n28228 & n28230 ;
  assign n28232 = ~n27436 & ~n28231 ;
  assign n28211 = ~n27391 & n27414 ;
  assign n28212 = ~n27448 & ~n28211 ;
  assign n28213 = n27411 & ~n28212 ;
  assign n28214 = ~n27411 & n27462 ;
  assign n28215 = n27468 & ~n28214 ;
  assign n28216 = ~n28213 & n28215 ;
  assign n28217 = n27436 & ~n28216 ;
  assign n28218 = ~n27411 & ~n27447 ;
  assign n28219 = n27411 & ~n27466 ;
  assign n28220 = n27399 & n27919 ;
  assign n28221 = ~n27423 & ~n28220 ;
  assign n28222 = n28219 & n28221 ;
  assign n28223 = ~n28218 & ~n28222 ;
  assign n28233 = ~n28217 & ~n28223 ;
  assign n28234 = ~n28232 & n28233 ;
  assign n28235 = ~\u2_desIn_r_reg[62]/NET0131  & ~n28234 ;
  assign n28236 = \u2_desIn_r_reg[62]/NET0131  & n28234 ;
  assign n28237 = ~n28235 & ~n28236 ;
  assign n28238 = n28122 & ~n28158 ;
  assign n28240 = n28144 & n28147 ;
  assign n28239 = n28106 & ~n28112 ;
  assign n28241 = ~n28122 & ~n28239 ;
  assign n28242 = n28154 & n28241 ;
  assign n28243 = ~n28240 & n28242 ;
  assign n28244 = ~n28238 & ~n28243 ;
  assign n28245 = n28114 & n28122 ;
  assign n28246 = ~n28105 & n28245 ;
  assign n28247 = n28144 & ~n28167 ;
  assign n28248 = ~n28246 & n28247 ;
  assign n28249 = n28112 & n28122 ;
  assign n28250 = ~n28099 & ~n28123 ;
  assign n28251 = ~n28249 & n28250 ;
  assign n28252 = ~n28248 & n28251 ;
  assign n28253 = ~n28244 & ~n28252 ;
  assign n28254 = n28132 & ~n28253 ;
  assign n28255 = ~n28105 & n28249 ;
  assign n28256 = ~n28144 & ~n28255 ;
  assign n28257 = ~n28248 & ~n28256 ;
  assign n28262 = n28114 & ~n28122 ;
  assign n28263 = ~n28153 & ~n28239 ;
  assign n28264 = ~n28262 & n28263 ;
  assign n28265 = ~n28144 & ~n28264 ;
  assign n28259 = ~n28114 & n28144 ;
  assign n28258 = ~n28105 & ~n28115 ;
  assign n28260 = ~n28153 & ~n28258 ;
  assign n28261 = n28259 & n28260 ;
  assign n28266 = ~n28135 & ~n28261 ;
  assign n28267 = ~n28265 & n28266 ;
  assign n28268 = ~n28132 & ~n28267 ;
  assign n28269 = ~n28257 & ~n28268 ;
  assign n28270 = ~n28254 & n28269 ;
  assign n28271 = ~\u2_desIn_r_reg[60]/NET0131  & ~n28270 ;
  assign n28272 = \u2_desIn_r_reg[60]/NET0131  & n28270 ;
  assign n28273 = ~n28271 & ~n28272 ;
  assign n28283 = ~n28122 & n28144 ;
  assign n28294 = ~n28105 & ~n28157 ;
  assign n28295 = n28283 & n28294 ;
  assign n28290 = ~n28134 & ~n28144 ;
  assign n28291 = ~n28116 & n28290 ;
  assign n28292 = ~n28113 & n28122 ;
  assign n28293 = n28259 & n28292 ;
  assign n28296 = ~n28291 & ~n28293 ;
  assign n28297 = ~n28295 & n28296 ;
  assign n28298 = ~n28164 & n28297 ;
  assign n28299 = n28132 & ~n28298 ;
  assign n28274 = n28099 & n28123 ;
  assign n28275 = ~n28245 & ~n28274 ;
  assign n28276 = ~n28147 & ~n28255 ;
  assign n28277 = n28275 & n28276 ;
  assign n28278 = n28144 & ~n28277 ;
  assign n28279 = ~n28099 & n28255 ;
  assign n28280 = ~n28278 & ~n28279 ;
  assign n28281 = ~n28132 & ~n28280 ;
  assign n28286 = ~n28116 & n28134 ;
  assign n28287 = ~n28125 & ~n28286 ;
  assign n28288 = ~n28132 & ~n28144 ;
  assign n28289 = ~n28287 & n28288 ;
  assign n28282 = n28153 & n28159 ;
  assign n28284 = ~n28152 & ~n28158 ;
  assign n28285 = n28283 & ~n28284 ;
  assign n28300 = ~n28282 & ~n28285 ;
  assign n28301 = ~n28289 & n28300 ;
  assign n28302 = ~n28281 & n28301 ;
  assign n28303 = ~n28299 & n28302 ;
  assign n28304 = ~\u2_desIn_r_reg[58]/NET0131  & ~n28303 ;
  assign n28305 = \u2_desIn_r_reg[58]/NET0131  & n28303 ;
  assign n28306 = ~n28304 & ~n28305 ;
  assign n28308 = ~n27543 & ~n27547 ;
  assign n28309 = n27481 & ~n28308 ;
  assign n28310 = ~n27665 & ~n27683 ;
  assign n28311 = n27965 & n28310 ;
  assign n28312 = ~n28309 & ~n28311 ;
  assign n28313 = ~n27661 & ~n27681 ;
  assign n28314 = ~n27967 & n28313 ;
  assign n28315 = ~n28312 & n28314 ;
  assign n28316 = n27520 & ~n28315 ;
  assign n28317 = ~n27507 & n27690 ;
  assign n28318 = n27481 & ~n27546 ;
  assign n28319 = ~n28317 & n28318 ;
  assign n28320 = n27536 & n27658 ;
  assign n28321 = ~n27662 & ~n28320 ;
  assign n28322 = ~n27975 & n28321 ;
  assign n28323 = ~n28319 & n28322 ;
  assign n28324 = ~n27520 & ~n28323 ;
  assign n28325 = ~n27481 & n27974 ;
  assign n28307 = n27529 & n27533 ;
  assign n28326 = ~n27972 & ~n28307 ;
  assign n28327 = ~n28325 & n28326 ;
  assign n28328 = ~n28324 & n28327 ;
  assign n28329 = ~n28316 & n28328 ;
  assign n28330 = ~\u2_desIn_r_reg[16]/NET0131  & ~n28329 ;
  assign n28331 = \u2_desIn_r_reg[16]/NET0131  & n28329 ;
  assign n28332 = ~n28330 & ~n28331 ;
  assign n28334 = ~n28122 & n28152 ;
  assign n28335 = n28275 & ~n28334 ;
  assign n28336 = n28132 & ~n28335 ;
  assign n28337 = ~n28165 & ~n28249 ;
  assign n28338 = ~n28132 & ~n28166 ;
  assign n28339 = ~n28337 & n28338 ;
  assign n28340 = ~n28336 & ~n28339 ;
  assign n28341 = n28144 & ~n28340 ;
  assign n28345 = n28122 & n28239 ;
  assign n28342 = ~n28105 & ~n28112 ;
  assign n28343 = ~n28144 & ~n28342 ;
  assign n28344 = n28337 & n28343 ;
  assign n28346 = ~n28286 & ~n28344 ;
  assign n28347 = ~n28345 & n28346 ;
  assign n28348 = ~n28132 & ~n28347 ;
  assign n28349 = ~n28147 & ~n28249 ;
  assign n28350 = n28149 & ~n28349 ;
  assign n28352 = n28105 & ~n28115 ;
  assign n28353 = n28146 & n28352 ;
  assign n28333 = n28159 & n28165 ;
  assign n28351 = n28161 & n28255 ;
  assign n28354 = ~n28333 & ~n28351 ;
  assign n28355 = ~n28353 & n28354 ;
  assign n28356 = ~n28350 & n28355 ;
  assign n28357 = ~n28348 & n28356 ;
  assign n28358 = ~n28341 & n28357 ;
  assign n28359 = \u2_desIn_r_reg[40]/NET0131  & ~n28358 ;
  assign n28360 = ~\u2_desIn_r_reg[40]/NET0131  & n28358 ;
  assign n28361 = ~n28359 & ~n28360 ;
  assign n28365 = n27436 & ~n27447 ;
  assign n28366 = ~n27421 & n28365 ;
  assign n28362 = ~n27422 & ~n27462 ;
  assign n28363 = ~n27385 & n27411 ;
  assign n28364 = ~n28362 & n28363 ;
  assign n28367 = ~n27451 & ~n28364 ;
  assign n28368 = n28366 & n28367 ;
  assign n28372 = ~n27441 & ~n27919 ;
  assign n28373 = n27411 & ~n28372 ;
  assign n28369 = n27411 & ~n27446 ;
  assign n28370 = ~n27393 & ~n27448 ;
  assign n28371 = ~n28369 & ~n28370 ;
  assign n28374 = ~n27436 & ~n28371 ;
  assign n28375 = ~n28373 & n28374 ;
  assign n28376 = ~n28368 & ~n28375 ;
  assign n28377 = ~n27419 & n28219 ;
  assign n28378 = n27404 & n27446 ;
  assign n28379 = ~n27411 & ~n27463 ;
  assign n28380 = ~n28378 & n28379 ;
  assign n28381 = ~n28211 & n28380 ;
  assign n28382 = ~n28377 & ~n28381 ;
  assign n28383 = ~n28376 & ~n28382 ;
  assign n28384 = ~\u2_desIn_r_reg[22]/NET0131  & ~n28383 ;
  assign n28385 = \u2_desIn_r_reg[22]/NET0131  & n28383 ;
  assign n28386 = ~n28384 & ~n28385 ;
  assign n28387 = n27024 & n27589 ;
  assign n28388 = ~n27024 & n27103 ;
  assign n28394 = ~n27070 & ~n28388 ;
  assign n28395 = ~n28387 & n28394 ;
  assign n28389 = ~n27051 & ~n28048 ;
  assign n28390 = ~n27037 & ~n28389 ;
  assign n28391 = ~n27072 & n27085 ;
  assign n28392 = ~n27056 & ~n28391 ;
  assign n28393 = n27037 & ~n28392 ;
  assign n28396 = ~n28390 & ~n28393 ;
  assign n28397 = n28395 & n28396 ;
  assign n28398 = n27599 & n28028 ;
  assign n28399 = n27024 & ~n28398 ;
  assign n28400 = n27054 & ~n28389 ;
  assign n28401 = n27070 & ~n27603 ;
  assign n28402 = ~n28400 & n28401 ;
  assign n28403 = ~n28399 & n28402 ;
  assign n28404 = ~n28397 & ~n28403 ;
  assign n28405 = ~n27037 & n27609 ;
  assign n28406 = ~n27073 & n28405 ;
  assign n28407 = ~n28404 & ~n28406 ;
  assign n28408 = ~\u2_desIn_r_reg[4]/NET0131  & ~n28407 ;
  assign n28409 = \u2_desIn_r_reg[4]/NET0131  & n28407 ;
  assign n28410 = ~n28408 & ~n28409 ;
  assign n28413 = n27766 & ~n27885 ;
  assign n28411 = ~n27779 & ~n28012 ;
  assign n28412 = ~n27766 & ~n28411 ;
  assign n28414 = ~n27864 & ~n28412 ;
  assign n28415 = ~n28413 & n28414 ;
  assign n28416 = n27773 & ~n28415 ;
  assign n28421 = ~n27861 & ~n27998 ;
  assign n28422 = ~n27759 & n28421 ;
  assign n28417 = n27766 & n27781 ;
  assign n28418 = n27742 & n27766 ;
  assign n28419 = ~n27749 & ~n28418 ;
  assign n28420 = n27871 & n28419 ;
  assign n28423 = ~n28417 & ~n28420 ;
  assign n28424 = n28422 & n28423 ;
  assign n28425 = ~n27773 & ~n28424 ;
  assign n28426 = ~n27766 & n27787 ;
  assign n28427 = n27742 & n27780 ;
  assign n28428 = ~n27995 & ~n28427 ;
  assign n28429 = n27766 & ~n28428 ;
  assign n28430 = ~n28426 & ~n28429 ;
  assign n28431 = ~n28425 & n28430 ;
  assign n28432 = ~n28416 & n28431 ;
  assign n28433 = ~\u2_desIn_r_reg[10]/P0001  & ~n28432 ;
  assign n28434 = \u2_desIn_r_reg[10]/P0001  & n28432 ;
  assign n28435 = ~n28433 & ~n28434 ;
  assign n28436 = decrypt_pad & ~\u1_uk_K_r14_reg[49]/NET0131  ;
  assign n28437 = ~decrypt_pad & ~\u1_uk_K_r14_reg[1]/NET0131  ;
  assign n28438 = ~n28436 & ~n28437 ;
  assign n28439 = \u1_R14_reg[31]/P0001  & ~n28438 ;
  assign n28440 = ~\u1_R14_reg[31]/P0001  & n28438 ;
  assign n28441 = ~n28439 & ~n28440 ;
  assign n28442 = decrypt_pad & ~\u1_uk_K_r14_reg[36]/NET0131  ;
  assign n28443 = ~decrypt_pad & ~\u1_uk_K_r14_reg[43]/NET0131  ;
  assign n28444 = ~n28442 & ~n28443 ;
  assign n28445 = \u1_R14_reg[29]/NET0131  & ~n28444 ;
  assign n28446 = ~\u1_R14_reg[29]/NET0131  & n28444 ;
  assign n28447 = ~n28445 & ~n28446 ;
  assign n28448 = decrypt_pad & ~\u1_uk_K_r14_reg[21]/NET0131  ;
  assign n28449 = ~decrypt_pad & ~\u1_uk_K_r14_reg[28]/NET0131  ;
  assign n28450 = ~n28448 & ~n28449 ;
  assign n28451 = \u1_R14_reg[1]/NET0131  & ~n28450 ;
  assign n28452 = ~\u1_R14_reg[1]/NET0131  & n28450 ;
  assign n28453 = ~n28451 & ~n28452 ;
  assign n28463 = n28447 & ~n28453 ;
  assign n28464 = decrypt_pad & ~\u1_uk_K_r14_reg[37]/NET0131  ;
  assign n28465 = ~decrypt_pad & ~\u1_uk_K_r14_reg[44]/NET0131  ;
  assign n28466 = ~n28464 & ~n28465 ;
  assign n28467 = \u1_R14_reg[30]/NET0131  & ~n28466 ;
  assign n28468 = ~\u1_R14_reg[30]/NET0131  & n28466 ;
  assign n28469 = ~n28467 & ~n28468 ;
  assign n28470 = n28463 & ~n28469 ;
  assign n28454 = ~n28447 & n28453 ;
  assign n28455 = decrypt_pad & ~\u1_uk_K_r14_reg[9]/NET0131  ;
  assign n28456 = ~decrypt_pad & ~\u1_uk_K_r14_reg[16]/NET0131  ;
  assign n28457 = ~n28455 & ~n28456 ;
  assign n28458 = \u1_R14_reg[28]/NET0131  & ~n28457 ;
  assign n28459 = ~\u1_R14_reg[28]/NET0131  & n28457 ;
  assign n28460 = ~n28458 & ~n28459 ;
  assign n28461 = n28454 & ~n28460 ;
  assign n28462 = n28447 & n28460 ;
  assign n28471 = ~n28461 & ~n28462 ;
  assign n28472 = ~n28470 & n28471 ;
  assign n28473 = n28441 & ~n28472 ;
  assign n28474 = n28460 & ~n28469 ;
  assign n28475 = ~n28453 & n28474 ;
  assign n28476 = ~n28447 & n28475 ;
  assign n28477 = decrypt_pad & ~\u1_uk_K_r14_reg[0]/P0001  ;
  assign n28478 = ~decrypt_pad & ~\u1_uk_K_r14_reg[7]/NET0131  ;
  assign n28479 = ~n28477 & ~n28478 ;
  assign n28480 = \u1_R14_reg[32]/NET0131  & ~n28479 ;
  assign n28481 = ~\u1_R14_reg[32]/NET0131  & n28479 ;
  assign n28482 = ~n28480 & ~n28481 ;
  assign n28483 = ~n28476 & ~n28482 ;
  assign n28484 = ~n28473 & n28483 ;
  assign n28488 = n28447 & ~n28469 ;
  assign n28489 = n28460 & n28488 ;
  assign n28498 = n28482 & ~n28489 ;
  assign n28493 = n28441 & ~n28447 ;
  assign n28494 = ~n28453 & ~n28460 ;
  assign n28495 = n28493 & n28494 ;
  assign n28496 = ~n28441 & n28469 ;
  assign n28497 = n28454 & n28496 ;
  assign n28499 = ~n28495 & ~n28497 ;
  assign n28500 = n28498 & n28499 ;
  assign n28485 = ~n28460 & n28469 ;
  assign n28486 = n28447 & n28485 ;
  assign n28487 = ~n28453 & n28486 ;
  assign n28490 = ~n28447 & n28460 ;
  assign n28491 = n28469 & n28490 ;
  assign n28492 = n28453 & n28491 ;
  assign n28501 = ~n28487 & ~n28492 ;
  assign n28502 = n28500 & n28501 ;
  assign n28503 = ~n28484 & ~n28502 ;
  assign n28510 = ~n28441 & ~n28491 ;
  assign n28511 = ~n28487 & n28510 ;
  assign n28504 = n28453 & ~n28460 ;
  assign n28505 = n28447 & n28504 ;
  assign n28506 = ~n28469 & n28505 ;
  assign n28507 = ~n28447 & ~n28460 ;
  assign n28508 = ~n28469 & n28507 ;
  assign n28509 = ~n28453 & n28508 ;
  assign n28512 = ~n28506 & ~n28509 ;
  assign n28513 = n28511 & n28512 ;
  assign n28515 = n28461 & ~n28469 ;
  assign n28514 = n28453 & n28486 ;
  assign n28516 = n28441 & ~n28514 ;
  assign n28517 = ~n28515 & n28516 ;
  assign n28518 = ~n28513 & ~n28517 ;
  assign n28519 = ~n28441 & ~n28482 ;
  assign n28520 = n28490 & n28519 ;
  assign n28521 = ~n28518 & ~n28520 ;
  assign n28522 = ~n28503 & n28521 ;
  assign n28523 = \u1_L14_reg[15]/P0001  & n28522 ;
  assign n28524 = ~\u1_L14_reg[15]/P0001  & ~n28522 ;
  assign n28525 = ~n28523 & ~n28524 ;
  assign n28526 = decrypt_pad & ~\u1_uk_K_r14_reg[53]/NET0131  ;
  assign n28527 = ~decrypt_pad & ~\u1_uk_K_r14_reg[3]/NET0131  ;
  assign n28528 = ~n28526 & ~n28527 ;
  assign n28529 = \u1_R14_reg[3]/NET0131  & ~n28528 ;
  assign n28530 = ~\u1_R14_reg[3]/NET0131  & n28528 ;
  assign n28531 = ~n28529 & ~n28530 ;
  assign n28532 = decrypt_pad & ~\u1_uk_K_r14_reg[19]/NET0131  ;
  assign n28533 = ~decrypt_pad & ~\u1_uk_K_r14_reg[26]/NET0131  ;
  assign n28534 = ~n28532 & ~n28533 ;
  assign n28535 = \u1_R14_reg[2]/NET0131  & ~n28534 ;
  assign n28536 = ~\u1_R14_reg[2]/NET0131  & n28534 ;
  assign n28537 = ~n28535 & ~n28536 ;
  assign n28552 = decrypt_pad & ~\u1_uk_K_r14_reg[40]/NET0131  ;
  assign n28553 = ~decrypt_pad & ~\u1_uk_K_r14_reg[47]/NET0131  ;
  assign n28554 = ~n28552 & ~n28553 ;
  assign n28555 = \u1_R14_reg[32]/NET0131  & ~n28554 ;
  assign n28556 = ~\u1_R14_reg[32]/NET0131  & n28554 ;
  assign n28557 = ~n28555 & ~n28556 ;
  assign n28538 = decrypt_pad & ~\u1_uk_K_r14_reg[34]/NET0131  ;
  assign n28539 = ~decrypt_pad & ~\u1_uk_K_r14_reg[41]/NET0131  ;
  assign n28540 = ~n28538 & ~n28539 ;
  assign n28541 = \u1_R14_reg[5]/NET0131  & ~n28540 ;
  assign n28542 = ~\u1_R14_reg[5]/NET0131  & n28540 ;
  assign n28543 = ~n28541 & ~n28542 ;
  assign n28545 = decrypt_pad & ~\u1_uk_K_r14_reg[4]/NET0131  ;
  assign n28546 = ~decrypt_pad & ~\u1_uk_K_r14_reg[11]/NET0131  ;
  assign n28547 = ~n28545 & ~n28546 ;
  assign n28548 = \u1_R14_reg[1]/NET0131  & ~n28547 ;
  assign n28549 = ~\u1_R14_reg[1]/NET0131  & n28547 ;
  assign n28550 = ~n28548 & ~n28549 ;
  assign n28562 = ~n28543 & ~n28550 ;
  assign n28563 = n28557 & n28562 ;
  assign n28564 = n28537 & n28563 ;
  assign n28565 = ~n28543 & ~n28557 ;
  assign n28566 = n28550 & n28565 ;
  assign n28567 = n28543 & ~n28550 ;
  assign n28568 = ~n28566 & ~n28567 ;
  assign n28569 = ~n28557 & ~n28568 ;
  assign n28570 = ~n28564 & ~n28569 ;
  assign n28571 = decrypt_pad & ~\u1_uk_K_r14_reg[6]/NET0131  ;
  assign n28572 = ~decrypt_pad & ~\u1_uk_K_r14_reg[13]/NET0131  ;
  assign n28573 = ~n28571 & ~n28572 ;
  assign n28574 = \u1_R14_reg[4]/NET0131  & ~n28573 ;
  assign n28575 = ~\u1_R14_reg[4]/NET0131  & n28573 ;
  assign n28576 = ~n28574 & ~n28575 ;
  assign n28577 = ~n28570 & n28576 ;
  assign n28544 = ~n28537 & ~n28543 ;
  assign n28551 = n28544 & n28550 ;
  assign n28558 = n28551 & n28557 ;
  assign n28559 = n28537 & n28550 ;
  assign n28560 = n28543 & n28557 ;
  assign n28561 = n28559 & n28560 ;
  assign n28578 = n28543 & ~n28557 ;
  assign n28579 = ~n28537 & ~n28550 ;
  assign n28580 = n28578 & n28579 ;
  assign n28581 = ~n28561 & ~n28580 ;
  assign n28582 = ~n28558 & n28581 ;
  assign n28583 = ~n28577 & n28582 ;
  assign n28584 = ~n28531 & ~n28583 ;
  assign n28585 = ~n28531 & n28557 ;
  assign n28586 = n28537 & n28585 ;
  assign n28587 = n28537 & ~n28557 ;
  assign n28588 = n28531 & n28587 ;
  assign n28589 = ~n28586 & ~n28588 ;
  assign n28590 = n28543 & ~n28589 ;
  assign n28593 = n28531 & n28566 ;
  assign n28591 = n28543 & n28559 ;
  assign n28595 = ~n28576 & ~n28591 ;
  assign n28592 = ~n28543 & n28579 ;
  assign n28594 = n28550 & n28585 ;
  assign n28596 = ~n28592 & ~n28594 ;
  assign n28597 = n28595 & n28596 ;
  assign n28598 = ~n28593 & n28597 ;
  assign n28599 = ~n28590 & n28598 ;
  assign n28602 = ~n28543 & n28559 ;
  assign n28603 = n28557 & n28602 ;
  assign n28604 = n28550 & n28578 ;
  assign n28605 = ~n28603 & ~n28604 ;
  assign n28606 = n28531 & ~n28605 ;
  assign n28607 = n28562 & n28588 ;
  assign n28600 = ~n28537 & n28560 ;
  assign n28601 = ~n28550 & n28600 ;
  assign n28608 = n28576 & ~n28601 ;
  assign n28609 = ~n28607 & n28608 ;
  assign n28610 = ~n28606 & n28609 ;
  assign n28611 = ~n28599 & ~n28610 ;
  assign n28612 = n28531 & n28557 ;
  assign n28613 = n28579 & n28612 ;
  assign n28614 = n28531 & ~n28537 ;
  assign n28615 = n28566 & n28614 ;
  assign n28616 = ~n28613 & ~n28615 ;
  assign n28617 = ~n28611 & n28616 ;
  assign n28618 = ~n28584 & n28617 ;
  assign n28619 = ~\u1_L14_reg[23]/P0001  & n28618 ;
  assign n28620 = \u1_L14_reg[23]/P0001  & ~n28618 ;
  assign n28621 = ~n28619 & ~n28620 ;
  assign n28622 = decrypt_pad & ~\u1_uk_K_r14_reg[10]/P0001  ;
  assign n28623 = ~decrypt_pad & ~\u1_uk_K_r14_reg[17]/NET0131  ;
  assign n28624 = ~n28622 & ~n28623 ;
  assign n28625 = \u1_R14_reg[12]/NET0131  & ~n28624 ;
  assign n28626 = ~\u1_R14_reg[12]/NET0131  & n28624 ;
  assign n28627 = ~n28625 & ~n28626 ;
  assign n28648 = decrypt_pad & ~\u1_uk_K_r14_reg[26]/NET0131  ;
  assign n28649 = ~decrypt_pad & ~\u1_uk_K_r14_reg[33]/NET0131  ;
  assign n28650 = ~n28648 & ~n28649 ;
  assign n28651 = \u1_R14_reg[10]/P0001  & ~n28650 ;
  assign n28652 = ~\u1_R14_reg[10]/P0001  & n28650 ;
  assign n28653 = ~n28651 & ~n28652 ;
  assign n28634 = decrypt_pad & ~\u1_uk_K_r14_reg[46]/NET0131  ;
  assign n28635 = ~decrypt_pad & ~\u1_uk_K_r14_reg[53]/NET0131  ;
  assign n28636 = ~n28634 & ~n28635 ;
  assign n28637 = \u1_R14_reg[8]/NET0131  & ~n28636 ;
  assign n28638 = ~\u1_R14_reg[8]/NET0131  & n28636 ;
  assign n28639 = ~n28637 & ~n28638 ;
  assign n28641 = decrypt_pad & ~\u1_uk_K_r14_reg[55]/NET0131  ;
  assign n28642 = ~decrypt_pad & ~\u1_uk_K_r14_reg[5]/NET0131  ;
  assign n28643 = ~n28641 & ~n28642 ;
  assign n28644 = \u1_R14_reg[13]/NET0131  & ~n28643 ;
  assign n28645 = ~\u1_R14_reg[13]/NET0131  & n28643 ;
  assign n28646 = ~n28644 & ~n28645 ;
  assign n28655 = ~n28639 & n28646 ;
  assign n28656 = ~n28653 & n28655 ;
  assign n28657 = ~n28639 & n28653 ;
  assign n28658 = ~n28646 & n28657 ;
  assign n28659 = ~n28656 & ~n28658 ;
  assign n28628 = decrypt_pad & ~\u1_uk_K_r14_reg[18]/NET0131  ;
  assign n28629 = ~decrypt_pad & ~\u1_uk_K_r14_reg[25]/NET0131  ;
  assign n28630 = ~n28628 & ~n28629 ;
  assign n28631 = \u1_R14_reg[9]/NET0131  & ~n28630 ;
  assign n28632 = ~\u1_R14_reg[9]/NET0131  & n28630 ;
  assign n28633 = ~n28631 & ~n28632 ;
  assign n28640 = ~n28633 & n28639 ;
  assign n28647 = n28640 & ~n28646 ;
  assign n28654 = n28647 & ~n28653 ;
  assign n28660 = decrypt_pad & ~\u1_uk_K_r14_reg[27]/NET0131  ;
  assign n28661 = ~decrypt_pad & ~\u1_uk_K_r14_reg[34]/NET0131  ;
  assign n28662 = ~n28660 & ~n28661 ;
  assign n28663 = \u1_R14_reg[11]/P0001  & ~n28662 ;
  assign n28664 = ~\u1_R14_reg[11]/P0001  & n28662 ;
  assign n28665 = ~n28663 & ~n28664 ;
  assign n28666 = ~n28654 & n28665 ;
  assign n28667 = n28659 & n28666 ;
  assign n28669 = n28633 & ~n28646 ;
  assign n28670 = ~n28639 & n28669 ;
  assign n28668 = n28639 & n28653 ;
  assign n28671 = ~n28665 & ~n28668 ;
  assign n28672 = ~n28670 & n28671 ;
  assign n28673 = ~n28667 & ~n28672 ;
  assign n28674 = n28627 & ~n28673 ;
  assign n28685 = n28668 & ~n28669 ;
  assign n28683 = n28633 & ~n28653 ;
  assign n28684 = ~n28646 & n28683 ;
  assign n28686 = n28665 & ~n28684 ;
  assign n28687 = ~n28685 & n28686 ;
  assign n28689 = n28639 & ~n28653 ;
  assign n28690 = ~n28669 & n28689 ;
  assign n28688 = n28633 & n28655 ;
  assign n28691 = ~n28665 & ~n28688 ;
  assign n28692 = ~n28690 & n28691 ;
  assign n28693 = ~n28687 & ~n28692 ;
  assign n28678 = ~n28633 & ~n28653 ;
  assign n28679 = n28639 & n28646 ;
  assign n28680 = ~n28639 & ~n28646 ;
  assign n28681 = ~n28679 & ~n28680 ;
  assign n28682 = n28678 & ~n28681 ;
  assign n28675 = ~n28633 & n28646 ;
  assign n28676 = n28653 & n28675 ;
  assign n28677 = ~n28639 & n28676 ;
  assign n28694 = ~n28627 & ~n28677 ;
  assign n28695 = ~n28682 & n28694 ;
  assign n28696 = ~n28693 & n28695 ;
  assign n28697 = ~n28674 & ~n28696 ;
  assign n28703 = n28665 & n28668 ;
  assign n28704 = n28675 & n28703 ;
  assign n28698 = n28653 & ~n28665 ;
  assign n28699 = n28669 & n28698 ;
  assign n28700 = n28633 & ~n28679 ;
  assign n28701 = n28627 & n28653 ;
  assign n28702 = n28700 & n28701 ;
  assign n28705 = ~n28699 & ~n28702 ;
  assign n28706 = ~n28704 & n28705 ;
  assign n28707 = ~n28697 & n28706 ;
  assign n28708 = ~\u1_L14_reg[30]/P0001  & n28707 ;
  assign n28709 = \u1_L14_reg[30]/P0001  & ~n28707 ;
  assign n28710 = ~n28708 & ~n28709 ;
  assign n28711 = decrypt_pad & ~\u1_uk_K_r14_reg[32]/NET0131  ;
  assign n28712 = ~decrypt_pad & ~\u1_uk_K_r14_reg[39]/P0001  ;
  assign n28713 = ~n28711 & ~n28712 ;
  assign n28714 = \u1_R14_reg[8]/NET0131  & ~n28713 ;
  assign n28715 = ~\u1_R14_reg[8]/NET0131  & n28713 ;
  assign n28716 = ~n28714 & ~n28715 ;
  assign n28723 = decrypt_pad & ~\u1_uk_K_r14_reg[20]/NET0131  ;
  assign n28724 = ~decrypt_pad & ~\u1_uk_K_r14_reg[27]/NET0131  ;
  assign n28725 = ~n28723 & ~n28724 ;
  assign n28726 = \u1_R14_reg[4]/NET0131  & ~n28725 ;
  assign n28727 = ~\u1_R14_reg[4]/NET0131  & n28725 ;
  assign n28728 = ~n28726 & ~n28727 ;
  assign n28729 = decrypt_pad & ~\u1_uk_K_r14_reg[12]/NET0131  ;
  assign n28730 = ~decrypt_pad & ~\u1_uk_K_r14_reg[19]/NET0131  ;
  assign n28731 = ~n28729 & ~n28730 ;
  assign n28732 = \u1_R14_reg[9]/NET0131  & ~n28731 ;
  assign n28733 = ~\u1_R14_reg[9]/NET0131  & n28731 ;
  assign n28734 = ~n28732 & ~n28733 ;
  assign n28752 = n28728 & n28734 ;
  assign n28735 = decrypt_pad & ~\u1_uk_K_r14_reg[24]/NET0131  ;
  assign n28736 = ~decrypt_pad & ~\u1_uk_K_r14_reg[6]/NET0131  ;
  assign n28737 = ~n28735 & ~n28736 ;
  assign n28738 = \u1_R14_reg[5]/NET0131  & ~n28737 ;
  assign n28739 = ~\u1_R14_reg[5]/NET0131  & n28737 ;
  assign n28740 = ~n28738 & ~n28739 ;
  assign n28742 = decrypt_pad & ~\u1_uk_K_r14_reg[47]/NET0131  ;
  assign n28743 = ~decrypt_pad & ~\u1_uk_K_r14_reg[54]/NET0131  ;
  assign n28744 = ~n28742 & ~n28743 ;
  assign n28745 = \u1_R14_reg[6]/NET0131  & ~n28744 ;
  assign n28746 = ~\u1_R14_reg[6]/NET0131  & n28744 ;
  assign n28747 = ~n28745 & ~n28746 ;
  assign n28770 = ~n28740 & n28747 ;
  assign n28717 = decrypt_pad & ~\u1_uk_K_r14_reg[41]/NET0131  ;
  assign n28718 = ~decrypt_pad & ~\u1_uk_K_r14_reg[48]/NET0131  ;
  assign n28719 = ~n28717 & ~n28718 ;
  assign n28720 = \u1_R14_reg[7]/P0001  & ~n28719 ;
  assign n28721 = ~\u1_R14_reg[7]/P0001  & n28719 ;
  assign n28722 = ~n28720 & ~n28721 ;
  assign n28771 = n28722 & n28740 ;
  assign n28772 = ~n28770 & ~n28771 ;
  assign n28777 = n28752 & ~n28772 ;
  assign n28764 = n28740 & ~n28747 ;
  assign n28773 = ~n28728 & ~n28764 ;
  assign n28774 = n28772 & n28773 ;
  assign n28757 = ~n28734 & ~n28740 ;
  assign n28775 = ~n28747 & n28757 ;
  assign n28741 = ~n28734 & n28740 ;
  assign n28766 = n28728 & n28747 ;
  assign n28776 = n28741 & n28766 ;
  assign n28778 = ~n28775 & ~n28776 ;
  assign n28779 = ~n28774 & n28778 ;
  assign n28780 = ~n28777 & n28779 ;
  assign n28781 = ~n28716 & ~n28780 ;
  assign n28753 = n28734 & ~n28740 ;
  assign n28754 = ~n28741 & ~n28753 ;
  assign n28755 = ~n28752 & ~n28754 ;
  assign n28756 = n28722 & n28755 ;
  assign n28748 = n28734 & n28747 ;
  assign n28749 = ~n28722 & n28728 ;
  assign n28750 = ~n28741 & n28749 ;
  assign n28751 = ~n28748 & n28750 ;
  assign n28758 = ~n28728 & n28747 ;
  assign n28759 = n28757 & n28758 ;
  assign n28760 = ~n28751 & ~n28759 ;
  assign n28761 = ~n28756 & n28760 ;
  assign n28762 = n28716 & ~n28761 ;
  assign n28763 = ~n28728 & ~n28734 ;
  assign n28765 = n28763 & n28764 ;
  assign n28767 = n28734 & n28766 ;
  assign n28768 = ~n28765 & ~n28767 ;
  assign n28769 = n28722 & ~n28768 ;
  assign n28782 = ~n28728 & n28740 ;
  assign n28783 = ~n28722 & n28734 ;
  assign n28784 = n28782 & n28783 ;
  assign n28785 = ~n28769 & ~n28784 ;
  assign n28786 = ~n28762 & n28785 ;
  assign n28787 = ~n28781 & n28786 ;
  assign n28788 = ~\u1_L14_reg[18]/P0001  & ~n28787 ;
  assign n28789 = \u1_L14_reg[18]/P0001  & n28787 ;
  assign n28790 = ~n28788 & ~n28789 ;
  assign n28837 = decrypt_pad & ~\u1_uk_K_r13_reg[24]/NET0131  ;
  assign n28838 = ~decrypt_pad & ~\u1_uk_K_r13_reg[20]/NET0131  ;
  assign n28839 = ~n28837 & ~n28838 ;
  assign n28840 = \u1_R13_reg[4]/NET0131  & ~n28839 ;
  assign n28841 = ~\u1_R13_reg[4]/NET0131  & n28839 ;
  assign n28842 = ~n28840 & ~n28841 ;
  assign n28791 = decrypt_pad & ~\u1_uk_K_r13_reg[46]/NET0131  ;
  assign n28792 = ~decrypt_pad & ~\u1_uk_K_r13_reg[10]/NET0131  ;
  assign n28793 = ~n28791 & ~n28792 ;
  assign n28794 = \u1_R13_reg[3]/NET0131  & ~n28793 ;
  assign n28795 = ~\u1_R13_reg[3]/NET0131  & n28793 ;
  assign n28796 = ~n28794 & ~n28795 ;
  assign n28819 = decrypt_pad & ~\u1_uk_K_r13_reg[33]/NET0131  ;
  assign n28820 = ~decrypt_pad & ~\u1_uk_K_r13_reg[54]/NET0131  ;
  assign n28821 = ~n28819 & ~n28820 ;
  assign n28822 = \u1_R13_reg[32]/NET0131  & ~n28821 ;
  assign n28823 = ~\u1_R13_reg[32]/NET0131  & n28821 ;
  assign n28824 = ~n28822 & ~n28823 ;
  assign n28804 = decrypt_pad & ~\u1_uk_K_r13_reg[27]/NET0131  ;
  assign n28805 = ~decrypt_pad & ~\u1_uk_K_r13_reg[48]/NET0131  ;
  assign n28806 = ~n28804 & ~n28805 ;
  assign n28807 = \u1_R13_reg[5]/NET0131  & ~n28806 ;
  assign n28808 = ~\u1_R13_reg[5]/NET0131  & n28806 ;
  assign n28809 = ~n28807 & ~n28808 ;
  assign n28797 = decrypt_pad & ~\u1_uk_K_r13_reg[54]/NET0131  ;
  assign n28798 = ~decrypt_pad & ~\u1_uk_K_r13_reg[18]/NET0131  ;
  assign n28799 = ~n28797 & ~n28798 ;
  assign n28800 = \u1_R13_reg[1]/NET0131  & ~n28799 ;
  assign n28801 = ~\u1_R13_reg[1]/NET0131  & n28799 ;
  assign n28802 = ~n28800 & ~n28801 ;
  assign n28810 = decrypt_pad & ~\u1_uk_K_r13_reg[12]/NET0131  ;
  assign n28811 = ~decrypt_pad & ~\u1_uk_K_r13_reg[33]/NET0131  ;
  assign n28812 = ~n28810 & ~n28811 ;
  assign n28813 = \u1_R13_reg[2]/NET0131  & ~n28812 ;
  assign n28814 = ~\u1_R13_reg[2]/NET0131  & n28812 ;
  assign n28815 = ~n28813 & ~n28814 ;
  assign n28844 = n28802 & n28815 ;
  assign n28845 = ~n28809 & n28844 ;
  assign n28846 = n28824 & n28845 ;
  assign n28847 = n28796 & n28846 ;
  assign n28848 = ~n28815 & n28824 ;
  assign n28803 = ~n28796 & n28802 ;
  assign n28849 = ~n28803 & n28809 ;
  assign n28850 = n28848 & n28849 ;
  assign n28862 = ~n28847 & ~n28850 ;
  assign n28851 = n28809 & ~n28824 ;
  assign n28852 = n28796 & n28815 ;
  assign n28853 = n28851 & n28852 ;
  assign n28816 = ~n28809 & ~n28815 ;
  assign n28854 = n28816 & ~n28824 ;
  assign n28855 = ~n28853 & ~n28854 ;
  assign n28856 = n28802 & ~n28855 ;
  assign n28858 = ~n28802 & n28824 ;
  assign n28859 = n28815 & ~n28858 ;
  assign n28826 = ~n28802 & n28809 ;
  assign n28857 = ~n28796 & ~n28848 ;
  assign n28860 = ~n28826 & n28857 ;
  assign n28861 = ~n28859 & n28860 ;
  assign n28863 = ~n28856 & ~n28861 ;
  assign n28864 = n28862 & n28863 ;
  assign n28865 = ~n28842 & ~n28864 ;
  assign n28827 = ~n28809 & ~n28824 ;
  assign n28828 = n28815 & n28827 ;
  assign n28829 = ~n28826 & ~n28828 ;
  assign n28830 = n28796 & ~n28829 ;
  assign n28817 = ~n28802 & n28816 ;
  assign n28818 = ~n28803 & ~n28817 ;
  assign n28825 = ~n28818 & n28824 ;
  assign n28831 = n28796 & ~n28815 ;
  assign n28832 = n28802 & ~n28831 ;
  assign n28833 = ~n28816 & ~n28824 ;
  assign n28834 = ~n28832 & n28833 ;
  assign n28835 = ~n28825 & ~n28834 ;
  assign n28836 = ~n28830 & n28835 ;
  assign n28843 = ~n28836 & n28842 ;
  assign n28866 = ~n28802 & ~n28815 ;
  assign n28867 = ~n28802 & n28851 ;
  assign n28868 = ~n28816 & ~n28867 ;
  assign n28869 = ~n28866 & ~n28868 ;
  assign n28870 = n28809 & n28844 ;
  assign n28871 = n28824 & n28870 ;
  assign n28872 = ~n28869 & ~n28871 ;
  assign n28873 = ~n28796 & ~n28872 ;
  assign n28874 = n28796 & ~n28802 ;
  assign n28875 = ~n28828 & ~n28848 ;
  assign n28876 = n28874 & ~n28875 ;
  assign n28877 = ~n28873 & ~n28876 ;
  assign n28878 = ~n28843 & n28877 ;
  assign n28879 = ~n28865 & n28878 ;
  assign n28880 = ~\u1_L13_reg[31]/NET0131  & ~n28879 ;
  assign n28881 = \u1_L13_reg[31]/NET0131  & n28879 ;
  assign n28882 = ~n28880 & ~n28881 ;
  assign n28883 = decrypt_pad & ~\u1_uk_K_r13_reg[28]/NET0131  ;
  assign n28884 = ~decrypt_pad & ~\u1_uk_K_r13_reg[49]/NET0131  ;
  assign n28885 = ~n28883 & ~n28884 ;
  assign n28886 = \u1_R13_reg[28]/NET0131  & ~n28885 ;
  assign n28887 = ~\u1_R13_reg[28]/NET0131  & n28885 ;
  assign n28888 = ~n28886 & ~n28887 ;
  assign n28918 = decrypt_pad & ~\u1_uk_K_r13_reg[45]/NET0131  ;
  assign n28919 = ~decrypt_pad & ~\u1_uk_K_r13_reg[7]/NET0131  ;
  assign n28920 = ~n28918 & ~n28919 ;
  assign n28921 = \u1_R13_reg[27]/P0001  & ~n28920 ;
  assign n28922 = ~\u1_R13_reg[27]/P0001  & n28920 ;
  assign n28923 = ~n28921 & ~n28922 ;
  assign n28902 = decrypt_pad & ~\u1_uk_K_r13_reg[8]/NET0131  ;
  assign n28903 = ~decrypt_pad & ~\u1_uk_K_r13_reg[29]/NET0131  ;
  assign n28904 = ~n28902 & ~n28903 ;
  assign n28905 = \u1_R13_reg[26]/NET0131  & ~n28904 ;
  assign n28906 = ~\u1_R13_reg[26]/NET0131  & n28904 ;
  assign n28907 = ~n28905 & ~n28906 ;
  assign n28889 = decrypt_pad & ~\u1_uk_K_r13_reg[51]/NET0131  ;
  assign n28890 = ~decrypt_pad & ~\u1_uk_K_r13_reg[45]/NET0131  ;
  assign n28891 = ~n28889 & ~n28890 ;
  assign n28892 = \u1_R13_reg[29]/NET0131  & ~n28891 ;
  assign n28893 = ~\u1_R13_reg[29]/NET0131  & n28891 ;
  assign n28894 = ~n28892 & ~n28893 ;
  assign n28908 = decrypt_pad & ~\u1_uk_K_r13_reg[43]/NET0131  ;
  assign n28909 = ~decrypt_pad & ~\u1_uk_K_r13_reg[9]/NET0131  ;
  assign n28910 = ~n28908 & ~n28909 ;
  assign n28911 = \u1_R13_reg[24]/NET0131  & ~n28910 ;
  assign n28912 = ~\u1_R13_reg[24]/NET0131  & n28910 ;
  assign n28913 = ~n28911 & ~n28912 ;
  assign n28924 = n28894 & n28913 ;
  assign n28895 = decrypt_pad & ~\u1_uk_K_r13_reg[23]/NET0131  ;
  assign n28896 = ~decrypt_pad & ~\u1_uk_K_r13_reg[44]/NET0131  ;
  assign n28897 = ~n28895 & ~n28896 ;
  assign n28898 = \u1_R13_reg[25]/NET0131  & ~n28897 ;
  assign n28899 = ~\u1_R13_reg[25]/NET0131  & n28897 ;
  assign n28900 = ~n28898 & ~n28899 ;
  assign n28925 = ~n28894 & ~n28900 ;
  assign n28926 = ~n28913 & n28925 ;
  assign n28927 = ~n28924 & ~n28926 ;
  assign n28928 = n28907 & ~n28927 ;
  assign n28929 = ~n28894 & n28913 ;
  assign n28930 = n28900 & n28929 ;
  assign n28931 = ~n28928 & ~n28930 ;
  assign n28932 = ~n28923 & ~n28931 ;
  assign n28933 = n28894 & ~n28913 ;
  assign n28934 = ~n28923 & n28933 ;
  assign n28935 = n28913 & n28925 ;
  assign n28936 = ~n28934 & ~n28935 ;
  assign n28937 = ~n28907 & ~n28936 ;
  assign n28901 = n28894 & n28900 ;
  assign n28914 = ~n28907 & ~n28913 ;
  assign n28915 = n28907 & n28913 ;
  assign n28916 = ~n28914 & ~n28915 ;
  assign n28917 = n28901 & ~n28916 ;
  assign n28938 = n28913 & n28923 ;
  assign n28939 = ~n28900 & ~n28907 ;
  assign n28940 = n28938 & n28939 ;
  assign n28941 = ~n28917 & ~n28940 ;
  assign n28942 = ~n28937 & n28941 ;
  assign n28943 = ~n28932 & n28942 ;
  assign n28944 = ~n28888 & ~n28943 ;
  assign n28958 = ~n28900 & n28907 ;
  assign n28960 = n28901 & ~n28907 ;
  assign n28961 = ~n28958 & ~n28960 ;
  assign n28962 = n28938 & ~n28961 ;
  assign n28959 = n28933 & n28958 ;
  assign n28963 = n28914 & n28925 ;
  assign n28964 = ~n28959 & ~n28963 ;
  assign n28965 = ~n28962 & n28964 ;
  assign n28966 = n28888 & ~n28965 ;
  assign n28945 = n28900 & ~n28916 ;
  assign n28946 = n28924 & n28939 ;
  assign n28947 = n28901 & ~n28913 ;
  assign n28948 = ~n28946 & ~n28947 ;
  assign n28949 = n28888 & ~n28948 ;
  assign n28950 = ~n28945 & ~n28949 ;
  assign n28951 = ~n28923 & ~n28950 ;
  assign n28952 = n28907 & ~n28913 ;
  assign n28953 = ~n28901 & ~n28925 ;
  assign n28954 = n28952 & n28953 ;
  assign n28955 = n28925 & ~n28952 ;
  assign n28956 = ~n28954 & ~n28955 ;
  assign n28957 = n28923 & ~n28956 ;
  assign n28967 = ~n28951 & ~n28957 ;
  assign n28968 = ~n28966 & n28967 ;
  assign n28969 = ~n28944 & n28968 ;
  assign n28970 = \u1_L13_reg[22]/NET0131  & n28969 ;
  assign n28971 = ~\u1_L13_reg[22]/NET0131  & ~n28969 ;
  assign n28972 = ~n28970 & ~n28971 ;
  assign n28986 = decrypt_pad & ~\u1_uk_K_r13_reg[50]/NET0131  ;
  assign n28987 = ~decrypt_pad & ~\u1_uk_K_r13_reg[16]/NET0131  ;
  assign n28988 = ~n28986 & ~n28987 ;
  assign n28989 = \u1_R13_reg[23]/P0001  & ~n28988 ;
  assign n28990 = ~\u1_R13_reg[23]/P0001  & n28988 ;
  assign n28991 = ~n28989 & ~n28990 ;
  assign n28994 = decrypt_pad & ~\u1_uk_K_r13_reg[37]/NET0131  ;
  assign n28995 = ~decrypt_pad & ~\u1_uk_K_r13_reg[31]/NET0131  ;
  assign n28996 = ~n28994 & ~n28995 ;
  assign n28997 = \u1_R13_reg[22]/NET0131  & ~n28996 ;
  assign n28998 = ~\u1_R13_reg[22]/NET0131  & n28996 ;
  assign n28999 = ~n28997 & ~n28998 ;
  assign n28973 = decrypt_pad & ~\u1_uk_K_r13_reg[0]/NET0131  ;
  assign n28974 = ~decrypt_pad & ~\u1_uk_K_r13_reg[21]/NET0131  ;
  assign n28975 = ~n28973 & ~n28974 ;
  assign n28976 = \u1_R13_reg[20]/NET0131  & ~n28975 ;
  assign n28977 = ~\u1_R13_reg[20]/NET0131  & n28975 ;
  assign n28978 = ~n28976 & ~n28977 ;
  assign n28979 = decrypt_pad & ~\u1_uk_K_r13_reg[15]/NET0131  ;
  assign n28980 = ~decrypt_pad & ~\u1_uk_K_r13_reg[36]/NET0131  ;
  assign n28981 = ~n28979 & ~n28980 ;
  assign n28982 = \u1_R13_reg[21]/NET0131  & ~n28981 ;
  assign n28983 = ~\u1_R13_reg[21]/NET0131  & n28981 ;
  assign n28984 = ~n28982 & ~n28983 ;
  assign n28993 = ~n28978 & n28984 ;
  assign n29000 = decrypt_pad & ~\u1_uk_K_r13_reg[16]/NET0131  ;
  assign n29001 = ~decrypt_pad & ~\u1_uk_K_r13_reg[37]/NET0131  ;
  assign n29002 = ~n29000 & ~n29001 ;
  assign n29003 = \u1_R13_reg[25]/NET0131  & ~n29002 ;
  assign n29004 = ~\u1_R13_reg[25]/NET0131  & n29002 ;
  assign n29005 = ~n29003 & ~n29004 ;
  assign n29009 = n28978 & n29005 ;
  assign n29050 = ~n28993 & ~n29009 ;
  assign n29051 = n28999 & ~n29050 ;
  assign n29016 = ~n28984 & n29005 ;
  assign n29053 = n28978 & n29016 ;
  assign n29052 = n28993 & n29005 ;
  assign n29054 = ~n28999 & ~n29052 ;
  assign n29055 = ~n29053 & n29054 ;
  assign n29056 = ~n29051 & ~n29055 ;
  assign n29057 = ~n28991 & ~n29056 ;
  assign n29020 = decrypt_pad & ~\u1_uk_K_r13_reg[21]/NET0131  ;
  assign n29021 = ~decrypt_pad & ~\u1_uk_K_r13_reg[42]/NET0131  ;
  assign n29022 = ~n29020 & ~n29021 ;
  assign n29023 = \u1_R13_reg[24]/NET0131  & ~n29022 ;
  assign n29024 = ~\u1_R13_reg[24]/NET0131  & n29022 ;
  assign n29025 = ~n29023 & ~n29024 ;
  assign n29037 = ~n28978 & n28999 ;
  assign n29011 = n28984 & ~n29005 ;
  assign n29045 = n28978 & ~n29011 ;
  assign n29046 = ~n29037 & ~n29045 ;
  assign n29006 = ~n28999 & ~n29005 ;
  assign n29047 = ~n28984 & ~n29006 ;
  assign n29048 = ~n29046 & ~n29047 ;
  assign n29049 = n28991 & ~n29048 ;
  assign n29058 = n29025 & ~n29049 ;
  assign n29059 = ~n29057 & n29058 ;
  assign n29026 = n28978 & ~n28999 ;
  assign n29027 = n28984 & n29026 ;
  assign n29028 = ~n28991 & ~n28999 ;
  assign n29029 = n28978 & n29028 ;
  assign n29030 = ~n29027 & ~n29029 ;
  assign n29031 = ~n29005 & ~n29030 ;
  assign n29038 = ~n29026 & ~n29037 ;
  assign n29039 = n28984 & ~n28991 ;
  assign n29040 = ~n29038 & n29039 ;
  assign n29017 = n28991 & ~n28999 ;
  assign n29018 = ~n28978 & n29017 ;
  assign n29034 = ~n28991 & ~n29009 ;
  assign n29032 = ~n28984 & n28999 ;
  assign n29033 = ~n28978 & ~n29005 ;
  assign n29035 = n29032 & ~n29033 ;
  assign n29036 = ~n29034 & n29035 ;
  assign n29041 = ~n29018 & ~n29036 ;
  assign n29042 = ~n29040 & n29041 ;
  assign n29043 = ~n29031 & n29042 ;
  assign n29044 = ~n29025 & ~n29043 ;
  assign n29012 = ~n28978 & n29011 ;
  assign n29013 = ~n28999 & ~n29012 ;
  assign n29010 = n28999 & ~n29009 ;
  assign n29014 = n28991 & ~n29010 ;
  assign n29015 = ~n29013 & n29014 ;
  assign n28985 = n28978 & ~n28984 ;
  assign n28992 = ~n28985 & ~n28991 ;
  assign n29007 = ~n28993 & n29006 ;
  assign n29008 = n28992 & n29007 ;
  assign n29019 = n29016 & n29018 ;
  assign n29060 = ~n29008 & ~n29019 ;
  assign n29061 = ~n29015 & n29060 ;
  assign n29062 = ~n29044 & n29061 ;
  assign n29063 = ~n29059 & n29062 ;
  assign n29064 = ~\u1_L13_reg[11]/NET0131  & n29063 ;
  assign n29065 = \u1_L13_reg[11]/NET0131  & ~n29063 ;
  assign n29066 = ~n29064 & ~n29065 ;
  assign n29067 = n29005 & n29026 ;
  assign n29068 = n29025 & n29067 ;
  assign n29069 = n28978 & n29011 ;
  assign n29070 = ~n28978 & ~n29011 ;
  assign n29071 = ~n29016 & n29070 ;
  assign n29072 = ~n29069 & ~n29071 ;
  assign n29073 = n28999 & ~n29072 ;
  assign n29074 = ~n29068 & ~n29073 ;
  assign n29075 = n28991 & ~n29074 ;
  assign n29076 = n28984 & n29005 ;
  assign n29077 = n28999 & n29076 ;
  assign n29078 = n28991 & ~n29012 ;
  assign n29079 = ~n28999 & ~n29045 ;
  assign n29080 = ~n29078 & n29079 ;
  assign n29081 = ~n29077 & ~n29080 ;
  assign n29082 = n29025 & ~n29081 ;
  assign n29103 = ~n29075 & ~n29082 ;
  assign n29083 = ~n28978 & n29016 ;
  assign n29084 = n28999 & n29083 ;
  assign n29085 = ~n29012 & ~n29084 ;
  assign n29086 = ~n29025 & ~n29085 ;
  assign n29087 = ~n29011 & ~n29016 ;
  assign n29088 = n28978 & n29087 ;
  assign n29089 = ~n29006 & ~n29088 ;
  assign n29090 = ~n29026 & ~n29089 ;
  assign n29091 = ~n29086 & ~n29090 ;
  assign n29092 = ~n28991 & ~n29091 ;
  assign n29093 = n28985 & n29006 ;
  assign n29094 = ~n28991 & ~n29067 ;
  assign n29095 = n28984 & n28999 ;
  assign n29096 = n29005 & ~n29095 ;
  assign n29097 = n29038 & n29096 ;
  assign n29098 = ~n29028 & ~n29069 ;
  assign n29099 = ~n29097 & n29098 ;
  assign n29100 = ~n29094 & ~n29099 ;
  assign n29101 = ~n29093 & ~n29100 ;
  assign n29102 = ~n29025 & ~n29101 ;
  assign n29104 = ~n29092 & ~n29102 ;
  assign n29105 = n29103 & n29104 ;
  assign n29106 = ~\u1_L13_reg[4]/NET0131  & ~n29105 ;
  assign n29107 = \u1_L13_reg[4]/NET0131  & n29105 ;
  assign n29108 = ~n29106 & ~n29107 ;
  assign n29121 = n28809 & n28824 ;
  assign n29130 = ~n28827 & ~n29121 ;
  assign n29131 = ~n28802 & ~n29130 ;
  assign n29132 = ~n28854 & ~n29131 ;
  assign n29133 = ~n28796 & ~n29132 ;
  assign n29134 = n28815 & n28867 ;
  assign n29135 = ~n28846 & ~n29134 ;
  assign n29136 = ~n29133 & n29135 ;
  assign n29137 = ~n28842 & ~n29136 ;
  assign n29109 = ~n28815 & n28851 ;
  assign n29110 = ~n28828 & ~n29109 ;
  assign n29111 = n28802 & ~n29110 ;
  assign n29112 = ~n28809 & n28858 ;
  assign n29113 = n28802 & n28824 ;
  assign n29114 = n28809 & n29113 ;
  assign n29115 = ~n29112 & ~n29114 ;
  assign n29116 = ~n28842 & ~n29115 ;
  assign n29117 = ~n29111 & ~n29116 ;
  assign n29118 = n28796 & ~n29117 ;
  assign n29120 = ~n28824 & ~n28866 ;
  assign n29122 = n28866 & n29121 ;
  assign n29123 = ~n29120 & ~n29122 ;
  assign n29124 = n28796 & ~n29123 ;
  assign n29125 = n28857 & ~n29120 ;
  assign n29119 = n28816 & n29113 ;
  assign n29126 = ~n28870 & ~n29119 ;
  assign n29127 = ~n29125 & n29126 ;
  assign n29128 = ~n29124 & n29127 ;
  assign n29129 = n28842 & ~n29128 ;
  assign n29138 = ~n29118 & ~n29129 ;
  assign n29139 = ~n29137 & n29138 ;
  assign n29140 = ~\u1_L13_reg[17]/NET0131  & ~n29139 ;
  assign n29141 = \u1_L13_reg[17]/NET0131  & n29139 ;
  assign n29142 = ~n29140 & ~n29141 ;
  assign n29156 = decrypt_pad & ~\u1_uk_K_r13_reg[18]/NET0131  ;
  assign n29157 = ~decrypt_pad & ~\u1_uk_K_r13_reg[39]/NET0131  ;
  assign n29158 = ~n29156 & ~n29157 ;
  assign n29159 = \u1_R13_reg[15]/NET0131  & ~n29158 ;
  assign n29160 = ~\u1_R13_reg[15]/NET0131  & n29158 ;
  assign n29161 = ~n29159 & ~n29160 ;
  assign n29179 = decrypt_pad & ~\u1_uk_K_r13_reg[10]/NET0131  ;
  assign n29180 = ~decrypt_pad & ~\u1_uk_K_r13_reg[6]/NET0131  ;
  assign n29181 = ~n29179 & ~n29180 ;
  assign n29182 = \u1_R13_reg[14]/NET0131  & ~n29181 ;
  assign n29183 = ~\u1_R13_reg[14]/NET0131  & n29181 ;
  assign n29184 = ~n29182 & ~n29183 ;
  assign n29195 = ~n29161 & ~n29184 ;
  assign n29143 = decrypt_pad & ~\u1_uk_K_r13_reg[47]/NET0131  ;
  assign n29144 = ~decrypt_pad & ~\u1_uk_K_r13_reg[11]/NET0131  ;
  assign n29145 = ~n29143 & ~n29144 ;
  assign n29146 = \u1_R13_reg[12]/NET0131  & ~n29145 ;
  assign n29147 = ~\u1_R13_reg[12]/NET0131  & n29145 ;
  assign n29148 = ~n29146 & ~n29147 ;
  assign n29162 = decrypt_pad & ~\u1_uk_K_r13_reg[41]/NET0131  ;
  assign n29163 = ~decrypt_pad & ~\u1_uk_K_r13_reg[5]/NET0131  ;
  assign n29164 = ~n29162 & ~n29163 ;
  assign n29165 = \u1_R13_reg[13]/NET0131  & ~n29164 ;
  assign n29166 = ~\u1_R13_reg[13]/NET0131  & n29164 ;
  assign n29167 = ~n29165 & ~n29166 ;
  assign n29196 = ~n29148 & n29167 ;
  assign n29197 = n29148 & ~n29167 ;
  assign n29198 = ~n29196 & ~n29197 ;
  assign n29199 = n29195 & ~n29198 ;
  assign n29149 = decrypt_pad & ~\u1_uk_K_r13_reg[6]/NET0131  ;
  assign n29150 = ~decrypt_pad & ~\u1_uk_K_r13_reg[27]/NET0131  ;
  assign n29151 = ~n29149 & ~n29150 ;
  assign n29152 = \u1_R13_reg[17]/NET0131  & ~n29151 ;
  assign n29153 = ~\u1_R13_reg[17]/NET0131  & n29151 ;
  assign n29154 = ~n29152 & ~n29153 ;
  assign n29186 = ~n29148 & n29154 ;
  assign n29193 = n29161 & n29186 ;
  assign n29194 = ~n29167 & n29193 ;
  assign n29155 = n29148 & ~n29154 ;
  assign n29168 = n29161 & n29167 ;
  assign n29169 = n29155 & n29168 ;
  assign n29170 = decrypt_pad & ~\u1_uk_K_r13_reg[26]/NET0131  ;
  assign n29171 = ~decrypt_pad & ~\u1_uk_K_r13_reg[47]/NET0131  ;
  assign n29172 = ~n29170 & ~n29171 ;
  assign n29173 = \u1_R13_reg[16]/NET0131  & ~n29172 ;
  assign n29174 = ~\u1_R13_reg[16]/NET0131  & n29172 ;
  assign n29175 = ~n29173 & ~n29174 ;
  assign n29200 = ~n29169 & n29175 ;
  assign n29201 = ~n29194 & n29200 ;
  assign n29202 = ~n29199 & n29201 ;
  assign n29176 = ~n29154 & ~n29167 ;
  assign n29177 = ~n29148 & n29176 ;
  assign n29178 = ~n29161 & n29177 ;
  assign n29185 = n29178 & n29184 ;
  assign n29187 = n29167 & ~n29184 ;
  assign n29188 = n29186 & n29187 ;
  assign n29189 = n29148 & n29154 ;
  assign n29190 = n29167 & n29189 ;
  assign n29191 = n29184 & n29190 ;
  assign n29192 = ~n29188 & ~n29191 ;
  assign n29203 = ~n29185 & n29192 ;
  assign n29204 = n29202 & n29203 ;
  assign n29206 = n29161 & n29177 ;
  assign n29205 = n29168 & n29189 ;
  assign n29219 = ~n29175 & ~n29205 ;
  assign n29220 = ~n29206 & n29219 ;
  assign n29207 = ~n29167 & n29189 ;
  assign n29208 = ~n29184 & n29207 ;
  assign n29209 = n29168 & n29184 ;
  assign n29210 = ~n29148 & n29209 ;
  assign n29221 = ~n29208 & ~n29210 ;
  assign n29222 = n29220 & n29221 ;
  assign n29211 = ~n29154 & n29196 ;
  assign n29212 = n29184 & n29211 ;
  assign n29213 = n29177 & ~n29184 ;
  assign n29214 = ~n29212 & ~n29213 ;
  assign n29215 = n29155 & n29184 ;
  assign n29216 = n29154 & ~n29167 ;
  assign n29217 = ~n29215 & ~n29216 ;
  assign n29218 = ~n29161 & ~n29217 ;
  assign n29223 = n29214 & ~n29218 ;
  assign n29224 = n29222 & n29223 ;
  assign n29225 = ~n29204 & ~n29224 ;
  assign n29226 = ~n29161 & ~n29188 ;
  assign n29227 = ~n29167 & n29184 ;
  assign n29228 = n29155 & n29227 ;
  assign n29229 = n29161 & ~n29228 ;
  assign n29230 = ~n29213 & n29229 ;
  assign n29231 = ~n29226 & ~n29230 ;
  assign n29232 = n29155 & ~n29184 ;
  assign n29233 = n29168 & n29232 ;
  assign n29234 = ~n29231 & ~n29233 ;
  assign n29235 = ~n29225 & n29234 ;
  assign n29236 = ~\u1_L13_reg[20]/NET0131  & ~n29235 ;
  assign n29237 = \u1_L13_reg[20]/NET0131  & n29235 ;
  assign n29238 = ~n29236 & ~n29237 ;
  assign n29275 = decrypt_pad & ~\u1_uk_K_r13_reg[25]/P0001  ;
  assign n29276 = ~decrypt_pad & ~\u1_uk_K_r13_reg[46]/NET0131  ;
  assign n29277 = ~n29275 & ~n29276 ;
  assign n29278 = \u1_R13_reg[8]/NET0131  & ~n29277 ;
  assign n29279 = ~\u1_R13_reg[8]/NET0131  & n29277 ;
  assign n29280 = ~n29278 & ~n29279 ;
  assign n29245 = decrypt_pad & ~\u1_uk_K_r13_reg[40]/NET0131  ;
  assign n29246 = ~decrypt_pad & ~\u1_uk_K_r13_reg[4]/NET0131  ;
  assign n29247 = ~n29245 & ~n29246 ;
  assign n29248 = \u1_R13_reg[6]/NET0131  & ~n29247 ;
  assign n29249 = ~\u1_R13_reg[6]/NET0131  & n29247 ;
  assign n29250 = ~n29248 & ~n29249 ;
  assign n29260 = decrypt_pad & ~\u1_uk_K_r13_reg[13]/NET0131  ;
  assign n29261 = ~decrypt_pad & ~\u1_uk_K_r13_reg[34]/NET0131  ;
  assign n29262 = ~n29260 & ~n29261 ;
  assign n29263 = \u1_R13_reg[4]/NET0131  & ~n29262 ;
  assign n29264 = ~\u1_R13_reg[4]/NET0131  & n29262 ;
  assign n29265 = ~n29263 & ~n29264 ;
  assign n29239 = decrypt_pad & ~\u1_uk_K_r13_reg[17]/NET0131  ;
  assign n29240 = ~decrypt_pad & ~\u1_uk_K_r13_reg[13]/NET0131  ;
  assign n29241 = ~n29239 & ~n29240 ;
  assign n29242 = \u1_R13_reg[5]/NET0131  & ~n29241 ;
  assign n29243 = ~\u1_R13_reg[5]/NET0131  & n29241 ;
  assign n29244 = ~n29242 & ~n29243 ;
  assign n29254 = decrypt_pad & ~\u1_uk_K_r13_reg[5]/NET0131  ;
  assign n29255 = ~decrypt_pad & ~\u1_uk_K_r13_reg[26]/NET0131  ;
  assign n29256 = ~n29254 & ~n29255 ;
  assign n29257 = \u1_R13_reg[9]/NET0131  & ~n29256 ;
  assign n29258 = ~\u1_R13_reg[9]/NET0131  & n29256 ;
  assign n29259 = ~n29257 & ~n29258 ;
  assign n29284 = ~n29244 & n29259 ;
  assign n29306 = ~n29265 & n29284 ;
  assign n29309 = n29244 & ~n29259 ;
  assign n29310 = ~n29306 & ~n29309 ;
  assign n29311 = ~n29250 & ~n29310 ;
  assign n29291 = n29250 & ~n29265 ;
  assign n29267 = decrypt_pad & ~\u1_uk_K_r13_reg[34]/NET0131  ;
  assign n29268 = ~decrypt_pad & ~\u1_uk_K_r13_reg[55]/NET0131  ;
  assign n29269 = ~n29267 & ~n29268 ;
  assign n29270 = \u1_R13_reg[7]/NET0131  & ~n29269 ;
  assign n29271 = ~\u1_R13_reg[7]/NET0131  & n29269 ;
  assign n29272 = ~n29270 & ~n29271 ;
  assign n29301 = ~n29244 & ~n29272 ;
  assign n29302 = ~n29291 & ~n29301 ;
  assign n29252 = ~n29244 & n29250 ;
  assign n29303 = ~n29252 & n29259 ;
  assign n29304 = ~n29302 & n29303 ;
  assign n29285 = n29250 & n29265 ;
  assign n29305 = ~n29284 & n29285 ;
  assign n29307 = ~n29305 & ~n29306 ;
  assign n29308 = ~n29272 & ~n29307 ;
  assign n29312 = ~n29304 & ~n29308 ;
  assign n29313 = ~n29311 & n29312 ;
  assign n29314 = ~n29280 & ~n29313 ;
  assign n29286 = n29284 & n29285 ;
  assign n29251 = n29244 & ~n29250 ;
  assign n29287 = ~n29259 & ~n29265 ;
  assign n29288 = ~n29251 & n29287 ;
  assign n29289 = ~n29286 & ~n29288 ;
  assign n29290 = ~n29272 & ~n29289 ;
  assign n29294 = ~n29259 & n29265 ;
  assign n29295 = ~n29250 & n29294 ;
  assign n29296 = ~n29244 & n29295 ;
  assign n29281 = n29244 & n29265 ;
  assign n29282 = ~n29250 & n29281 ;
  assign n29283 = n29259 & n29282 ;
  assign n29292 = n29244 & n29272 ;
  assign n29293 = ~n29291 & n29292 ;
  assign n29297 = ~n29283 & ~n29293 ;
  assign n29298 = ~n29296 & n29297 ;
  assign n29299 = ~n29290 & n29298 ;
  assign n29300 = n29280 & ~n29299 ;
  assign n29253 = ~n29251 & ~n29252 ;
  assign n29266 = n29259 & ~n29265 ;
  assign n29273 = n29266 & ~n29272 ;
  assign n29274 = n29253 & n29273 ;
  assign n29317 = ~n29280 & n29286 ;
  assign n29315 = n29252 & ~n29265 ;
  assign n29316 = ~n29259 & n29315 ;
  assign n29318 = ~n29282 & ~n29316 ;
  assign n29319 = ~n29317 & n29318 ;
  assign n29320 = n29272 & ~n29319 ;
  assign n29321 = ~n29274 & ~n29320 ;
  assign n29322 = ~n29300 & n29321 ;
  assign n29323 = ~n29314 & n29322 ;
  assign n29324 = \u1_L13_reg[2]/NET0131  & n29323 ;
  assign n29325 = ~\u1_L13_reg[2]/NET0131  & ~n29323 ;
  assign n29326 = ~n29324 & ~n29325 ;
  assign n29327 = n28984 & ~n29037 ;
  assign n29328 = ~n29009 & ~n29026 ;
  assign n29329 = n29327 & n29328 ;
  assign n29330 = n29094 & ~n29329 ;
  assign n29331 = ~n29005 & ~n29032 ;
  assign n29332 = ~n29327 & n29331 ;
  assign n29333 = n28991 & ~n29088 ;
  assign n29334 = ~n29332 & n29333 ;
  assign n29335 = ~n29330 & ~n29334 ;
  assign n29336 = ~n29025 & ~n29084 ;
  assign n29337 = ~n29335 & n29336 ;
  assign n29343 = ~n29052 & ~n29329 ;
  assign n29344 = n28991 & ~n29343 ;
  assign n29340 = n29010 & ~n29033 ;
  assign n29338 = ~n28999 & ~n29050 ;
  assign n29339 = n28991 & ~n29047 ;
  assign n29341 = ~n29338 & ~n29339 ;
  assign n29342 = ~n29340 & n29341 ;
  assign n29345 = n29025 & ~n29342 ;
  assign n29346 = ~n29344 & n29345 ;
  assign n29347 = ~n29337 & ~n29346 ;
  assign n29348 = n29017 & n29076 ;
  assign n29349 = ~n29093 & ~n29348 ;
  assign n29350 = ~n29347 & n29349 ;
  assign n29351 = \u1_L13_reg[29]/NET0131  & ~n29350 ;
  assign n29352 = ~\u1_L13_reg[29]/NET0131  & n29350 ;
  assign n29353 = ~n29351 & ~n29352 ;
  assign n29408 = decrypt_pad & ~\u1_uk_K_r13_reg[52]/P0001  ;
  assign n29409 = ~decrypt_pad & ~\u1_uk_K_r13_reg[14]/NET0131  ;
  assign n29410 = ~n29408 & ~n29409 ;
  assign n29411 = \u1_R13_reg[32]/NET0131  & ~n29410 ;
  assign n29412 = ~\u1_R13_reg[32]/NET0131  & n29410 ;
  assign n29413 = ~n29411 & ~n29412 ;
  assign n29354 = decrypt_pad & ~\u1_uk_K_r13_reg[42]/NET0131  ;
  assign n29355 = ~decrypt_pad & ~\u1_uk_K_r13_reg[8]/NET0131  ;
  assign n29356 = ~n29354 & ~n29355 ;
  assign n29357 = \u1_R13_reg[31]/P0001  & ~n29356 ;
  assign n29358 = ~\u1_R13_reg[31]/P0001  & n29356 ;
  assign n29359 = ~n29357 & ~n29358 ;
  assign n29360 = decrypt_pad & ~\u1_uk_K_r13_reg[30]/NET0131  ;
  assign n29361 = ~decrypt_pad & ~\u1_uk_K_r13_reg[51]/NET0131  ;
  assign n29362 = ~n29360 & ~n29361 ;
  assign n29363 = \u1_R13_reg[30]/NET0131  & ~n29362 ;
  assign n29364 = ~\u1_R13_reg[30]/NET0131  & n29362 ;
  assign n29365 = ~n29363 & ~n29364 ;
  assign n29367 = decrypt_pad & ~\u1_uk_K_r13_reg[29]/NET0131  ;
  assign n29368 = ~decrypt_pad & ~\u1_uk_K_r13_reg[50]/NET0131  ;
  assign n29369 = ~n29367 & ~n29368 ;
  assign n29370 = \u1_R13_reg[29]/NET0131  & ~n29369 ;
  assign n29371 = ~\u1_R13_reg[29]/NET0131  & n29369 ;
  assign n29372 = ~n29370 & ~n29371 ;
  assign n29382 = decrypt_pad & ~\u1_uk_K_r13_reg[2]/NET0131  ;
  assign n29383 = ~decrypt_pad & ~\u1_uk_K_r13_reg[23]/NET0131  ;
  assign n29384 = ~n29382 & ~n29383 ;
  assign n29385 = \u1_R13_reg[28]/NET0131  & ~n29384 ;
  assign n29386 = ~\u1_R13_reg[28]/NET0131  & n29384 ;
  assign n29387 = ~n29385 & ~n29386 ;
  assign n29389 = ~n29372 & n29387 ;
  assign n29374 = decrypt_pad & ~\u1_uk_K_r13_reg[14]/NET0131  ;
  assign n29375 = ~decrypt_pad & ~\u1_uk_K_r13_reg[35]/NET0131  ;
  assign n29376 = ~n29374 & ~n29375 ;
  assign n29377 = \u1_R13_reg[1]/NET0131  & ~n29376 ;
  assign n29378 = ~\u1_R13_reg[1]/NET0131  & n29376 ;
  assign n29379 = ~n29377 & ~n29378 ;
  assign n29396 = n29379 & n29387 ;
  assign n29436 = ~n29389 & ~n29396 ;
  assign n29437 = ~n29365 & ~n29436 ;
  assign n29397 = n29365 & n29372 ;
  assign n29435 = ~n29379 & n29397 ;
  assign n29428 = ~n29379 & ~n29387 ;
  assign n29438 = n29372 & n29428 ;
  assign n29439 = ~n29435 & ~n29438 ;
  assign n29440 = ~n29437 & n29439 ;
  assign n29441 = n29359 & ~n29440 ;
  assign n29421 = ~n29387 & n29397 ;
  assign n29434 = n29379 & n29421 ;
  assign n29423 = ~n29365 & ~n29372 ;
  assign n29442 = ~n29387 & n29423 ;
  assign n29443 = ~n29359 & n29442 ;
  assign n29444 = ~n29434 & ~n29443 ;
  assign n29445 = ~n29441 & n29444 ;
  assign n29446 = n29413 & ~n29445 ;
  assign n29390 = n29365 & n29389 ;
  assign n29391 = ~n29379 & n29390 ;
  assign n29392 = n29379 & ~n29387 ;
  assign n29393 = ~n29372 & n29392 ;
  assign n29394 = ~n29391 & ~n29393 ;
  assign n29395 = n29359 & ~n29394 ;
  assign n29366 = ~n29359 & ~n29365 ;
  assign n29373 = ~n29365 & n29372 ;
  assign n29380 = n29373 & ~n29379 ;
  assign n29381 = ~n29366 & ~n29380 ;
  assign n29388 = ~n29381 & n29387 ;
  assign n29398 = n29396 & n29397 ;
  assign n29399 = ~n29379 & n29387 ;
  assign n29402 = ~n29359 & ~n29399 ;
  assign n29400 = ~n29365 & ~n29379 ;
  assign n29401 = ~n29372 & n29379 ;
  assign n29403 = ~n29400 & ~n29401 ;
  assign n29404 = n29402 & n29403 ;
  assign n29405 = ~n29398 & ~n29404 ;
  assign n29406 = ~n29388 & n29405 ;
  assign n29407 = ~n29395 & n29406 ;
  assign n29414 = ~n29407 & ~n29413 ;
  assign n29422 = ~n29379 & n29421 ;
  assign n29424 = n29379 & n29423 ;
  assign n29425 = n29387 & n29424 ;
  assign n29426 = ~n29422 & ~n29425 ;
  assign n29427 = n29365 & n29393 ;
  assign n29429 = ~n29372 & n29428 ;
  assign n29430 = ~n29365 & n29429 ;
  assign n29431 = ~n29427 & ~n29430 ;
  assign n29432 = n29426 & n29431 ;
  assign n29433 = n29359 & ~n29432 ;
  assign n29415 = ~n29359 & n29365 ;
  assign n29416 = n29389 & n29413 ;
  assign n29417 = n29415 & n29416 ;
  assign n29418 = n29372 & n29387 ;
  assign n29419 = ~n29379 & n29418 ;
  assign n29420 = n29366 & n29419 ;
  assign n29447 = ~n29417 & ~n29420 ;
  assign n29448 = ~n29433 & n29447 ;
  assign n29449 = ~n29414 & n29448 ;
  assign n29450 = ~n29446 & n29449 ;
  assign n29451 = \u1_L13_reg[5]/NET0131  & ~n29450 ;
  assign n29452 = ~\u1_L13_reg[5]/NET0131  & n29450 ;
  assign n29453 = ~n29451 & ~n29452 ;
  assign n29454 = n29285 & n29309 ;
  assign n29455 = ~n29283 & ~n29454 ;
  assign n29456 = ~n29265 & n29309 ;
  assign n29457 = n29284 & n29291 ;
  assign n29458 = ~n29456 & ~n29457 ;
  assign n29459 = ~n29296 & n29458 ;
  assign n29460 = ~n29280 & ~n29459 ;
  assign n29461 = n29455 & ~n29460 ;
  assign n29462 = ~n29272 & ~n29461 ;
  assign n29464 = ~n29250 & ~n29259 ;
  assign n29465 = ~n29244 & ~n29266 ;
  assign n29466 = ~n29464 & n29465 ;
  assign n29467 = ~n29272 & ~n29466 ;
  assign n29469 = n29250 & n29266 ;
  assign n29468 = ~n29244 & n29464 ;
  assign n29470 = n29272 & ~n29468 ;
  assign n29471 = ~n29469 & n29470 ;
  assign n29472 = ~n29467 & ~n29471 ;
  assign n29463 = ~n29250 & n29456 ;
  assign n29473 = n29280 & ~n29304 ;
  assign n29474 = ~n29463 & n29473 ;
  assign n29475 = n29455 & n29474 ;
  assign n29476 = ~n29472 & n29475 ;
  assign n29480 = ~n29294 & ~n29465 ;
  assign n29479 = ~n29251 & n29294 ;
  assign n29481 = n29272 & ~n29479 ;
  assign n29482 = ~n29480 & n29481 ;
  assign n29483 = n29272 & n29285 ;
  assign n29484 = ~n29309 & n29483 ;
  assign n29477 = ~n29250 & n29266 ;
  assign n29478 = ~n29301 & n29477 ;
  assign n29485 = ~n29280 & ~n29478 ;
  assign n29486 = ~n29484 & n29485 ;
  assign n29487 = ~n29482 & n29486 ;
  assign n29488 = ~n29476 & ~n29487 ;
  assign n29489 = ~n29462 & ~n29488 ;
  assign n29490 = ~\u1_L13_reg[13]/NET0131  & n29489 ;
  assign n29491 = \u1_L13_reg[13]/NET0131  & ~n29489 ;
  assign n29492 = ~n29490 & ~n29491 ;
  assign n29493 = decrypt_pad & ~\u1_uk_K_r13_reg[49]/NET0131  ;
  assign n29494 = ~decrypt_pad & ~\u1_uk_K_r13_reg[15]/NET0131  ;
  assign n29495 = ~n29493 & ~n29494 ;
  assign n29496 = \u1_R13_reg[19]/NET0131  & ~n29495 ;
  assign n29497 = ~\u1_R13_reg[19]/NET0131  & n29495 ;
  assign n29498 = ~n29496 & ~n29497 ;
  assign n29499 = decrypt_pad & ~\u1_uk_K_r13_reg[22]/NET0131  ;
  assign n29500 = ~decrypt_pad & ~\u1_uk_K_r13_reg[43]/NET0131  ;
  assign n29501 = ~n29499 & ~n29500 ;
  assign n29502 = \u1_R13_reg[16]/NET0131  & ~n29501 ;
  assign n29503 = ~\u1_R13_reg[16]/NET0131  & n29501 ;
  assign n29504 = ~n29502 & ~n29503 ;
  assign n29505 = decrypt_pad & ~\u1_uk_K_r13_reg[38]/NET0131  ;
  assign n29506 = ~decrypt_pad & ~\u1_uk_K_r13_reg[0]/NET0131  ;
  assign n29507 = ~n29505 & ~n29506 ;
  assign n29508 = \u1_R13_reg[21]/NET0131  & ~n29507 ;
  assign n29509 = ~\u1_R13_reg[21]/NET0131  & n29507 ;
  assign n29510 = ~n29508 & ~n29509 ;
  assign n29512 = decrypt_pad & ~\u1_uk_K_r13_reg[44]/NET0131  ;
  assign n29513 = ~decrypt_pad & ~\u1_uk_K_r13_reg[38]/NET0131  ;
  assign n29514 = ~n29512 & ~n29513 ;
  assign n29515 = \u1_R13_reg[17]/NET0131  & ~n29514 ;
  assign n29516 = ~\u1_R13_reg[17]/NET0131  & n29514 ;
  assign n29517 = ~n29515 & ~n29516 ;
  assign n29519 = decrypt_pad & ~\u1_uk_K_r13_reg[7]/NET0131  ;
  assign n29520 = ~decrypt_pad & ~\u1_uk_K_r13_reg[28]/NET0131  ;
  assign n29521 = ~n29519 & ~n29520 ;
  assign n29522 = \u1_R13_reg[18]/NET0131  & ~n29521 ;
  assign n29523 = ~\u1_R13_reg[18]/NET0131  & n29521 ;
  assign n29524 = ~n29522 & ~n29523 ;
  assign n29530 = n29517 & ~n29524 ;
  assign n29531 = n29510 & n29530 ;
  assign n29532 = n29504 & n29531 ;
  assign n29511 = n29504 & ~n29510 ;
  assign n29518 = n29511 & ~n29517 ;
  assign n29525 = n29518 & ~n29524 ;
  assign n29526 = ~n29504 & n29510 ;
  assign n29527 = ~n29517 & n29526 ;
  assign n29528 = ~n29510 & n29517 ;
  assign n29529 = n29524 & n29528 ;
  assign n29533 = ~n29527 & ~n29529 ;
  assign n29534 = ~n29525 & n29533 ;
  assign n29535 = ~n29532 & n29534 ;
  assign n29536 = ~n29498 & ~n29535 ;
  assign n29544 = n29510 & n29524 ;
  assign n29545 = n29504 & n29544 ;
  assign n29540 = ~n29504 & n29530 ;
  assign n29542 = ~n29504 & ~n29510 ;
  assign n29543 = ~n29517 & n29542 ;
  assign n29546 = ~n29540 & ~n29543 ;
  assign n29547 = ~n29545 & n29546 ;
  assign n29548 = n29498 & ~n29547 ;
  assign n29537 = n29504 & n29510 ;
  assign n29538 = ~n29517 & n29524 ;
  assign n29539 = n29537 & n29538 ;
  assign n29541 = ~n29510 & n29540 ;
  assign n29549 = ~n29539 & ~n29541 ;
  assign n29550 = ~n29548 & n29549 ;
  assign n29551 = ~n29536 & n29550 ;
  assign n29552 = decrypt_pad & ~\u1_uk_K_r13_reg[9]/NET0131  ;
  assign n29553 = ~decrypt_pad & ~\u1_uk_K_r13_reg[30]/NET0131  ;
  assign n29554 = ~n29552 & ~n29553 ;
  assign n29555 = \u1_R13_reg[20]/NET0131  & ~n29554 ;
  assign n29556 = ~\u1_R13_reg[20]/NET0131  & n29554 ;
  assign n29557 = ~n29555 & ~n29556 ;
  assign n29558 = ~n29551 & ~n29557 ;
  assign n29563 = n29504 & n29528 ;
  assign n29561 = ~n29524 & n29537 ;
  assign n29562 = n29526 & ~n29530 ;
  assign n29564 = ~n29561 & ~n29562 ;
  assign n29565 = ~n29563 & n29564 ;
  assign n29566 = n29498 & ~n29565 ;
  assign n29567 = ~n29498 & ~n29524 ;
  assign n29568 = n29517 & n29526 ;
  assign n29569 = ~n29543 & ~n29568 ;
  assign n29570 = n29567 & ~n29569 ;
  assign n29559 = ~n29530 & ~n29538 ;
  assign n29560 = n29511 & ~n29559 ;
  assign n29571 = n29498 & n29517 ;
  assign n29572 = n29537 & ~n29571 ;
  assign n29573 = n29559 & n29572 ;
  assign n29574 = ~n29560 & ~n29573 ;
  assign n29575 = ~n29570 & n29574 ;
  assign n29576 = ~n29566 & n29575 ;
  assign n29577 = n29557 & ~n29576 ;
  assign n29578 = ~n29524 & n29563 ;
  assign n29579 = n29524 & n29543 ;
  assign n29580 = ~n29578 & ~n29579 ;
  assign n29581 = n29498 & ~n29580 ;
  assign n29582 = n29526 & n29538 ;
  assign n29583 = ~n29504 & n29524 ;
  assign n29584 = n29528 & n29583 ;
  assign n29585 = ~n29582 & ~n29584 ;
  assign n29586 = ~n29498 & ~n29585 ;
  assign n29587 = ~n29581 & ~n29586 ;
  assign n29588 = ~n29577 & n29587 ;
  assign n29589 = ~n29558 & n29588 ;
  assign n29590 = ~\u1_L13_reg[14]/NET0131  & ~n29589 ;
  assign n29591 = \u1_L13_reg[14]/NET0131  & n29589 ;
  assign n29592 = ~n29590 & ~n29591 ;
  assign n29616 = n29365 & n29418 ;
  assign n29615 = n29372 & n29392 ;
  assign n29617 = ~n29424 & ~n29615 ;
  assign n29618 = ~n29616 & n29617 ;
  assign n29619 = n29359 & ~n29618 ;
  assign n29609 = n29379 & n29390 ;
  assign n29610 = n29387 & n29400 ;
  assign n29611 = ~n29609 & ~n29610 ;
  assign n29612 = ~n29359 & ~n29611 ;
  assign n29613 = ~n29419 & ~n29429 ;
  assign n29614 = n29365 & ~n29613 ;
  assign n29620 = ~n29365 & n29393 ;
  assign n29621 = ~n29614 & ~n29620 ;
  assign n29622 = ~n29612 & n29621 ;
  assign n29623 = ~n29619 & n29622 ;
  assign n29624 = n29413 & ~n29623 ;
  assign n29598 = ~n29359 & n29438 ;
  assign n29596 = ~n29366 & ~n29373 ;
  assign n29597 = n29396 & ~n29596 ;
  assign n29601 = ~n29430 & ~n29597 ;
  assign n29602 = ~n29598 & n29601 ;
  assign n29593 = ~n29390 & ~n29419 ;
  assign n29594 = n29359 & ~n29593 ;
  assign n29595 = n29392 & n29415 ;
  assign n29599 = ~n29421 & ~n29595 ;
  assign n29600 = ~n29391 & n29599 ;
  assign n29603 = ~n29594 & n29600 ;
  assign n29604 = n29602 & n29603 ;
  assign n29605 = ~n29413 & ~n29604 ;
  assign n29606 = n29359 & n29442 ;
  assign n29607 = n29372 & n29396 ;
  assign n29608 = n29366 & n29607 ;
  assign n29625 = ~n29606 & ~n29608 ;
  assign n29626 = ~n29605 & n29625 ;
  assign n29627 = ~n29624 & n29626 ;
  assign n29628 = ~\u1_L13_reg[21]/NET0131  & ~n29627 ;
  assign n29629 = \u1_L13_reg[21]/NET0131  & n29627 ;
  assign n29630 = ~n29628 & ~n29629 ;
  assign n29641 = ~n29176 & ~n29227 ;
  assign n29642 = n29161 & ~n29641 ;
  assign n29643 = n29154 & n29195 ;
  assign n29644 = ~n29187 & ~n29643 ;
  assign n29645 = ~n29642 & n29644 ;
  assign n29646 = n29148 & ~n29645 ;
  assign n29647 = ~n29184 & n29193 ;
  assign n29648 = ~n29178 & ~n29647 ;
  assign n29649 = n29214 & n29648 ;
  assign n29650 = ~n29646 & n29649 ;
  assign n29651 = ~n29175 & ~n29650 ;
  assign n29631 = ~n29148 & n29227 ;
  assign n29632 = n29154 & n29631 ;
  assign n29633 = ~n29191 & ~n29632 ;
  assign n29634 = n29155 & ~n29187 ;
  assign n29635 = n29226 & ~n29634 ;
  assign n29636 = n29161 & ~n29211 ;
  assign n29637 = ~n29208 & n29636 ;
  assign n29638 = ~n29635 & ~n29637 ;
  assign n29639 = n29633 & ~n29638 ;
  assign n29640 = n29175 & ~n29639 ;
  assign n29652 = ~n29213 & n29633 ;
  assign n29653 = ~n29161 & ~n29652 ;
  assign n29654 = ~n29210 & ~n29233 ;
  assign n29655 = ~n29653 & n29654 ;
  assign n29656 = ~n29640 & n29655 ;
  assign n29657 = ~n29651 & n29656 ;
  assign n29658 = \u1_L13_reg[10]/NET0131  & n29657 ;
  assign n29659 = ~\u1_L13_reg[10]/NET0131  & ~n29657 ;
  assign n29660 = ~n29658 & ~n29659 ;
  assign n29661 = n28929 & n28939 ;
  assign n29672 = ~n28888 & ~n29661 ;
  assign n29662 = n28915 & ~n28923 ;
  assign n29663 = ~n28894 & ~n28913 ;
  assign n29664 = n28900 & ~n28907 ;
  assign n29665 = n29663 & n29664 ;
  assign n29673 = ~n29662 & ~n29665 ;
  assign n29674 = n29672 & n29673 ;
  assign n29669 = ~n28900 & ~n28923 ;
  assign n29670 = n28933 & ~n29664 ;
  assign n29671 = ~n29669 & n29670 ;
  assign n29666 = ~n28929 & ~n28933 ;
  assign n29667 = n28958 & n29666 ;
  assign n29668 = ~n28923 & ~n28953 ;
  assign n29675 = ~n29667 & ~n29668 ;
  assign n29676 = ~n29671 & n29675 ;
  assign n29677 = n29674 & n29676 ;
  assign n29684 = n28900 & n28952 ;
  assign n29685 = ~n28894 & n29684 ;
  assign n29678 = n28901 & n28914 ;
  assign n29686 = n28888 & ~n28946 ;
  assign n29687 = ~n29678 & n29686 ;
  assign n29688 = ~n29685 & n29687 ;
  assign n29679 = ~n28929 & ~n28934 ;
  assign n29680 = n28958 & ~n29679 ;
  assign n29681 = n28900 & n28913 ;
  assign n29682 = ~n28963 & ~n29681 ;
  assign n29683 = n28923 & ~n29682 ;
  assign n29689 = ~n29680 & ~n29683 ;
  assign n29690 = n29688 & n29689 ;
  assign n29691 = ~n29677 & ~n29690 ;
  assign n29692 = \u1_L13_reg[12]/NET0131  & n29691 ;
  assign n29693 = ~\u1_L13_reg[12]/NET0131  & ~n29691 ;
  assign n29694 = ~n29692 & ~n29693 ;
  assign n29695 = ~n29380 & ~n29418 ;
  assign n29696 = ~n29393 & n29695 ;
  assign n29697 = n29359 & ~n29696 ;
  assign n29698 = ~n29372 & n29610 ;
  assign n29699 = ~n29697 & ~n29698 ;
  assign n29700 = ~n29413 & ~n29699 ;
  assign n29701 = ~n29365 & n29418 ;
  assign n29703 = n29401 & n29415 ;
  assign n29704 = ~n29701 & ~n29703 ;
  assign n29705 = ~n29422 & n29704 ;
  assign n29702 = n29359 & n29429 ;
  assign n29706 = ~n29609 & ~n29702 ;
  assign n29707 = n29705 & n29706 ;
  assign n29708 = n29413 & ~n29707 ;
  assign n29711 = ~n29359 & ~n29390 ;
  assign n29709 = n29373 & n29392 ;
  assign n29710 = n29389 & ~n29413 ;
  assign n29712 = ~n29709 & ~n29710 ;
  assign n29713 = n29711 & n29712 ;
  assign n29714 = ~n29422 & ~n29430 ;
  assign n29715 = n29713 & n29714 ;
  assign n29716 = n29359 & ~n29434 ;
  assign n29717 = ~n29620 & n29716 ;
  assign n29718 = ~n29715 & ~n29717 ;
  assign n29719 = ~n29708 & ~n29718 ;
  assign n29720 = ~n29700 & n29719 ;
  assign n29721 = ~\u1_L13_reg[15]/P0001  & ~n29720 ;
  assign n29722 = \u1_L13_reg[15]/P0001  & n29720 ;
  assign n29723 = ~n29721 & ~n29722 ;
  assign n29724 = n28991 & ~n29027 ;
  assign n29725 = ~n29083 & n29724 ;
  assign n29726 = ~n28992 & ~n29725 ;
  assign n29728 = ~n28999 & ~n29009 ;
  assign n29729 = ~n29087 & n29728 ;
  assign n29727 = n29037 & n29087 ;
  assign n29730 = n29025 & ~n29727 ;
  assign n29731 = ~n29729 & n29730 ;
  assign n29732 = ~n29726 & n29731 ;
  assign n29734 = ~n28991 & n29071 ;
  assign n29733 = ~n29070 & n29724 ;
  assign n29735 = n29009 & n29095 ;
  assign n29736 = ~n29025 & ~n29735 ;
  assign n29737 = ~n29733 & n29736 ;
  assign n29738 = ~n29734 & n29737 ;
  assign n29739 = ~n29732 & ~n29738 ;
  assign n29740 = n29029 & ~n29087 ;
  assign n29741 = ~n29019 & ~n29740 ;
  assign n29742 = ~n29739 & n29741 ;
  assign n29743 = \u1_L13_reg[19]/P0001  & n29742 ;
  assign n29744 = ~\u1_L13_reg[19]/P0001  & ~n29742 ;
  assign n29745 = ~n29743 & ~n29744 ;
  assign n29766 = ~n29184 & n29197 ;
  assign n29767 = ~n29216 & ~n29766 ;
  assign n29768 = n29175 & ~n29767 ;
  assign n29769 = ~n29212 & n29633 ;
  assign n29770 = ~n29768 & n29769 ;
  assign n29771 = n29161 & ~n29770 ;
  assign n29746 = ~n29148 & ~n29184 ;
  assign n29747 = ~n29154 & n29746 ;
  assign n29748 = n29229 & ~n29747 ;
  assign n29749 = ~n29161 & ~n29207 ;
  assign n29750 = ~n29232 & n29749 ;
  assign n29751 = ~n29748 & ~n29750 ;
  assign n29752 = n29167 & n29232 ;
  assign n29753 = n29192 & ~n29752 ;
  assign n29754 = ~n29751 & n29753 ;
  assign n29755 = ~n29175 & ~n29754 ;
  assign n29756 = ~n29155 & n29187 ;
  assign n29757 = n29154 & n29196 ;
  assign n29758 = ~n29756 & ~n29757 ;
  assign n29759 = ~n29161 & ~n29758 ;
  assign n29760 = n29184 & ~n29189 ;
  assign n29761 = n29198 & n29760 ;
  assign n29762 = ~n29759 & ~n29761 ;
  assign n29763 = n29175 & ~n29762 ;
  assign n29764 = ~n29154 & ~n29161 ;
  assign n29765 = n29761 & n29764 ;
  assign n29772 = ~n29763 & ~n29765 ;
  assign n29773 = ~n29755 & n29772 ;
  assign n29774 = ~n29771 & n29773 ;
  assign n29775 = ~\u1_L13_reg[1]/NET0131  & ~n29774 ;
  assign n29776 = \u1_L13_reg[1]/NET0131  & n29774 ;
  assign n29777 = ~n29775 & ~n29776 ;
  assign n29798 = n28815 & n29121 ;
  assign n29799 = ~n29113 & ~n29798 ;
  assign n29800 = ~n28796 & ~n29799 ;
  assign n29779 = n28802 & n28827 ;
  assign n29801 = n28796 & n29779 ;
  assign n29802 = ~n28817 & ~n28853 ;
  assign n29803 = ~n28870 & n29802 ;
  assign n29804 = ~n29801 & n29803 ;
  assign n29805 = ~n29800 & n29804 ;
  assign n29806 = ~n28842 & ~n29805 ;
  assign n29782 = ~n28842 & ~n29114 ;
  assign n29783 = n28815 & ~n29115 ;
  assign n29784 = ~n29782 & n29783 ;
  assign n29780 = ~n28867 & ~n29779 ;
  assign n29781 = n28842 & ~n29780 ;
  assign n29778 = n28851 & n28866 ;
  assign n29785 = ~n29119 & ~n29778 ;
  assign n29786 = ~n29781 & n29785 ;
  assign n29787 = ~n29784 & n29786 ;
  assign n29788 = ~n28796 & ~n29787 ;
  assign n29789 = ~n28858 & ~n29779 ;
  assign n29790 = n28831 & ~n29789 ;
  assign n29792 = n28802 & n29130 ;
  assign n29793 = n28796 & ~n28816 ;
  assign n29794 = n29792 & n29793 ;
  assign n29791 = n28828 & n28874 ;
  assign n29795 = ~n29122 & ~n29791 ;
  assign n29796 = ~n29794 & n29795 ;
  assign n29797 = n28842 & ~n29796 ;
  assign n29807 = ~n29790 & ~n29797 ;
  assign n29808 = ~n29788 & n29807 ;
  assign n29809 = ~n29806 & n29808 ;
  assign n29810 = ~\u1_L13_reg[23]/P0001  & n29809 ;
  assign n29811 = \u1_L13_reg[23]/P0001  & ~n29809 ;
  assign n29812 = ~n29810 & ~n29811 ;
  assign n29813 = ~n29517 & ~n29524 ;
  assign n29814 = ~n29583 & ~n29813 ;
  assign n29815 = ~n29510 & ~n29814 ;
  assign n29816 = ~n29504 & ~n29517 ;
  assign n29817 = n29517 & n29537 ;
  assign n29818 = ~n29816 & ~n29817 ;
  assign n29819 = ~n29815 & n29818 ;
  assign n29820 = n29498 & ~n29819 ;
  assign n29821 = ~n29517 & n29537 ;
  assign n29822 = ~n29540 & ~n29821 ;
  assign n29823 = ~n29498 & ~n29822 ;
  assign n29824 = n29504 & n29529 ;
  assign n29825 = ~n29531 & ~n29824 ;
  assign n29826 = ~n29823 & n29825 ;
  assign n29827 = ~n29820 & n29826 ;
  assign n29828 = n29557 & ~n29827 ;
  assign n29838 = n29498 & ~n29528 ;
  assign n29837 = ~n29498 & ~n29816 ;
  assign n29839 = ~n29524 & ~n29837 ;
  assign n29840 = ~n29838 & n29839 ;
  assign n29833 = ~n29498 & n29518 ;
  assign n29834 = n29498 & ~n29510 ;
  assign n29835 = n29517 & n29583 ;
  assign n29836 = ~n29834 & n29835 ;
  assign n29841 = ~n29833 & ~n29836 ;
  assign n29842 = ~n29840 & n29841 ;
  assign n29843 = ~n29557 & ~n29842 ;
  assign n29829 = ~n29579 & ~n29824 ;
  assign n29830 = n29526 & n29813 ;
  assign n29831 = n29829 & ~n29830 ;
  assign n29832 = n29498 & ~n29831 ;
  assign n29844 = ~n29498 & n29504 ;
  assign n29845 = n29538 & n29844 ;
  assign n29846 = ~n29532 & ~n29845 ;
  assign n29847 = ~n29832 & n29846 ;
  assign n29848 = ~n29843 & n29847 ;
  assign n29849 = ~n29828 & n29848 ;
  assign n29850 = ~\u1_L13_reg[25]/NET0131  & ~n29849 ;
  assign n29851 = \u1_L13_reg[25]/NET0131  & n29849 ;
  assign n29852 = ~n29850 & ~n29851 ;
  assign n29867 = n29184 & n29189 ;
  assign n29868 = n29216 & n29746 ;
  assign n29869 = ~n29867 & ~n29868 ;
  assign n29870 = ~n29161 & ~n29869 ;
  assign n29875 = ~n29206 & ~n29870 ;
  assign n29871 = ~n29215 & ~n29747 ;
  assign n29872 = n29167 & ~n29871 ;
  assign n29873 = ~n29193 & ~n29757 ;
  assign n29874 = n29184 & ~n29873 ;
  assign n29876 = ~n29872 & ~n29874 ;
  assign n29877 = n29875 & n29876 ;
  assign n29878 = n29175 & ~n29877 ;
  assign n29855 = ~n29176 & ~n29631 ;
  assign n29856 = ~n29175 & ~n29855 ;
  assign n29857 = ~n29154 & ~n29198 ;
  assign n29858 = ~n29190 & ~n29857 ;
  assign n29859 = ~n29184 & ~n29858 ;
  assign n29860 = ~n29856 & ~n29859 ;
  assign n29861 = ~n29161 & ~n29860 ;
  assign n29853 = ~n29188 & ~n29208 ;
  assign n29854 = n29161 & ~n29853 ;
  assign n29862 = ~n29186 & n29209 ;
  assign n29863 = ~n29169 & ~n29188 ;
  assign n29864 = ~n29766 & n29863 ;
  assign n29865 = ~n29862 & n29864 ;
  assign n29866 = ~n29175 & ~n29865 ;
  assign n29879 = ~n29854 & ~n29866 ;
  assign n29880 = ~n29861 & n29879 ;
  assign n29881 = ~n29878 & n29880 ;
  assign n29882 = ~\u1_L13_reg[26]/NET0131  & ~n29881 ;
  assign n29883 = \u1_L13_reg[26]/NET0131  & n29881 ;
  assign n29884 = ~n29882 & ~n29883 ;
  assign n29888 = n29250 & n29456 ;
  assign n29890 = n29259 & n29281 ;
  assign n29889 = ~n29244 & n29294 ;
  assign n29885 = ~n29250 & n29265 ;
  assign n29891 = n29272 & ~n29885 ;
  assign n29892 = ~n29889 & n29891 ;
  assign n29893 = ~n29890 & n29892 ;
  assign n29894 = ~n29888 & n29893 ;
  assign n29896 = n29250 & ~n29259 ;
  assign n29897 = ~n29265 & ~n29284 ;
  assign n29898 = ~n29896 & n29897 ;
  assign n29895 = ~n29272 & ~n29315 ;
  assign n29899 = ~n29454 & n29895 ;
  assign n29900 = ~n29898 & n29899 ;
  assign n29901 = ~n29894 & ~n29900 ;
  assign n29886 = ~n29291 & ~n29885 ;
  assign n29887 = n29284 & ~n29886 ;
  assign n29902 = n29280 & ~n29887 ;
  assign n29903 = ~n29901 & n29902 ;
  assign n29906 = n29272 & ~n29898 ;
  assign n29907 = ~n29281 & ~n29295 ;
  assign n29908 = ~n29306 & n29907 ;
  assign n29909 = n29895 & n29908 ;
  assign n29910 = ~n29906 & ~n29909 ;
  assign n29904 = n29250 & ~n29889 ;
  assign n29905 = ~n29480 & n29904 ;
  assign n29911 = ~n29280 & ~n29905 ;
  assign n29912 = ~n29910 & n29911 ;
  assign n29913 = ~n29903 & ~n29912 ;
  assign n29914 = ~\u1_L13_reg[28]/NET0131  & n29913 ;
  assign n29915 = \u1_L13_reg[28]/NET0131  & ~n29913 ;
  assign n29916 = ~n29914 & ~n29915 ;
  assign n29918 = n29498 & ~n29525 ;
  assign n29919 = ~n29817 & n29918 ;
  assign n29920 = n29526 & ~n29538 ;
  assign n29921 = ~n29498 & ~n29821 ;
  assign n29922 = ~n29920 & n29921 ;
  assign n29923 = ~n29919 & ~n29922 ;
  assign n29924 = ~n29540 & n29829 ;
  assign n29925 = ~n29923 & n29924 ;
  assign n29926 = ~n29557 & ~n29925 ;
  assign n29930 = n29542 & n29813 ;
  assign n29931 = ~n29821 & ~n29930 ;
  assign n29932 = n29498 & ~n29931 ;
  assign n29933 = n29504 & n29567 ;
  assign n29934 = n29585 & ~n29933 ;
  assign n29935 = ~n29932 & n29934 ;
  assign n29936 = n29557 & ~n29935 ;
  assign n29917 = ~n29510 & n29845 ;
  assign n29927 = n29526 & ~n29559 ;
  assign n29928 = ~n29529 & ~n29927 ;
  assign n29929 = n29498 & ~n29928 ;
  assign n29937 = ~n29917 & ~n29929 ;
  assign n29938 = ~n29936 & n29937 ;
  assign n29939 = ~n29926 & n29938 ;
  assign n29940 = ~\u1_L13_reg[8]/NET0131  & ~n29939 ;
  assign n29941 = \u1_L13_reg[8]/NET0131  & n29939 ;
  assign n29942 = ~n29940 & ~n29941 ;
  assign n29944 = ~n28826 & ~n28845 ;
  assign n29945 = ~n29779 & n29944 ;
  assign n29946 = n28796 & ~n29945 ;
  assign n29947 = n28802 & ~n28851 ;
  assign n29948 = ~n28826 & ~n29947 ;
  assign n29949 = ~n28796 & n29948 ;
  assign n29943 = n28815 & n29131 ;
  assign n29950 = ~n28815 & n29114 ;
  assign n29951 = ~n29943 & ~n29950 ;
  assign n29952 = ~n29949 & n29951 ;
  assign n29953 = ~n29946 & n29952 ;
  assign n29954 = ~n28842 & ~n29953 ;
  assign n29955 = ~n28824 & n28870 ;
  assign n29956 = ~n29950 & ~n29955 ;
  assign n29957 = ~n28796 & ~n29956 ;
  assign n29959 = n28815 & ~n29131 ;
  assign n29960 = ~n29792 & n29959 ;
  assign n29958 = n28831 & n29948 ;
  assign n29961 = ~n29119 & ~n29958 ;
  assign n29962 = ~n29960 & n29961 ;
  assign n29963 = n28842 & ~n29962 ;
  assign n29964 = ~n29957 & ~n29963 ;
  assign n29965 = ~n29954 & n29964 ;
  assign n29966 = ~\u1_L13_reg[9]/NET0131  & ~n29965 ;
  assign n29967 = \u1_L13_reg[9]/NET0131  & n29965 ;
  assign n29968 = ~n29966 & ~n29967 ;
  assign n29971 = ~n28939 & ~n29663 ;
  assign n29972 = n28927 & ~n29971 ;
  assign n29973 = n28924 & n28958 ;
  assign n29974 = ~n29972 & ~n29973 ;
  assign n29975 = ~n28923 & ~n29974 ;
  assign n29969 = n28907 & n28929 ;
  assign n29970 = ~n29669 & n29969 ;
  assign n29976 = ~n28926 & ~n28960 ;
  assign n29977 = n28923 & ~n29976 ;
  assign n29978 = ~n29970 & ~n29977 ;
  assign n29979 = ~n29975 & n29978 ;
  assign n29980 = n28888 & ~n29979 ;
  assign n29981 = n28923 & ~n28959 ;
  assign n29982 = ~n28923 & ~n29684 ;
  assign n29983 = n28913 & n28960 ;
  assign n29984 = n29982 & ~n29983 ;
  assign n29985 = ~n29981 & ~n29984 ;
  assign n29986 = ~n28907 & n28929 ;
  assign n29990 = n29668 & ~n29986 ;
  assign n29987 = n28924 & ~n29664 ;
  assign n29988 = ~n29986 & ~n29987 ;
  assign n29989 = ~n29669 & ~n29988 ;
  assign n29991 = ~n28954 & ~n29989 ;
  assign n29992 = ~n29990 & n29991 ;
  assign n29993 = ~n28888 & ~n29992 ;
  assign n29994 = ~n29985 & ~n29993 ;
  assign n29995 = ~n29980 & n29994 ;
  assign n29996 = \u1_L13_reg[32]/NET0131  & n29995 ;
  assign n29997 = ~\u1_L13_reg[32]/NET0131  & ~n29995 ;
  assign n29998 = ~n29996 & ~n29997 ;
  assign n30015 = ~n29365 & n29438 ;
  assign n30016 = ~n29607 & ~n30015 ;
  assign n30017 = n29359 & ~n30016 ;
  assign n30012 = ~n29419 & ~n29442 ;
  assign n30013 = ~n29615 & n30012 ;
  assign n30014 = ~n29359 & ~n30013 ;
  assign n30018 = ~n29391 & ~n29424 ;
  assign n30019 = ~n29434 & n30018 ;
  assign n30020 = ~n30014 & n30019 ;
  assign n30021 = ~n30017 & n30020 ;
  assign n30022 = n29413 & ~n30021 ;
  assign n30000 = n29359 & ~n29380 ;
  assign n29999 = ~n29373 & n29379 ;
  assign n30001 = ~n29421 & ~n29999 ;
  assign n30002 = n30000 & n30001 ;
  assign n30003 = n29396 & n29415 ;
  assign n30004 = ~n29427 & ~n30003 ;
  assign n30005 = ~n29598 & n30004 ;
  assign n30006 = ~n30002 & n30005 ;
  assign n30007 = ~n29413 & ~n30006 ;
  assign n30011 = ~n29359 & ~n29426 ;
  assign n30008 = n29359 & n29365 ;
  assign n30009 = ~n29372 & ~n29379 ;
  assign n30010 = n30008 & n30009 ;
  assign n30023 = ~n29420 & ~n30010 ;
  assign n30024 = ~n30011 & n30023 ;
  assign n30025 = ~n30007 & n30024 ;
  assign n30026 = ~n30022 & n30025 ;
  assign n30027 = \u1_L13_reg[27]/NET0131  & n30026 ;
  assign n30028 = ~\u1_L13_reg[27]/NET0131  & ~n30026 ;
  assign n30029 = ~n30027 & ~n30028 ;
  assign n30031 = ~n29542 & ~n29544 ;
  assign n30032 = n29921 & n30031 ;
  assign n30033 = ~n29524 & n29526 ;
  assign n30034 = n29498 & ~n29563 ;
  assign n30035 = ~n30033 & n30034 ;
  assign n30036 = ~n30032 & ~n30035 ;
  assign n30030 = ~n29511 & n29538 ;
  assign n30037 = ~n29557 & ~n30030 ;
  assign n30038 = ~n30036 & n30037 ;
  assign n30040 = ~n29504 & n29528 ;
  assign n30041 = ~n29561 & ~n30040 ;
  assign n30042 = n29498 & ~n30041 ;
  assign n30044 = ~n29532 & n29557 ;
  assign n30039 = n29518 & n29524 ;
  assign n30043 = ~n29498 & n29568 ;
  assign n30045 = ~n30039 & ~n30043 ;
  assign n30046 = n30044 & n30045 ;
  assign n30047 = ~n30042 & n30046 ;
  assign n30048 = ~n30038 & ~n30047 ;
  assign n30049 = ~n29582 & n29918 ;
  assign n30050 = ~n29498 & ~n29539 ;
  assign n30051 = ~n29930 & n30050 ;
  assign n30052 = ~n29578 & n30051 ;
  assign n30053 = ~n30049 & ~n30052 ;
  assign n30054 = ~n30048 & ~n30053 ;
  assign n30055 = ~\u1_L13_reg[3]/NET0131  & ~n30054 ;
  assign n30056 = \u1_L13_reg[3]/NET0131  & n30054 ;
  assign n30057 = ~n30055 & ~n30056 ;
  assign n30092 = decrypt_pad & ~\u1_uk_K_r13_reg[20]/NET0131  ;
  assign n30093 = ~decrypt_pad & ~\u1_uk_K_r13_reg[41]/NET0131  ;
  assign n30094 = ~n30092 & ~n30093 ;
  assign n30095 = \u1_R13_reg[11]/P0001  & ~n30094 ;
  assign n30096 = ~\u1_R13_reg[11]/P0001  & n30094 ;
  assign n30097 = ~n30095 & ~n30096 ;
  assign n30084 = decrypt_pad & ~\u1_uk_K_r13_reg[3]/NET0131  ;
  assign n30085 = ~decrypt_pad & ~\u1_uk_K_r13_reg[24]/NET0131  ;
  assign n30086 = ~n30084 & ~n30085 ;
  assign n30087 = \u1_R13_reg[12]/NET0131  & ~n30086 ;
  assign n30088 = ~\u1_R13_reg[12]/NET0131  & n30086 ;
  assign n30089 = ~n30087 & ~n30088 ;
  assign n30058 = decrypt_pad & ~\u1_uk_K_r13_reg[48]/NET0131  ;
  assign n30059 = ~decrypt_pad & ~\u1_uk_K_r13_reg[12]/NET0131  ;
  assign n30060 = ~n30058 & ~n30059 ;
  assign n30061 = \u1_R13_reg[13]/NET0131  & ~n30060 ;
  assign n30062 = ~\u1_R13_reg[13]/NET0131  & n30060 ;
  assign n30063 = ~n30061 & ~n30062 ;
  assign n30071 = decrypt_pad & ~\u1_uk_K_r13_reg[11]/NET0131  ;
  assign n30072 = ~decrypt_pad & ~\u1_uk_K_r13_reg[32]/NET0131  ;
  assign n30073 = ~n30071 & ~n30072 ;
  assign n30074 = \u1_R13_reg[9]/NET0131  & ~n30073 ;
  assign n30075 = ~\u1_R13_reg[9]/NET0131  & n30073 ;
  assign n30076 = ~n30074 & ~n30075 ;
  assign n30098 = n30063 & ~n30076 ;
  assign n30077 = decrypt_pad & ~\u1_uk_K_r13_reg[19]/NET0131  ;
  assign n30078 = ~decrypt_pad & ~\u1_uk_K_r13_reg[40]/NET0131  ;
  assign n30079 = ~n30077 & ~n30078 ;
  assign n30080 = \u1_R13_reg[10]/NET0131  & ~n30079 ;
  assign n30081 = ~\u1_R13_reg[10]/NET0131  & n30079 ;
  assign n30082 = ~n30080 & ~n30081 ;
  assign n30064 = decrypt_pad & ~\u1_uk_K_r13_reg[39]/NET0131  ;
  assign n30065 = ~decrypt_pad & ~\u1_uk_K_r13_reg[3]/NET0131  ;
  assign n30066 = ~n30064 & ~n30065 ;
  assign n30067 = \u1_R13_reg[8]/NET0131  & ~n30066 ;
  assign n30068 = ~\u1_R13_reg[8]/NET0131  & n30066 ;
  assign n30069 = ~n30067 & ~n30068 ;
  assign n30100 = n30063 & ~n30069 ;
  assign n30101 = n30082 & n30100 ;
  assign n30102 = ~n30063 & n30069 ;
  assign n30103 = n30076 & n30102 ;
  assign n30104 = ~n30101 & ~n30103 ;
  assign n30105 = ~n30098 & n30104 ;
  assign n30106 = n30089 & ~n30105 ;
  assign n30099 = n30082 & n30098 ;
  assign n30070 = ~n30063 & ~n30069 ;
  assign n30107 = n30070 & ~n30076 ;
  assign n30108 = ~n30082 & n30107 ;
  assign n30109 = ~n30099 & ~n30108 ;
  assign n30110 = ~n30106 & n30109 ;
  assign n30111 = n30097 & ~n30110 ;
  assign n30083 = n30076 & n30082 ;
  assign n30119 = ~n30076 & ~n30082 ;
  assign n30120 = ~n30083 & ~n30119 ;
  assign n30121 = ~n30069 & n30097 ;
  assign n30123 = ~n30100 & ~n30102 ;
  assign n30126 = ~n30121 & ~n30123 ;
  assign n30127 = ~n30120 & ~n30126 ;
  assign n30122 = n30076 & n30121 ;
  assign n30124 = n30120 & ~n30122 ;
  assign n30125 = ~n30123 & n30124 ;
  assign n30128 = ~n30089 & ~n30125 ;
  assign n30129 = ~n30127 & n30128 ;
  assign n30090 = n30083 & n30089 ;
  assign n30091 = n30070 & n30090 ;
  assign n30113 = n30076 & ~n30082 ;
  assign n30114 = ~n30069 & ~n30113 ;
  assign n30115 = n30089 & ~n30097 ;
  assign n30112 = ~n30063 & n30076 ;
  assign n30116 = ~n30098 & ~n30112 ;
  assign n30117 = n30115 & n30116 ;
  assign n30118 = ~n30114 & n30117 ;
  assign n30130 = ~n30091 & ~n30118 ;
  assign n30131 = ~n30129 & n30130 ;
  assign n30132 = ~n30111 & n30131 ;
  assign n30133 = ~\u1_L13_reg[6]/NET0131  & ~n30132 ;
  assign n30134 = \u1_L13_reg[6]/NET0131  & n30132 ;
  assign n30135 = ~n30133 & ~n30134 ;
  assign n30136 = n28900 & ~n29666 ;
  assign n30137 = n28907 & n30136 ;
  assign n30138 = ~n29973 & ~n30137 ;
  assign n30139 = ~n28907 & n29666 ;
  assign n30140 = ~n28925 & n30139 ;
  assign n30141 = n28923 & ~n30140 ;
  assign n30142 = ~n28900 & n28914 ;
  assign n30143 = ~n29969 & ~n30142 ;
  assign n30144 = n29982 & n30143 ;
  assign n30145 = ~n30136 & n30144 ;
  assign n30146 = ~n30141 & ~n30145 ;
  assign n30147 = n30138 & ~n30146 ;
  assign n30148 = n28888 & ~n30147 ;
  assign n30150 = ~n28923 & n30140 ;
  assign n30151 = n28925 & n28952 ;
  assign n30152 = ~n30150 & ~n30151 ;
  assign n30153 = ~n28888 & ~n30152 ;
  assign n30149 = ~n28923 & ~n30138 ;
  assign n30154 = n28888 & ~n30151 ;
  assign n30155 = ~n28900 & n28924 ;
  assign n30156 = n28923 & ~n30155 ;
  assign n30157 = ~n30139 & n30156 ;
  assign n30158 = ~n30154 & n30157 ;
  assign n30159 = ~n30137 & n30158 ;
  assign n30160 = ~n30149 & ~n30159 ;
  assign n30161 = ~n30153 & n30160 ;
  assign n30162 = ~n30148 & n30161 ;
  assign n30163 = \u1_L13_reg[7]/NET0131  & n30162 ;
  assign n30164 = ~\u1_L13_reg[7]/NET0131  & ~n30162 ;
  assign n30165 = ~n30163 & ~n30164 ;
  assign n30177 = n30070 & n30082 ;
  assign n30178 = ~n30082 & n30100 ;
  assign n30179 = ~n30177 & ~n30178 ;
  assign n30180 = n30102 & n30119 ;
  assign n30181 = n30179 & ~n30180 ;
  assign n30182 = n30097 & ~n30181 ;
  assign n30183 = n30089 & ~n30182 ;
  assign n30166 = n30069 & n30082 ;
  assign n30186 = ~n30112 & n30166 ;
  assign n30185 = ~n30063 & n30113 ;
  assign n30187 = ~n30089 & n30097 ;
  assign n30188 = ~n30185 & n30187 ;
  assign n30189 = ~n30186 & n30188 ;
  assign n30191 = n30069 & ~n30082 ;
  assign n30192 = ~n30112 & n30191 ;
  assign n30190 = n30076 & n30100 ;
  assign n30193 = ~n30097 & ~n30190 ;
  assign n30194 = ~n30192 & n30193 ;
  assign n30195 = ~n30189 & ~n30194 ;
  assign n30184 = n30119 & n30123 ;
  assign n30196 = ~n30076 & n30100 ;
  assign n30197 = n30082 & n30196 ;
  assign n30198 = ~n30184 & ~n30197 ;
  assign n30199 = ~n30195 & n30198 ;
  assign n30200 = ~n30183 & ~n30199 ;
  assign n30167 = n30070 & n30076 ;
  assign n30168 = ~n30166 & ~n30167 ;
  assign n30169 = n30115 & ~n30168 ;
  assign n30174 = n30082 & n30097 ;
  assign n30170 = n30063 & n30069 ;
  assign n30175 = ~n30076 & n30170 ;
  assign n30176 = n30174 & n30175 ;
  assign n30171 = n30090 & ~n30170 ;
  assign n30172 = n30082 & ~n30097 ;
  assign n30173 = n30112 & n30172 ;
  assign n30201 = ~n30171 & ~n30173 ;
  assign n30202 = ~n30176 & n30201 ;
  assign n30203 = ~n30169 & n30202 ;
  assign n30204 = ~n30200 & n30203 ;
  assign n30205 = \u1_L13_reg[30]/NET0131  & ~n30204 ;
  assign n30206 = ~\u1_L13_reg[30]/NET0131  & n30204 ;
  assign n30207 = ~n30205 & ~n30206 ;
  assign n30208 = ~n30103 & ~n30107 ;
  assign n30209 = n30174 & ~n30208 ;
  assign n30215 = n30082 & ~n30190 ;
  assign n30216 = n30076 & n30170 ;
  assign n30217 = ~n30196 & ~n30216 ;
  assign n30219 = n30112 & n30121 ;
  assign n30218 = ~n30076 & n30102 ;
  assign n30220 = ~n30082 & ~n30218 ;
  assign n30221 = ~n30219 & n30220 ;
  assign n30222 = n30217 & n30221 ;
  assign n30223 = ~n30215 & ~n30222 ;
  assign n30211 = ~n30076 & n30166 ;
  assign n30210 = ~n30082 & n30102 ;
  assign n30212 = ~n30177 & ~n30210 ;
  assign n30213 = ~n30211 & n30212 ;
  assign n30214 = ~n30097 & ~n30213 ;
  assign n30224 = n30089 & ~n30214 ;
  assign n30225 = ~n30223 & n30224 ;
  assign n30230 = n30070 & ~n30082 ;
  assign n30231 = ~n30211 & ~n30230 ;
  assign n30232 = n30217 & n30231 ;
  assign n30233 = ~n30097 & ~n30232 ;
  assign n30226 = ~n30076 & ~n30170 ;
  assign n30227 = ~n30070 & n30097 ;
  assign n30228 = ~n30216 & n30227 ;
  assign n30229 = ~n30226 & n30228 ;
  assign n30234 = ~n30089 & ~n30108 ;
  assign n30235 = ~n30229 & n30234 ;
  assign n30236 = ~n30233 & n30235 ;
  assign n30237 = ~n30225 & ~n30236 ;
  assign n30238 = ~n30209 & ~n30237 ;
  assign n30239 = ~\u1_L13_reg[16]/NET0131  & ~n30238 ;
  assign n30240 = \u1_L13_reg[16]/NET0131  & n30238 ;
  assign n30241 = ~n30239 & ~n30240 ;
  assign n30246 = n29272 & ~n29310 ;
  assign n30243 = n29259 & n29885 ;
  assign n30244 = ~n29889 & ~n30243 ;
  assign n30245 = ~n29272 & ~n30244 ;
  assign n30247 = ~n29316 & ~n30245 ;
  assign n30248 = ~n30246 & n30247 ;
  assign n30249 = n29280 & ~n30248 ;
  assign n30253 = ~n29265 & ~n29292 ;
  assign n30254 = n29253 & n30253 ;
  assign n30250 = n29259 & ~n29272 ;
  assign n30251 = n29281 & ~n29464 ;
  assign n30252 = ~n30250 & n30251 ;
  assign n30255 = ~n29286 & ~n29468 ;
  assign n30256 = ~n30252 & n30255 ;
  assign n30257 = ~n30254 & n30256 ;
  assign n30258 = ~n29280 & ~n30257 ;
  assign n30242 = n29244 & n29273 ;
  assign n30259 = ~n29285 & ~n29456 ;
  assign n30260 = n29272 & ~n29896 ;
  assign n30261 = ~n30259 & n30260 ;
  assign n30262 = ~n30242 & ~n30261 ;
  assign n30263 = ~n30258 & n30262 ;
  assign n30264 = ~n30249 & n30263 ;
  assign n30265 = ~\u1_L13_reg[18]/P0001  & ~n30264 ;
  assign n30266 = \u1_L13_reg[18]/P0001  & n30264 ;
  assign n30267 = ~n30265 & ~n30266 ;
  assign n30282 = ~n30167 & ~n30211 ;
  assign n30283 = n30179 & n30282 ;
  assign n30284 = n30097 & ~n30283 ;
  assign n30285 = n30082 & n30218 ;
  assign n30286 = ~n30284 & ~n30285 ;
  assign n30287 = ~n30089 & ~n30286 ;
  assign n30272 = n30119 & n30126 ;
  assign n30269 = n30076 & n30166 ;
  assign n30270 = ~n30101 & ~n30269 ;
  assign n30271 = n30097 & ~n30270 ;
  assign n30273 = ~n30097 & ~n30119 ;
  assign n30274 = n30123 & n30273 ;
  assign n30275 = ~n30082 & n30097 ;
  assign n30276 = ~n30076 & ~n30100 ;
  assign n30277 = n30275 & n30276 ;
  assign n30278 = ~n30274 & ~n30277 ;
  assign n30279 = ~n30271 & n30278 ;
  assign n30280 = ~n30272 & n30279 ;
  assign n30281 = n30089 & ~n30280 ;
  assign n30290 = n30104 & ~n30184 ;
  assign n30291 = ~n30089 & ~n30097 ;
  assign n30292 = ~n30290 & n30291 ;
  assign n30268 = n30172 & n30216 ;
  assign n30288 = ~n30190 & ~n30218 ;
  assign n30289 = n30275 & ~n30288 ;
  assign n30293 = ~n30268 & ~n30289 ;
  assign n30294 = ~n30292 & n30293 ;
  assign n30295 = ~n30281 & n30294 ;
  assign n30296 = ~n30287 & n30295 ;
  assign n30297 = ~\u1_L13_reg[24]/NET0131  & ~n30296 ;
  assign n30298 = \u1_L13_reg[24]/NET0131  & n30296 ;
  assign n30299 = ~n30297 & ~n30298 ;
  assign n30349 = decrypt_pad & ~\u1_uk_K_r12_reg[14]/NET0131  ;
  assign n30350 = ~decrypt_pad & ~\u1_uk_K_r12_reg[8]/NET0131  ;
  assign n30351 = ~n30349 & ~n30350 ;
  assign n30352 = \u1_R12_reg[28]/NET0131  & ~n30351 ;
  assign n30353 = ~\u1_R12_reg[28]/NET0131  & n30351 ;
  assign n30354 = ~n30352 & ~n30353 ;
  assign n30300 = decrypt_pad & ~\u1_uk_K_r12_reg[31]/NET0131  ;
  assign n30301 = ~decrypt_pad & ~\u1_uk_K_r12_reg[21]/NET0131  ;
  assign n30302 = ~n30300 & ~n30301 ;
  assign n30303 = \u1_R12_reg[27]/NET0131  & ~n30302 ;
  assign n30304 = ~\u1_R12_reg[27]/NET0131  & n30302 ;
  assign n30305 = ~n30303 & ~n30304 ;
  assign n30312 = decrypt_pad & ~\u1_uk_K_r12_reg[29]/NET0131  ;
  assign n30313 = ~decrypt_pad & ~\u1_uk_K_r12_reg[23]/NET0131  ;
  assign n30314 = ~n30312 & ~n30313 ;
  assign n30315 = \u1_R12_reg[24]/NET0131  & ~n30314 ;
  assign n30316 = ~\u1_R12_reg[24]/NET0131  & n30314 ;
  assign n30317 = ~n30315 & ~n30316 ;
  assign n30326 = decrypt_pad & ~\u1_uk_K_r12_reg[49]/NET0131  ;
  assign n30327 = ~decrypt_pad & ~\u1_uk_K_r12_reg[43]/NET0131  ;
  assign n30328 = ~n30326 & ~n30327 ;
  assign n30329 = \u1_R12_reg[26]/NET0131  & ~n30328 ;
  assign n30330 = ~\u1_R12_reg[26]/NET0131  & n30328 ;
  assign n30331 = ~n30329 & ~n30330 ;
  assign n30306 = decrypt_pad & ~\u1_uk_K_r12_reg[37]/NET0131  ;
  assign n30307 = ~decrypt_pad & ~\u1_uk_K_r12_reg[0]/NET0131  ;
  assign n30308 = ~n30306 & ~n30307 ;
  assign n30309 = \u1_R12_reg[29]/NET0131  & ~n30308 ;
  assign n30310 = ~\u1_R12_reg[29]/NET0131  & n30308 ;
  assign n30311 = ~n30309 & ~n30310 ;
  assign n30319 = decrypt_pad & ~\u1_uk_K_r12_reg[9]/NET0131  ;
  assign n30320 = ~decrypt_pad & ~\u1_uk_K_r12_reg[31]/NET0131  ;
  assign n30321 = ~n30319 & ~n30320 ;
  assign n30322 = \u1_R12_reg[25]/NET0131  & ~n30321 ;
  assign n30323 = ~\u1_R12_reg[25]/NET0131  & n30321 ;
  assign n30324 = ~n30322 & ~n30323 ;
  assign n30355 = n30311 & n30324 ;
  assign n30382 = ~n30331 & n30355 ;
  assign n30383 = n30317 & n30382 ;
  assign n30333 = n30317 & ~n30324 ;
  assign n30384 = n30331 & n30333 ;
  assign n30385 = ~n30383 & ~n30384 ;
  assign n30386 = n30305 & ~n30385 ;
  assign n30377 = n30311 & n30333 ;
  assign n30378 = ~n30331 & n30377 ;
  assign n30318 = n30311 & ~n30317 ;
  assign n30379 = n30318 & n30324 ;
  assign n30380 = ~n30378 & ~n30379 ;
  assign n30381 = ~n30305 & ~n30380 ;
  assign n30325 = n30318 & ~n30324 ;
  assign n30332 = n30325 & n30331 ;
  assign n30341 = ~n30311 & ~n30324 ;
  assign n30345 = ~n30317 & ~n30331 ;
  assign n30376 = n30341 & n30345 ;
  assign n30387 = ~n30332 & ~n30376 ;
  assign n30388 = ~n30381 & n30387 ;
  assign n30389 = ~n30386 & n30388 ;
  assign n30390 = n30354 & ~n30389 ;
  assign n30335 = ~n30311 & ~n30317 ;
  assign n30361 = ~n30324 & n30335 ;
  assign n30362 = n30331 & n30361 ;
  assign n30344 = n30317 & n30331 ;
  assign n30363 = n30311 & n30344 ;
  assign n30364 = n30317 & n30324 ;
  assign n30365 = ~n30311 & n30364 ;
  assign n30366 = ~n30363 & ~n30365 ;
  assign n30367 = ~n30362 & n30366 ;
  assign n30368 = ~n30305 & ~n30367 ;
  assign n30358 = ~n30305 & ~n30318 ;
  assign n30357 = n30305 & ~n30333 ;
  assign n30359 = ~n30331 & ~n30357 ;
  assign n30360 = ~n30358 & n30359 ;
  assign n30346 = ~n30344 & ~n30345 ;
  assign n30356 = ~n30346 & n30355 ;
  assign n30369 = ~n30311 & n30317 ;
  assign n30370 = ~n30331 & n30369 ;
  assign n30371 = ~n30324 & n30370 ;
  assign n30372 = ~n30356 & ~n30371 ;
  assign n30373 = ~n30360 & n30372 ;
  assign n30374 = ~n30368 & n30373 ;
  assign n30375 = ~n30354 & ~n30374 ;
  assign n30334 = ~n30311 & n30333 ;
  assign n30336 = n30324 & n30331 ;
  assign n30337 = n30335 & n30336 ;
  assign n30338 = ~n30334 & ~n30337 ;
  assign n30339 = ~n30332 & n30338 ;
  assign n30340 = n30305 & ~n30339 ;
  assign n30342 = n30305 & ~n30331 ;
  assign n30343 = n30341 & n30342 ;
  assign n30347 = ~n30305 & n30324 ;
  assign n30348 = ~n30346 & n30347 ;
  assign n30391 = ~n30343 & ~n30348 ;
  assign n30392 = ~n30340 & n30391 ;
  assign n30393 = ~n30375 & n30392 ;
  assign n30394 = ~n30390 & n30393 ;
  assign n30395 = ~\u1_L12_reg[22]/NET0131  & ~n30394 ;
  assign n30396 = \u1_L12_reg[22]/NET0131  & n30394 ;
  assign n30397 = ~n30395 & ~n30396 ;
  assign n30398 = decrypt_pad & ~\u1_uk_K_r12_reg[10]/P0001  ;
  assign n30399 = ~decrypt_pad & ~\u1_uk_K_r12_reg[34]/NET0131  ;
  assign n30400 = ~n30398 & ~n30399 ;
  assign n30401 = \u1_R12_reg[4]/NET0131  & ~n30400 ;
  assign n30402 = ~\u1_R12_reg[4]/NET0131  & n30400 ;
  assign n30403 = ~n30401 & ~n30402 ;
  assign n30404 = decrypt_pad & ~\u1_uk_K_r12_reg[40]/NET0131  ;
  assign n30405 = ~decrypt_pad & ~\u1_uk_K_r12_reg[32]/NET0131  ;
  assign n30406 = ~n30404 & ~n30405 ;
  assign n30407 = \u1_R12_reg[1]/NET0131  & ~n30406 ;
  assign n30408 = ~\u1_R12_reg[1]/NET0131  & n30406 ;
  assign n30409 = ~n30407 & ~n30408 ;
  assign n30410 = decrypt_pad & ~\u1_uk_K_r12_reg[13]/NET0131  ;
  assign n30411 = ~decrypt_pad & ~\u1_uk_K_r12_reg[5]/NET0131  ;
  assign n30412 = ~n30410 & ~n30411 ;
  assign n30413 = \u1_R12_reg[5]/NET0131  & ~n30412 ;
  assign n30414 = ~\u1_R12_reg[5]/NET0131  & n30412 ;
  assign n30415 = ~n30413 & ~n30414 ;
  assign n30416 = ~n30409 & ~n30415 ;
  assign n30417 = decrypt_pad & ~\u1_uk_K_r12_reg[19]/NET0131  ;
  assign n30418 = ~decrypt_pad & ~\u1_uk_K_r12_reg[11]/NET0131  ;
  assign n30419 = ~n30417 & ~n30418 ;
  assign n30420 = \u1_R12_reg[32]/NET0131  & ~n30419 ;
  assign n30421 = ~\u1_R12_reg[32]/NET0131  & n30419 ;
  assign n30422 = ~n30420 & ~n30421 ;
  assign n30423 = n30416 & n30422 ;
  assign n30424 = decrypt_pad & ~\u1_uk_K_r12_reg[55]/NET0131  ;
  assign n30425 = ~decrypt_pad & ~\u1_uk_K_r12_reg[47]/NET0131  ;
  assign n30426 = ~n30424 & ~n30425 ;
  assign n30427 = \u1_R12_reg[2]/NET0131  & ~n30426 ;
  assign n30428 = ~\u1_R12_reg[2]/NET0131  & n30426 ;
  assign n30429 = ~n30427 & ~n30428 ;
  assign n30430 = n30423 & n30429 ;
  assign n30431 = ~n30409 & n30415 ;
  assign n30432 = ~n30422 & ~n30429 ;
  assign n30433 = ~n30431 & n30432 ;
  assign n30434 = ~n30430 & ~n30433 ;
  assign n30435 = decrypt_pad & ~\u1_uk_K_r12_reg[32]/NET0131  ;
  assign n30436 = ~decrypt_pad & ~\u1_uk_K_r12_reg[24]/NET0131  ;
  assign n30437 = ~n30435 & ~n30436 ;
  assign n30438 = \u1_R12_reg[3]/NET0131  & ~n30437 ;
  assign n30439 = ~\u1_R12_reg[3]/NET0131  & n30437 ;
  assign n30440 = ~n30438 & ~n30439 ;
  assign n30441 = ~n30434 & ~n30440 ;
  assign n30442 = n30415 & n30422 ;
  assign n30449 = n30409 & ~n30440 ;
  assign n30450 = n30442 & ~n30449 ;
  assign n30443 = ~n30415 & ~n30422 ;
  assign n30448 = n30409 & n30443 ;
  assign n30451 = ~n30429 & ~n30448 ;
  assign n30452 = ~n30450 & n30451 ;
  assign n30444 = ~n30442 & ~n30443 ;
  assign n30445 = n30409 & n30444 ;
  assign n30446 = n30429 & ~n30445 ;
  assign n30447 = n30429 & ~n30440 ;
  assign n30453 = ~n30446 & ~n30447 ;
  assign n30454 = ~n30452 & n30453 ;
  assign n30455 = ~n30441 & ~n30454 ;
  assign n30456 = ~n30403 & ~n30455 ;
  assign n30466 = n30429 & n30443 ;
  assign n30469 = ~n30431 & ~n30466 ;
  assign n30470 = n30440 & ~n30469 ;
  assign n30457 = ~n30415 & ~n30429 ;
  assign n30475 = n30422 & ~n30457 ;
  assign n30476 = ~n30409 & ~n30432 ;
  assign n30477 = ~n30475 & n30476 ;
  assign n30460 = n30415 & ~n30422 ;
  assign n30471 = ~n30429 & n30440 ;
  assign n30472 = n30409 & ~n30471 ;
  assign n30473 = n30460 & ~n30472 ;
  assign n30474 = n30422 & n30449 ;
  assign n30478 = ~n30473 & ~n30474 ;
  assign n30479 = ~n30477 & n30478 ;
  assign n30480 = ~n30470 & n30479 ;
  assign n30481 = n30403 & ~n30480 ;
  assign n30458 = n30409 & n30457 ;
  assign n30459 = n30409 & n30442 ;
  assign n30461 = ~n30409 & n30460 ;
  assign n30462 = ~n30459 & ~n30461 ;
  assign n30463 = n30429 & ~n30462 ;
  assign n30464 = ~n30458 & ~n30463 ;
  assign n30465 = ~n30440 & ~n30464 ;
  assign n30467 = ~n30409 & n30440 ;
  assign n30468 = n30466 & n30467 ;
  assign n30482 = n30422 & ~n30429 ;
  assign n30483 = n30467 & n30482 ;
  assign n30484 = ~n30468 & ~n30483 ;
  assign n30485 = ~n30465 & n30484 ;
  assign n30486 = ~n30481 & n30485 ;
  assign n30487 = ~n30456 & n30486 ;
  assign n30488 = ~\u1_L12_reg[31]/NET0131  & ~n30487 ;
  assign n30489 = \u1_L12_reg[31]/NET0131  & n30487 ;
  assign n30490 = ~n30488 & ~n30489 ;
  assign n30547 = decrypt_pad & ~\u1_uk_K_r12_reg[7]/P0001  ;
  assign n30548 = ~decrypt_pad & ~\u1_uk_K_r12_reg[1]/NET0131  ;
  assign n30549 = ~n30547 & ~n30548 ;
  assign n30550 = \u1_R12_reg[24]/NET0131  & ~n30549 ;
  assign n30551 = ~\u1_R12_reg[24]/NET0131  & n30549 ;
  assign n30552 = ~n30550 & ~n30551 ;
  assign n30514 = decrypt_pad & ~\u1_uk_K_r12_reg[36]/NET0131  ;
  assign n30515 = ~decrypt_pad & ~\u1_uk_K_r12_reg[30]/NET0131  ;
  assign n30516 = ~n30514 & ~n30515 ;
  assign n30517 = \u1_R12_reg[23]/NET0131  & ~n30516 ;
  assign n30518 = ~\u1_R12_reg[23]/NET0131  & n30516 ;
  assign n30519 = ~n30517 & ~n30518 ;
  assign n30497 = decrypt_pad & ~\u1_uk_K_r12_reg[1]/NET0131  ;
  assign n30498 = ~decrypt_pad & ~\u1_uk_K_r12_reg[50]/NET0131  ;
  assign n30499 = ~n30497 & ~n30498 ;
  assign n30500 = \u1_R12_reg[21]/NET0131  & ~n30499 ;
  assign n30501 = ~\u1_R12_reg[21]/NET0131  & n30499 ;
  assign n30502 = ~n30500 & ~n30501 ;
  assign n30504 = decrypt_pad & ~\u1_uk_K_r12_reg[45]/NET0131  ;
  assign n30505 = ~decrypt_pad & ~\u1_uk_K_r12_reg[35]/NET0131  ;
  assign n30506 = ~n30504 & ~n30505 ;
  assign n30507 = \u1_R12_reg[20]/NET0131  & ~n30506 ;
  assign n30508 = ~\u1_R12_reg[20]/NET0131  & n30506 ;
  assign n30509 = ~n30507 & ~n30508 ;
  assign n30525 = decrypt_pad & ~\u1_uk_K_r12_reg[2]/NET0131  ;
  assign n30526 = ~decrypt_pad & ~\u1_uk_K_r12_reg[51]/NET0131  ;
  assign n30527 = ~n30525 & ~n30526 ;
  assign n30528 = \u1_R12_reg[25]/NET0131  & ~n30527 ;
  assign n30529 = ~\u1_R12_reg[25]/NET0131  & n30527 ;
  assign n30530 = ~n30528 & ~n30529 ;
  assign n30537 = n30509 & n30530 ;
  assign n30556 = n30502 & n30537 ;
  assign n30491 = decrypt_pad & ~\u1_uk_K_r12_reg[23]/NET0131  ;
  assign n30492 = ~decrypt_pad & ~\u1_uk_K_r12_reg[45]/NET0131  ;
  assign n30493 = ~n30491 & ~n30492 ;
  assign n30494 = \u1_R12_reg[22]/NET0131  & ~n30493 ;
  assign n30495 = ~\u1_R12_reg[22]/NET0131  & n30493 ;
  assign n30496 = ~n30494 & ~n30495 ;
  assign n30503 = n30496 & n30502 ;
  assign n30510 = n30503 & ~n30509 ;
  assign n30535 = n30509 & ~n30530 ;
  assign n30554 = ~n30496 & ~n30502 ;
  assign n30555 = n30535 & n30554 ;
  assign n30557 = ~n30510 & ~n30555 ;
  assign n30558 = ~n30556 & n30557 ;
  assign n30559 = n30519 & ~n30558 ;
  assign n30534 = ~n30496 & ~n30519 ;
  assign n30560 = n30534 & n30537 ;
  assign n30561 = ~n30502 & n30560 ;
  assign n30562 = n30502 & n30530 ;
  assign n30563 = ~n30496 & ~n30562 ;
  assign n30564 = ~n30519 & ~n30537 ;
  assign n30565 = ~n30510 & n30564 ;
  assign n30566 = ~n30563 & n30565 ;
  assign n30567 = ~n30561 & ~n30566 ;
  assign n30568 = ~n30559 & n30567 ;
  assign n30569 = n30552 & ~n30568 ;
  assign n30511 = ~n30496 & n30509 ;
  assign n30512 = n30502 & n30511 ;
  assign n30513 = ~n30510 & ~n30512 ;
  assign n30520 = ~n30513 & ~n30519 ;
  assign n30536 = n30534 & n30535 ;
  assign n30538 = n30496 & ~n30502 ;
  assign n30539 = n30537 & n30538 ;
  assign n30540 = ~n30536 & ~n30539 ;
  assign n30521 = ~n30502 & n30509 ;
  assign n30522 = n30496 & ~n30521 ;
  assign n30523 = ~n30511 & n30519 ;
  assign n30524 = ~n30522 & n30523 ;
  assign n30531 = ~n30509 & n30530 ;
  assign n30532 = ~n30502 & n30519 ;
  assign n30533 = n30531 & n30532 ;
  assign n30541 = n30502 & ~n30530 ;
  assign n30542 = n30511 & n30541 ;
  assign n30543 = ~n30533 & ~n30542 ;
  assign n30544 = ~n30524 & n30543 ;
  assign n30545 = n30540 & n30544 ;
  assign n30546 = ~n30520 & n30545 ;
  assign n30553 = ~n30546 & ~n30552 ;
  assign n30576 = n30502 & n30535 ;
  assign n30577 = ~n30519 & n30576 ;
  assign n30578 = ~n30533 & ~n30577 ;
  assign n30579 = ~n30496 & ~n30578 ;
  assign n30570 = ~n30509 & ~n30530 ;
  assign n30571 = ~n30502 & n30570 ;
  assign n30572 = n30534 & n30571 ;
  assign n30573 = ~n30496 & n30541 ;
  assign n30574 = ~n30537 & ~n30573 ;
  assign n30575 = n30523 & ~n30574 ;
  assign n30580 = ~n30572 & ~n30575 ;
  assign n30581 = ~n30579 & n30580 ;
  assign n30582 = ~n30553 & n30581 ;
  assign n30583 = ~n30569 & n30582 ;
  assign n30584 = ~\u1_L12_reg[11]/NET0131  & n30583 ;
  assign n30585 = \u1_L12_reg[11]/NET0131  & ~n30583 ;
  assign n30586 = ~n30584 & ~n30585 ;
  assign n30587 = decrypt_pad & ~\u1_uk_K_r12_reg[27]/NET0131  ;
  assign n30588 = ~decrypt_pad & ~\u1_uk_K_r12_reg[19]/NET0131  ;
  assign n30589 = ~n30587 & ~n30588 ;
  assign n30590 = \u1_R12_reg[13]/NET0131  & ~n30589 ;
  assign n30591 = ~\u1_R12_reg[13]/NET0131  & n30589 ;
  assign n30592 = ~n30590 & ~n30591 ;
  assign n30600 = decrypt_pad & ~\u1_uk_K_r12_reg[33]/NET0131  ;
  assign n30601 = ~decrypt_pad & ~\u1_uk_K_r12_reg[25]/NET0131  ;
  assign n30602 = ~n30600 & ~n30601 ;
  assign n30603 = \u1_R12_reg[12]/NET0131  & ~n30602 ;
  assign n30604 = ~\u1_R12_reg[12]/NET0131  & n30602 ;
  assign n30605 = ~n30603 & ~n30604 ;
  assign n30606 = decrypt_pad & ~\u1_uk_K_r12_reg[17]/NET0131  ;
  assign n30607 = ~decrypt_pad & ~\u1_uk_K_r12_reg[41]/NET0131  ;
  assign n30608 = ~n30606 & ~n30607 ;
  assign n30609 = \u1_R12_reg[17]/NET0131  & ~n30608 ;
  assign n30610 = ~\u1_R12_reg[17]/NET0131  & n30608 ;
  assign n30611 = ~n30609 & ~n30610 ;
  assign n30612 = ~n30605 & ~n30611 ;
  assign n30613 = decrypt_pad & ~\u1_uk_K_r12_reg[53]/NET0131  ;
  assign n30614 = ~decrypt_pad & ~\u1_uk_K_r12_reg[20]/NET0131  ;
  assign n30615 = ~n30613 & ~n30614 ;
  assign n30616 = \u1_R12_reg[14]/NET0131  & ~n30615 ;
  assign n30617 = ~\u1_R12_reg[14]/NET0131  & n30615 ;
  assign n30618 = ~n30616 & ~n30617 ;
  assign n30619 = n30612 & ~n30618 ;
  assign n30631 = ~n30592 & n30619 ;
  assign n30632 = n30592 & n30612 ;
  assign n30633 = n30618 & n30632 ;
  assign n30634 = ~n30631 & ~n30633 ;
  assign n30593 = decrypt_pad & ~\u1_uk_K_r12_reg[4]/NET0131  ;
  assign n30594 = ~decrypt_pad & ~\u1_uk_K_r12_reg[53]/NET0131  ;
  assign n30595 = ~n30593 & ~n30594 ;
  assign n30596 = \u1_R12_reg[15]/NET0131  & ~n30595 ;
  assign n30597 = ~\u1_R12_reg[15]/NET0131  & n30595 ;
  assign n30598 = ~n30596 & ~n30597 ;
  assign n30624 = n30592 & n30598 ;
  assign n30638 = n30618 & n30624 ;
  assign n30639 = ~n30605 & n30638 ;
  assign n30635 = ~n30592 & n30605 ;
  assign n30636 = n30611 & ~n30618 ;
  assign n30637 = n30635 & n30636 ;
  assign n30640 = decrypt_pad & ~\u1_uk_K_r12_reg[12]/NET0131  ;
  assign n30641 = ~decrypt_pad & ~\u1_uk_K_r12_reg[4]/NET0131  ;
  assign n30642 = ~n30640 & ~n30641 ;
  assign n30643 = \u1_R12_reg[16]/NET0131  & ~n30642 ;
  assign n30644 = ~\u1_R12_reg[16]/NET0131  & n30642 ;
  assign n30645 = ~n30643 & ~n30644 ;
  assign n30656 = ~n30637 & ~n30645 ;
  assign n30657 = ~n30639 & n30656 ;
  assign n30658 = n30634 & n30657 ;
  assign n30620 = n30605 & ~n30611 ;
  assign n30621 = n30618 & n30620 ;
  assign n30646 = ~n30592 & n30611 ;
  assign n30647 = ~n30621 & ~n30646 ;
  assign n30648 = ~n30598 & ~n30647 ;
  assign n30652 = n30605 & n30611 ;
  assign n30653 = ~n30612 & ~n30652 ;
  assign n30649 = n30592 & n30605 ;
  assign n30650 = ~n30592 & ~n30605 ;
  assign n30651 = ~n30649 & ~n30650 ;
  assign n30654 = n30598 & ~n30651 ;
  assign n30655 = ~n30653 & n30654 ;
  assign n30659 = ~n30648 & ~n30655 ;
  assign n30660 = n30658 & n30659 ;
  assign n30625 = n30620 & n30624 ;
  assign n30627 = ~n30605 & n30611 ;
  assign n30628 = n30592 & n30627 ;
  assign n30661 = ~n30618 & n30628 ;
  assign n30662 = ~n30625 & ~n30661 ;
  assign n30663 = ~n30598 & ~n30611 ;
  assign n30664 = n30618 & n30650 ;
  assign n30665 = n30663 & n30664 ;
  assign n30670 = n30611 & n30618 ;
  assign n30671 = n30649 & n30670 ;
  assign n30672 = n30645 & ~n30671 ;
  assign n30673 = ~n30665 & n30672 ;
  assign n30629 = ~n30598 & ~n30618 ;
  assign n30666 = n30629 & n30651 ;
  assign n30667 = n30598 & n30611 ;
  assign n30668 = ~n30605 & n30667 ;
  assign n30669 = ~n30592 & n30668 ;
  assign n30674 = ~n30666 & ~n30669 ;
  assign n30675 = n30673 & n30674 ;
  assign n30676 = n30662 & n30675 ;
  assign n30677 = ~n30660 & ~n30676 ;
  assign n30599 = ~n30592 & n30598 ;
  assign n30622 = ~n30619 & ~n30621 ;
  assign n30623 = n30599 & ~n30622 ;
  assign n30626 = ~n30618 & n30625 ;
  assign n30630 = n30628 & n30629 ;
  assign n30678 = ~n30626 & ~n30630 ;
  assign n30679 = ~n30623 & n30678 ;
  assign n30680 = ~n30677 & n30679 ;
  assign n30681 = ~\u1_L12_reg[20]/NET0131  & ~n30680 ;
  assign n30682 = \u1_L12_reg[20]/NET0131  & n30680 ;
  assign n30683 = ~n30681 & ~n30682 ;
  assign n30705 = ~n30409 & ~n30429 ;
  assign n30706 = ~n30422 & ~n30705 ;
  assign n30707 = n30442 & n30705 ;
  assign n30708 = ~n30706 & ~n30707 ;
  assign n30709 = n30440 & ~n30708 ;
  assign n30710 = ~n30440 & ~n30482 ;
  assign n30711 = ~n30706 & n30710 ;
  assign n30684 = n30409 & n30429 ;
  assign n30703 = n30415 & n30684 ;
  assign n30704 = n30422 & n30458 ;
  assign n30712 = ~n30703 & ~n30704 ;
  assign n30713 = ~n30711 & n30712 ;
  assign n30714 = ~n30709 & n30713 ;
  assign n30715 = n30403 & ~n30714 ;
  assign n30687 = ~n30409 & ~n30444 ;
  assign n30688 = ~n30422 & n30457 ;
  assign n30689 = ~n30687 & ~n30688 ;
  assign n30690 = ~n30440 & ~n30689 ;
  assign n30691 = ~n30423 & ~n30459 ;
  assign n30692 = n30440 & ~n30691 ;
  assign n30685 = ~n30415 & n30684 ;
  assign n30686 = n30422 & n30685 ;
  assign n30693 = n30429 & n30461 ;
  assign n30694 = ~n30686 & ~n30693 ;
  assign n30695 = ~n30692 & n30694 ;
  assign n30696 = ~n30690 & n30695 ;
  assign n30697 = ~n30403 & ~n30696 ;
  assign n30700 = n30429 & ~n30448 ;
  assign n30698 = n30409 & n30460 ;
  assign n30699 = ~n30429 & ~n30698 ;
  assign n30701 = n30440 & ~n30699 ;
  assign n30702 = ~n30700 & n30701 ;
  assign n30716 = ~n30697 & ~n30702 ;
  assign n30717 = ~n30715 & n30716 ;
  assign n30718 = ~\u1_L12_reg[17]/NET0131  & ~n30717 ;
  assign n30719 = \u1_L12_reg[17]/NET0131  & n30717 ;
  assign n30720 = ~n30718 & ~n30719 ;
  assign n30729 = n30311 & n30384 ;
  assign n30726 = n30305 & n30325 ;
  assign n30727 = ~n30341 & ~n30355 ;
  assign n30728 = ~n30305 & ~n30727 ;
  assign n30733 = ~n30726 & ~n30728 ;
  assign n30734 = ~n30729 & n30733 ;
  assign n30722 = ~n30305 & n30344 ;
  assign n30721 = n30318 & n30336 ;
  assign n30730 = ~n30354 & ~n30721 ;
  assign n30731 = ~n30722 & n30730 ;
  assign n30723 = ~n30324 & ~n30331 ;
  assign n30724 = n30335 & ~n30336 ;
  assign n30725 = ~n30723 & n30724 ;
  assign n30732 = ~n30371 & ~n30725 ;
  assign n30735 = n30731 & n30732 ;
  assign n30736 = n30734 & n30735 ;
  assign n30740 = ~n30341 & ~n30345 ;
  assign n30741 = ~n30344 & ~n30355 ;
  assign n30742 = ~n30740 & ~n30741 ;
  assign n30743 = ~n30337 & n30354 ;
  assign n30744 = ~n30378 & n30743 ;
  assign n30745 = ~n30742 & n30744 ;
  assign n30737 = ~n30305 & n30332 ;
  assign n30738 = ~n30364 & ~n30376 ;
  assign n30739 = n30305 & ~n30738 ;
  assign n30746 = ~n30737 & ~n30739 ;
  assign n30747 = n30745 & n30746 ;
  assign n30748 = ~n30736 & ~n30747 ;
  assign n30749 = \u1_L12_reg[12]/NET0131  & n30748 ;
  assign n30750 = ~\u1_L12_reg[12]/NET0131  & ~n30748 ;
  assign n30751 = ~n30749 & ~n30750 ;
  assign n30752 = decrypt_pad & ~\u1_uk_K_r12_reg[43]/NET0131  ;
  assign n30753 = ~decrypt_pad & ~\u1_uk_K_r12_reg[37]/NET0131  ;
  assign n30754 = ~n30752 & ~n30753 ;
  assign n30755 = \u1_R12_reg[28]/NET0131  & ~n30754 ;
  assign n30756 = ~\u1_R12_reg[28]/NET0131  & n30754 ;
  assign n30757 = ~n30755 & ~n30756 ;
  assign n30758 = decrypt_pad & ~\u1_uk_K_r12_reg[15]/NET0131  ;
  assign n30759 = ~decrypt_pad & ~\u1_uk_K_r12_reg[9]/NET0131  ;
  assign n30760 = ~n30758 & ~n30759 ;
  assign n30761 = \u1_R12_reg[29]/NET0131  & ~n30760 ;
  assign n30762 = ~\u1_R12_reg[29]/NET0131  & n30760 ;
  assign n30763 = ~n30761 & ~n30762 ;
  assign n30764 = n30757 & ~n30763 ;
  assign n30765 = decrypt_pad & ~\u1_uk_K_r12_reg[0]/NET0131  ;
  assign n30766 = ~decrypt_pad & ~\u1_uk_K_r12_reg[49]/NET0131  ;
  assign n30767 = ~n30765 & ~n30766 ;
  assign n30768 = \u1_R12_reg[1]/NET0131  & ~n30767 ;
  assign n30769 = ~\u1_R12_reg[1]/NET0131  & n30767 ;
  assign n30770 = ~n30768 & ~n30769 ;
  assign n30773 = decrypt_pad & ~\u1_uk_K_r12_reg[16]/NET0131  ;
  assign n30774 = ~decrypt_pad & ~\u1_uk_K_r12_reg[38]/NET0131  ;
  assign n30775 = ~n30773 & ~n30774 ;
  assign n30776 = \u1_R12_reg[30]/NET0131  & ~n30775 ;
  assign n30777 = ~\u1_R12_reg[30]/NET0131  & n30775 ;
  assign n30778 = ~n30776 & ~n30777 ;
  assign n30786 = ~n30757 & n30778 ;
  assign n30787 = ~n30770 & n30786 ;
  assign n30788 = n30763 & n30787 ;
  assign n30789 = ~n30757 & ~n30763 ;
  assign n30790 = ~n30778 & n30789 ;
  assign n30791 = ~n30770 & n30790 ;
  assign n30792 = ~n30788 & ~n30791 ;
  assign n30771 = n30763 & n30770 ;
  assign n30772 = ~n30757 & n30771 ;
  assign n30779 = n30772 & ~n30778 ;
  assign n30780 = decrypt_pad & ~\u1_uk_K_r12_reg[28]/NET0131  ;
  assign n30781 = ~decrypt_pad & ~\u1_uk_K_r12_reg[22]/NET0131  ;
  assign n30782 = ~n30780 & ~n30781 ;
  assign n30783 = \u1_R12_reg[31]/NET0131  & ~n30782 ;
  assign n30784 = ~\u1_R12_reg[31]/NET0131  & n30782 ;
  assign n30785 = ~n30783 & ~n30784 ;
  assign n30793 = n30757 & n30778 ;
  assign n30794 = ~n30763 & n30793 ;
  assign n30795 = ~n30785 & ~n30794 ;
  assign n30796 = ~n30779 & n30795 ;
  assign n30797 = n30792 & n30796 ;
  assign n30798 = ~n30764 & n30797 ;
  assign n30803 = n30770 & n30789 ;
  assign n30804 = ~n30778 & n30803 ;
  assign n30805 = n30771 & n30786 ;
  assign n30806 = n30785 & ~n30805 ;
  assign n30807 = ~n30804 & n30806 ;
  assign n30799 = n30757 & n30763 ;
  assign n30800 = n30763 & ~n30778 ;
  assign n30801 = ~n30770 & n30800 ;
  assign n30802 = ~n30799 & ~n30801 ;
  assign n30808 = n30802 & ~n30803 ;
  assign n30809 = n30807 & n30808 ;
  assign n30810 = ~n30798 & ~n30809 ;
  assign n30811 = decrypt_pad & ~\u1_uk_K_r12_reg[38]/NET0131  ;
  assign n30812 = ~decrypt_pad & ~\u1_uk_K_r12_reg[28]/NET0131  ;
  assign n30813 = ~n30811 & ~n30812 ;
  assign n30814 = \u1_R12_reg[32]/NET0131  & ~n30813 ;
  assign n30815 = ~\u1_R12_reg[32]/NET0131  & n30813 ;
  assign n30816 = ~n30814 & ~n30815 ;
  assign n30817 = ~n30763 & ~n30770 ;
  assign n30818 = n30757 & ~n30778 ;
  assign n30819 = n30817 & n30818 ;
  assign n30820 = ~n30816 & ~n30819 ;
  assign n30821 = ~n30810 & n30820 ;
  assign n30822 = ~n30770 & n30789 ;
  assign n30823 = n30807 & ~n30822 ;
  assign n30824 = ~n30797 & ~n30823 ;
  assign n30829 = ~n30778 & n30799 ;
  assign n30825 = n30770 & ~n30785 ;
  assign n30826 = ~n30763 & n30778 ;
  assign n30827 = n30825 & n30826 ;
  assign n30830 = n30816 & ~n30827 ;
  assign n30831 = ~n30829 & n30830 ;
  assign n30828 = n30770 & n30794 ;
  assign n30832 = ~n30788 & ~n30828 ;
  assign n30833 = n30831 & n30832 ;
  assign n30834 = ~n30824 & n30833 ;
  assign n30835 = ~n30821 & ~n30834 ;
  assign n30836 = ~\u1_L12_reg[15]/P0001  & n30835 ;
  assign n30837 = \u1_L12_reg[15]/P0001  & ~n30835 ;
  assign n30838 = ~n30836 & ~n30837 ;
  assign n30840 = n30592 & ~n30618 ;
  assign n30855 = ~n30605 & ~n30840 ;
  assign n30856 = ~n30618 & n30649 ;
  assign n30857 = ~n30855 & ~n30856 ;
  assign n30858 = ~n30620 & ~n30857 ;
  assign n30850 = n30605 & ~n30618 ;
  assign n30851 = ~n30611 & ~n30850 ;
  assign n30859 = ~n30599 & ~n30851 ;
  assign n30860 = ~n30858 & n30859 ;
  assign n30852 = n30618 & ~n30635 ;
  assign n30853 = n30598 & n30851 ;
  assign n30854 = ~n30852 & n30853 ;
  assign n30861 = ~n30645 & ~n30854 ;
  assign n30862 = ~n30860 & n30861 ;
  assign n30839 = n30592 & n30621 ;
  assign n30863 = n30645 & ~n30839 ;
  assign n30864 = n30599 & ~n30851 ;
  assign n30865 = ~n30664 & ~n30864 ;
  assign n30866 = n30863 & n30865 ;
  assign n30867 = ~n30862 & ~n30866 ;
  assign n30841 = ~n30620 & n30840 ;
  assign n30842 = ~n30628 & ~n30841 ;
  assign n30843 = n30645 & ~n30842 ;
  assign n30844 = ~n30598 & ~n30839 ;
  assign n30845 = ~n30843 & n30844 ;
  assign n30846 = ~n30651 & n30670 ;
  assign n30847 = n30598 & ~n30633 ;
  assign n30848 = ~n30846 & n30847 ;
  assign n30849 = ~n30845 & ~n30848 ;
  assign n30868 = ~n30665 & ~n30849 ;
  assign n30869 = ~n30867 & n30868 ;
  assign n30870 = ~\u1_L12_reg[1]/NET0131  & ~n30869 ;
  assign n30871 = \u1_L12_reg[1]/NET0131  & n30869 ;
  assign n30872 = ~n30870 & ~n30871 ;
  assign n30899 = n30763 & n30793 ;
  assign n30897 = ~n30763 & n30770 ;
  assign n30898 = ~n30778 & n30897 ;
  assign n30900 = ~n30772 & ~n30898 ;
  assign n30901 = ~n30899 & n30900 ;
  assign n30902 = n30785 & ~n30901 ;
  assign n30894 = ~n30770 & n30818 ;
  assign n30895 = ~n30828 & ~n30894 ;
  assign n30896 = ~n30785 & ~n30895 ;
  assign n30884 = ~n30770 & n30799 ;
  assign n30892 = ~n30822 & ~n30884 ;
  assign n30893 = n30778 & ~n30892 ;
  assign n30903 = ~n30804 & ~n30893 ;
  assign n30904 = ~n30896 & n30903 ;
  assign n30905 = ~n30902 & n30904 ;
  assign n30906 = n30816 & ~n30905 ;
  assign n30885 = ~n30794 & ~n30884 ;
  assign n30886 = n30785 & ~n30885 ;
  assign n30875 = ~n30786 & ~n30818 ;
  assign n30876 = n30757 & ~n30770 ;
  assign n30877 = n30763 & ~n30876 ;
  assign n30878 = ~n30825 & ~n30877 ;
  assign n30879 = ~n30875 & ~n30878 ;
  assign n30880 = n30793 & n30817 ;
  assign n30881 = n30763 & ~n30770 ;
  assign n30882 = ~n30757 & ~n30785 ;
  assign n30883 = n30881 & n30882 ;
  assign n30887 = ~n30880 & ~n30883 ;
  assign n30888 = ~n30791 & n30887 ;
  assign n30889 = ~n30879 & n30888 ;
  assign n30890 = ~n30886 & n30889 ;
  assign n30891 = ~n30816 & ~n30890 ;
  assign n30873 = n30825 & n30829 ;
  assign n30874 = n30785 & n30790 ;
  assign n30907 = ~n30873 & ~n30874 ;
  assign n30908 = ~n30891 & n30907 ;
  assign n30909 = ~n30906 & n30908 ;
  assign n30910 = ~\u1_L12_reg[21]/NET0131  & ~n30909 ;
  assign n30911 = \u1_L12_reg[21]/NET0131  & n30909 ;
  assign n30912 = ~n30910 & ~n30911 ;
  assign n30913 = ~n30599 & ~n30840 ;
  assign n30914 = n30612 & ~n30913 ;
  assign n30921 = n30863 & ~n30914 ;
  assign n30915 = ~n30628 & ~n30668 ;
  assign n30916 = n30618 & ~n30915 ;
  assign n30917 = ~n30592 & n30636 ;
  assign n30918 = ~n30652 & ~n30917 ;
  assign n30919 = ~n30598 & ~n30850 ;
  assign n30920 = ~n30918 & n30919 ;
  assign n30922 = ~n30916 & ~n30920 ;
  assign n30923 = n30921 & n30922 ;
  assign n30924 = ~n30627 & n30638 ;
  assign n30928 = ~n30645 & ~n30924 ;
  assign n30925 = ~n30598 & n30664 ;
  assign n30926 = ~n30663 & ~n30850 ;
  assign n30927 = ~n30592 & ~n30926 ;
  assign n30929 = ~n30925 & ~n30927 ;
  assign n30930 = n30928 & n30929 ;
  assign n30931 = n30662 & n30930 ;
  assign n30932 = ~n30923 & ~n30931 ;
  assign n30933 = ~n30663 & ~n30667 ;
  assign n30936 = ~n30651 & ~n30933 ;
  assign n30934 = ~n30598 & n30649 ;
  assign n30935 = n30933 & ~n30934 ;
  assign n30937 = ~n30618 & ~n30935 ;
  assign n30938 = ~n30936 & n30937 ;
  assign n30939 = ~n30932 & ~n30938 ;
  assign n30940 = ~\u1_L12_reg[26]/NET0131  & ~n30939 ;
  assign n30941 = \u1_L12_reg[26]/NET0131  & n30939 ;
  assign n30942 = ~n30940 & ~n30941 ;
  assign n30959 = ~n30502 & n30535 ;
  assign n30960 = ~n30556 & ~n30959 ;
  assign n30961 = ~n30510 & ~n30554 ;
  assign n30962 = ~n30530 & ~n30961 ;
  assign n30963 = n30960 & ~n30962 ;
  assign n30964 = n30519 & ~n30963 ;
  assign n30943 = n30496 & ~n30535 ;
  assign n30947 = n30502 & ~n30511 ;
  assign n30948 = ~n30943 & n30947 ;
  assign n30965 = ~n30519 & n30948 ;
  assign n30966 = n30531 & n30538 ;
  assign n30967 = ~n30560 & ~n30966 ;
  assign n30968 = ~n30965 & n30967 ;
  assign n30969 = ~n30964 & n30968 ;
  assign n30970 = ~n30552 & ~n30969 ;
  assign n30949 = n30502 & n30531 ;
  assign n30950 = ~n30948 & ~n30949 ;
  assign n30951 = n30519 & ~n30950 ;
  assign n30944 = ~n30531 & n30943 ;
  assign n30945 = ~n30571 & ~n30944 ;
  assign n30946 = ~n30519 & ~n30945 ;
  assign n30953 = n30496 & n30571 ;
  assign n30952 = n30531 & n30554 ;
  assign n30954 = n30540 & ~n30952 ;
  assign n30955 = ~n30953 & n30954 ;
  assign n30956 = ~n30946 & n30955 ;
  assign n30957 = ~n30951 & n30956 ;
  assign n30958 = n30552 & ~n30957 ;
  assign n30971 = ~n30496 & n30519 ;
  assign n30972 = n30562 & n30971 ;
  assign n30973 = ~n30555 & ~n30972 ;
  assign n30974 = ~n30958 & n30973 ;
  assign n30975 = ~n30970 & n30974 ;
  assign n30976 = \u1_L12_reg[29]/NET0131  & ~n30975 ;
  assign n30977 = ~\u1_L12_reg[29]/NET0131  & n30975 ;
  assign n30978 = ~n30976 & ~n30977 ;
  assign n30979 = decrypt_pad & ~\u1_uk_K_r12_reg[24]/NET0131  ;
  assign n30980 = ~decrypt_pad & ~\u1_uk_K_r12_reg[48]/NET0131  ;
  assign n30981 = ~n30979 & ~n30980 ;
  assign n30982 = \u1_R12_reg[4]/NET0131  & ~n30981 ;
  assign n30983 = ~\u1_R12_reg[4]/NET0131  & n30981 ;
  assign n30984 = ~n30982 & ~n30983 ;
  assign n30985 = decrypt_pad & ~\u1_uk_K_r12_reg[48]/NET0131  ;
  assign n30986 = ~decrypt_pad & ~\u1_uk_K_r12_reg[40]/NET0131  ;
  assign n30987 = ~n30985 & ~n30986 ;
  assign n30988 = \u1_R12_reg[9]/NET0131  & ~n30987 ;
  assign n30989 = ~\u1_R12_reg[9]/NET0131  & n30987 ;
  assign n30990 = ~n30988 & ~n30989 ;
  assign n30991 = n30984 & ~n30990 ;
  assign n30992 = ~n30984 & n30990 ;
  assign n30993 = decrypt_pad & ~\u1_uk_K_r12_reg[3]/NET0131  ;
  assign n30994 = ~decrypt_pad & ~\u1_uk_K_r12_reg[27]/NET0131  ;
  assign n30995 = ~n30993 & ~n30994 ;
  assign n30996 = \u1_R12_reg[5]/NET0131  & ~n30995 ;
  assign n30997 = ~\u1_R12_reg[5]/NET0131  & n30995 ;
  assign n30998 = ~n30996 & ~n30997 ;
  assign n30999 = n30992 & ~n30998 ;
  assign n31000 = n30984 & n30998 ;
  assign n31001 = ~n30999 & ~n31000 ;
  assign n31002 = ~n30991 & n31001 ;
  assign n31003 = decrypt_pad & ~\u1_uk_K_r12_reg[26]/NET0131  ;
  assign n31004 = ~decrypt_pad & ~\u1_uk_K_r12_reg[18]/NET0131  ;
  assign n31005 = ~n31003 & ~n31004 ;
  assign n31006 = \u1_R12_reg[6]/NET0131  & ~n31005 ;
  assign n31007 = ~\u1_R12_reg[6]/NET0131  & n31005 ;
  assign n31008 = ~n31006 & ~n31007 ;
  assign n31009 = decrypt_pad & ~\u1_uk_K_r12_reg[20]/NET0131  ;
  assign n31010 = ~decrypt_pad & ~\u1_uk_K_r12_reg[12]/NET0131  ;
  assign n31011 = ~n31009 & ~n31010 ;
  assign n31012 = \u1_R12_reg[7]/NET0131  & ~n31011 ;
  assign n31013 = ~\u1_R12_reg[7]/NET0131  & n31011 ;
  assign n31014 = ~n31012 & ~n31013 ;
  assign n31015 = n31008 & ~n31014 ;
  assign n31016 = ~n31002 & n31015 ;
  assign n31017 = ~n30990 & n30998 ;
  assign n31018 = ~n30999 & ~n31017 ;
  assign n31019 = ~n31008 & ~n31018 ;
  assign n31020 = decrypt_pad & ~\u1_uk_K_r12_reg[11]/NET0131  ;
  assign n31021 = ~decrypt_pad & ~\u1_uk_K_r12_reg[3]/NET0131  ;
  assign n31022 = ~n31020 & ~n31021 ;
  assign n31023 = \u1_R12_reg[8]/NET0131  & ~n31022 ;
  assign n31024 = ~\u1_R12_reg[8]/NET0131  & n31022 ;
  assign n31025 = ~n31023 & ~n31024 ;
  assign n31037 = ~n31019 & ~n31025 ;
  assign n31026 = n30984 & n30990 ;
  assign n31027 = n31008 & n31026 ;
  assign n31028 = ~n30998 & n31027 ;
  assign n31029 = n31014 & n31028 ;
  assign n31030 = ~n30984 & n31008 ;
  assign n31032 = n30998 & ~n31030 ;
  assign n31031 = n31014 & ~n31030 ;
  assign n31033 = ~n30998 & n31008 ;
  assign n31034 = n30990 & ~n31033 ;
  assign n31035 = ~n31031 & n31034 ;
  assign n31036 = ~n31032 & n31035 ;
  assign n31038 = ~n31029 & ~n31036 ;
  assign n31039 = n31037 & n31038 ;
  assign n31040 = ~n31016 & n31039 ;
  assign n31042 = n30991 & ~n30998 ;
  assign n31043 = n30998 & n31026 ;
  assign n31044 = ~n31042 & ~n31043 ;
  assign n31045 = ~n31008 & ~n31044 ;
  assign n31041 = n31014 & n31032 ;
  assign n31046 = n31025 & ~n31041 ;
  assign n31047 = ~n31045 & n31046 ;
  assign n31048 = ~n31040 & ~n31047 ;
  assign n31049 = n30998 & ~n31008 ;
  assign n31050 = ~n30984 & ~n30990 ;
  assign n31051 = ~n31028 & ~n31050 ;
  assign n31052 = n31025 & ~n31051 ;
  assign n31053 = ~n30984 & ~n31033 ;
  assign n31054 = n30990 & n31053 ;
  assign n31055 = ~n31052 & ~n31054 ;
  assign n31056 = ~n31049 & ~n31055 ;
  assign n31057 = ~n31014 & ~n31056 ;
  assign n31058 = ~n30998 & n31030 ;
  assign n31059 = ~n30990 & n31058 ;
  assign n31060 = n30984 & ~n31008 ;
  assign n31061 = n30998 & n31060 ;
  assign n31062 = n31014 & ~n31061 ;
  assign n31063 = ~n31059 & n31062 ;
  assign n31064 = ~n31057 & ~n31063 ;
  assign n31065 = ~n31048 & ~n31064 ;
  assign n31066 = \u1_L12_reg[2]/NET0131  & n31065 ;
  assign n31067 = ~\u1_L12_reg[2]/NET0131  & ~n31065 ;
  assign n31068 = ~n31066 & ~n31067 ;
  assign n31073 = n30992 & n30998 ;
  assign n31074 = ~n31008 & n31050 ;
  assign n31075 = ~n31073 & ~n31074 ;
  assign n31076 = ~n30990 & n31008 ;
  assign n31077 = n31000 & n31076 ;
  assign n31078 = ~n31014 & ~n31058 ;
  assign n31079 = ~n31077 & n31078 ;
  assign n31080 = n31075 & n31079 ;
  assign n31081 = ~n30984 & n31017 ;
  assign n31082 = n31008 & n31081 ;
  assign n31083 = n31014 & n31044 ;
  assign n31084 = ~n31082 & n31083 ;
  assign n31085 = ~n31080 & ~n31084 ;
  assign n31069 = ~n30998 & n31026 ;
  assign n31070 = ~n31014 & ~n31069 ;
  assign n31071 = n31060 & ~n31070 ;
  assign n31072 = n30992 & n31033 ;
  assign n31086 = n31025 & ~n31072 ;
  assign n31087 = ~n31071 & n31086 ;
  assign n31088 = ~n31085 & n31087 ;
  assign n31089 = n31014 & n31075 ;
  assign n31090 = n30991 & ~n31008 ;
  assign n31091 = n31001 & ~n31090 ;
  assign n31092 = n31079 & n31091 ;
  assign n31093 = ~n31089 & ~n31092 ;
  assign n31094 = ~n30992 & n31008 ;
  assign n31095 = ~n30991 & n30998 ;
  assign n31096 = ~n31042 & ~n31095 ;
  assign n31097 = n31094 & n31096 ;
  assign n31098 = ~n31025 & ~n31097 ;
  assign n31099 = ~n31093 & n31098 ;
  assign n31100 = ~n31088 & ~n31099 ;
  assign n31101 = ~\u1_L12_reg[28]/NET0131  & n31100 ;
  assign n31102 = \u1_L12_reg[28]/NET0131  & ~n31100 ;
  assign n31103 = ~n31101 & ~n31102 ;
  assign n31114 = n30509 & n30971 ;
  assign n31115 = ~n30503 & ~n31114 ;
  assign n31116 = n30530 & ~n31115 ;
  assign n31112 = ~n30534 & ~n30573 ;
  assign n31113 = ~n30509 & ~n31112 ;
  assign n31111 = n30534 & n30541 ;
  assign n31117 = n30552 & ~n31111 ;
  assign n31118 = ~n31113 & n31117 ;
  assign n31119 = ~n31116 & n31118 ;
  assign n31105 = n30519 & ~n30576 ;
  assign n31120 = ~n30511 & n30530 ;
  assign n31121 = ~n30522 & n31120 ;
  assign n31122 = n31105 & ~n31121 ;
  assign n31123 = n30502 & n30570 ;
  assign n31124 = ~n30519 & ~n30966 ;
  assign n31125 = ~n31123 & n31124 ;
  assign n31126 = ~n31122 & ~n31125 ;
  assign n31127 = ~n30552 & ~n30555 ;
  assign n31128 = ~n30560 & n31127 ;
  assign n31129 = ~n31126 & n31128 ;
  assign n31130 = ~n31119 & ~n31129 ;
  assign n31104 = n30534 & n30570 ;
  assign n31108 = ~n30519 & n30960 ;
  assign n31106 = ~n30571 & ~n30949 ;
  assign n31107 = n31105 & n31106 ;
  assign n31109 = n30496 & ~n31107 ;
  assign n31110 = ~n31108 & n31109 ;
  assign n31131 = ~n31104 & ~n31110 ;
  assign n31132 = ~n31130 & n31131 ;
  assign n31133 = ~\u1_L12_reg[4]/NET0131  & ~n31132 ;
  assign n31134 = \u1_L12_reg[4]/NET0131  & n31132 ;
  assign n31135 = ~n31133 & ~n31134 ;
  assign n31149 = ~n30598 & n30653 ;
  assign n31150 = n30857 & n31149 ;
  assign n31147 = ~n30632 & ~n30637 ;
  assign n31148 = n30598 & ~n31147 ;
  assign n31151 = ~n30846 & ~n31148 ;
  assign n31152 = ~n31150 & n31151 ;
  assign n31153 = n30645 & ~n31152 ;
  assign n31137 = n30629 & n30652 ;
  assign n31136 = n30650 & n30663 ;
  assign n31141 = ~n30856 & ~n31136 ;
  assign n31142 = ~n31137 & n31141 ;
  assign n31138 = n30599 & n30605 ;
  assign n31139 = ~n30636 & n31138 ;
  assign n31140 = ~n30618 & n30668 ;
  assign n31143 = ~n31139 & ~n31140 ;
  assign n31144 = n31142 & n31143 ;
  assign n31145 = n30634 & n31144 ;
  assign n31146 = ~n30645 & ~n31145 ;
  assign n31154 = ~n30631 & ~n30846 ;
  assign n31155 = ~n30598 & ~n31154 ;
  assign n31156 = ~n30626 & ~n30639 ;
  assign n31157 = ~n31155 & n31156 ;
  assign n31158 = ~n31146 & n31157 ;
  assign n31159 = ~n31153 & n31158 ;
  assign n31160 = ~\u1_L12_reg[10]/NET0131  & ~n31159 ;
  assign n31161 = \u1_L12_reg[10]/NET0131  & n31159 ;
  assign n31162 = ~n31160 & ~n31161 ;
  assign n31163 = decrypt_pad & ~\u1_uk_K_r12_reg[51]/NET0131  ;
  assign n31164 = ~decrypt_pad & ~\u1_uk_K_r12_reg[14]/NET0131  ;
  assign n31165 = ~n31163 & ~n31164 ;
  assign n31166 = \u1_R12_reg[21]/NET0131  & ~n31165 ;
  assign n31167 = ~\u1_R12_reg[21]/NET0131  & n31165 ;
  assign n31168 = ~n31166 & ~n31167 ;
  assign n31169 = decrypt_pad & ~\u1_uk_K_r12_reg[52]/NET0131  ;
  assign n31170 = ~decrypt_pad & ~\u1_uk_K_r12_reg[42]/NET0131  ;
  assign n31171 = ~n31169 & ~n31170 ;
  assign n31172 = \u1_R12_reg[18]/NET0131  & ~n31171 ;
  assign n31173 = ~\u1_R12_reg[18]/NET0131  & n31171 ;
  assign n31174 = ~n31172 & ~n31173 ;
  assign n31175 = n31168 & n31174 ;
  assign n31176 = decrypt_pad & ~\u1_uk_K_r12_reg[8]/NET0131  ;
  assign n31177 = ~decrypt_pad & ~\u1_uk_K_r12_reg[2]/NET0131  ;
  assign n31178 = ~n31176 & ~n31177 ;
  assign n31179 = \u1_R12_reg[16]/NET0131  & ~n31178 ;
  assign n31180 = ~\u1_R12_reg[16]/NET0131  & n31178 ;
  assign n31181 = ~n31179 & ~n31180 ;
  assign n31182 = ~n31168 & ~n31181 ;
  assign n31183 = ~n31175 & ~n31182 ;
  assign n31184 = decrypt_pad & ~\u1_uk_K_r12_reg[30]/NET0131  ;
  assign n31185 = ~decrypt_pad & ~\u1_uk_K_r12_reg[52]/NET0131  ;
  assign n31186 = ~n31184 & ~n31185 ;
  assign n31187 = \u1_R12_reg[17]/NET0131  & ~n31186 ;
  assign n31188 = ~\u1_R12_reg[17]/NET0131  & n31186 ;
  assign n31189 = ~n31187 & ~n31188 ;
  assign n31190 = n31181 & ~n31189 ;
  assign n31191 = ~n31174 & n31189 ;
  assign n31192 = ~n31190 & ~n31191 ;
  assign n31193 = ~n31183 & ~n31192 ;
  assign n31204 = ~n31181 & ~n31189 ;
  assign n31205 = n31168 & n31204 ;
  assign n31196 = ~n31168 & n31189 ;
  assign n31197 = n31174 & n31196 ;
  assign n31198 = decrypt_pad & ~\u1_uk_K_r12_reg[35]/NET0131  ;
  assign n31199 = ~decrypt_pad & ~\u1_uk_K_r12_reg[29]/NET0131  ;
  assign n31200 = ~n31198 & ~n31199 ;
  assign n31201 = \u1_R12_reg[19]/NET0131  & ~n31200 ;
  assign n31202 = ~\u1_R12_reg[19]/NET0131  & n31200 ;
  assign n31203 = ~n31201 & ~n31202 ;
  assign n31209 = ~n31197 & ~n31203 ;
  assign n31210 = ~n31205 & n31209 ;
  assign n31194 = ~n31168 & n31190 ;
  assign n31195 = ~n31174 & n31194 ;
  assign n31206 = ~n31174 & n31181 ;
  assign n31207 = n31168 & n31206 ;
  assign n31208 = n31189 & n31207 ;
  assign n31211 = ~n31195 & ~n31208 ;
  assign n31212 = n31210 & n31211 ;
  assign n31213 = n31174 & n31181 ;
  assign n31214 = n31168 & n31213 ;
  assign n31217 = n31203 & ~n31214 ;
  assign n31215 = n31182 & ~n31189 ;
  assign n31216 = ~n31181 & n31191 ;
  assign n31218 = ~n31215 & ~n31216 ;
  assign n31219 = n31217 & n31218 ;
  assign n31220 = ~n31212 & ~n31219 ;
  assign n31221 = ~n31193 & ~n31220 ;
  assign n31222 = decrypt_pad & ~\u1_uk_K_r12_reg[50]/NET0131  ;
  assign n31223 = ~decrypt_pad & ~\u1_uk_K_r12_reg[44]/P0001  ;
  assign n31224 = ~n31222 & ~n31223 ;
  assign n31225 = \u1_R12_reg[20]/NET0131  & ~n31224 ;
  assign n31226 = ~\u1_R12_reg[20]/NET0131  & n31224 ;
  assign n31227 = ~n31225 & ~n31226 ;
  assign n31228 = ~n31221 & ~n31227 ;
  assign n31229 = n31181 & n31196 ;
  assign n31230 = n31168 & ~n31213 ;
  assign n31231 = ~n31216 & n31230 ;
  assign n31232 = ~n31229 & ~n31231 ;
  assign n31233 = n31203 & ~n31232 ;
  assign n31238 = ~n31174 & ~n31181 ;
  assign n31239 = ~n31214 & ~n31238 ;
  assign n31234 = n31168 & ~n31189 ;
  assign n31235 = ~n31196 & ~n31234 ;
  assign n31240 = ~n31203 & n31235 ;
  assign n31241 = ~n31239 & n31240 ;
  assign n31236 = n31206 & ~n31235 ;
  assign n31237 = n31174 & n31194 ;
  assign n31242 = ~n31236 & ~n31237 ;
  assign n31243 = ~n31241 & n31242 ;
  assign n31244 = ~n31233 & n31243 ;
  assign n31245 = n31227 & ~n31244 ;
  assign n31246 = n31174 & ~n31181 ;
  assign n31247 = ~n31235 & n31246 ;
  assign n31248 = ~n31203 & n31247 ;
  assign n31249 = n31174 & n31215 ;
  assign n31250 = ~n31174 & n31229 ;
  assign n31251 = ~n31249 & ~n31250 ;
  assign n31252 = n31203 & ~n31251 ;
  assign n31253 = ~n31248 & ~n31252 ;
  assign n31254 = ~n31245 & n31253 ;
  assign n31255 = ~n31228 & n31254 ;
  assign n31256 = ~\u1_L12_reg[14]/NET0131  & ~n31255 ;
  assign n31257 = \u1_L12_reg[14]/NET0131  & n31255 ;
  assign n31258 = ~n31256 & ~n31257 ;
  assign n31272 = ~n31168 & ~n31191 ;
  assign n31273 = ~n31213 & n31272 ;
  assign n31260 = n31168 & n31189 ;
  assign n31271 = n31181 & n31260 ;
  assign n31274 = ~n31204 & ~n31271 ;
  assign n31275 = ~n31273 & n31274 ;
  assign n31276 = n31203 & ~n31275 ;
  assign n31278 = n31181 & n31234 ;
  assign n31279 = ~n31216 & ~n31278 ;
  assign n31280 = ~n31203 & ~n31279 ;
  assign n31277 = n31168 & n31191 ;
  assign n31281 = n31181 & n31197 ;
  assign n31282 = ~n31277 & ~n31281 ;
  assign n31283 = ~n31280 & n31282 ;
  assign n31284 = ~n31276 & n31283 ;
  assign n31285 = n31227 & ~n31284 ;
  assign n31259 = n31189 & ~n31246 ;
  assign n31261 = ~n31204 & ~n31234 ;
  assign n31262 = ~n31203 & n31261 ;
  assign n31263 = ~n31260 & ~n31262 ;
  assign n31264 = ~n31259 & ~n31263 ;
  assign n31266 = ~n31203 & ~n31204 ;
  assign n31265 = ~n31196 & n31203 ;
  assign n31267 = ~n31174 & ~n31265 ;
  assign n31268 = ~n31266 & n31267 ;
  assign n31269 = ~n31264 & ~n31268 ;
  assign n31270 = ~n31227 & ~n31269 ;
  assign n31288 = ~n31249 & ~n31281 ;
  assign n31289 = n31168 & n31238 ;
  assign n31290 = ~n31189 & n31289 ;
  assign n31291 = n31288 & ~n31290 ;
  assign n31292 = n31203 & ~n31291 ;
  assign n31286 = n31174 & ~n31203 ;
  assign n31287 = n31190 & n31286 ;
  assign n31293 = ~n31208 & ~n31287 ;
  assign n31294 = ~n31292 & n31293 ;
  assign n31295 = ~n31270 & n31294 ;
  assign n31296 = ~n31285 & n31295 ;
  assign n31297 = ~\u1_L12_reg[25]/NET0131  & ~n31296 ;
  assign n31298 = \u1_L12_reg[25]/NET0131  & n31296 ;
  assign n31299 = ~n31297 & ~n31298 ;
  assign n31305 = ~n31014 & ~n31072 ;
  assign n31306 = ~n31081 & n31305 ;
  assign n31300 = ~n30990 & ~n30998 ;
  assign n31301 = ~n31008 & n31300 ;
  assign n31302 = n30984 & n31301 ;
  assign n31303 = n30992 & n31049 ;
  assign n31304 = ~n31025 & ~n31303 ;
  assign n31307 = ~n31302 & n31304 ;
  assign n31308 = n31306 & n31307 ;
  assign n31309 = n31008 & n31300 ;
  assign n31310 = n31070 & ~n31309 ;
  assign n31311 = n30990 & n31030 ;
  assign n31312 = n31014 & ~n31301 ;
  assign n31313 = ~n31311 & n31312 ;
  assign n31314 = ~n31310 & ~n31313 ;
  assign n31315 = ~n31008 & n31081 ;
  assign n31316 = n31025 & ~n31315 ;
  assign n31317 = ~n31036 & n31316 ;
  assign n31318 = ~n31314 & n31317 ;
  assign n31319 = ~n31308 & ~n31318 ;
  assign n31320 = n30990 & n31060 ;
  assign n31321 = n30998 & n31320 ;
  assign n31322 = ~n31077 & ~n31321 ;
  assign n31323 = ~n31319 & n31322 ;
  assign n31325 = ~n31008 & n31096 ;
  assign n31324 = ~n31017 & n31094 ;
  assign n31326 = n31014 & n31304 ;
  assign n31327 = ~n31324 & n31326 ;
  assign n31328 = ~n31325 & n31327 ;
  assign n31329 = ~n31323 & ~n31328 ;
  assign n31330 = ~\u1_L12_reg[13]/NET0131  & ~n31329 ;
  assign n31331 = \u1_L12_reg[13]/NET0131  & n31329 ;
  assign n31332 = ~n31330 & ~n31331 ;
  assign n31335 = ~n30512 & n30519 ;
  assign n31336 = ~n30509 & ~n30541 ;
  assign n31337 = n31335 & ~n31336 ;
  assign n31334 = ~n30519 & ~n31106 ;
  assign n31333 = n30496 & n30556 ;
  assign n31338 = ~n30552 & ~n31333 ;
  assign n31339 = ~n31334 & n31338 ;
  assign n31340 = ~n31337 & n31339 ;
  assign n31343 = n30496 & ~n31106 ;
  assign n31341 = ~n30519 & ~n30521 ;
  assign n31342 = ~n31335 & ~n31341 ;
  assign n31344 = ~n30533 & n30552 ;
  assign n31345 = ~n30573 & ~n30952 ;
  assign n31346 = n31344 & n31345 ;
  assign n31347 = ~n31342 & n31346 ;
  assign n31348 = ~n31343 & n31347 ;
  assign n31349 = ~n31340 & ~n31348 ;
  assign n31350 = ~n30561 & ~n30579 ;
  assign n31351 = ~n31349 & n31350 ;
  assign n31352 = ~\u1_L12_reg[19]/NET0131  & ~n31351 ;
  assign n31353 = \u1_L12_reg[19]/NET0131  & n31351 ;
  assign n31354 = ~n31352 & ~n31353 ;
  assign n31373 = ~n30448 & ~n30461 ;
  assign n31374 = ~n30430 & n31373 ;
  assign n31375 = n30403 & ~n31374 ;
  assign n31376 = ~n30429 & n30461 ;
  assign n31377 = ~n30704 & ~n31376 ;
  assign n31378 = ~n31375 & n31377 ;
  assign n31379 = ~n30440 & ~n31378 ;
  assign n31356 = n30440 & ~n30457 ;
  assign n31357 = n30445 & n31356 ;
  assign n31358 = n30403 & ~n30707 ;
  assign n31359 = ~n30468 & n31358 ;
  assign n31360 = ~n31357 & n31359 ;
  assign n31361 = n30429 & n30440 ;
  assign n31362 = n30460 & n31361 ;
  assign n31367 = ~n30703 & ~n31362 ;
  assign n31363 = n30442 & n30447 ;
  assign n31364 = ~n30409 & n30457 ;
  assign n31368 = ~n31363 & ~n31364 ;
  assign n31369 = n31367 & n31368 ;
  assign n31365 = n30440 & n30448 ;
  assign n31366 = ~n30403 & ~n30474 ;
  assign n31370 = ~n31365 & n31366 ;
  assign n31371 = n31369 & n31370 ;
  assign n31372 = ~n31360 & ~n31371 ;
  assign n31380 = n30448 & n30471 ;
  assign n31355 = n30447 & n30459 ;
  assign n31381 = ~n30483 & ~n31355 ;
  assign n31382 = ~n31380 & n31381 ;
  assign n31383 = ~n31372 & n31382 ;
  assign n31384 = ~n31379 & n31383 ;
  assign n31385 = ~\u1_L12_reg[23]/P0001  & n31384 ;
  assign n31386 = \u1_L12_reg[23]/P0001  & ~n31384 ;
  assign n31387 = ~n31385 & ~n31386 ;
  assign n31405 = ~n30802 & ~n30876 ;
  assign n31406 = n30785 & ~n31405 ;
  assign n31407 = ~n30785 & ~n30790 ;
  assign n31408 = ~n30772 & ~n30884 ;
  assign n31409 = n31407 & n31408 ;
  assign n31410 = ~n31406 & ~n31409 ;
  assign n31411 = ~n30805 & ~n30880 ;
  assign n31412 = ~n30898 & n31411 ;
  assign n31413 = ~n31410 & n31412 ;
  assign n31414 = n30816 & ~n31413 ;
  assign n31390 = ~n30800 & ~n30876 ;
  assign n31391 = ~n30817 & n31390 ;
  assign n31392 = n30785 & ~n30801 ;
  assign n31393 = ~n31391 & n31392 ;
  assign n31388 = n30778 & n30803 ;
  assign n31389 = n30793 & n30825 ;
  assign n31394 = ~n30883 & ~n31389 ;
  assign n31395 = ~n31388 & n31394 ;
  assign n31396 = ~n31393 & n31395 ;
  assign n31397 = ~n30816 & ~n31396 ;
  assign n31398 = ~n30770 & n30785 ;
  assign n31399 = n30826 & n31398 ;
  assign n31400 = n30800 & n30876 ;
  assign n31401 = ~n31390 & ~n31400 ;
  assign n31402 = ~n30818 & ~n30881 ;
  assign n31403 = ~n30785 & ~n31402 ;
  assign n31404 = ~n31401 & n31403 ;
  assign n31415 = ~n31399 & ~n31404 ;
  assign n31416 = ~n31397 & n31415 ;
  assign n31417 = ~n31414 & n31416 ;
  assign n31418 = \u1_L12_reg[27]/NET0131  & n31417 ;
  assign n31419 = ~\u1_L12_reg[27]/NET0131  & ~n31417 ;
  assign n31420 = ~n31418 & ~n31419 ;
  assign n31421 = n30305 & ~n30332 ;
  assign n31422 = ~n30317 & n30336 ;
  assign n31423 = ~n30305 & ~n31422 ;
  assign n31424 = ~n30383 & n31423 ;
  assign n31425 = ~n31421 & ~n31424 ;
  assign n31427 = ~n30335 & ~n30723 ;
  assign n31428 = ~n30318 & ~n30369 ;
  assign n31429 = ~n30324 & n31428 ;
  assign n31430 = ~n31427 & ~n31429 ;
  assign n31431 = ~n30305 & ~n30729 ;
  assign n31432 = ~n31430 & n31431 ;
  assign n31434 = n30305 & ~n30361 ;
  assign n31433 = n30331 & n30369 ;
  assign n31435 = ~n30382 & ~n31433 ;
  assign n31436 = n31434 & n31435 ;
  assign n31437 = ~n31432 & ~n31436 ;
  assign n31426 = n30336 & n30369 ;
  assign n31438 = n30354 & ~n31426 ;
  assign n31439 = ~n31437 & n31438 ;
  assign n31442 = n30741 & n31427 ;
  assign n31440 = n30336 & n31428 ;
  assign n31445 = ~n30354 & ~n31440 ;
  assign n31446 = ~n31442 & n31445 ;
  assign n31441 = ~n30370 & n30728 ;
  assign n31443 = ~n30370 & ~n30377 ;
  assign n31444 = n30305 & ~n31443 ;
  assign n31447 = ~n31441 & ~n31444 ;
  assign n31448 = n31446 & n31447 ;
  assign n31449 = ~n31439 & ~n31448 ;
  assign n31450 = ~n31425 & ~n31449 ;
  assign n31451 = \u1_L12_reg[32]/NET0131  & n31450 ;
  assign n31452 = ~\u1_L12_reg[32]/NET0131  & ~n31450 ;
  assign n31453 = ~n31451 & ~n31452 ;
  assign n31491 = decrypt_pad & ~\u1_uk_K_r12_reg[6]/NET0131  ;
  assign n31492 = ~decrypt_pad & ~\u1_uk_K_r12_reg[55]/NET0131  ;
  assign n31493 = ~n31491 & ~n31492 ;
  assign n31494 = \u1_R12_reg[11]/NET0131  & ~n31493 ;
  assign n31495 = ~\u1_R12_reg[11]/NET0131  & n31493 ;
  assign n31496 = ~n31494 & ~n31495 ;
  assign n31480 = decrypt_pad & ~\u1_uk_K_r12_reg[46]/NET0131  ;
  assign n31481 = ~decrypt_pad & ~\u1_uk_K_r12_reg[13]/NET0131  ;
  assign n31482 = ~n31480 & ~n31481 ;
  assign n31483 = \u1_R12_reg[12]/NET0131  & ~n31482 ;
  assign n31484 = ~\u1_R12_reg[12]/NET0131  & n31482 ;
  assign n31485 = ~n31483 & ~n31484 ;
  assign n31460 = decrypt_pad & ~\u1_uk_K_r12_reg[34]/NET0131  ;
  assign n31461 = ~decrypt_pad & ~\u1_uk_K_r12_reg[26]/NET0131  ;
  assign n31462 = ~n31460 & ~n31461 ;
  assign n31463 = \u1_R12_reg[13]/NET0131  & ~n31462 ;
  assign n31464 = ~\u1_R12_reg[13]/NET0131  & n31462 ;
  assign n31465 = ~n31463 & ~n31464 ;
  assign n31467 = decrypt_pad & ~\u1_uk_K_r12_reg[54]/NET0131  ;
  assign n31468 = ~decrypt_pad & ~\u1_uk_K_r12_reg[46]/NET0131  ;
  assign n31469 = ~n31467 & ~n31468 ;
  assign n31470 = \u1_R12_reg[9]/NET0131  & ~n31469 ;
  assign n31471 = ~\u1_R12_reg[9]/NET0131  & n31469 ;
  assign n31472 = ~n31470 & ~n31471 ;
  assign n31514 = n31465 & ~n31472 ;
  assign n31454 = decrypt_pad & ~\u1_uk_K_r12_reg[25]/NET0131  ;
  assign n31455 = ~decrypt_pad & ~\u1_uk_K_r12_reg[17]/NET0131  ;
  assign n31456 = ~n31454 & ~n31455 ;
  assign n31457 = \u1_R12_reg[8]/NET0131  & ~n31456 ;
  assign n31458 = ~\u1_R12_reg[8]/NET0131  & n31456 ;
  assign n31459 = ~n31457 & ~n31458 ;
  assign n31466 = ~n31459 & ~n31465 ;
  assign n31515 = ~n31465 & n31472 ;
  assign n31473 = decrypt_pad & ~\u1_uk_K_r12_reg[5]/NET0131  ;
  assign n31474 = ~decrypt_pad & ~\u1_uk_K_r12_reg[54]/NET0131  ;
  assign n31475 = ~n31473 & ~n31474 ;
  assign n31476 = \u1_R12_reg[10]/NET0131  & ~n31475 ;
  assign n31477 = ~\u1_R12_reg[10]/NET0131  & n31475 ;
  assign n31478 = ~n31476 & ~n31477 ;
  assign n31516 = ~n31459 & n31478 ;
  assign n31517 = ~n31515 & ~n31516 ;
  assign n31518 = ~n31466 & ~n31517 ;
  assign n31519 = ~n31514 & ~n31518 ;
  assign n31520 = n31485 & ~n31519 ;
  assign n31498 = n31465 & n31478 ;
  assign n31521 = ~n31465 & ~n31478 ;
  assign n31522 = ~n31498 & ~n31521 ;
  assign n31523 = ~n31459 & ~n31472 ;
  assign n31524 = ~n31514 & ~n31523 ;
  assign n31525 = ~n31522 & ~n31524 ;
  assign n31526 = ~n31520 & ~n31525 ;
  assign n31527 = n31496 & ~n31526 ;
  assign n31479 = n31472 & n31478 ;
  assign n31502 = ~n31472 & ~n31478 ;
  assign n31503 = n31459 & n31465 ;
  assign n31504 = ~n31466 & ~n31503 ;
  assign n31505 = ~n31502 & ~n31504 ;
  assign n31506 = ~n31479 & n31505 ;
  assign n31490 = ~n31459 & n31472 ;
  assign n31497 = ~n31478 & n31496 ;
  assign n31499 = ~n31496 & n31498 ;
  assign n31500 = ~n31497 & ~n31499 ;
  assign n31501 = n31490 & ~n31500 ;
  assign n31488 = ~n31465 & n31479 ;
  assign n31489 = n31459 & n31488 ;
  assign n31507 = n31465 & n31496 ;
  assign n31508 = n31502 & ~n31507 ;
  assign n31509 = n31504 & n31508 ;
  assign n31510 = ~n31489 & ~n31509 ;
  assign n31511 = ~n31501 & n31510 ;
  assign n31512 = ~n31506 & n31511 ;
  assign n31513 = ~n31485 & ~n31512 ;
  assign n31486 = n31479 & n31485 ;
  assign n31487 = n31466 & n31486 ;
  assign n31528 = n31485 & ~n31496 ;
  assign n31529 = n31517 & n31528 ;
  assign n31530 = n31524 & n31529 ;
  assign n31531 = ~n31487 & ~n31530 ;
  assign n31532 = ~n31513 & n31531 ;
  assign n31533 = ~n31527 & n31532 ;
  assign n31534 = ~\u1_L12_reg[6]/NET0131  & ~n31533 ;
  assign n31535 = \u1_L12_reg[6]/NET0131  & n31533 ;
  assign n31536 = ~n31534 & ~n31535 ;
  assign n31537 = n30324 & ~n31428 ;
  assign n31538 = n30331 & n31537 ;
  assign n31539 = ~n30729 & ~n31538 ;
  assign n31540 = ~n30331 & ~n30341 ;
  assign n31541 = n31428 & n31540 ;
  assign n31542 = n30305 & ~n31541 ;
  assign n31543 = ~n30324 & n30345 ;
  assign n31544 = ~n31433 & ~n31543 ;
  assign n31545 = n31423 & n31544 ;
  assign n31546 = ~n31537 & n31545 ;
  assign n31547 = ~n31542 & ~n31546 ;
  assign n31548 = n31539 & ~n31547 ;
  assign n31549 = n30354 & ~n31548 ;
  assign n31550 = n30331 & ~n30333 ;
  assign n31551 = n31428 & ~n31550 ;
  assign n31552 = ~n30354 & ~n31551 ;
  assign n31553 = ~n31538 & n31552 ;
  assign n31554 = ~n30362 & ~n31553 ;
  assign n31555 = n30305 & ~n31554 ;
  assign n31556 = ~n30305 & ~n31539 ;
  assign n31557 = ~n30305 & n31541 ;
  assign n31558 = ~n30362 & ~n31557 ;
  assign n31559 = ~n30354 & ~n31558 ;
  assign n31560 = ~n31556 & ~n31559 ;
  assign n31561 = ~n31555 & n31560 ;
  assign n31562 = ~n31549 & n31561 ;
  assign n31563 = ~\u1_L12_reg[7]/NET0131  & ~n31562 ;
  assign n31564 = \u1_L12_reg[7]/NET0131  & n31562 ;
  assign n31565 = ~n31563 & ~n31564 ;
  assign n31579 = ~n31195 & n31203 ;
  assign n31581 = ~n31203 & ~n31278 ;
  assign n31580 = ~n31181 & n31260 ;
  assign n31582 = ~n31289 & ~n31580 ;
  assign n31583 = n31581 & n31582 ;
  assign n31584 = ~n31579 & ~n31583 ;
  assign n31585 = n31203 & n31271 ;
  assign n31586 = ~n31216 & ~n31585 ;
  assign n31587 = n31288 & n31586 ;
  assign n31588 = ~n31584 & n31587 ;
  assign n31589 = ~n31227 & ~n31588 ;
  assign n31567 = ~n31174 & n31215 ;
  assign n31568 = ~n31278 & ~n31567 ;
  assign n31569 = n31227 & ~n31568 ;
  assign n31566 = n31189 & n31289 ;
  assign n31570 = n31175 & n31204 ;
  assign n31571 = ~n31197 & ~n31570 ;
  assign n31572 = ~n31566 & n31571 ;
  assign n31573 = ~n31569 & n31572 ;
  assign n31574 = n31203 & ~n31573 ;
  assign n31575 = n31227 & n31247 ;
  assign n31576 = n31206 & n31227 ;
  assign n31577 = ~n31237 & ~n31576 ;
  assign n31578 = ~n31203 & ~n31577 ;
  assign n31590 = ~n31575 & ~n31578 ;
  assign n31591 = ~n31574 & n31590 ;
  assign n31592 = ~n31589 & n31591 ;
  assign n31593 = ~\u1_L12_reg[8]/NET0131  & ~n31592 ;
  assign n31594 = \u1_L12_reg[8]/NET0131  & n31592 ;
  assign n31595 = ~n31593 & ~n31594 ;
  assign n31606 = n31459 & n31472 ;
  assign n31607 = ~n31523 & ~n31606 ;
  assign n31608 = n31465 & ~n31607 ;
  assign n31615 = ~n31496 & n31608 ;
  assign n31616 = n31466 & ~n31478 ;
  assign n31617 = ~n31615 & ~n31616 ;
  assign n31604 = n31472 & n31496 ;
  assign n31618 = ~n31485 & ~n31604 ;
  assign n31619 = ~n31617 & n31618 ;
  assign n31609 = n31466 & n31604 ;
  assign n31603 = n31459 & ~n31465 ;
  assign n31605 = n31603 & ~n31604 ;
  assign n31610 = ~n31478 & ~n31605 ;
  assign n31611 = ~n31609 & n31610 ;
  assign n31612 = ~n31608 & n31611 ;
  assign n31600 = n31465 & n31490 ;
  assign n31599 = n31466 & ~n31496 ;
  assign n31601 = n31478 & ~n31599 ;
  assign n31602 = ~n31600 & n31601 ;
  assign n31613 = n31485 & ~n31602 ;
  assign n31614 = ~n31612 & n31613 ;
  assign n31596 = n31459 & n31478 ;
  assign n31597 = ~n31472 & n31596 ;
  assign n31598 = ~n31496 & n31597 ;
  assign n31620 = ~n31465 & ~n31606 ;
  assign n31621 = ~n31485 & ~n31620 ;
  assign n31622 = n31478 & ~n31607 ;
  assign n31623 = ~n31621 & ~n31622 ;
  assign n31624 = n31496 & ~n31608 ;
  assign n31625 = ~n31623 & n31624 ;
  assign n31626 = ~n31598 & ~n31625 ;
  assign n31627 = ~n31614 & n31626 ;
  assign n31628 = ~n31619 & n31627 ;
  assign n31629 = ~\u1_L12_reg[16]/NET0131  & ~n31628 ;
  assign n31630 = \u1_L12_reg[16]/NET0131  & n31628 ;
  assign n31631 = ~n31629 & ~n31630 ;
  assign n31647 = ~n31459 & n31465 ;
  assign n31648 = n31502 & ~n31647 ;
  assign n31649 = ~n31606 & ~n31647 ;
  assign n31650 = n31478 & ~n31649 ;
  assign n31651 = ~n31648 & ~n31650 ;
  assign n31652 = n31496 & ~n31651 ;
  assign n31653 = ~n31496 & n31505 ;
  assign n31654 = ~n31509 & ~n31653 ;
  assign n31655 = ~n31652 & n31654 ;
  assign n31656 = n31485 & ~n31655 ;
  assign n31632 = ~n31465 & n31597 ;
  assign n31633 = ~n31459 & n31522 ;
  assign n31634 = ~n31515 & ~n31596 ;
  assign n31635 = ~n31633 & n31634 ;
  assign n31636 = n31496 & ~n31606 ;
  assign n31637 = ~n31635 & n31636 ;
  assign n31638 = ~n31632 & ~n31637 ;
  assign n31639 = ~n31485 & ~n31638 ;
  assign n31641 = n31502 & ~n31504 ;
  assign n31642 = ~n31518 & ~n31641 ;
  assign n31643 = ~n31485 & ~n31496 ;
  assign n31644 = ~n31642 & n31643 ;
  assign n31640 = n31499 & n31606 ;
  assign n31645 = n31497 & n31504 ;
  assign n31646 = n31607 & n31645 ;
  assign n31657 = ~n31640 & ~n31646 ;
  assign n31658 = ~n31644 & n31657 ;
  assign n31659 = ~n31639 & n31658 ;
  assign n31660 = ~n31656 & n31659 ;
  assign n31661 = ~\u1_L12_reg[24]/NET0131  & ~n31660 ;
  assign n31662 = \u1_L12_reg[24]/NET0131  & n31660 ;
  assign n31663 = ~n31661 & ~n31662 ;
  assign n31674 = ~n31488 & ~n31634 ;
  assign n31675 = ~n31485 & ~n31674 ;
  assign n31671 = n31502 & n31603 ;
  assign n31672 = n31485 & ~n31671 ;
  assign n31673 = ~n31633 & n31672 ;
  assign n31676 = n31496 & ~n31673 ;
  assign n31677 = ~n31675 & n31676 ;
  assign n31666 = ~n31496 & ~n31523 ;
  assign n31667 = n31634 & n31666 ;
  assign n31665 = n31498 & n31523 ;
  assign n31668 = ~n31641 & ~n31665 ;
  assign n31669 = ~n31667 & n31668 ;
  assign n31670 = ~n31485 & ~n31669 ;
  assign n31678 = n31466 & n31472 ;
  assign n31679 = ~n31596 & ~n31678 ;
  assign n31680 = n31528 & ~n31679 ;
  assign n31682 = n31507 & n31597 ;
  assign n31664 = n31488 & ~n31496 ;
  assign n31681 = n31486 & ~n31503 ;
  assign n31683 = ~n31664 & ~n31681 ;
  assign n31684 = ~n31682 & n31683 ;
  assign n31685 = ~n31680 & n31684 ;
  assign n31686 = ~n31670 & n31685 ;
  assign n31687 = ~n31677 & n31686 ;
  assign n31688 = \u1_L12_reg[30]/NET0131  & ~n31687 ;
  assign n31689 = ~\u1_L12_reg[30]/NET0131  & n31687 ;
  assign n31690 = ~n31688 & ~n31689 ;
  assign n31692 = ~n30431 & ~n30448 ;
  assign n31693 = ~n30685 & n31692 ;
  assign n31694 = n30440 & ~n31693 ;
  assign n31695 = ~n30416 & ~n30698 ;
  assign n31696 = ~n30440 & ~n31695 ;
  assign n31691 = n30429 & n30687 ;
  assign n31697 = ~n30429 & n30459 ;
  assign n31698 = ~n31691 & ~n31697 ;
  assign n31699 = ~n31696 & n31698 ;
  assign n31700 = ~n31694 & n31699 ;
  assign n31701 = ~n30403 & ~n31700 ;
  assign n31702 = n30429 & n30698 ;
  assign n31703 = ~n31697 & ~n31702 ;
  assign n31704 = ~n30440 & ~n31703 ;
  assign n31705 = n30446 & ~n30687 ;
  assign n31706 = n30471 & ~n31695 ;
  assign n31707 = ~n30704 & ~n31706 ;
  assign n31708 = ~n31705 & n31707 ;
  assign n31709 = n30403 & ~n31708 ;
  assign n31710 = ~n31704 & ~n31709 ;
  assign n31711 = ~n31701 & n31710 ;
  assign n31712 = ~\u1_L12_reg[9]/NET0131  & ~n31711 ;
  assign n31713 = \u1_L12_reg[9]/NET0131  & n31711 ;
  assign n31714 = ~n31712 & ~n31713 ;
  assign n31715 = n31227 & ~n31237 ;
  assign n31716 = ~n31213 & n31260 ;
  assign n31717 = n31715 & ~n31716 ;
  assign n31718 = n31174 & ~n31261 ;
  assign n31719 = ~n31227 & ~n31718 ;
  assign n31720 = n31183 & ~n31278 ;
  assign n31721 = n31719 & n31720 ;
  assign n31722 = ~n31717 & ~n31721 ;
  assign n31723 = ~n31189 & ~n31246 ;
  assign n31724 = ~n31183 & n31723 ;
  assign n31725 = ~n31203 & ~n31250 ;
  assign n31726 = ~n31724 & n31725 ;
  assign n31727 = ~n31722 & n31726 ;
  assign n31728 = ~n31181 & n31196 ;
  assign n31729 = ~n31207 & ~n31728 ;
  assign n31730 = n31715 & n31729 ;
  assign n31731 = ~n31229 & ~n31289 ;
  assign n31732 = n31719 & n31731 ;
  assign n31733 = ~n31730 & ~n31732 ;
  assign n31734 = ~n31570 & n31579 ;
  assign n31735 = ~n31733 & n31734 ;
  assign n31736 = ~n31727 & ~n31735 ;
  assign n31737 = ~\u1_L12_reg[3]/NET0131  & n31736 ;
  assign n31738 = \u1_L12_reg[3]/NET0131  & ~n31736 ;
  assign n31739 = ~n31737 & ~n31738 ;
  assign n31743 = n31014 & ~n31018 ;
  assign n31741 = ~n31042 & ~n31320 ;
  assign n31742 = ~n31014 & ~n31741 ;
  assign n31744 = ~n31059 & ~n31742 ;
  assign n31745 = ~n31743 & n31744 ;
  assign n31746 = n31025 & ~n31745 ;
  assign n31750 = ~n31077 & ~n31301 ;
  assign n31751 = ~n31028 & n31750 ;
  assign n31747 = n31014 & n31043 ;
  assign n31748 = n30998 & ~n31015 ;
  assign n31749 = n31053 & ~n31748 ;
  assign n31752 = ~n31747 & ~n31749 ;
  assign n31753 = n31751 & n31752 ;
  assign n31754 = ~n31025 & ~n31753 ;
  assign n31740 = ~n31014 & n31073 ;
  assign n31755 = ~n31027 & ~n31315 ;
  assign n31756 = n31014 & ~n31755 ;
  assign n31757 = ~n31740 & ~n31756 ;
  assign n31758 = ~n31754 & n31757 ;
  assign n31759 = ~n31746 & n31758 ;
  assign n31760 = ~\u1_L12_reg[18]/P0001  & ~n31759 ;
  assign n31761 = \u1_L12_reg[18]/P0001  & n31759 ;
  assign n31762 = ~n31760 & ~n31761 ;
  assign n31763 = decrypt_pad & ~\u1_uk_K_r11_reg[18]/NET0131  ;
  assign n31764 = ~decrypt_pad & ~\u1_uk_K_r11_reg[13]/NET0131  ;
  assign n31765 = ~n31763 & ~n31764 ;
  assign n31766 = \u1_R11_reg[3]/NET0131  & ~n31765 ;
  assign n31767 = ~\u1_R11_reg[3]/NET0131  & n31765 ;
  assign n31768 = ~n31766 & ~n31767 ;
  assign n31769 = decrypt_pad & ~\u1_uk_K_r11_reg[26]/NET0131  ;
  assign n31770 = ~decrypt_pad & ~\u1_uk_K_r11_reg[46]/NET0131  ;
  assign n31771 = ~n31769 & ~n31770 ;
  assign n31772 = \u1_R11_reg[1]/NET0131  & ~n31771 ;
  assign n31773 = ~\u1_R11_reg[1]/NET0131  & n31771 ;
  assign n31774 = ~n31772 & ~n31773 ;
  assign n31783 = decrypt_pad & ~\u1_uk_K_r11_reg[24]/NET0131  ;
  assign n31784 = ~decrypt_pad & ~\u1_uk_K_r11_reg[19]/NET0131  ;
  assign n31785 = ~n31783 & ~n31784 ;
  assign n31786 = \u1_R11_reg[5]/NET0131  & ~n31785 ;
  assign n31787 = ~\u1_R11_reg[5]/NET0131  & n31785 ;
  assign n31788 = ~n31786 & ~n31787 ;
  assign n31803 = ~n31774 & n31788 ;
  assign n31776 = decrypt_pad & ~\u1_uk_K_r11_reg[41]/NET0131  ;
  assign n31777 = ~decrypt_pad & ~\u1_uk_K_r11_reg[4]/NET0131  ;
  assign n31778 = ~n31776 & ~n31777 ;
  assign n31779 = \u1_R11_reg[2]/NET0131  & ~n31778 ;
  assign n31780 = ~\u1_R11_reg[2]/NET0131  & n31778 ;
  assign n31781 = ~n31779 & ~n31780 ;
  assign n31791 = decrypt_pad & ~\u1_uk_K_r11_reg[5]/NET0131  ;
  assign n31792 = ~decrypt_pad & ~\u1_uk_K_r11_reg[25]/NET0131  ;
  assign n31793 = ~n31791 & ~n31792 ;
  assign n31794 = \u1_R11_reg[32]/NET0131  & ~n31793 ;
  assign n31795 = ~\u1_R11_reg[32]/NET0131  & n31793 ;
  assign n31796 = ~n31794 & ~n31795 ;
  assign n31804 = ~n31788 & ~n31796 ;
  assign n31805 = n31781 & n31804 ;
  assign n31806 = ~n31803 & ~n31805 ;
  assign n31807 = n31768 & ~n31806 ;
  assign n31775 = ~n31768 & n31774 ;
  assign n31782 = ~n31774 & ~n31781 ;
  assign n31789 = n31782 & ~n31788 ;
  assign n31790 = ~n31775 & ~n31789 ;
  assign n31797 = ~n31790 & n31796 ;
  assign n31798 = n31768 & ~n31781 ;
  assign n31799 = n31774 & ~n31798 ;
  assign n31800 = ~n31781 & ~n31788 ;
  assign n31801 = ~n31796 & ~n31800 ;
  assign n31802 = ~n31799 & n31801 ;
  assign n31808 = decrypt_pad & ~\u1_uk_K_r11_reg[53]/P0001  ;
  assign n31809 = ~decrypt_pad & ~\u1_uk_K_r11_reg[48]/NET0131  ;
  assign n31810 = ~n31808 & ~n31809 ;
  assign n31811 = \u1_R11_reg[4]/NET0131  & ~n31810 ;
  assign n31812 = ~\u1_R11_reg[4]/NET0131  & n31810 ;
  assign n31813 = ~n31811 & ~n31812 ;
  assign n31814 = ~n31802 & n31813 ;
  assign n31815 = ~n31797 & n31814 ;
  assign n31816 = ~n31807 & n31815 ;
  assign n31820 = n31768 & ~n31796 ;
  assign n31821 = n31781 & n31820 ;
  assign n31822 = n31788 & n31821 ;
  assign n31823 = ~n31796 & n31800 ;
  assign n31824 = ~n31822 & ~n31823 ;
  assign n31825 = n31774 & ~n31824 ;
  assign n31828 = ~n31781 & n31796 ;
  assign n31829 = ~n31768 & ~n31828 ;
  assign n31826 = ~n31774 & n31796 ;
  assign n31827 = n31781 & ~n31826 ;
  assign n31830 = ~n31803 & ~n31827 ;
  assign n31831 = n31829 & n31830 ;
  assign n31832 = n31768 & n31796 ;
  assign n31833 = n31774 & ~n31788 ;
  assign n31834 = n31781 & n31833 ;
  assign n31835 = n31832 & n31834 ;
  assign n31817 = n31788 & n31796 ;
  assign n31818 = ~n31775 & ~n31781 ;
  assign n31819 = n31817 & n31818 ;
  assign n31836 = ~n31813 & ~n31819 ;
  assign n31837 = ~n31835 & n31836 ;
  assign n31838 = ~n31831 & n31837 ;
  assign n31839 = ~n31825 & n31838 ;
  assign n31840 = ~n31816 & ~n31839 ;
  assign n31843 = n31774 & n31788 ;
  assign n31844 = n31781 & n31843 ;
  assign n31845 = n31796 & n31844 ;
  assign n31846 = ~n31774 & n31781 ;
  assign n31847 = ~n31800 & ~n31846 ;
  assign n31841 = ~n31774 & ~n31788 ;
  assign n31848 = ~n31826 & ~n31841 ;
  assign n31849 = ~n31847 & n31848 ;
  assign n31850 = ~n31845 & ~n31849 ;
  assign n31851 = ~n31768 & ~n31850 ;
  assign n31842 = n31821 & n31841 ;
  assign n31852 = n31798 & n31826 ;
  assign n31853 = ~n31842 & ~n31852 ;
  assign n31854 = ~n31851 & n31853 ;
  assign n31855 = ~n31840 & n31854 ;
  assign n31856 = ~\u1_L11_reg[31]/NET0131  & ~n31855 ;
  assign n31857 = \u1_L11_reg[31]/NET0131  & n31855 ;
  assign n31858 = ~n31856 & ~n31857 ;
  assign n31913 = decrypt_pad & ~\u1_uk_K_r11_reg[52]/NET0131  ;
  assign n31914 = ~decrypt_pad & ~\u1_uk_K_r11_reg[15]/NET0131  ;
  assign n31915 = ~n31913 & ~n31914 ;
  assign n31916 = \u1_R11_reg[24]/NET0131  & ~n31915 ;
  assign n31917 = ~\u1_R11_reg[24]/NET0131  & n31915 ;
  assign n31918 = ~n31916 & ~n31917 ;
  assign n31882 = decrypt_pad & ~\u1_uk_K_r11_reg[22]/NET0131  ;
  assign n31883 = ~decrypt_pad & ~\u1_uk_K_r11_reg[44]/NET0131  ;
  assign n31884 = ~n31882 & ~n31883 ;
  assign n31885 = \u1_R11_reg[23]/NET0131  & ~n31884 ;
  assign n31886 = ~\u1_R11_reg[23]/NET0131  & n31884 ;
  assign n31887 = ~n31885 & ~n31886 ;
  assign n31859 = decrypt_pad & ~\u1_uk_K_r11_reg[42]/NET0131  ;
  assign n31860 = ~decrypt_pad & ~\u1_uk_K_r11_reg[9]/NET0131  ;
  assign n31861 = ~n31859 & ~n31860 ;
  assign n31862 = \u1_R11_reg[21]/NET0131  & ~n31861 ;
  assign n31863 = ~\u1_R11_reg[21]/NET0131  & n31861 ;
  assign n31864 = ~n31862 & ~n31863 ;
  assign n31865 = decrypt_pad & ~\u1_uk_K_r11_reg[31]/NET0131  ;
  assign n31866 = ~decrypt_pad & ~\u1_uk_K_r11_reg[49]/NET0131  ;
  assign n31867 = ~n31865 & ~n31866 ;
  assign n31868 = \u1_R11_reg[20]/NET0131  & ~n31867 ;
  assign n31869 = ~\u1_R11_reg[20]/NET0131  & n31867 ;
  assign n31870 = ~n31868 & ~n31869 ;
  assign n31871 = n31864 & ~n31870 ;
  assign n31872 = decrypt_pad & ~\u1_uk_K_r11_reg[9]/NET0131  ;
  assign n31873 = ~decrypt_pad & ~\u1_uk_K_r11_reg[0]/NET0131  ;
  assign n31874 = ~n31872 & ~n31873 ;
  assign n31875 = \u1_R11_reg[22]/NET0131  & ~n31874 ;
  assign n31876 = ~\u1_R11_reg[22]/NET0131  & n31874 ;
  assign n31877 = ~n31875 & ~n31876 ;
  assign n31878 = n31871 & n31877 ;
  assign n31890 = decrypt_pad & ~\u1_uk_K_r11_reg[43]/NET0131  ;
  assign n31891 = ~decrypt_pad & ~\u1_uk_K_r11_reg[38]/NET0131  ;
  assign n31892 = ~n31890 & ~n31891 ;
  assign n31893 = \u1_R11_reg[25]/NET0131  & ~n31892 ;
  assign n31894 = ~\u1_R11_reg[25]/NET0131  & n31892 ;
  assign n31895 = ~n31893 & ~n31894 ;
  assign n31938 = n31864 & ~n31895 ;
  assign n31939 = n31870 & ~n31938 ;
  assign n31896 = ~n31877 & ~n31895 ;
  assign n31940 = ~n31864 & ~n31896 ;
  assign n31941 = n31939 & ~n31940 ;
  assign n31942 = ~n31878 & ~n31941 ;
  assign n31943 = n31887 & ~n31942 ;
  assign n31901 = n31870 & n31895 ;
  assign n31934 = ~n31871 & ~n31901 ;
  assign n31935 = n31877 & ~n31934 ;
  assign n31906 = ~n31870 & n31895 ;
  assign n31932 = n31864 & n31906 ;
  assign n31933 = ~n31877 & ~n31932 ;
  assign n31936 = ~n31887 & ~n31933 ;
  assign n31937 = ~n31935 & n31936 ;
  assign n31928 = ~n31877 & ~n31887 ;
  assign n31944 = n31901 & n31928 ;
  assign n31945 = ~n31864 & n31944 ;
  assign n31946 = ~n31937 & ~n31945 ;
  assign n31947 = ~n31943 & n31946 ;
  assign n31948 = n31918 & ~n31947 ;
  assign n31879 = n31864 & n31870 ;
  assign n31880 = ~n31877 & n31879 ;
  assign n31881 = ~n31878 & ~n31880 ;
  assign n31888 = ~n31881 & ~n31887 ;
  assign n31897 = ~n31864 & n31887 ;
  assign n31907 = n31897 & n31906 ;
  assign n31904 = n31879 & n31896 ;
  assign n31889 = ~n31877 & n31887 ;
  assign n31905 = ~n31870 & n31889 ;
  assign n31908 = ~n31904 & ~n31905 ;
  assign n31909 = ~n31907 & n31908 ;
  assign n31898 = ~n31896 & ~n31897 ;
  assign n31899 = n31870 & ~n31889 ;
  assign n31900 = ~n31898 & n31899 ;
  assign n31902 = n31877 & n31901 ;
  assign n31903 = ~n31864 & n31902 ;
  assign n31910 = ~n31900 & ~n31903 ;
  assign n31911 = n31909 & n31910 ;
  assign n31912 = ~n31888 & n31911 ;
  assign n31919 = ~n31912 & ~n31918 ;
  assign n31924 = n31879 & ~n31895 ;
  assign n31925 = ~n31887 & n31924 ;
  assign n31926 = ~n31907 & ~n31925 ;
  assign n31927 = ~n31877 & ~n31926 ;
  assign n31920 = n31871 & ~n31895 ;
  assign n31921 = ~n31877 & n31920 ;
  assign n31922 = ~n31902 & ~n31921 ;
  assign n31923 = n31887 & ~n31922 ;
  assign n31929 = ~n31870 & ~n31895 ;
  assign n31930 = n31928 & n31929 ;
  assign n31931 = ~n31864 & n31930 ;
  assign n31949 = ~n31923 & ~n31931 ;
  assign n31950 = ~n31927 & n31949 ;
  assign n31951 = ~n31919 & n31950 ;
  assign n31952 = ~n31948 & n31951 ;
  assign n31953 = \u1_L11_reg[11]/NET0131  & ~n31952 ;
  assign n31954 = ~\u1_L11_reg[11]/NET0131  & n31952 ;
  assign n31955 = ~n31953 & ~n31954 ;
  assign n31971 = decrypt_pad & ~\u1_uk_K_r11_reg[44]/NET0131  ;
  assign n31972 = ~decrypt_pad & ~\u1_uk_K_r11_reg[35]/NET0131  ;
  assign n31973 = ~n31971 & ~n31972 ;
  assign n31974 = \u1_R11_reg[27]/NET0131  & ~n31973 ;
  assign n31975 = ~\u1_R11_reg[27]/NET0131  & n31973 ;
  assign n31976 = ~n31974 & ~n31975 ;
  assign n31956 = decrypt_pad & ~\u1_uk_K_r11_reg[15]/NET0131  ;
  assign n31957 = ~decrypt_pad & ~\u1_uk_K_r11_reg[37]/NET0131  ;
  assign n31958 = ~n31956 & ~n31957 ;
  assign n31959 = \u1_R11_reg[24]/NET0131  & ~n31958 ;
  assign n31960 = ~\u1_R11_reg[24]/NET0131  & n31958 ;
  assign n31961 = ~n31959 & ~n31960 ;
  assign n31977 = decrypt_pad & ~\u1_uk_K_r11_reg[50]/NET0131  ;
  assign n31978 = ~decrypt_pad & ~\u1_uk_K_r11_reg[45]/NET0131  ;
  assign n31979 = ~n31977 & ~n31978 ;
  assign n31980 = \u1_R11_reg[25]/NET0131  & ~n31979 ;
  assign n31981 = ~\u1_R11_reg[25]/NET0131  & n31979 ;
  assign n31982 = ~n31980 & ~n31981 ;
  assign n32003 = n31961 & n31982 ;
  assign n31962 = decrypt_pad & ~\u1_uk_K_r11_reg[35]/NET0131  ;
  assign n31963 = ~decrypt_pad & ~\u1_uk_K_r11_reg[2]/NET0131  ;
  assign n31964 = ~n31962 & ~n31963 ;
  assign n31965 = \u1_R11_reg[26]/NET0131  & ~n31964 ;
  assign n31966 = ~\u1_R11_reg[26]/NET0131  & n31964 ;
  assign n31967 = ~n31965 & ~n31966 ;
  assign n31985 = decrypt_pad & ~\u1_uk_K_r11_reg[23]/NET0131  ;
  assign n31986 = ~decrypt_pad & ~\u1_uk_K_r11_reg[14]/NET0131  ;
  assign n31987 = ~n31985 & ~n31986 ;
  assign n31988 = \u1_R11_reg[29]/NET0131  & ~n31987 ;
  assign n31989 = ~\u1_R11_reg[29]/NET0131  & n31987 ;
  assign n31990 = ~n31988 & ~n31989 ;
  assign n32004 = ~n31967 & n31990 ;
  assign n32005 = n32003 & n32004 ;
  assign n31994 = n31967 & ~n31982 ;
  assign n32006 = n31961 & n31994 ;
  assign n32007 = ~n32005 & ~n32006 ;
  assign n32008 = n31976 & ~n32007 ;
  assign n32017 = ~n31961 & ~n31982 ;
  assign n32018 = ~n32003 & ~n32017 ;
  assign n32019 = ~n31976 & n31990 ;
  assign n32020 = ~n31994 & n32019 ;
  assign n32021 = n32018 & n32020 ;
  assign n31997 = ~n31961 & ~n31990 ;
  assign n32015 = ~n31967 & ~n31982 ;
  assign n32016 = n31997 & n32015 ;
  assign n31995 = ~n31961 & n31990 ;
  assign n31996 = n31994 & n31995 ;
  assign n32009 = decrypt_pad & ~\u1_uk_K_r11_reg[0]/NET0131  ;
  assign n32010 = ~decrypt_pad & ~\u1_uk_K_r11_reg[22]/NET0131  ;
  assign n32011 = ~n32009 & ~n32010 ;
  assign n32012 = \u1_R11_reg[28]/NET0131  & ~n32011 ;
  assign n32013 = ~\u1_R11_reg[28]/NET0131  & n32011 ;
  assign n32014 = ~n32012 & ~n32013 ;
  assign n32022 = ~n31996 & n32014 ;
  assign n32023 = ~n32016 & n32022 ;
  assign n32024 = ~n32021 & n32023 ;
  assign n32025 = ~n32008 & n32024 ;
  assign n31968 = ~n31961 & ~n31967 ;
  assign n31969 = n31961 & n31967 ;
  assign n31970 = ~n31968 & ~n31969 ;
  assign n32026 = n31976 & ~n31982 ;
  assign n32027 = n31990 & ~n32026 ;
  assign n32028 = ~n31970 & n32027 ;
  assign n32034 = ~n32014 & ~n32028 ;
  assign n32029 = n31994 & n31997 ;
  assign n32030 = ~n31976 & n32029 ;
  assign n31983 = ~n31976 & n31982 ;
  assign n32031 = ~n31983 & ~n32015 ;
  assign n32032 = n31961 & ~n32019 ;
  assign n32033 = ~n32031 & n32032 ;
  assign n32035 = ~n32030 & ~n32033 ;
  assign n32036 = n32034 & n32035 ;
  assign n32037 = ~n32025 & ~n32036 ;
  assign n31984 = ~n31970 & n31983 ;
  assign n31991 = ~n31982 & ~n31990 ;
  assign n31992 = ~n31961 & n31967 ;
  assign n31993 = n31991 & ~n31992 ;
  assign n31998 = n31967 & n31982 ;
  assign n31999 = n31997 & n31998 ;
  assign n32000 = ~n31996 & ~n31999 ;
  assign n32001 = ~n31993 & n32000 ;
  assign n32002 = n31976 & ~n32001 ;
  assign n32038 = ~n31984 & ~n32002 ;
  assign n32039 = ~n32037 & n32038 ;
  assign n32040 = \u1_L11_reg[22]/NET0131  & n32039 ;
  assign n32041 = ~\u1_L11_reg[22]/NET0131  & ~n32039 ;
  assign n32042 = ~n32040 & ~n32041 ;
  assign n32055 = decrypt_pad & ~\u1_uk_K_r11_reg[13]/NET0131  ;
  assign n32056 = ~decrypt_pad & ~\u1_uk_K_r11_reg[33]/NET0131  ;
  assign n32057 = ~n32055 & ~n32056 ;
  assign n32058 = \u1_R11_reg[13]/NET0131  & ~n32057 ;
  assign n32059 = ~\u1_R11_reg[13]/NET0131  & n32057 ;
  assign n32060 = ~n32058 & ~n32059 ;
  assign n32049 = decrypt_pad & ~\u1_uk_K_r11_reg[19]/NET0131  ;
  assign n32050 = ~decrypt_pad & ~\u1_uk_K_r11_reg[39]/NET0131  ;
  assign n32051 = ~n32049 & ~n32050 ;
  assign n32052 = \u1_R11_reg[12]/NET0131  & ~n32051 ;
  assign n32053 = ~\u1_R11_reg[12]/NET0131  & n32051 ;
  assign n32054 = ~n32052 & ~n32053 ;
  assign n32068 = decrypt_pad & ~\u1_uk_K_r11_reg[3]/NET0131  ;
  assign n32069 = ~decrypt_pad & ~\u1_uk_K_r11_reg[55]/NET0131  ;
  assign n32070 = ~n32068 & ~n32069 ;
  assign n32071 = \u1_R11_reg[17]/NET0131  & ~n32070 ;
  assign n32072 = ~\u1_R11_reg[17]/NET0131  & n32070 ;
  assign n32073 = ~n32071 & ~n32072 ;
  assign n32100 = n32054 & n32073 ;
  assign n32101 = n32060 & n32100 ;
  assign n32043 = decrypt_pad & ~\u1_uk_K_r11_reg[47]/NET0131  ;
  assign n32044 = ~decrypt_pad & ~\u1_uk_K_r11_reg[10]/NET0131  ;
  assign n32045 = ~n32043 & ~n32044 ;
  assign n32046 = \u1_R11_reg[15]/NET0131  & ~n32045 ;
  assign n32047 = ~\u1_R11_reg[15]/NET0131  & n32045 ;
  assign n32048 = ~n32046 & ~n32047 ;
  assign n32098 = ~n32060 & ~n32073 ;
  assign n32099 = ~n32054 & n32098 ;
  assign n32102 = n32048 & ~n32099 ;
  assign n32103 = ~n32101 & n32102 ;
  assign n32062 = decrypt_pad & ~\u1_uk_K_r11_reg[39]/NET0131  ;
  assign n32063 = ~decrypt_pad & ~\u1_uk_K_r11_reg[34]/NET0131  ;
  assign n32064 = ~n32062 & ~n32063 ;
  assign n32065 = \u1_R11_reg[14]/NET0131  & ~n32064 ;
  assign n32066 = ~\u1_R11_reg[14]/NET0131  & n32064 ;
  assign n32067 = ~n32065 & ~n32066 ;
  assign n32080 = n32054 & ~n32073 ;
  assign n32104 = n32067 & n32080 ;
  assign n32105 = ~n32060 & n32073 ;
  assign n32106 = ~n32048 & ~n32105 ;
  assign n32107 = ~n32104 & n32106 ;
  assign n32108 = ~n32103 & ~n32107 ;
  assign n32077 = ~n32067 & ~n32073 ;
  assign n32078 = ~n32054 & n32077 ;
  assign n32079 = ~n32060 & n32078 ;
  assign n32061 = ~n32054 & n32060 ;
  assign n32089 = n32061 & ~n32073 ;
  assign n32090 = n32067 & n32089 ;
  assign n32091 = ~n32079 & ~n32090 ;
  assign n32111 = n32054 & ~n32067 ;
  assign n32112 = ~n32060 & n32111 ;
  assign n32113 = n32073 & n32112 ;
  assign n32092 = decrypt_pad & ~\u1_uk_K_r11_reg[55]/NET0131  ;
  assign n32093 = ~decrypt_pad & ~\u1_uk_K_r11_reg[18]/NET0131  ;
  assign n32094 = ~n32092 & ~n32093 ;
  assign n32095 = \u1_R11_reg[16]/NET0131  & ~n32094 ;
  assign n32096 = ~\u1_R11_reg[16]/NET0131  & n32094 ;
  assign n32097 = ~n32095 & ~n32096 ;
  assign n32086 = n32048 & n32060 ;
  assign n32109 = n32067 & n32086 ;
  assign n32110 = ~n32054 & n32109 ;
  assign n32114 = ~n32097 & ~n32110 ;
  assign n32115 = ~n32113 & n32114 ;
  assign n32116 = n32091 & n32115 ;
  assign n32117 = ~n32108 & n32116 ;
  assign n32118 = ~n32048 & n32099 ;
  assign n32119 = ~n32101 & ~n32118 ;
  assign n32120 = n32067 & ~n32119 ;
  assign n32121 = ~n32048 & ~n32067 ;
  assign n32122 = n32054 & ~n32060 ;
  assign n32123 = ~n32061 & ~n32122 ;
  assign n32124 = n32121 & ~n32123 ;
  assign n32129 = n32097 & ~n32124 ;
  assign n32074 = ~n32067 & n32073 ;
  assign n32075 = n32061 & n32074 ;
  assign n32087 = n32080 & n32086 ;
  assign n32125 = ~n32075 & ~n32087 ;
  assign n32126 = ~n32054 & n32073 ;
  assign n32127 = n32048 & n32126 ;
  assign n32128 = ~n32060 & n32127 ;
  assign n32130 = n32125 & ~n32128 ;
  assign n32131 = n32129 & n32130 ;
  assign n32132 = ~n32120 & n32131 ;
  assign n32133 = ~n32117 & ~n32132 ;
  assign n32076 = ~n32048 & ~n32075 ;
  assign n32081 = ~n32060 & n32067 ;
  assign n32082 = n32080 & n32081 ;
  assign n32083 = n32048 & ~n32082 ;
  assign n32084 = ~n32079 & n32083 ;
  assign n32085 = ~n32076 & ~n32084 ;
  assign n32088 = ~n32067 & n32087 ;
  assign n32134 = ~n32085 & ~n32088 ;
  assign n32135 = ~n32133 & n32134 ;
  assign n32136 = ~\u1_L11_reg[20]/NET0131  & ~n32135 ;
  assign n32137 = \u1_L11_reg[20]/NET0131  & n32135 ;
  assign n32138 = ~n32136 & ~n32137 ;
  assign n32144 = ~n31864 & n31895 ;
  assign n32145 = n31939 & ~n32144 ;
  assign n32146 = ~n31864 & ~n31877 ;
  assign n32147 = ~n31878 & ~n32146 ;
  assign n32148 = ~n31895 & ~n32147 ;
  assign n32149 = ~n32145 & ~n32148 ;
  assign n32150 = n31887 & ~n32149 ;
  assign n32139 = ~n31877 & ~n31934 ;
  assign n32140 = n31877 & ~n31895 ;
  assign n32141 = n31879 & n32140 ;
  assign n32142 = ~n32139 & ~n32141 ;
  assign n32143 = ~n31887 & ~n32142 ;
  assign n32151 = ~n31870 & n32144 ;
  assign n32152 = n31877 & n32151 ;
  assign n32153 = ~n32143 & ~n32152 ;
  assign n32154 = ~n32150 & n32153 ;
  assign n32155 = ~n31918 & ~n32154 ;
  assign n32160 = n31871 & ~n32140 ;
  assign n32161 = ~n32141 & ~n32160 ;
  assign n32162 = n31887 & ~n32161 ;
  assign n32164 = n31877 & ~n31901 ;
  assign n32165 = ~n31929 & n32164 ;
  assign n32163 = n31887 & ~n31940 ;
  assign n32166 = ~n32139 & ~n32163 ;
  assign n32167 = ~n32165 & n32166 ;
  assign n32168 = ~n32162 & ~n32167 ;
  assign n32169 = n31918 & ~n32168 ;
  assign n32156 = ~n31864 & n31870 ;
  assign n32157 = n31896 & n32156 ;
  assign n32158 = n31864 & n31895 ;
  assign n32159 = n31889 & n32158 ;
  assign n32170 = ~n32157 & ~n32159 ;
  assign n32171 = ~n32169 & n32170 ;
  assign n32172 = ~n32155 & n32171 ;
  assign n32173 = \u1_L11_reg[29]/NET0131  & ~n32172 ;
  assign n32174 = ~\u1_L11_reg[29]/NET0131  & n32172 ;
  assign n32175 = ~n32173 & ~n32174 ;
  assign n32176 = decrypt_pad & ~\u1_uk_K_r11_reg[51]/NET0131  ;
  assign n32177 = ~decrypt_pad & ~\u1_uk_K_r11_reg[42]/NET0131  ;
  assign n32178 = ~n32176 & ~n32177 ;
  assign n32179 = \u1_R11_reg[32]/NET0131  & ~n32178 ;
  assign n32180 = ~\u1_R11_reg[32]/NET0131  & n32178 ;
  assign n32181 = ~n32179 & ~n32180 ;
  assign n32202 = decrypt_pad & ~\u1_uk_K_r11_reg[1]/NET0131  ;
  assign n32203 = ~decrypt_pad & ~\u1_uk_K_r11_reg[23]/NET0131  ;
  assign n32204 = ~n32202 & ~n32203 ;
  assign n32205 = \u1_R11_reg[29]/NET0131  & ~n32204 ;
  assign n32206 = ~\u1_R11_reg[29]/NET0131  & n32204 ;
  assign n32207 = ~n32205 & ~n32206 ;
  assign n32188 = decrypt_pad & ~\u1_uk_K_r11_reg[45]/NET0131  ;
  assign n32189 = ~decrypt_pad & ~\u1_uk_K_r11_reg[8]/NET0131  ;
  assign n32190 = ~n32188 & ~n32189 ;
  assign n32191 = \u1_R11_reg[1]/NET0131  & ~n32190 ;
  assign n32192 = ~\u1_R11_reg[1]/NET0131  & n32190 ;
  assign n32193 = ~n32191 & ~n32192 ;
  assign n32182 = decrypt_pad & ~\u1_uk_K_r11_reg[29]/NET0131  ;
  assign n32183 = ~decrypt_pad & ~\u1_uk_K_r11_reg[51]/NET0131  ;
  assign n32184 = ~n32182 & ~n32183 ;
  assign n32185 = \u1_R11_reg[28]/NET0131  & ~n32184 ;
  assign n32186 = ~\u1_R11_reg[28]/NET0131  & n32184 ;
  assign n32187 = ~n32185 & ~n32186 ;
  assign n32195 = decrypt_pad & ~\u1_uk_K_r11_reg[2]/NET0131  ;
  assign n32196 = ~decrypt_pad & ~\u1_uk_K_r11_reg[52]/NET0131  ;
  assign n32197 = ~n32195 & ~n32196 ;
  assign n32198 = \u1_R11_reg[30]/NET0131  & ~n32197 ;
  assign n32199 = ~\u1_R11_reg[30]/NET0131  & n32197 ;
  assign n32200 = ~n32198 & ~n32199 ;
  assign n32225 = n32187 & ~n32200 ;
  assign n32230 = ~n32193 & n32225 ;
  assign n32231 = n32207 & n32230 ;
  assign n32209 = decrypt_pad & ~\u1_uk_K_r11_reg[14]/NET0131  ;
  assign n32210 = ~decrypt_pad & ~\u1_uk_K_r11_reg[36]/NET0131  ;
  assign n32211 = ~n32209 & ~n32210 ;
  assign n32212 = \u1_R11_reg[31]/NET0131  & ~n32211 ;
  assign n32213 = ~\u1_R11_reg[31]/NET0131  & n32211 ;
  assign n32214 = ~n32212 & ~n32213 ;
  assign n32240 = ~n32193 & n32207 ;
  assign n32256 = ~n32225 & ~n32240 ;
  assign n32257 = n32214 & ~n32256 ;
  assign n32258 = ~n32231 & n32257 ;
  assign n32217 = ~n32187 & n32193 ;
  assign n32249 = n32207 & n32217 ;
  assign n32250 = n32200 & n32249 ;
  assign n32237 = ~n32200 & ~n32207 ;
  assign n32251 = ~n32187 & n32237 ;
  assign n32252 = n32187 & ~n32207 ;
  assign n32253 = n32200 & n32252 ;
  assign n32254 = ~n32251 & ~n32253 ;
  assign n32255 = ~n32214 & ~n32254 ;
  assign n32259 = ~n32250 & ~n32255 ;
  assign n32260 = ~n32258 & n32259 ;
  assign n32261 = n32181 & ~n32260 ;
  assign n32194 = ~n32187 & ~n32193 ;
  assign n32201 = n32194 & n32200 ;
  assign n32208 = n32193 & n32207 ;
  assign n32215 = ~n32208 & ~n32214 ;
  assign n32216 = ~n32201 & n32215 ;
  assign n32219 = n32200 & ~n32207 ;
  assign n32220 = ~n32193 & n32219 ;
  assign n32221 = n32187 & n32220 ;
  assign n32218 = ~n32207 & n32217 ;
  assign n32222 = n32214 & ~n32218 ;
  assign n32223 = ~n32221 & n32222 ;
  assign n32224 = ~n32216 & ~n32223 ;
  assign n32226 = ~n32214 & n32225 ;
  assign n32227 = n32187 & n32207 ;
  assign n32228 = n32200 & n32227 ;
  assign n32229 = n32193 & n32228 ;
  assign n32232 = ~n32226 & ~n32229 ;
  assign n32233 = ~n32231 & n32232 ;
  assign n32234 = ~n32224 & n32233 ;
  assign n32235 = ~n32181 & ~n32234 ;
  assign n32241 = ~n32187 & n32200 ;
  assign n32242 = n32240 & n32241 ;
  assign n32243 = n32194 & n32237 ;
  assign n32244 = ~n32242 & ~n32243 ;
  assign n32236 = n32217 & n32219 ;
  assign n32238 = n32187 & n32193 ;
  assign n32239 = n32237 & n32238 ;
  assign n32245 = ~n32236 & ~n32239 ;
  assign n32246 = n32244 & n32245 ;
  assign n32247 = n32214 & ~n32246 ;
  assign n32248 = n32226 & n32240 ;
  assign n32262 = ~n32247 & ~n32248 ;
  assign n32263 = ~n32235 & n32262 ;
  assign n32264 = ~n32261 & n32263 ;
  assign n32265 = \u1_L11_reg[5]/NET0131  & ~n32264 ;
  assign n32266 = ~\u1_L11_reg[5]/NET0131  & n32264 ;
  assign n32267 = ~n32265 & ~n32266 ;
  assign n32270 = n31889 & n31901 ;
  assign n32268 = n31877 & n32158 ;
  assign n32271 = n31918 & ~n32268 ;
  assign n32272 = ~n32270 & n32271 ;
  assign n32269 = n31928 & ~n31939 ;
  assign n32273 = ~n31921 & ~n32269 ;
  assign n32274 = n32272 & n32273 ;
  assign n32276 = n31887 & ~n31924 ;
  assign n32275 = ~n31877 & n31906 ;
  assign n32277 = ~n31903 & ~n32275 ;
  assign n32278 = n32276 & n32277 ;
  assign n32279 = ~n31887 & ~n31920 ;
  assign n32280 = ~n32152 & n32279 ;
  assign n32281 = ~n32278 & ~n32280 ;
  assign n32282 = ~n31918 & ~n31944 ;
  assign n32283 = ~n32157 & n32282 ;
  assign n32284 = ~n32281 & n32283 ;
  assign n32285 = ~n32274 & ~n32284 ;
  assign n32287 = ~n31870 & ~n31938 ;
  assign n32288 = ~n32144 & n32287 ;
  assign n32289 = n32276 & ~n32288 ;
  assign n32286 = ~n31887 & ~n32145 ;
  assign n32290 = n31877 & ~n32286 ;
  assign n32291 = ~n32289 & n32290 ;
  assign n32292 = ~n31930 & ~n32291 ;
  assign n32293 = ~n32285 & n32292 ;
  assign n32294 = ~\u1_L11_reg[4]/NET0131  & ~n32293 ;
  assign n32295 = \u1_L11_reg[4]/NET0131  & n32293 ;
  assign n32296 = ~n32294 & ~n32295 ;
  assign n32309 = decrypt_pad & ~\u1_uk_K_r11_reg[12]/NET0131  ;
  assign n32310 = ~decrypt_pad & ~\u1_uk_K_r11_reg[32]/NET0131  ;
  assign n32311 = ~n32309 & ~n32310 ;
  assign n32312 = \u1_R11_reg[6]/NET0131  & ~n32311 ;
  assign n32313 = ~\u1_R11_reg[6]/NET0131  & n32311 ;
  assign n32314 = ~n32312 & ~n32313 ;
  assign n32303 = decrypt_pad & ~\u1_uk_K_r11_reg[34]/NET0131  ;
  assign n32304 = ~decrypt_pad & ~\u1_uk_K_r11_reg[54]/NET0131  ;
  assign n32305 = ~n32303 & ~n32304 ;
  assign n32306 = \u1_R11_reg[9]/NET0131  & ~n32305 ;
  assign n32307 = ~\u1_R11_reg[9]/NET0131  & n32305 ;
  assign n32308 = ~n32306 & ~n32307 ;
  assign n32315 = decrypt_pad & ~\u1_uk_K_r11_reg[46]/NET0131  ;
  assign n32316 = ~decrypt_pad & ~\u1_uk_K_r11_reg[41]/NET0131  ;
  assign n32317 = ~n32315 & ~n32316 ;
  assign n32318 = \u1_R11_reg[5]/NET0131  & ~n32317 ;
  assign n32319 = ~\u1_R11_reg[5]/NET0131  & n32317 ;
  assign n32320 = ~n32318 & ~n32319 ;
  assign n32334 = ~n32308 & n32320 ;
  assign n32322 = decrypt_pad & ~\u1_uk_K_r11_reg[10]/NET0131  ;
  assign n32323 = ~decrypt_pad & ~\u1_uk_K_r11_reg[5]/NET0131  ;
  assign n32324 = ~n32322 & ~n32323 ;
  assign n32325 = \u1_R11_reg[4]/NET0131  & ~n32324 ;
  assign n32326 = ~\u1_R11_reg[4]/NET0131  & n32324 ;
  assign n32327 = ~n32325 & ~n32326 ;
  assign n32335 = n32308 & ~n32320 ;
  assign n32336 = ~n32327 & n32335 ;
  assign n32337 = ~n32334 & ~n32336 ;
  assign n32338 = ~n32314 & ~n32337 ;
  assign n32297 = decrypt_pad & ~\u1_uk_K_r11_reg[6]/NET0131  ;
  assign n32298 = ~decrypt_pad & ~\u1_uk_K_r11_reg[26]/NET0131  ;
  assign n32299 = ~n32297 & ~n32298 ;
  assign n32300 = \u1_R11_reg[7]/NET0131  & ~n32299 ;
  assign n32301 = ~\u1_R11_reg[7]/NET0131  & n32299 ;
  assign n32302 = ~n32300 & ~n32301 ;
  assign n32339 = n32314 & n32327 ;
  assign n32340 = n32302 & n32339 ;
  assign n32341 = n32335 & n32340 ;
  assign n32352 = decrypt_pad & ~\u1_uk_K_r11_reg[54]/NET0131  ;
  assign n32353 = ~decrypt_pad & ~\u1_uk_K_r11_reg[17]/NET0131  ;
  assign n32354 = ~n32352 & ~n32353 ;
  assign n32355 = \u1_R11_reg[8]/NET0131  & ~n32354 ;
  assign n32356 = ~\u1_R11_reg[8]/NET0131  & n32354 ;
  assign n32357 = ~n32355 & ~n32356 ;
  assign n32358 = ~n32341 & ~n32357 ;
  assign n32359 = ~n32338 & n32358 ;
  assign n32342 = ~n32302 & ~n32320 ;
  assign n32343 = n32308 & ~n32314 ;
  assign n32344 = n32342 & n32343 ;
  assign n32345 = n32308 & ~n32327 ;
  assign n32346 = n32320 & n32345 ;
  assign n32347 = n32314 & n32346 ;
  assign n32348 = ~n32344 & ~n32347 ;
  assign n32349 = ~n32335 & n32339 ;
  assign n32350 = ~n32336 & ~n32349 ;
  assign n32351 = ~n32302 & ~n32350 ;
  assign n32360 = n32348 & ~n32351 ;
  assign n32361 = n32359 & n32360 ;
  assign n32363 = n32308 & n32327 ;
  assign n32366 = ~n32308 & ~n32327 ;
  assign n32370 = ~n32363 & ~n32366 ;
  assign n32368 = n32320 & n32327 ;
  assign n32369 = ~n32302 & ~n32368 ;
  assign n32371 = n32314 & n32369 ;
  assign n32372 = ~n32370 & n32371 ;
  assign n32330 = ~n32314 & n32327 ;
  assign n32376 = ~n32308 & n32330 ;
  assign n32377 = ~n32320 & n32376 ;
  assign n32362 = ~n32314 & n32320 ;
  assign n32364 = n32362 & n32363 ;
  assign n32365 = n32357 & ~n32364 ;
  assign n32367 = n32342 & n32366 ;
  assign n32373 = n32314 & ~n32327 ;
  assign n32374 = n32302 & n32320 ;
  assign n32375 = ~n32373 & n32374 ;
  assign n32378 = ~n32367 & ~n32375 ;
  assign n32379 = n32365 & n32378 ;
  assign n32380 = ~n32377 & n32379 ;
  assign n32381 = ~n32372 & n32380 ;
  assign n32382 = ~n32361 & ~n32381 ;
  assign n32321 = n32314 & ~n32320 ;
  assign n32328 = n32321 & ~n32327 ;
  assign n32329 = ~n32308 & n32328 ;
  assign n32331 = n32320 & n32330 ;
  assign n32332 = ~n32329 & ~n32331 ;
  assign n32333 = n32302 & ~n32332 ;
  assign n32383 = ~n32321 & ~n32362 ;
  assign n32384 = ~n32302 & n32345 ;
  assign n32385 = n32383 & n32384 ;
  assign n32386 = ~n32333 & ~n32385 ;
  assign n32387 = ~n32382 & n32386 ;
  assign n32388 = \u1_L11_reg[2]/NET0131  & n32387 ;
  assign n32389 = ~\u1_L11_reg[2]/NET0131  & ~n32387 ;
  assign n32390 = ~n32388 & ~n32389 ;
  assign n32402 = n32048 & ~n32113 ;
  assign n32403 = ~n32089 & n32402 ;
  assign n32404 = n32060 & ~n32067 ;
  assign n32405 = n32080 & ~n32404 ;
  assign n32406 = n32076 & ~n32405 ;
  assign n32407 = ~n32403 & ~n32406 ;
  assign n32408 = n32067 & n32101 ;
  assign n32409 = ~n32054 & n32081 ;
  assign n32410 = n32073 & n32409 ;
  assign n32411 = ~n32408 & ~n32410 ;
  assign n32412 = ~n32407 & n32411 ;
  assign n32413 = n32097 & ~n32412 ;
  assign n32391 = n32060 & n32111 ;
  assign n32392 = n32100 & n32121 ;
  assign n32396 = ~n32391 & ~n32392 ;
  assign n32397 = ~n32118 & n32396 ;
  assign n32393 = n32048 & ~n32074 ;
  assign n32394 = n32122 & n32393 ;
  assign n32395 = ~n32067 & n32127 ;
  assign n32398 = ~n32394 & ~n32395 ;
  assign n32399 = n32397 & n32398 ;
  assign n32400 = n32091 & n32399 ;
  assign n32401 = ~n32097 & ~n32400 ;
  assign n32414 = ~n32079 & n32411 ;
  assign n32415 = ~n32048 & ~n32414 ;
  assign n32416 = ~n32088 & ~n32110 ;
  assign n32417 = ~n32415 & n32416 ;
  assign n32418 = ~n32401 & n32417 ;
  assign n32419 = ~n32413 & n32418 ;
  assign n32420 = ~\u1_L11_reg[10]/NET0131  & ~n32419 ;
  assign n32421 = \u1_L11_reg[10]/NET0131  & n32419 ;
  assign n32422 = ~n32420 & ~n32421 ;
  assign n32429 = ~n31961 & ~n32015 ;
  assign n32430 = n31967 & ~n31990 ;
  assign n32431 = n31961 & ~n32430 ;
  assign n32432 = ~n32429 & ~n32431 ;
  assign n32428 = ~n31968 & n31982 ;
  assign n32433 = ~n31969 & n31990 ;
  assign n32434 = ~n32428 & ~n32433 ;
  assign n32435 = ~n32432 & n32434 ;
  assign n32425 = n31982 & n31990 ;
  assign n32426 = ~n31991 & ~n32425 ;
  assign n32427 = ~n31976 & ~n32426 ;
  assign n32423 = ~n31998 & ~n32026 ;
  assign n32424 = n31995 & ~n32423 ;
  assign n32436 = n31969 & ~n31976 ;
  assign n32437 = ~n32014 & ~n32436 ;
  assign n32438 = ~n32424 & n32437 ;
  assign n32439 = ~n32427 & n32438 ;
  assign n32440 = ~n32435 & n32439 ;
  assign n32441 = ~n31982 & ~n31997 ;
  assign n32442 = n31976 & ~n32441 ;
  assign n32443 = ~n32429 & n32442 ;
  assign n32445 = ~n32004 & ~n32430 ;
  assign n32446 = n32018 & ~n32445 ;
  assign n32444 = ~n31976 & n31996 ;
  assign n32447 = n32014 & ~n32444 ;
  assign n32448 = ~n32446 & n32447 ;
  assign n32449 = ~n32443 & n32448 ;
  assign n32450 = ~n32440 & ~n32449 ;
  assign n32451 = \u1_L11_reg[12]/NET0131  & n32450 ;
  assign n32452 = ~\u1_L11_reg[12]/NET0131  & ~n32450 ;
  assign n32453 = ~n32451 & ~n32452 ;
  assign n32456 = n32320 & n32366 ;
  assign n32457 = n32335 & n32373 ;
  assign n32458 = ~n32456 & ~n32457 ;
  assign n32459 = ~n32377 & n32458 ;
  assign n32460 = ~n32357 & ~n32459 ;
  assign n32454 = ~n32308 & n32368 ;
  assign n32455 = n32314 & n32454 ;
  assign n32461 = ~n32364 & ~n32455 ;
  assign n32462 = ~n32460 & n32461 ;
  assign n32463 = ~n32302 & ~n32462 ;
  assign n32464 = ~n32320 & ~n32370 ;
  assign n32465 = ~n32314 & n32454 ;
  assign n32466 = ~n32464 & ~n32465 ;
  assign n32467 = n32302 & ~n32466 ;
  assign n32469 = ~n32327 & ~n32342 ;
  assign n32470 = n32343 & n32469 ;
  assign n32468 = ~n32334 & n32340 ;
  assign n32471 = ~n32357 & ~n32468 ;
  assign n32472 = ~n32470 & n32471 ;
  assign n32473 = ~n32467 & n32472 ;
  assign n32482 = n32362 & n32366 ;
  assign n32483 = n32365 & ~n32482 ;
  assign n32479 = ~n32308 & ~n32314 ;
  assign n32480 = n32342 & ~n32345 ;
  assign n32481 = ~n32479 & n32480 ;
  assign n32484 = ~n32455 & ~n32481 ;
  assign n32485 = n32483 & n32484 ;
  assign n32474 = ~n32308 & ~n32320 ;
  assign n32475 = ~n32314 & n32474 ;
  assign n32476 = n32314 & n32345 ;
  assign n32477 = ~n32475 & ~n32476 ;
  assign n32478 = n32302 & ~n32477 ;
  assign n32486 = n32348 & ~n32478 ;
  assign n32487 = n32485 & n32486 ;
  assign n32488 = ~n32473 & ~n32487 ;
  assign n32489 = ~n32463 & ~n32488 ;
  assign n32490 = ~\u1_L11_reg[13]/NET0131  & n32489 ;
  assign n32491 = \u1_L11_reg[13]/NET0131  & ~n32489 ;
  assign n32492 = ~n32490 & ~n32491 ;
  assign n32493 = ~n32207 & n32230 ;
  assign n32494 = ~n32200 & n32207 ;
  assign n32495 = ~n32193 & n32494 ;
  assign n32496 = ~n32218 & ~n32227 ;
  assign n32497 = ~n32495 & n32496 ;
  assign n32498 = n32214 & ~n32497 ;
  assign n32499 = ~n32493 & ~n32498 ;
  assign n32500 = ~n32181 & ~n32499 ;
  assign n32508 = ~n32187 & n32214 ;
  assign n32509 = n32193 & n32219 ;
  assign n32510 = ~n32508 & n32509 ;
  assign n32507 = ~n32200 & n32227 ;
  assign n32505 = ~n32207 & n32214 ;
  assign n32506 = n32194 & n32505 ;
  assign n32511 = ~n32242 & ~n32506 ;
  assign n32512 = ~n32507 & n32511 ;
  assign n32513 = ~n32510 & n32512 ;
  assign n32514 = n32181 & ~n32513 ;
  assign n32501 = ~n32219 & ~n32249 ;
  assign n32502 = ~n32241 & ~n32501 ;
  assign n32503 = n32244 & ~n32502 ;
  assign n32504 = ~n32214 & ~n32503 ;
  assign n32515 = n32193 & n32251 ;
  assign n32516 = ~n32250 & ~n32515 ;
  assign n32517 = n32214 & ~n32516 ;
  assign n32518 = ~n32181 & ~n32214 ;
  assign n32519 = n32252 & n32518 ;
  assign n32520 = ~n32517 & ~n32519 ;
  assign n32521 = ~n32504 & n32520 ;
  assign n32522 = ~n32514 & n32521 ;
  assign n32523 = ~n32500 & n32522 ;
  assign n32524 = ~\u1_L11_reg[15]/P0001  & ~n32523 ;
  assign n32525 = \u1_L11_reg[15]/P0001  & n32523 ;
  assign n32526 = ~n32524 & ~n32525 ;
  assign n32529 = ~n31887 & n32288 ;
  assign n32527 = ~n31880 & n31887 ;
  assign n32528 = ~n32287 & n32527 ;
  assign n32530 = n31870 & n32268 ;
  assign n32531 = ~n31918 & ~n32530 ;
  assign n32532 = ~n32528 & n32531 ;
  assign n32533 = ~n32529 & n32532 ;
  assign n32534 = n31877 & n32288 ;
  assign n32539 = ~n31907 & n31918 ;
  assign n32540 = ~n32534 & n32539 ;
  assign n32535 = ~n31938 & ~n32151 ;
  assign n32536 = ~n31877 & ~n32535 ;
  assign n32537 = ~n31887 & ~n32156 ;
  assign n32538 = ~n32527 & ~n32537 ;
  assign n32541 = ~n32536 & ~n32538 ;
  assign n32542 = n32540 & n32541 ;
  assign n32543 = ~n32533 & ~n32542 ;
  assign n32544 = ~n31927 & ~n31945 ;
  assign n32545 = ~n32543 & n32544 ;
  assign n32546 = ~\u1_L11_reg[19]/P0001  & ~n32545 ;
  assign n32547 = \u1_L11_reg[19]/P0001  & n32545 ;
  assign n32548 = ~n32546 & ~n32547 ;
  assign n32558 = n32193 & n32225 ;
  assign n32559 = ~n32505 & n32558 ;
  assign n32553 = n32207 & n32241 ;
  assign n32560 = ~n32181 & ~n32553 ;
  assign n32554 = n32200 & ~n32214 ;
  assign n32555 = n32217 & n32554 ;
  assign n32556 = ~n32187 & ~n32214 ;
  assign n32557 = n32240 & n32556 ;
  assign n32561 = ~n32555 & ~n32557 ;
  assign n32562 = n32560 & n32561 ;
  assign n32563 = ~n32559 & n32562 ;
  assign n32549 = ~n32193 & ~n32254 ;
  assign n32550 = n32187 & n32240 ;
  assign n32551 = ~n32253 & ~n32550 ;
  assign n32552 = n32214 & ~n32551 ;
  assign n32564 = ~n32549 & ~n32552 ;
  assign n32565 = n32563 & n32564 ;
  assign n32567 = n32214 & ~n32228 ;
  assign n32566 = n32193 & n32237 ;
  assign n32568 = ~n32249 & ~n32566 ;
  assign n32569 = n32567 & n32568 ;
  assign n32570 = n32219 & n32238 ;
  assign n32571 = ~n32214 & ~n32230 ;
  assign n32572 = ~n32570 & n32571 ;
  assign n32573 = ~n32569 & ~n32572 ;
  assign n32574 = n32194 & ~n32207 ;
  assign n32575 = ~n32550 & ~n32574 ;
  assign n32576 = n32200 & ~n32575 ;
  assign n32577 = n32181 & ~n32515 ;
  assign n32578 = ~n32576 & n32577 ;
  assign n32579 = ~n32573 & n32578 ;
  assign n32580 = ~n32565 & ~n32579 ;
  assign n32581 = n32208 & n32226 ;
  assign n32582 = n32214 & n32251 ;
  assign n32583 = ~n32581 & ~n32582 ;
  assign n32584 = ~n32580 & n32583 ;
  assign n32585 = ~\u1_L11_reg[21]/NET0131  & ~n32584 ;
  assign n32586 = \u1_L11_reg[21]/NET0131  & n32584 ;
  assign n32587 = ~n32585 & ~n32586 ;
  assign n32608 = ~n32105 & ~n32112 ;
  assign n32609 = n32097 & ~n32608 ;
  assign n32610 = ~n32090 & n32411 ;
  assign n32611 = ~n32609 & n32610 ;
  assign n32612 = n32048 & ~n32611 ;
  assign n32588 = ~n32077 & ~n32105 ;
  assign n32589 = n32054 & ~n32588 ;
  assign n32590 = ~n32048 & ~n32589 ;
  assign n32591 = ~n32078 & n32083 ;
  assign n32592 = ~n32590 & ~n32591 ;
  assign n32593 = ~n32080 & ~n32126 ;
  assign n32594 = n32404 & ~n32593 ;
  assign n32595 = ~n32408 & ~n32594 ;
  assign n32596 = ~n32592 & n32595 ;
  assign n32597 = ~n32097 & ~n32596 ;
  assign n32598 = ~n32080 & n32404 ;
  assign n32599 = n32060 & n32126 ;
  assign n32600 = ~n32598 & ~n32599 ;
  assign n32601 = ~n32048 & ~n32600 ;
  assign n32602 = n32060 & n32104 ;
  assign n32603 = ~n32409 & ~n32602 ;
  assign n32604 = ~n32601 & n32603 ;
  assign n32605 = n32097 & ~n32604 ;
  assign n32606 = ~n32048 & ~n32073 ;
  assign n32607 = ~n32603 & n32606 ;
  assign n32613 = ~n32605 & ~n32607 ;
  assign n32614 = ~n32597 & n32613 ;
  assign n32615 = ~n32612 & n32614 ;
  assign n32616 = ~\u1_L11_reg[1]/NET0131  & ~n32615 ;
  assign n32617 = \u1_L11_reg[1]/NET0131  & n32615 ;
  assign n32618 = ~n32616 & ~n32617 ;
  assign n32634 = ~n31804 & ~n31817 ;
  assign n32635 = ~n31774 & ~n32634 ;
  assign n32636 = n31774 & n32634 ;
  assign n32637 = ~n32635 & ~n32636 ;
  assign n32638 = n31796 & ~n31846 ;
  assign n32639 = ~n31768 & ~n32638 ;
  assign n32640 = n32637 & n32639 ;
  assign n32641 = n31782 & n31817 ;
  assign n32642 = n31820 & n31843 ;
  assign n32643 = ~n32641 & ~n32642 ;
  assign n32644 = ~n31835 & n32643 ;
  assign n32645 = ~n31842 & n32644 ;
  assign n32646 = ~n32640 & n32645 ;
  assign n32647 = n31813 & ~n32646 ;
  assign n32619 = ~n31768 & n31796 ;
  assign n32620 = ~n31782 & n32619 ;
  assign n32621 = ~n31841 & n32620 ;
  assign n32622 = ~n31789 & ~n31844 ;
  assign n32623 = ~n31822 & n32622 ;
  assign n32624 = ~n32621 & n32623 ;
  assign n32625 = ~n31813 & ~n32624 ;
  assign n32629 = ~n31804 & ~n31843 ;
  assign n32630 = ~n31781 & ~n31826 ;
  assign n32631 = n32629 & n32630 ;
  assign n32632 = ~n31845 & ~n32631 ;
  assign n32633 = ~n31768 & ~n32632 ;
  assign n32626 = n31781 & n31813 ;
  assign n32627 = n31820 & n31833 ;
  assign n32628 = ~n32626 & n32627 ;
  assign n32648 = ~n31852 & ~n32628 ;
  assign n32649 = ~n32633 & n32648 ;
  assign n32650 = ~n32625 & n32649 ;
  assign n32651 = ~n32647 & n32650 ;
  assign n32652 = \u1_L11_reg[23]/NET0131  & ~n32651 ;
  assign n32653 = ~\u1_L11_reg[23]/NET0131  & n32651 ;
  assign n32654 = ~n32652 & ~n32653 ;
  assign n32684 = decrypt_pad & ~\u1_uk_K_r11_reg[21]/NET0131  ;
  assign n32685 = ~decrypt_pad & ~\u1_uk_K_r11_reg[43]/NET0131  ;
  assign n32686 = ~n32684 & ~n32685 ;
  assign n32687 = \u1_R11_reg[19]/NET0131  & ~n32686 ;
  assign n32688 = ~\u1_R11_reg[19]/NET0131  & n32686 ;
  assign n32689 = ~n32687 & ~n32688 ;
  assign n32655 = decrypt_pad & ~\u1_uk_K_r11_reg[16]/NET0131  ;
  assign n32656 = ~decrypt_pad & ~\u1_uk_K_r11_reg[7]/NET0131  ;
  assign n32657 = ~n32655 & ~n32656 ;
  assign n32658 = \u1_R11_reg[17]/NET0131  & ~n32657 ;
  assign n32659 = ~\u1_R11_reg[17]/NET0131  & n32657 ;
  assign n32660 = ~n32658 & ~n32659 ;
  assign n32668 = decrypt_pad & ~\u1_uk_K_r11_reg[37]/NET0131  ;
  assign n32669 = ~decrypt_pad & ~\u1_uk_K_r11_reg[28]/NET0131  ;
  assign n32670 = ~n32668 & ~n32669 ;
  assign n32671 = \u1_R11_reg[21]/NET0131  & ~n32670 ;
  assign n32672 = ~\u1_R11_reg[21]/NET0131  & n32670 ;
  assign n32673 = ~n32671 & ~n32672 ;
  assign n32675 = decrypt_pad & ~\u1_uk_K_r11_reg[49]/NET0131  ;
  assign n32676 = ~decrypt_pad & ~\u1_uk_K_r11_reg[16]/NET0131  ;
  assign n32677 = ~n32675 & ~n32676 ;
  assign n32678 = \u1_R11_reg[16]/NET0131  & ~n32677 ;
  assign n32679 = ~\u1_R11_reg[16]/NET0131  & n32677 ;
  assign n32680 = ~n32678 & ~n32679 ;
  assign n32690 = n32673 & n32680 ;
  assign n32691 = ~n32660 & n32690 ;
  assign n32692 = ~n32689 & ~n32691 ;
  assign n32661 = decrypt_pad & ~\u1_uk_K_r11_reg[38]/NET0131  ;
  assign n32662 = ~decrypt_pad & ~\u1_uk_K_r11_reg[1]/NET0131  ;
  assign n32663 = ~n32661 & ~n32662 ;
  assign n32664 = \u1_R11_reg[18]/NET0131  & ~n32663 ;
  assign n32665 = ~\u1_R11_reg[18]/NET0131  & n32663 ;
  assign n32666 = ~n32664 & ~n32665 ;
  assign n32667 = n32660 & ~n32666 ;
  assign n32693 = n32667 & ~n32680 ;
  assign n32694 = n32692 & ~n32693 ;
  assign n32696 = ~n32660 & ~n32666 ;
  assign n32697 = n32666 & ~n32680 ;
  assign n32698 = ~n32696 & ~n32697 ;
  assign n32699 = ~n32673 & ~n32698 ;
  assign n32700 = n32660 & n32690 ;
  assign n32695 = ~n32660 & ~n32680 ;
  assign n32701 = n32689 & ~n32695 ;
  assign n32702 = ~n32700 & n32701 ;
  assign n32703 = ~n32699 & n32702 ;
  assign n32704 = ~n32694 & ~n32703 ;
  assign n32674 = n32667 & n32673 ;
  assign n32681 = ~n32673 & n32680 ;
  assign n32682 = n32660 & n32681 ;
  assign n32683 = n32666 & n32682 ;
  assign n32705 = ~n32674 & ~n32683 ;
  assign n32706 = ~n32704 & n32705 ;
  assign n32707 = decrypt_pad & ~\u1_uk_K_r11_reg[36]/NET0131  ;
  assign n32708 = ~decrypt_pad & ~\u1_uk_K_r11_reg[31]/NET0131  ;
  assign n32709 = ~n32707 & ~n32708 ;
  assign n32710 = \u1_R11_reg[20]/NET0131  & ~n32709 ;
  assign n32711 = ~\u1_R11_reg[20]/NET0131  & n32709 ;
  assign n32712 = ~n32710 & ~n32711 ;
  assign n32713 = ~n32706 & n32712 ;
  assign n32729 = ~n32673 & ~n32680 ;
  assign n32730 = ~n32660 & n32729 ;
  assign n32731 = n32666 & n32730 ;
  assign n32732 = ~n32683 & ~n32731 ;
  assign n32733 = n32673 & ~n32680 ;
  assign n32734 = n32696 & n32733 ;
  assign n32735 = n32732 & ~n32734 ;
  assign n32736 = n32689 & ~n32735 ;
  assign n32714 = ~n32673 & n32689 ;
  assign n32716 = n32666 & n32714 ;
  assign n32715 = ~n32697 & ~n32714 ;
  assign n32717 = n32660 & ~n32715 ;
  assign n32718 = ~n32716 & n32717 ;
  assign n32719 = ~n32660 & ~n32689 ;
  assign n32720 = ~n32690 & n32719 ;
  assign n32721 = ~n32697 & n32720 ;
  assign n32722 = ~n32718 & ~n32721 ;
  assign n32723 = ~n32712 & ~n32722 ;
  assign n32724 = ~n32666 & n32690 ;
  assign n32725 = n32660 & n32724 ;
  assign n32726 = ~n32660 & n32680 ;
  assign n32727 = n32666 & ~n32689 ;
  assign n32728 = n32726 & n32727 ;
  assign n32737 = ~n32725 & ~n32728 ;
  assign n32738 = ~n32723 & n32737 ;
  assign n32739 = ~n32736 & n32738 ;
  assign n32740 = ~n32713 & n32739 ;
  assign n32741 = ~\u1_L11_reg[25]/NET0131  & ~n32740 ;
  assign n32742 = \u1_L11_reg[25]/NET0131  & n32740 ;
  assign n32743 = ~n32741 & ~n32742 ;
  assign n32746 = n32320 & ~n32479 ;
  assign n32747 = ~n32370 & n32746 ;
  assign n32744 = n32314 & ~n32474 ;
  assign n32745 = n32327 & ~n32744 ;
  assign n32748 = n32302 & ~n32457 ;
  assign n32749 = ~n32745 & n32748 ;
  assign n32750 = ~n32747 & n32749 ;
  assign n32753 = ~n32328 & ~n32455 ;
  assign n32751 = ~n32302 & ~n32346 ;
  assign n32752 = ~n32314 & n32366 ;
  assign n32754 = n32330 & n32335 ;
  assign n32755 = ~n32752 & ~n32754 ;
  assign n32756 = n32751 & n32755 ;
  assign n32757 = n32753 & n32756 ;
  assign n32758 = ~n32750 & ~n32757 ;
  assign n32759 = n32357 & ~n32758 ;
  assign n32760 = ~n32336 & n32369 ;
  assign n32761 = ~n32376 & n32760 ;
  assign n32762 = n32753 & n32761 ;
  assign n32763 = n32302 & ~n32346 ;
  assign n32764 = ~n32752 & n32763 ;
  assign n32765 = ~n32762 & ~n32764 ;
  assign n32766 = ~n32454 & ~n32464 ;
  assign n32767 = n32314 & ~n32766 ;
  assign n32768 = ~n32357 & ~n32767 ;
  assign n32769 = ~n32765 & n32768 ;
  assign n32770 = ~n32759 & ~n32769 ;
  assign n32771 = \u1_L11_reg[28]/NET0131  & n32770 ;
  assign n32772 = ~\u1_L11_reg[28]/NET0131  & ~n32770 ;
  assign n32773 = ~n32771 & ~n32772 ;
  assign n32776 = n32689 & ~n32693 ;
  assign n32775 = n32666 & n32690 ;
  assign n32777 = ~n32730 & ~n32775 ;
  assign n32778 = n32776 & n32777 ;
  assign n32779 = n32681 & n32696 ;
  assign n32783 = ~n32689 & ~n32779 ;
  assign n32780 = n32660 & n32666 ;
  assign n32781 = ~n32673 & n32780 ;
  assign n32782 = n32673 & n32695 ;
  assign n32784 = ~n32781 & ~n32782 ;
  assign n32785 = n32783 & n32784 ;
  assign n32786 = ~n32725 & n32785 ;
  assign n32787 = ~n32778 & ~n32786 ;
  assign n32774 = n32666 & n32691 ;
  assign n32788 = n32667 & n32729 ;
  assign n32789 = ~n32774 & ~n32788 ;
  assign n32790 = ~n32787 & n32789 ;
  assign n32791 = ~n32712 & ~n32790 ;
  assign n32795 = ~n32667 & n32733 ;
  assign n32796 = ~n32682 & ~n32724 ;
  assign n32797 = ~n32795 & n32796 ;
  assign n32798 = n32689 & ~n32797 ;
  assign n32799 = ~n32666 & ~n32689 ;
  assign n32800 = n32660 & n32733 ;
  assign n32801 = ~n32730 & ~n32800 ;
  assign n32802 = n32799 & ~n32801 ;
  assign n32792 = ~n32660 & n32666 ;
  assign n32793 = ~n32667 & ~n32792 ;
  assign n32794 = n32681 & ~n32793 ;
  assign n32803 = n32660 & ~n32727 ;
  assign n32804 = n32690 & ~n32792 ;
  assign n32805 = ~n32803 & n32804 ;
  assign n32806 = ~n32794 & ~n32805 ;
  assign n32807 = ~n32802 & n32806 ;
  assign n32808 = ~n32798 & n32807 ;
  assign n32809 = n32712 & ~n32808 ;
  assign n32810 = ~n32666 & n32682 ;
  assign n32811 = ~n32731 & ~n32810 ;
  assign n32812 = n32689 & ~n32811 ;
  assign n32813 = n32733 & n32792 ;
  assign n32814 = ~n32680 & n32781 ;
  assign n32815 = ~n32813 & ~n32814 ;
  assign n32816 = ~n32689 & ~n32815 ;
  assign n32817 = ~n32812 & ~n32816 ;
  assign n32818 = ~n32809 & n32817 ;
  assign n32819 = ~n32791 & n32818 ;
  assign n32820 = ~\u1_L11_reg[14]/NET0131  & ~n32819 ;
  assign n32821 = \u1_L11_reg[14]/NET0131  & n32819 ;
  assign n32822 = ~n32820 & ~n32821 ;
  assign n32823 = ~n32075 & n32402 ;
  assign n32824 = ~n32073 & ~n32123 ;
  assign n32825 = ~n32101 & ~n32824 ;
  assign n32826 = ~n32067 & ~n32825 ;
  assign n32827 = ~n32098 & ~n32409 ;
  assign n32828 = ~n32097 & ~n32827 ;
  assign n32829 = ~n32048 & ~n32828 ;
  assign n32830 = ~n32826 & n32829 ;
  assign n32831 = ~n32823 & ~n32830 ;
  assign n32840 = n32097 & ~n32602 ;
  assign n32836 = n32048 & n32099 ;
  assign n32839 = ~n32067 & n32089 ;
  assign n32841 = ~n32836 & ~n32839 ;
  assign n32842 = n32840 & n32841 ;
  assign n32832 = ~n32060 & n32074 ;
  assign n32833 = ~n32100 & ~n32832 ;
  assign n32834 = ~n32048 & ~n32111 ;
  assign n32835 = ~n32833 & n32834 ;
  assign n32837 = ~n32127 & ~n32599 ;
  assign n32838 = n32067 & ~n32837 ;
  assign n32843 = ~n32835 & ~n32838 ;
  assign n32844 = n32842 & n32843 ;
  assign n32845 = n32109 & ~n32126 ;
  assign n32846 = ~n32097 & ~n32112 ;
  assign n32847 = n32125 & n32846 ;
  assign n32848 = ~n32845 & n32847 ;
  assign n32849 = ~n32844 & ~n32848 ;
  assign n32850 = ~n32831 & ~n32849 ;
  assign n32851 = ~\u1_L11_reg[26]/NET0131  & ~n32850 ;
  assign n32852 = \u1_L11_reg[26]/NET0131  & n32850 ;
  assign n32853 = ~n32851 & ~n32852 ;
  assign n32854 = n32681 & n32792 ;
  assign n32855 = ~n32689 & ~n32854 ;
  assign n32856 = n32689 & ~n32733 ;
  assign n32857 = ~n32793 & ~n32856 ;
  assign n32858 = ~n32781 & ~n32857 ;
  assign n32859 = ~n32855 & ~n32858 ;
  assign n32861 = ~n32666 & n32730 ;
  assign n32862 = ~n32691 & ~n32861 ;
  assign n32863 = n32689 & ~n32862 ;
  assign n32860 = n32680 & n32799 ;
  assign n32864 = n32712 & ~n32860 ;
  assign n32865 = n32815 & n32864 ;
  assign n32866 = ~n32863 & n32865 ;
  assign n32867 = n32733 & ~n32792 ;
  assign n32868 = n32692 & ~n32867 ;
  assign n32869 = n32689 & ~n32779 ;
  assign n32870 = ~n32700 & n32869 ;
  assign n32871 = ~n32868 & ~n32870 ;
  assign n32872 = ~n32693 & ~n32712 ;
  assign n32873 = n32732 & n32872 ;
  assign n32874 = ~n32871 & n32873 ;
  assign n32875 = ~n32866 & ~n32874 ;
  assign n32876 = ~n32859 & ~n32875 ;
  assign n32877 = ~\u1_L11_reg[8]/NET0131  & ~n32876 ;
  assign n32878 = \u1_L11_reg[8]/NET0131  & n32876 ;
  assign n32879 = ~n32877 & ~n32878 ;
  assign n32887 = ~n32221 & ~n32566 ;
  assign n32888 = ~n32250 & n32887 ;
  assign n32880 = ~n32194 & ~n32238 ;
  assign n32881 = n32207 & ~n32880 ;
  assign n32882 = n32214 & ~n32241 ;
  assign n32883 = n32881 & n32882 ;
  assign n32884 = ~n32214 & ~n32219 ;
  assign n32885 = ~n32252 & n32884 ;
  assign n32886 = ~n32881 & n32885 ;
  assign n32889 = ~n32883 & ~n32886 ;
  assign n32890 = n32888 & n32889 ;
  assign n32891 = n32181 & ~n32890 ;
  assign n32894 = n32214 & ~n32495 ;
  assign n32893 = n32193 & ~n32494 ;
  assign n32895 = ~n32553 & ~n32893 ;
  assign n32896 = n32894 & n32895 ;
  assign n32892 = n32238 & n32554 ;
  assign n32897 = ~n32236 & ~n32557 ;
  assign n32898 = ~n32892 & n32897 ;
  assign n32899 = ~n32896 & n32898 ;
  assign n32900 = ~n32181 & ~n32899 ;
  assign n32901 = ~n32239 & ~n32242 ;
  assign n32902 = ~n32214 & ~n32901 ;
  assign n32903 = n32214 & n32220 ;
  assign n32904 = ~n32248 & ~n32903 ;
  assign n32905 = ~n32902 & n32904 ;
  assign n32906 = ~n32900 & n32905 ;
  assign n32907 = ~n32891 & n32906 ;
  assign n32908 = ~\u1_L11_reg[27]/NET0131  & ~n32907 ;
  assign n32909 = \u1_L11_reg[27]/NET0131  & n32907 ;
  assign n32910 = ~n32908 & ~n32909 ;
  assign n32911 = n31976 & ~n31996 ;
  assign n32912 = ~n31961 & n31998 ;
  assign n32913 = ~n31976 & ~n32912 ;
  assign n32914 = ~n32005 & n32913 ;
  assign n32915 = ~n32911 & ~n32914 ;
  assign n32921 = n31961 & n31990 ;
  assign n32922 = ~n31997 & ~n32921 ;
  assign n32923 = ~n32004 & n32426 ;
  assign n32924 = ~n32922 & ~n32923 ;
  assign n32925 = ~n32015 & n32922 ;
  assign n32926 = ~n31976 & ~n32925 ;
  assign n32927 = ~n32924 & n32926 ;
  assign n32919 = n31982 & ~n32004 ;
  assign n32920 = n32442 & ~n32919 ;
  assign n32916 = ~n31976 & ~n31982 ;
  assign n32917 = n31969 & ~n31990 ;
  assign n32918 = ~n32916 & n32917 ;
  assign n32928 = n32014 & ~n32918 ;
  assign n32929 = ~n32920 & n32928 ;
  assign n32930 = ~n32927 & n32929 ;
  assign n32933 = ~n32026 & ~n32919 ;
  assign n32934 = n32431 & ~n32933 ;
  assign n32931 = n31961 & n32015 ;
  assign n32932 = n32427 & ~n32931 ;
  assign n32935 = n32000 & ~n32014 ;
  assign n32936 = ~n32932 & n32935 ;
  assign n32937 = ~n32934 & n32936 ;
  assign n32938 = ~n32930 & ~n32937 ;
  assign n32939 = ~n32915 & ~n32938 ;
  assign n32940 = \u1_L11_reg[32]/NET0131  & n32939 ;
  assign n32941 = ~\u1_L11_reg[32]/NET0131  & ~n32939 ;
  assign n32942 = ~n32940 & ~n32941 ;
  assign n32943 = n32712 & ~n32854 ;
  assign n32944 = ~n32725 & n32943 ;
  assign n32945 = ~n32800 & n32944 ;
  assign n32946 = ~n32666 & ~n32726 ;
  assign n32947 = n32673 & ~n32946 ;
  assign n32948 = ~n32712 & ~n32729 ;
  assign n32949 = ~n32947 & n32948 ;
  assign n32950 = ~n32945 & ~n32949 ;
  assign n32951 = ~n32689 & ~n32774 ;
  assign n32952 = ~n32810 & ~n32861 ;
  assign n32953 = n32951 & n32952 ;
  assign n32954 = ~n32950 & n32953 ;
  assign n32957 = ~n32682 & ~n32712 ;
  assign n32955 = ~n32666 & n32733 ;
  assign n32956 = ~n32681 & n32792 ;
  assign n32958 = ~n32955 & ~n32956 ;
  assign n32959 = n32957 & n32958 ;
  assign n32960 = n32660 & n32729 ;
  assign n32961 = ~n32724 & ~n32960 ;
  assign n32962 = n32944 & n32961 ;
  assign n32963 = ~n32959 & ~n32962 ;
  assign n32964 = ~n32813 & n32869 ;
  assign n32965 = ~n32963 & n32964 ;
  assign n32966 = ~n32954 & ~n32965 ;
  assign n32967 = ~\u1_L11_reg[3]/NET0131  & n32966 ;
  assign n32968 = \u1_L11_reg[3]/NET0131  & ~n32966 ;
  assign n32969 = ~n32967 & ~n32968 ;
  assign n33004 = decrypt_pad & ~\u1_uk_K_r11_reg[17]/NET0131  ;
  assign n33005 = ~decrypt_pad & ~\u1_uk_K_r11_reg[12]/NET0131  ;
  assign n33006 = ~n33004 & ~n33005 ;
  assign n33007 = \u1_R11_reg[11]/NET0131  & ~n33006 ;
  assign n33008 = ~\u1_R11_reg[11]/NET0131  & n33006 ;
  assign n33009 = ~n33007 & ~n33008 ;
  assign n32996 = decrypt_pad & ~\u1_uk_K_r11_reg[32]/NET0131  ;
  assign n32997 = ~decrypt_pad & ~\u1_uk_K_r11_reg[27]/P0001  ;
  assign n32998 = ~n32996 & ~n32997 ;
  assign n32999 = \u1_R11_reg[12]/NET0131  & ~n32998 ;
  assign n33000 = ~\u1_R11_reg[12]/NET0131  & n32998 ;
  assign n33001 = ~n32999 & ~n33000 ;
  assign n32970 = decrypt_pad & ~\u1_uk_K_r11_reg[20]/NET0131  ;
  assign n32971 = ~decrypt_pad & ~\u1_uk_K_r11_reg[40]/NET0131  ;
  assign n32972 = ~n32970 & ~n32971 ;
  assign n32973 = \u1_R11_reg[13]/NET0131  & ~n32972 ;
  assign n32974 = ~\u1_R11_reg[13]/NET0131  & n32972 ;
  assign n32975 = ~n32973 & ~n32974 ;
  assign n32983 = decrypt_pad & ~\u1_uk_K_r11_reg[40]/NET0131  ;
  assign n32984 = ~decrypt_pad & ~\u1_uk_K_r11_reg[3]/NET0131  ;
  assign n32985 = ~n32983 & ~n32984 ;
  assign n32986 = \u1_R11_reg[9]/NET0131  & ~n32985 ;
  assign n32987 = ~\u1_R11_reg[9]/NET0131  & n32985 ;
  assign n32988 = ~n32986 & ~n32987 ;
  assign n33010 = n32975 & ~n32988 ;
  assign n32989 = decrypt_pad & ~\u1_uk_K_r11_reg[48]/NET0131  ;
  assign n32990 = ~decrypt_pad & ~\u1_uk_K_r11_reg[11]/NET0131  ;
  assign n32991 = ~n32989 & ~n32990 ;
  assign n32992 = \u1_R11_reg[10]/NET0131  & ~n32991 ;
  assign n32993 = ~\u1_R11_reg[10]/NET0131  & n32991 ;
  assign n32994 = ~n32992 & ~n32993 ;
  assign n32976 = decrypt_pad & ~\u1_uk_K_r11_reg[11]/NET0131  ;
  assign n32977 = ~decrypt_pad & ~\u1_uk_K_r11_reg[6]/NET0131  ;
  assign n32978 = ~n32976 & ~n32977 ;
  assign n32979 = \u1_R11_reg[8]/NET0131  & ~n32978 ;
  assign n32980 = ~\u1_R11_reg[8]/NET0131  & n32978 ;
  assign n32981 = ~n32979 & ~n32980 ;
  assign n33012 = n32975 & ~n32981 ;
  assign n33013 = n32994 & n33012 ;
  assign n33014 = ~n32975 & n32988 ;
  assign n33015 = n32981 & n33014 ;
  assign n33016 = ~n33013 & ~n33015 ;
  assign n33017 = ~n33010 & n33016 ;
  assign n33018 = n33001 & ~n33017 ;
  assign n33011 = n32994 & n33010 ;
  assign n32982 = ~n32975 & ~n32981 ;
  assign n33019 = n32982 & ~n32988 ;
  assign n33020 = ~n32994 & n33019 ;
  assign n33021 = ~n33011 & ~n33020 ;
  assign n33022 = ~n33018 & n33021 ;
  assign n33023 = n33009 & ~n33022 ;
  assign n32995 = n32988 & n32994 ;
  assign n33032 = ~n32988 & ~n32994 ;
  assign n33033 = ~n32995 & ~n33032 ;
  assign n33030 = n32975 & n32981 ;
  assign n33031 = ~n32982 & ~n33030 ;
  assign n33034 = ~n32981 & n33009 ;
  assign n33038 = n33031 & ~n33034 ;
  assign n33039 = ~n33033 & ~n33038 ;
  assign n33035 = n32988 & n33034 ;
  assign n33036 = n33031 & n33033 ;
  assign n33037 = ~n33035 & n33036 ;
  assign n33040 = ~n33001 & ~n33037 ;
  assign n33041 = ~n33039 & n33040 ;
  assign n33002 = n32995 & n33001 ;
  assign n33003 = n32982 & n33002 ;
  assign n33026 = ~n33009 & ~n33014 ;
  assign n33024 = n32988 & ~n32994 ;
  assign n33025 = ~n32981 & ~n33024 ;
  assign n33027 = n33001 & ~n33010 ;
  assign n33028 = ~n33025 & n33027 ;
  assign n33029 = n33026 & n33028 ;
  assign n33042 = ~n33003 & ~n33029 ;
  assign n33043 = ~n33041 & n33042 ;
  assign n33044 = ~n33023 & n33043 ;
  assign n33045 = ~\u1_L11_reg[6]/NET0131  & ~n33044 ;
  assign n33046 = \u1_L11_reg[6]/NET0131  & n33044 ;
  assign n33047 = ~n33045 & ~n33046 ;
  assign n33049 = n31982 & n32922 ;
  assign n33059 = n31967 & n33049 ;
  assign n33053 = ~n31967 & ~n32922 ;
  assign n33048 = ~n31982 & n32921 ;
  assign n33060 = n31976 & ~n33048 ;
  assign n33061 = ~n33053 & n33060 ;
  assign n33062 = ~n33059 & n33061 ;
  assign n33063 = ~n32014 & ~n33062 ;
  assign n33054 = ~n31991 & n33053 ;
  assign n33064 = n31976 & ~n33054 ;
  assign n33065 = ~n32432 & n32913 ;
  assign n33066 = ~n33049 & n33065 ;
  assign n33067 = ~n33064 & ~n33066 ;
  assign n33050 = ~n33048 & ~n33049 ;
  assign n33051 = n31967 & ~n33050 ;
  assign n33068 = n32014 & ~n33051 ;
  assign n33069 = ~n33067 & n33068 ;
  assign n33070 = ~n33063 & ~n33069 ;
  assign n33052 = ~n31976 & n33051 ;
  assign n33055 = ~n31976 & n33054 ;
  assign n33056 = ~n32029 & ~n33055 ;
  assign n33057 = ~n31976 & n32014 ;
  assign n33058 = ~n33056 & ~n33057 ;
  assign n33071 = ~n33052 & ~n33058 ;
  assign n33072 = ~n33070 & n33071 ;
  assign n33073 = ~\u1_L11_reg[7]/NET0131  & ~n33072 ;
  assign n33074 = \u1_L11_reg[7]/NET0131  & n33072 ;
  assign n33075 = ~n33073 & ~n33074 ;
  assign n33093 = n31781 & n32637 ;
  assign n33077 = ~n31841 & ~n31843 ;
  assign n33078 = ~n31817 & ~n33077 ;
  assign n33092 = n31798 & n33078 ;
  assign n33082 = ~n31788 & n31828 ;
  assign n33094 = n31774 & n33082 ;
  assign n33095 = ~n33092 & ~n33094 ;
  assign n33096 = ~n33093 & n33095 ;
  assign n33097 = n31813 & ~n33096 ;
  assign n33083 = n31768 & n33077 ;
  assign n33084 = ~n33082 & n33083 ;
  assign n33079 = ~n31768 & n33078 ;
  assign n33076 = n31846 & ~n32634 ;
  assign n33080 = ~n31781 & n31843 ;
  assign n33081 = n31796 & n33080 ;
  assign n33085 = ~n33076 & ~n33081 ;
  assign n33086 = ~n33079 & n33085 ;
  assign n33087 = ~n33084 & n33086 ;
  assign n33088 = ~n31813 & ~n33087 ;
  assign n33089 = ~n31796 & n31844 ;
  assign n33090 = ~n33081 & ~n33089 ;
  assign n33091 = ~n31768 & ~n33090 ;
  assign n33098 = ~n33088 & ~n33091 ;
  assign n33099 = ~n33097 & n33098 ;
  assign n33100 = ~\u1_L11_reg[9]/NET0131  & ~n33099 ;
  assign n33101 = \u1_L11_reg[9]/NET0131  & n33099 ;
  assign n33102 = ~n33100 & ~n33101 ;
  assign n33103 = n32988 & n33030 ;
  assign n33104 = ~n32988 & ~n33030 ;
  assign n33105 = ~n33103 & ~n33104 ;
  assign n33106 = ~n32982 & ~n33105 ;
  assign n33107 = n33014 & n33034 ;
  assign n33108 = ~n33106 & ~n33107 ;
  assign n33109 = ~n32994 & ~n33108 ;
  assign n33110 = n32982 & n32994 ;
  assign n33111 = ~n32975 & n32981 ;
  assign n33112 = ~n32994 & n33111 ;
  assign n33113 = ~n33110 & ~n33112 ;
  assign n33114 = ~n33009 & ~n33113 ;
  assign n33115 = n32995 & n33012 ;
  assign n33116 = n33001 & ~n33115 ;
  assign n33117 = ~n33114 & n33116 ;
  assign n33118 = ~n33109 & n33117 ;
  assign n33120 = n32982 & ~n32994 ;
  assign n33119 = ~n32988 & n33012 ;
  assign n33121 = ~n33103 & ~n33119 ;
  assign n33122 = ~n33120 & n33121 ;
  assign n33123 = ~n33009 & ~n33122 ;
  assign n33124 = ~n32982 & n33009 ;
  assign n33125 = n33105 & n33124 ;
  assign n33126 = ~n33001 & ~n33020 ;
  assign n33127 = ~n33125 & n33126 ;
  assign n33128 = ~n33123 & n33127 ;
  assign n33129 = ~n33118 & ~n33128 ;
  assign n33130 = ~n33015 & ~n33019 ;
  assign n33131 = n32994 & ~n33130 ;
  assign n33132 = n33009 & ~n33131 ;
  assign n33133 = n32981 & n32994 ;
  assign n33134 = ~n32988 & n33133 ;
  assign n33135 = ~n33009 & ~n33134 ;
  assign n33136 = ~n33132 & ~n33135 ;
  assign n33137 = ~n33129 & ~n33136 ;
  assign n33138 = ~\u1_L11_reg[16]/NET0131  & ~n33137 ;
  assign n33139 = \u1_L11_reg[16]/NET0131  & n33137 ;
  assign n33140 = ~n33138 & ~n33139 ;
  assign n33143 = n33031 & ~n33032 ;
  assign n33144 = ~n33031 & n33032 ;
  assign n33145 = ~n33143 & ~n33144 ;
  assign n33146 = n33001 & ~n33145 ;
  assign n33147 = ~n33001 & n33016 ;
  assign n33148 = ~n33144 & n33147 ;
  assign n33149 = ~n33146 & ~n33148 ;
  assign n33150 = ~n33009 & ~n33149 ;
  assign n33154 = ~n33012 & n33032 ;
  assign n33153 = n32988 & n33133 ;
  assign n33155 = ~n33013 & ~n33153 ;
  assign n33156 = ~n33154 & n33155 ;
  assign n33157 = n33001 & ~n33156 ;
  assign n33151 = ~n32994 & n33012 ;
  assign n33152 = n32988 & n33151 ;
  assign n33158 = ~n32988 & n33112 ;
  assign n33159 = n33009 & ~n33158 ;
  assign n33160 = ~n33152 & n33159 ;
  assign n33161 = ~n33157 & n33160 ;
  assign n33162 = ~n33150 & ~n33161 ;
  assign n33141 = n32994 & ~n33009 ;
  assign n33142 = n33103 & n33141 ;
  assign n33163 = ~n32975 & n33134 ;
  assign n33164 = ~n33110 & ~n33151 ;
  assign n33165 = n32982 & n32988 ;
  assign n33166 = ~n33134 & ~n33165 ;
  assign n33167 = n33164 & n33166 ;
  assign n33168 = n33009 & ~n33167 ;
  assign n33169 = ~n33163 & ~n33168 ;
  assign n33170 = ~n33001 & ~n33169 ;
  assign n33171 = ~n33142 & ~n33170 ;
  assign n33172 = ~n33162 & n33171 ;
  assign n33173 = ~\u1_L11_reg[24]/NET0131  & ~n33172 ;
  assign n33174 = \u1_L11_reg[24]/NET0131  & n33172 ;
  assign n33175 = ~n33173 & ~n33174 ;
  assign n33178 = n33159 & n33164 ;
  assign n33179 = ~n33009 & ~n33133 ;
  assign n33180 = ~n33165 & n33179 ;
  assign n33181 = ~n33178 & ~n33180 ;
  assign n33182 = n33001 & ~n33181 ;
  assign n33183 = ~n32994 & ~n33119 ;
  assign n33184 = ~n33013 & ~n33183 ;
  assign n33185 = ~n32988 & ~n33111 ;
  assign n33186 = ~n33026 & ~n33185 ;
  assign n33187 = ~n33184 & ~n33186 ;
  assign n33188 = ~n33014 & n33133 ;
  assign n33189 = ~n32975 & n33024 ;
  assign n33190 = ~n33188 & ~n33189 ;
  assign n33191 = n33009 & ~n33190 ;
  assign n33192 = ~n33001 & ~n33191 ;
  assign n33193 = ~n33187 & n33192 ;
  assign n33194 = ~n33182 & ~n33193 ;
  assign n33195 = n33009 & n33010 ;
  assign n33196 = n33133 & n33195 ;
  assign n33176 = n33002 & ~n33030 ;
  assign n33177 = n33014 & n33141 ;
  assign n33197 = ~n33176 & ~n33177 ;
  assign n33198 = ~n33196 & n33197 ;
  assign n33199 = ~n33194 & n33198 ;
  assign n33200 = \u1_L11_reg[30]/NET0131  & ~n33199 ;
  assign n33201 = ~\u1_L11_reg[30]/NET0131  & n33199 ;
  assign n33202 = ~n33200 & ~n33201 ;
  assign n33218 = ~n32455 & ~n32475 ;
  assign n33214 = ~n32321 & ~n32374 ;
  assign n33215 = n32363 & ~n33214 ;
  assign n33216 = ~n32327 & ~n32374 ;
  assign n33217 = n32383 & n33216 ;
  assign n33219 = ~n33215 & ~n33217 ;
  assign n33220 = n33218 & n33219 ;
  assign n33221 = ~n32357 & ~n33220 ;
  assign n33203 = n32302 & ~n32337 ;
  assign n33204 = ~n32343 & ~n32474 ;
  assign n33205 = ~n32302 & n32327 ;
  assign n33206 = ~n33204 & n33205 ;
  assign n33207 = ~n32329 & ~n33206 ;
  assign n33208 = ~n33203 & n33207 ;
  assign n33209 = n32357 & ~n33208 ;
  assign n33210 = n32314 & n32363 ;
  assign n33211 = n32302 & ~n32482 ;
  assign n33212 = ~n33210 & n33211 ;
  assign n33213 = ~n32751 & ~n33212 ;
  assign n33222 = ~n33209 & ~n33213 ;
  assign n33223 = ~n33221 & n33222 ;
  assign n33224 = \u1_L11_reg[18]/P0001  & n33223 ;
  assign n33225 = ~\u1_L11_reg[18]/P0001  & ~n33223 ;
  assign n33226 = ~n33224 & ~n33225 ;
  assign n33227 = decrypt_pad & ~\u1_uk_K_r10_reg[45]/P0001  ;
  assign n33228 = ~decrypt_pad & ~\u1_uk_K_r10_reg[36]/NET0131  ;
  assign n33229 = ~n33227 & ~n33228 ;
  assign n33230 = \u1_R10_reg[28]/NET0131  & ~n33229 ;
  assign n33231 = ~\u1_R10_reg[28]/NET0131  & n33229 ;
  assign n33232 = ~n33230 & ~n33231 ;
  assign n33233 = decrypt_pad & ~\u1_uk_K_r10_reg[21]/NET0131  ;
  assign n33234 = ~decrypt_pad & ~\u1_uk_K_r10_reg[16]/NET0131  ;
  assign n33235 = ~n33233 & ~n33234 ;
  assign n33236 = \u1_R10_reg[26]/NET0131  & ~n33235 ;
  assign n33237 = ~\u1_R10_reg[26]/NET0131  & n33235 ;
  assign n33238 = ~n33236 & ~n33237 ;
  assign n33239 = decrypt_pad & ~\u1_uk_K_r10_reg[36]/NET0131  ;
  assign n33240 = ~decrypt_pad & ~\u1_uk_K_r10_reg[0]/NET0131  ;
  assign n33241 = ~n33239 & ~n33240 ;
  assign n33242 = \u1_R10_reg[25]/NET0131  & ~n33241 ;
  assign n33243 = ~\u1_R10_reg[25]/NET0131  & n33241 ;
  assign n33244 = ~n33242 & ~n33243 ;
  assign n33273 = ~n33238 & ~n33244 ;
  assign n33245 = decrypt_pad & ~\u1_uk_K_r10_reg[9]/NET0131  ;
  assign n33246 = ~decrypt_pad & ~\u1_uk_K_r10_reg[28]/NET0131  ;
  assign n33247 = ~n33245 & ~n33246 ;
  assign n33248 = \u1_R10_reg[29]/NET0131  & ~n33247 ;
  assign n33249 = ~\u1_R10_reg[29]/NET0131  & n33247 ;
  assign n33250 = ~n33248 & ~n33249 ;
  assign n33276 = ~n33238 & ~n33250 ;
  assign n33296 = ~n33273 & ~n33276 ;
  assign n33252 = decrypt_pad & ~\u1_uk_K_r10_reg[1]/NET0131  ;
  assign n33253 = ~decrypt_pad & ~\u1_uk_K_r10_reg[51]/NET0131  ;
  assign n33254 = ~n33252 & ~n33253 ;
  assign n33255 = \u1_R10_reg[24]/NET0131  & ~n33254 ;
  assign n33256 = ~\u1_R10_reg[24]/NET0131  & n33254 ;
  assign n33257 = ~n33255 & ~n33256 ;
  assign n33260 = decrypt_pad & ~\u1_uk_K_r10_reg[30]/NET0131  ;
  assign n33261 = ~decrypt_pad & ~\u1_uk_K_r10_reg[49]/NET0131  ;
  assign n33262 = ~n33260 & ~n33261 ;
  assign n33263 = \u1_R10_reg[27]/NET0131  & ~n33262 ;
  assign n33264 = ~\u1_R10_reg[27]/NET0131  & n33262 ;
  assign n33265 = ~n33263 & ~n33264 ;
  assign n33275 = n33238 & n33244 ;
  assign n33295 = n33265 & ~n33275 ;
  assign n33297 = n33257 & n33295 ;
  assign n33298 = n33296 & n33297 ;
  assign n33289 = n33250 & n33257 ;
  assign n33290 = n33273 & n33289 ;
  assign n33291 = n33244 & n33250 ;
  assign n33292 = ~n33257 & n33291 ;
  assign n33293 = ~n33290 & ~n33292 ;
  assign n33294 = ~n33265 & ~n33293 ;
  assign n33284 = ~n33250 & ~n33257 ;
  assign n33285 = n33273 & n33284 ;
  assign n33286 = n33250 & ~n33257 ;
  assign n33287 = n33238 & ~n33244 ;
  assign n33288 = n33286 & n33287 ;
  assign n33299 = ~n33285 & ~n33288 ;
  assign n33300 = ~n33294 & n33299 ;
  assign n33301 = ~n33298 & n33300 ;
  assign n33302 = n33232 & ~n33301 ;
  assign n33277 = ~n33265 & ~n33275 ;
  assign n33278 = ~n33276 & n33277 ;
  assign n33274 = n33265 & ~n33273 ;
  assign n33279 = n33257 & ~n33274 ;
  assign n33280 = ~n33278 & n33279 ;
  assign n33251 = ~n33244 & ~n33250 ;
  assign n33258 = n33251 & ~n33257 ;
  assign n33259 = n33238 & n33258 ;
  assign n33266 = n33259 & ~n33265 ;
  assign n33267 = ~n33238 & ~n33257 ;
  assign n33268 = n33238 & n33257 ;
  assign n33269 = ~n33267 & ~n33268 ;
  assign n33270 = ~n33244 & n33265 ;
  assign n33271 = n33250 & ~n33270 ;
  assign n33272 = ~n33269 & n33271 ;
  assign n33281 = ~n33266 & ~n33272 ;
  assign n33282 = ~n33280 & n33281 ;
  assign n33283 = ~n33232 & ~n33282 ;
  assign n33305 = n33275 & n33284 ;
  assign n33306 = ~n33288 & ~n33305 ;
  assign n33307 = ~n33250 & n33257 ;
  assign n33308 = ~n33244 & n33307 ;
  assign n33309 = n33306 & ~n33308 ;
  assign n33310 = n33265 & ~n33309 ;
  assign n33303 = n33244 & ~n33265 ;
  assign n33304 = ~n33269 & n33303 ;
  assign n33311 = n33270 & n33276 ;
  assign n33312 = ~n33304 & ~n33311 ;
  assign n33313 = ~n33310 & n33312 ;
  assign n33314 = ~n33283 & n33313 ;
  assign n33315 = ~n33302 & n33314 ;
  assign n33316 = ~\u1_L10_reg[22]/NET0131  & ~n33315 ;
  assign n33317 = \u1_L10_reg[22]/NET0131  & n33315 ;
  assign n33318 = ~n33316 & ~n33317 ;
  assign n33338 = decrypt_pad & ~\u1_uk_K_r10_reg[4]/NET0131  ;
  assign n33339 = ~decrypt_pad & ~\u1_uk_K_r10_reg[27]/NET0131  ;
  assign n33340 = ~n33338 & ~n33339 ;
  assign n33341 = \u1_R10_reg[3]/NET0131  & ~n33340 ;
  assign n33342 = ~\u1_R10_reg[3]/NET0131  & n33340 ;
  assign n33343 = ~n33341 & ~n33342 ;
  assign n33325 = decrypt_pad & ~\u1_uk_K_r10_reg[12]/NET0131  ;
  assign n33326 = ~decrypt_pad & ~\u1_uk_K_r10_reg[3]/NET0131  ;
  assign n33327 = ~n33325 & ~n33326 ;
  assign n33328 = \u1_R10_reg[1]/NET0131  & ~n33327 ;
  assign n33329 = ~\u1_R10_reg[1]/NET0131  & n33327 ;
  assign n33330 = ~n33328 & ~n33329 ;
  assign n33344 = decrypt_pad & ~\u1_uk_K_r10_reg[48]/NET0131  ;
  assign n33345 = ~decrypt_pad & ~\u1_uk_K_r10_reg[39]/NET0131  ;
  assign n33346 = ~n33344 & ~n33345 ;
  assign n33347 = \u1_R10_reg[32]/NET0131  & ~n33346 ;
  assign n33348 = ~\u1_R10_reg[32]/NET0131  & n33346 ;
  assign n33349 = ~n33347 & ~n33348 ;
  assign n33362 = n33330 & n33349 ;
  assign n33319 = decrypt_pad & ~\u1_uk_K_r10_reg[10]/NET0131  ;
  assign n33320 = ~decrypt_pad & ~\u1_uk_K_r10_reg[33]/NET0131  ;
  assign n33321 = ~n33319 & ~n33320 ;
  assign n33322 = \u1_R10_reg[5]/NET0131  & ~n33321 ;
  assign n33323 = ~\u1_R10_reg[5]/NET0131  & n33321 ;
  assign n33324 = ~n33322 & ~n33323 ;
  assign n33331 = decrypt_pad & ~\u1_uk_K_r10_reg[27]/NET0131  ;
  assign n33332 = ~decrypt_pad & ~\u1_uk_K_r10_reg[18]/NET0131  ;
  assign n33333 = ~n33331 & ~n33332 ;
  assign n33334 = \u1_R10_reg[2]/NET0131  & ~n33333 ;
  assign n33335 = ~\u1_R10_reg[2]/NET0131  & n33333 ;
  assign n33336 = ~n33334 & ~n33335 ;
  assign n33384 = ~n33324 & n33336 ;
  assign n33385 = n33362 & n33384 ;
  assign n33386 = n33343 & n33385 ;
  assign n33363 = decrypt_pad & ~\u1_uk_K_r10_reg[39]/NET0131  ;
  assign n33364 = ~decrypt_pad & ~\u1_uk_K_r10_reg[5]/NET0131  ;
  assign n33365 = ~n33363 & ~n33364 ;
  assign n33366 = \u1_R10_reg[4]/NET0131  & ~n33365 ;
  assign n33367 = ~\u1_R10_reg[4]/NET0131  & n33365 ;
  assign n33368 = ~n33366 & ~n33367 ;
  assign n33356 = n33336 & ~n33349 ;
  assign n33376 = n33324 & n33343 ;
  assign n33377 = n33356 & n33376 ;
  assign n33378 = n33330 & n33377 ;
  assign n33393 = ~n33368 & ~n33378 ;
  assign n33394 = ~n33386 & n33393 ;
  assign n33380 = ~n33336 & n33349 ;
  assign n33381 = ~n33356 & ~n33380 ;
  assign n33357 = n33324 & ~n33330 ;
  assign n33379 = ~n33343 & ~n33362 ;
  assign n33382 = ~n33357 & n33379 ;
  assign n33383 = n33381 & n33382 ;
  assign n33359 = n33324 & n33349 ;
  assign n33387 = n33330 & ~n33343 ;
  assign n33388 = n33359 & ~n33387 ;
  assign n33389 = ~n33324 & ~n33349 ;
  assign n33390 = n33330 & n33389 ;
  assign n33391 = ~n33388 & ~n33390 ;
  assign n33392 = ~n33336 & ~n33391 ;
  assign n33395 = ~n33383 & ~n33392 ;
  assign n33396 = n33394 & n33395 ;
  assign n33401 = ~n33324 & n33380 ;
  assign n33400 = n33324 & ~n33349 ;
  assign n33402 = ~n33356 & ~n33376 ;
  assign n33403 = ~n33400 & n33402 ;
  assign n33404 = ~n33401 & n33403 ;
  assign n33405 = ~n33330 & ~n33404 ;
  assign n33350 = n33343 & ~n33349 ;
  assign n33397 = n33324 & ~n33336 ;
  assign n33398 = ~n33384 & ~n33397 ;
  assign n33399 = n33350 & ~n33398 ;
  assign n33406 = n33368 & ~n33399 ;
  assign n33407 = ~n33405 & n33406 ;
  assign n33408 = ~n33396 & ~n33407 ;
  assign n33360 = n33336 & n33359 ;
  assign n33361 = n33330 & n33360 ;
  assign n33370 = ~n33324 & n33330 ;
  assign n33371 = ~n33336 & n33370 ;
  assign n33358 = n33356 & n33357 ;
  assign n33369 = n33362 & n33368 ;
  assign n33372 = ~n33358 & ~n33369 ;
  assign n33373 = ~n33371 & n33372 ;
  assign n33374 = ~n33361 & n33373 ;
  assign n33375 = ~n33343 & ~n33374 ;
  assign n33337 = ~n33330 & n33336 ;
  assign n33351 = ~n33324 & n33337 ;
  assign n33352 = n33350 & n33351 ;
  assign n33353 = ~n33330 & ~n33336 ;
  assign n33354 = n33343 & n33349 ;
  assign n33355 = n33353 & n33354 ;
  assign n33409 = ~n33352 & ~n33355 ;
  assign n33410 = ~n33375 & n33409 ;
  assign n33411 = ~n33408 & n33410 ;
  assign n33412 = ~\u1_L10_reg[31]/NET0131  & ~n33411 ;
  assign n33413 = \u1_L10_reg[31]/NET0131  & n33411 ;
  assign n33414 = ~n33412 & ~n33413 ;
  assign n33415 = decrypt_pad & ~\u1_uk_K_r10_reg[38]/NET0131  ;
  assign n33416 = ~decrypt_pad & ~\u1_uk_K_r10_reg[29]/NET0131  ;
  assign n33417 = ~n33415 & ~n33416 ;
  assign n33418 = \u1_R10_reg[24]/NET0131  & ~n33417 ;
  assign n33419 = ~\u1_R10_reg[24]/NET0131  & n33417 ;
  assign n33420 = ~n33418 & ~n33419 ;
  assign n33434 = decrypt_pad & ~\u1_uk_K_r10_reg[50]/NET0131  ;
  assign n33435 = ~decrypt_pad & ~\u1_uk_K_r10_reg[14]/NET0131  ;
  assign n33436 = ~n33434 & ~n33435 ;
  assign n33437 = \u1_R10_reg[22]/NET0131  & ~n33436 ;
  assign n33438 = ~\u1_R10_reg[22]/NET0131  & n33436 ;
  assign n33439 = ~n33437 & ~n33438 ;
  assign n33421 = decrypt_pad & ~\u1_uk_K_r10_reg[28]/NET0131  ;
  assign n33422 = ~decrypt_pad & ~\u1_uk_K_r10_reg[23]/NET0131  ;
  assign n33423 = ~n33421 & ~n33422 ;
  assign n33424 = \u1_R10_reg[21]/NET0131  & ~n33423 ;
  assign n33425 = ~\u1_R10_reg[21]/NET0131  & n33423 ;
  assign n33426 = ~n33424 & ~n33425 ;
  assign n33427 = decrypt_pad & ~\u1_uk_K_r10_reg[44]/NET0131  ;
  assign n33428 = ~decrypt_pad & ~\u1_uk_K_r10_reg[8]/NET0131  ;
  assign n33429 = ~n33427 & ~n33428 ;
  assign n33430 = \u1_R10_reg[20]/NET0131  & ~n33429 ;
  assign n33431 = ~\u1_R10_reg[20]/NET0131  & n33429 ;
  assign n33432 = ~n33430 & ~n33431 ;
  assign n33433 = n33426 & ~n33432 ;
  assign n33451 = decrypt_pad & ~\u1_uk_K_r10_reg[29]/NET0131  ;
  assign n33452 = ~decrypt_pad & ~\u1_uk_K_r10_reg[52]/NET0131  ;
  assign n33453 = ~n33451 & ~n33452 ;
  assign n33454 = \u1_R10_reg[25]/NET0131  & ~n33453 ;
  assign n33455 = ~\u1_R10_reg[25]/NET0131  & n33453 ;
  assign n33456 = ~n33454 & ~n33455 ;
  assign n33461 = n33432 & n33456 ;
  assign n33499 = ~n33433 & ~n33461 ;
  assign n33500 = n33439 & ~n33499 ;
  assign n33444 = decrypt_pad & ~\u1_uk_K_r10_reg[8]/NET0131  ;
  assign n33445 = ~decrypt_pad & ~\u1_uk_K_r10_reg[31]/NET0131  ;
  assign n33446 = ~n33444 & ~n33445 ;
  assign n33447 = \u1_R10_reg[23]/NET0131  & ~n33446 ;
  assign n33448 = ~\u1_R10_reg[23]/NET0131  & n33446 ;
  assign n33449 = ~n33447 & ~n33448 ;
  assign n33480 = ~n33432 & n33456 ;
  assign n33497 = n33426 & n33480 ;
  assign n33498 = ~n33439 & ~n33497 ;
  assign n33501 = ~n33449 & ~n33498 ;
  assign n33502 = ~n33500 & n33501 ;
  assign n33491 = n33426 & n33461 ;
  assign n33440 = n33433 & n33439 ;
  assign n33457 = n33432 & ~n33456 ;
  assign n33479 = ~n33426 & ~n33439 ;
  assign n33490 = n33457 & n33479 ;
  assign n33492 = ~n33440 & ~n33490 ;
  assign n33493 = ~n33491 & n33492 ;
  assign n33494 = n33449 & ~n33493 ;
  assign n33458 = ~n33439 & ~n33449 ;
  assign n33495 = n33458 & n33461 ;
  assign n33496 = ~n33426 & n33495 ;
  assign n33503 = ~n33494 & ~n33496 ;
  assign n33504 = ~n33502 & n33503 ;
  assign n33505 = n33420 & ~n33504 ;
  assign n33462 = ~n33426 & n33439 ;
  assign n33466 = ~n33432 & ~n33456 ;
  assign n33467 = n33462 & n33466 ;
  assign n33464 = ~n33432 & ~n33439 ;
  assign n33465 = ~n33462 & ~n33464 ;
  assign n33468 = n33449 & ~n33465 ;
  assign n33469 = ~n33467 & n33468 ;
  assign n33441 = n33426 & ~n33439 ;
  assign n33442 = n33432 & n33441 ;
  assign n33443 = ~n33440 & ~n33442 ;
  assign n33450 = ~n33443 & ~n33449 ;
  assign n33459 = ~n33441 & ~n33458 ;
  assign n33460 = n33457 & ~n33459 ;
  assign n33463 = n33461 & n33462 ;
  assign n33470 = ~n33460 & ~n33463 ;
  assign n33471 = ~n33450 & n33470 ;
  assign n33472 = ~n33469 & n33471 ;
  assign n33473 = ~n33420 & ~n33472 ;
  assign n33481 = n33449 & n33480 ;
  assign n33482 = n33479 & n33481 ;
  assign n33483 = n33432 & ~n33449 ;
  assign n33484 = ~n33439 & ~n33456 ;
  assign n33485 = n33426 & n33484 ;
  assign n33486 = n33483 & n33485 ;
  assign n33487 = ~n33482 & ~n33486 ;
  assign n33474 = n33426 & n33466 ;
  assign n33475 = ~n33439 & ~n33474 ;
  assign n33476 = n33439 & ~n33461 ;
  assign n33477 = n33449 & ~n33476 ;
  assign n33478 = ~n33475 & n33477 ;
  assign n33488 = ~n33426 & n33466 ;
  assign n33489 = n33458 & n33488 ;
  assign n33506 = ~n33478 & ~n33489 ;
  assign n33507 = n33487 & n33506 ;
  assign n33508 = ~n33473 & n33507 ;
  assign n33509 = ~n33505 & n33508 ;
  assign n33510 = \u1_L10_reg[11]/NET0131  & ~n33509 ;
  assign n33511 = ~\u1_L10_reg[11]/NET0131  & n33509 ;
  assign n33512 = ~n33510 & ~n33511 ;
  assign n33525 = decrypt_pad & ~\u1_uk_K_r10_reg[24]/NET0131  ;
  assign n33526 = ~decrypt_pad & ~\u1_uk_K_r10_reg[47]/NET0131  ;
  assign n33527 = ~n33525 & ~n33526 ;
  assign n33528 = \u1_R10_reg[13]/NET0131  & ~n33527 ;
  assign n33529 = ~\u1_R10_reg[13]/NET0131  & n33527 ;
  assign n33530 = ~n33528 & ~n33529 ;
  assign n33519 = decrypt_pad & ~\u1_uk_K_r10_reg[5]/NET0131  ;
  assign n33520 = ~decrypt_pad & ~\u1_uk_K_r10_reg[53]/NET0131  ;
  assign n33521 = ~n33519 & ~n33520 ;
  assign n33522 = \u1_R10_reg[12]/NET0131  & ~n33521 ;
  assign n33523 = ~\u1_R10_reg[12]/NET0131  & n33521 ;
  assign n33524 = ~n33522 & ~n33523 ;
  assign n33538 = decrypt_pad & ~\u1_uk_K_r10_reg[46]/NET0131  ;
  assign n33539 = ~decrypt_pad & ~\u1_uk_K_r10_reg[12]/NET0131  ;
  assign n33540 = ~n33538 & ~n33539 ;
  assign n33541 = \u1_R10_reg[17]/NET0131  & ~n33540 ;
  assign n33542 = ~\u1_R10_reg[17]/NET0131  & n33540 ;
  assign n33543 = ~n33541 & ~n33542 ;
  assign n33568 = n33524 & n33543 ;
  assign n33569 = n33530 & n33568 ;
  assign n33513 = decrypt_pad & ~\u1_uk_K_r10_reg[33]/NET0131  ;
  assign n33514 = ~decrypt_pad & ~\u1_uk_K_r10_reg[24]/NET0131  ;
  assign n33515 = ~n33513 & ~n33514 ;
  assign n33516 = \u1_R10_reg[15]/NET0131  & ~n33515 ;
  assign n33517 = ~\u1_R10_reg[15]/NET0131  & n33515 ;
  assign n33518 = ~n33516 & ~n33517 ;
  assign n33551 = ~n33530 & ~n33543 ;
  assign n33552 = ~n33524 & n33551 ;
  assign n33570 = n33518 & ~n33552 ;
  assign n33571 = ~n33569 & n33570 ;
  assign n33532 = decrypt_pad & ~\u1_uk_K_r10_reg[25]/NET0131  ;
  assign n33533 = ~decrypt_pad & ~\u1_uk_K_r10_reg[48]/NET0131  ;
  assign n33534 = ~n33532 & ~n33533 ;
  assign n33535 = \u1_R10_reg[14]/NET0131  & ~n33534 ;
  assign n33536 = ~\u1_R10_reg[14]/NET0131  & n33534 ;
  assign n33537 = ~n33535 & ~n33536 ;
  assign n33547 = n33524 & ~n33543 ;
  assign n33573 = n33537 & n33547 ;
  assign n33572 = ~n33530 & n33543 ;
  assign n33574 = ~n33518 & ~n33572 ;
  assign n33575 = ~n33573 & n33574 ;
  assign n33576 = ~n33571 & ~n33575 ;
  assign n33553 = ~n33537 & n33552 ;
  assign n33531 = ~n33524 & n33530 ;
  assign n33559 = n33531 & ~n33543 ;
  assign n33560 = n33537 & n33559 ;
  assign n33561 = ~n33553 & ~n33560 ;
  assign n33556 = n33518 & n33530 ;
  assign n33577 = n33537 & n33556 ;
  assign n33578 = ~n33524 & n33577 ;
  assign n33562 = decrypt_pad & ~\u1_uk_K_r10_reg[41]/P0001  ;
  assign n33563 = ~decrypt_pad & ~\u1_uk_K_r10_reg[32]/NET0131  ;
  assign n33564 = ~n33562 & ~n33563 ;
  assign n33565 = \u1_R10_reg[16]/NET0131  & ~n33564 ;
  assign n33566 = ~\u1_R10_reg[16]/NET0131  & n33564 ;
  assign n33567 = ~n33565 & ~n33566 ;
  assign n33544 = ~n33537 & n33543 ;
  assign n33579 = n33524 & ~n33530 ;
  assign n33580 = n33544 & n33579 ;
  assign n33581 = ~n33567 & ~n33580 ;
  assign n33582 = ~n33578 & n33581 ;
  assign n33583 = n33561 & n33582 ;
  assign n33584 = ~n33576 & n33583 ;
  assign n33585 = ~n33524 & n33543 ;
  assign n33586 = n33518 & n33585 ;
  assign n33587 = ~n33530 & n33586 ;
  assign n33595 = n33567 & ~n33587 ;
  assign n33545 = n33531 & n33544 ;
  assign n33557 = n33547 & n33556 ;
  assign n33588 = ~n33545 & ~n33557 ;
  assign n33589 = n33537 & n33569 ;
  assign n33596 = n33588 & ~n33589 ;
  assign n33590 = ~n33531 & ~n33579 ;
  assign n33591 = ~n33518 & ~n33537 ;
  assign n33592 = ~n33590 & n33591 ;
  assign n33593 = ~n33518 & n33537 ;
  assign n33594 = n33552 & n33593 ;
  assign n33597 = ~n33592 & ~n33594 ;
  assign n33598 = n33596 & n33597 ;
  assign n33599 = n33595 & n33598 ;
  assign n33600 = ~n33584 & ~n33599 ;
  assign n33546 = ~n33518 & ~n33545 ;
  assign n33548 = ~n33530 & n33537 ;
  assign n33549 = n33547 & n33548 ;
  assign n33550 = n33518 & ~n33549 ;
  assign n33554 = n33550 & ~n33553 ;
  assign n33555 = ~n33546 & ~n33554 ;
  assign n33558 = ~n33537 & n33557 ;
  assign n33601 = ~n33555 & ~n33558 ;
  assign n33602 = ~n33600 & n33601 ;
  assign n33603 = ~\u1_L10_reg[20]/NET0131  & ~n33602 ;
  assign n33604 = \u1_L10_reg[20]/NET0131  & n33602 ;
  assign n33605 = ~n33603 & ~n33604 ;
  assign n33618 = n33548 & n33585 ;
  assign n33619 = ~n33589 & ~n33618 ;
  assign n33622 = n33518 & ~n33580 ;
  assign n33623 = ~n33559 & n33622 ;
  assign n33624 = n33530 & ~n33537 ;
  assign n33625 = n33547 & ~n33624 ;
  assign n33626 = n33546 & ~n33625 ;
  assign n33627 = ~n33623 & ~n33626 ;
  assign n33628 = n33619 & ~n33627 ;
  assign n33629 = n33567 & ~n33628 ;
  assign n33612 = n33518 & ~n33544 ;
  assign n33613 = n33579 & n33612 ;
  assign n33614 = n33561 & ~n33613 ;
  assign n33606 = n33524 & n33530 ;
  assign n33607 = ~n33586 & ~n33606 ;
  assign n33608 = ~n33537 & ~n33607 ;
  assign n33609 = n33524 & n33544 ;
  assign n33610 = ~n33552 & ~n33609 ;
  assign n33611 = ~n33518 & ~n33610 ;
  assign n33615 = ~n33608 & ~n33611 ;
  assign n33616 = n33614 & n33615 ;
  assign n33617 = ~n33567 & ~n33616 ;
  assign n33620 = ~n33553 & n33619 ;
  assign n33621 = ~n33518 & ~n33620 ;
  assign n33630 = ~n33558 & ~n33578 ;
  assign n33631 = ~n33621 & n33630 ;
  assign n33632 = ~n33617 & n33631 ;
  assign n33633 = ~n33629 & n33632 ;
  assign n33634 = ~\u1_L10_reg[10]/NET0131  & ~n33633 ;
  assign n33635 = \u1_L10_reg[10]/NET0131  & n33633 ;
  assign n33636 = ~n33634 & ~n33635 ;
  assign n33643 = ~n33273 & ~n33275 ;
  assign n33644 = n33284 & n33643 ;
  assign n33641 = ~n33270 & ~n33275 ;
  assign n33642 = n33286 & ~n33641 ;
  assign n33648 = ~n33232 & ~n33642 ;
  assign n33649 = ~n33644 & n33648 ;
  assign n33637 = n33257 & n33276 ;
  assign n33638 = n33250 & n33268 ;
  assign n33639 = ~n33637 & ~n33638 ;
  assign n33640 = ~n33244 & ~n33639 ;
  assign n33645 = ~n33251 & ~n33291 ;
  assign n33646 = ~n33268 & n33645 ;
  assign n33647 = ~n33265 & ~n33646 ;
  assign n33650 = ~n33640 & ~n33647 ;
  assign n33651 = n33649 & n33650 ;
  assign n33652 = ~n33265 & n33288 ;
  assign n33658 = n33232 & ~n33290 ;
  assign n33659 = ~n33305 & n33658 ;
  assign n33660 = ~n33652 & n33659 ;
  assign n33653 = ~n33267 & ~n33308 ;
  assign n33654 = n33296 & ~n33653 ;
  assign n33655 = n33244 & n33257 ;
  assign n33656 = ~n33285 & ~n33655 ;
  assign n33657 = n33265 & ~n33656 ;
  assign n33661 = ~n33654 & ~n33657 ;
  assign n33662 = n33660 & n33661 ;
  assign n33663 = ~n33651 & ~n33662 ;
  assign n33664 = \u1_L10_reg[12]/NET0131  & n33663 ;
  assign n33665 = ~\u1_L10_reg[12]/NET0131  & ~n33663 ;
  assign n33666 = ~n33664 & ~n33665 ;
  assign n33725 = decrypt_pad & ~\u1_uk_K_r10_reg[22]/NET0131  ;
  assign n33726 = ~decrypt_pad & ~\u1_uk_K_r10_reg[45]/P0001  ;
  assign n33727 = ~n33725 & ~n33726 ;
  assign n33728 = \u1_R10_reg[20]/NET0131  & ~n33727 ;
  assign n33729 = ~\u1_R10_reg[20]/NET0131  & n33727 ;
  assign n33730 = ~n33728 & ~n33729 ;
  assign n33695 = decrypt_pad & ~\u1_uk_K_r10_reg[7]/NET0131  ;
  assign n33696 = ~decrypt_pad & ~\u1_uk_K_r10_reg[2]/NET0131  ;
  assign n33697 = ~n33695 & ~n33696 ;
  assign n33698 = \u1_R10_reg[19]/NET0131  & ~n33697 ;
  assign n33699 = ~\u1_R10_reg[19]/NET0131  & n33697 ;
  assign n33700 = ~n33698 & ~n33699 ;
  assign n33687 = decrypt_pad & ~\u1_uk_K_r10_reg[2]/NET0131  ;
  assign n33688 = ~decrypt_pad & ~\u1_uk_K_r10_reg[21]/NET0131  ;
  assign n33689 = ~n33687 & ~n33688 ;
  assign n33690 = \u1_R10_reg[17]/NET0131  & ~n33689 ;
  assign n33691 = ~\u1_R10_reg[17]/NET0131  & n33689 ;
  assign n33692 = ~n33690 & ~n33691 ;
  assign n33673 = decrypt_pad & ~\u1_uk_K_r10_reg[35]/NET0131  ;
  assign n33674 = ~decrypt_pad & ~\u1_uk_K_r10_reg[30]/NET0131  ;
  assign n33675 = ~n33673 & ~n33674 ;
  assign n33676 = \u1_R10_reg[16]/NET0131  & ~n33675 ;
  assign n33677 = ~\u1_R10_reg[16]/NET0131  & n33675 ;
  assign n33678 = ~n33676 & ~n33677 ;
  assign n33680 = decrypt_pad & ~\u1_uk_K_r10_reg[23]/NET0131  ;
  assign n33681 = ~decrypt_pad & ~\u1_uk_K_r10_reg[42]/NET0131  ;
  assign n33682 = ~n33680 & ~n33681 ;
  assign n33683 = \u1_R10_reg[21]/NET0131  & ~n33682 ;
  assign n33684 = ~\u1_R10_reg[21]/NET0131  & n33682 ;
  assign n33685 = ~n33683 & ~n33684 ;
  assign n33732 = n33678 & ~n33685 ;
  assign n33733 = n33692 & n33732 ;
  assign n33667 = decrypt_pad & ~\u1_uk_K_r10_reg[51]/NET0131  ;
  assign n33668 = ~decrypt_pad & ~\u1_uk_K_r10_reg[15]/NET0131  ;
  assign n33669 = ~n33667 & ~n33668 ;
  assign n33670 = \u1_R10_reg[18]/NET0131  & ~n33669 ;
  assign n33671 = ~\u1_R10_reg[18]/NET0131  & n33669 ;
  assign n33672 = ~n33670 & ~n33671 ;
  assign n33693 = ~n33672 & n33692 ;
  assign n33694 = ~n33678 & n33693 ;
  assign n33679 = n33672 & n33678 ;
  assign n33734 = ~n33679 & n33685 ;
  assign n33735 = ~n33694 & n33734 ;
  assign n33736 = ~n33733 & ~n33735 ;
  assign n33737 = n33700 & ~n33736 ;
  assign n33701 = ~n33678 & ~n33685 ;
  assign n33702 = ~n33692 & n33701 ;
  assign n33714 = ~n33678 & n33685 ;
  assign n33740 = n33692 & n33714 ;
  assign n33741 = ~n33702 & ~n33740 ;
  assign n33742 = ~n33672 & ~n33700 ;
  assign n33743 = ~n33741 & n33742 ;
  assign n33711 = n33678 & n33685 ;
  assign n33712 = n33692 & n33711 ;
  assign n33744 = n33672 & ~n33700 ;
  assign n33745 = n33712 & n33744 ;
  assign n33738 = ~n33672 & n33711 ;
  assign n33739 = ~n33692 & n33738 ;
  assign n33746 = n33693 & n33732 ;
  assign n33747 = n33672 & ~n33692 ;
  assign n33748 = n33732 & n33747 ;
  assign n33749 = ~n33746 & ~n33748 ;
  assign n33750 = ~n33739 & n33749 ;
  assign n33751 = ~n33745 & n33750 ;
  assign n33752 = ~n33743 & n33751 ;
  assign n33753 = ~n33737 & n33752 ;
  assign n33754 = n33730 & ~n33753 ;
  assign n33686 = n33679 & n33685 ;
  assign n33703 = ~n33686 & n33700 ;
  assign n33704 = ~n33694 & ~n33702 ;
  assign n33705 = n33703 & n33704 ;
  assign n33715 = ~n33692 & n33714 ;
  assign n33706 = n33672 & n33692 ;
  assign n33707 = ~n33685 & n33706 ;
  assign n33716 = ~n33700 & ~n33707 ;
  assign n33717 = ~n33715 & n33716 ;
  assign n33708 = n33678 & ~n33692 ;
  assign n33709 = ~n33685 & n33708 ;
  assign n33710 = ~n33672 & n33709 ;
  assign n33713 = ~n33672 & n33712 ;
  assign n33718 = ~n33710 & ~n33713 ;
  assign n33719 = n33717 & n33718 ;
  assign n33720 = ~n33705 & ~n33719 ;
  assign n33721 = n33686 & ~n33692 ;
  assign n33722 = ~n33685 & n33694 ;
  assign n33723 = ~n33721 & ~n33722 ;
  assign n33724 = ~n33720 & n33723 ;
  assign n33731 = ~n33724 & ~n33730 ;
  assign n33755 = n33672 & n33702 ;
  assign n33756 = ~n33746 & ~n33755 ;
  assign n33757 = n33700 & ~n33756 ;
  assign n33758 = n33714 & n33747 ;
  assign n33759 = n33701 & n33706 ;
  assign n33760 = ~n33758 & ~n33759 ;
  assign n33761 = ~n33700 & ~n33760 ;
  assign n33762 = ~n33757 & ~n33761 ;
  assign n33763 = ~n33731 & n33762 ;
  assign n33764 = ~n33754 & n33763 ;
  assign n33765 = ~\u1_L10_reg[14]/NET0131  & ~n33764 ;
  assign n33766 = \u1_L10_reg[14]/NET0131  & n33764 ;
  assign n33767 = ~n33765 & ~n33766 ;
  assign n33782 = ~n33336 & n33389 ;
  assign n33783 = ~n33359 & ~n33389 ;
  assign n33784 = ~n33330 & ~n33783 ;
  assign n33785 = ~n33782 & ~n33784 ;
  assign n33786 = ~n33343 & ~n33785 ;
  assign n33780 = ~n33357 & ~n33370 ;
  assign n33781 = n33354 & n33780 ;
  assign n33787 = ~n33358 & ~n33385 ;
  assign n33788 = ~n33781 & n33787 ;
  assign n33789 = ~n33786 & n33788 ;
  assign n33790 = ~n33368 & ~n33789 ;
  assign n33768 = n33330 & n33399 ;
  assign n33771 = ~n33349 & ~n33353 ;
  assign n33772 = n33353 & n33359 ;
  assign n33773 = ~n33771 & ~n33772 ;
  assign n33774 = n33343 & ~n33773 ;
  assign n33769 = n33330 & ~n33389 ;
  assign n33770 = n33398 & n33769 ;
  assign n33775 = ~n33343 & ~n33380 ;
  assign n33776 = ~n33771 & n33775 ;
  assign n33777 = ~n33770 & ~n33776 ;
  assign n33778 = ~n33774 & n33777 ;
  assign n33779 = n33368 & ~n33778 ;
  assign n33791 = ~n33768 & ~n33779 ;
  assign n33792 = ~n33790 & n33791 ;
  assign n33793 = ~\u1_L10_reg[17]/NET0131  & ~n33792 ;
  assign n33794 = \u1_L10_reg[17]/NET0131  & n33792 ;
  assign n33795 = ~n33793 & ~n33794 ;
  assign n33796 = decrypt_pad & ~\u1_uk_K_r10_reg[43]/NET0131  ;
  assign n33797 = ~decrypt_pad & ~\u1_uk_K_r10_reg[7]/NET0131  ;
  assign n33798 = ~n33796 & ~n33797 ;
  assign n33799 = \u1_R10_reg[30]/NET0131  & ~n33798 ;
  assign n33800 = ~\u1_R10_reg[30]/NET0131  & n33798 ;
  assign n33801 = ~n33799 & ~n33800 ;
  assign n33802 = decrypt_pad & ~\u1_uk_K_r10_reg[31]/NET0131  ;
  assign n33803 = ~decrypt_pad & ~\u1_uk_K_r10_reg[22]/NET0131  ;
  assign n33804 = ~n33802 & ~n33803 ;
  assign n33805 = \u1_R10_reg[1]/NET0131  & ~n33804 ;
  assign n33806 = ~\u1_R10_reg[1]/NET0131  & n33804 ;
  assign n33807 = ~n33805 & ~n33806 ;
  assign n33808 = ~n33801 & ~n33807 ;
  assign n33809 = decrypt_pad & ~\u1_uk_K_r10_reg[15]/NET0131  ;
  assign n33810 = ~decrypt_pad & ~\u1_uk_K_r10_reg[38]/NET0131  ;
  assign n33811 = ~n33809 & ~n33810 ;
  assign n33812 = \u1_R10_reg[28]/NET0131  & ~n33811 ;
  assign n33813 = ~\u1_R10_reg[28]/NET0131  & n33811 ;
  assign n33814 = ~n33812 & ~n33813 ;
  assign n33815 = ~n33808 & ~n33814 ;
  assign n33816 = decrypt_pad & ~\u1_uk_K_r10_reg[42]/NET0131  ;
  assign n33817 = ~decrypt_pad & ~\u1_uk_K_r10_reg[37]/NET0131  ;
  assign n33818 = ~n33816 & ~n33817 ;
  assign n33819 = \u1_R10_reg[29]/NET0131  & ~n33818 ;
  assign n33820 = ~\u1_R10_reg[29]/NET0131  & n33818 ;
  assign n33821 = ~n33819 & ~n33820 ;
  assign n33822 = ~n33815 & n33821 ;
  assign n33823 = n33807 & ~n33814 ;
  assign n33824 = ~n33821 & n33823 ;
  assign n33825 = ~n33822 & ~n33824 ;
  assign n33826 = decrypt_pad & ~\u1_uk_K_r10_reg[0]/NET0131  ;
  assign n33827 = ~decrypt_pad & ~\u1_uk_K_r10_reg[50]/NET0131  ;
  assign n33828 = ~n33826 & ~n33827 ;
  assign n33829 = \u1_R10_reg[31]/P0001  & ~n33828 ;
  assign n33830 = ~\u1_R10_reg[31]/P0001  & n33828 ;
  assign n33831 = ~n33829 & ~n33830 ;
  assign n33832 = ~n33825 & n33831 ;
  assign n33833 = ~n33801 & ~n33821 ;
  assign n33834 = ~n33807 & n33814 ;
  assign n33835 = n33833 & n33834 ;
  assign n33836 = ~n33832 & ~n33835 ;
  assign n33837 = decrypt_pad & ~\u1_uk_K_r10_reg[37]/NET0131  ;
  assign n33838 = ~decrypt_pad & ~\u1_uk_K_r10_reg[1]/NET0131  ;
  assign n33839 = ~n33837 & ~n33838 ;
  assign n33840 = \u1_R10_reg[32]/NET0131  & ~n33839 ;
  assign n33841 = ~\u1_R10_reg[32]/NET0131  & n33839 ;
  assign n33842 = ~n33840 & ~n33841 ;
  assign n33843 = ~n33836 & ~n33842 ;
  assign n33853 = n33801 & n33821 ;
  assign n33854 = ~n33814 & n33853 ;
  assign n33855 = ~n33807 & n33854 ;
  assign n33850 = ~n33807 & ~n33814 ;
  assign n33867 = n33833 & n33850 ;
  assign n33868 = ~n33855 & ~n33867 ;
  assign n33847 = n33801 & ~n33821 ;
  assign n33869 = n33814 & n33847 ;
  assign n33844 = ~n33801 & n33821 ;
  assign n33870 = n33823 & n33844 ;
  assign n33871 = ~n33869 & ~n33870 ;
  assign n33872 = n33868 & n33871 ;
  assign n33873 = ~n33831 & ~n33872 ;
  assign n33845 = n33814 & n33844 ;
  assign n33846 = ~n33814 & n33831 ;
  assign n33848 = n33807 & n33847 ;
  assign n33849 = ~n33846 & n33848 ;
  assign n33856 = ~n33845 & ~n33849 ;
  assign n33851 = ~n33821 & n33850 ;
  assign n33852 = n33831 & n33851 ;
  assign n33857 = ~n33852 & ~n33855 ;
  assign n33858 = n33856 & n33857 ;
  assign n33859 = n33842 & ~n33858 ;
  assign n33860 = ~n33801 & n33824 ;
  assign n33861 = n33807 & n33854 ;
  assign n33862 = ~n33860 & ~n33861 ;
  assign n33863 = n33831 & ~n33862 ;
  assign n33864 = n33814 & ~n33821 ;
  assign n33865 = ~n33831 & ~n33842 ;
  assign n33866 = n33864 & n33865 ;
  assign n33874 = ~n33863 & ~n33866 ;
  assign n33875 = ~n33859 & n33874 ;
  assign n33876 = ~n33873 & n33875 ;
  assign n33877 = ~n33843 & n33876 ;
  assign n33878 = ~\u1_L10_reg[15]/P0001  & ~n33877 ;
  assign n33879 = \u1_L10_reg[15]/P0001  & n33877 ;
  assign n33880 = ~n33878 & ~n33879 ;
  assign n33903 = n33524 & ~n33537 ;
  assign n33904 = ~n33530 & n33903 ;
  assign n33905 = ~n33572 & ~n33904 ;
  assign n33906 = n33567 & ~n33905 ;
  assign n33907 = ~n33560 & n33619 ;
  assign n33908 = ~n33906 & n33907 ;
  assign n33909 = n33518 & ~n33908 ;
  assign n33889 = ~n33537 & ~n33543 ;
  assign n33890 = ~n33524 & n33889 ;
  assign n33891 = n33550 & ~n33890 ;
  assign n33892 = ~n33572 & ~n33889 ;
  assign n33893 = n33524 & ~n33892 ;
  assign n33894 = ~n33518 & ~n33893 ;
  assign n33895 = ~n33891 & ~n33894 ;
  assign n33896 = ~n33547 & ~n33585 ;
  assign n33897 = n33624 & ~n33896 ;
  assign n33898 = ~n33589 & ~n33897 ;
  assign n33899 = ~n33895 & n33898 ;
  assign n33900 = ~n33567 & ~n33899 ;
  assign n33881 = ~n33547 & n33624 ;
  assign n33882 = n33530 & n33585 ;
  assign n33883 = ~n33881 & ~n33882 ;
  assign n33884 = ~n33518 & ~n33883 ;
  assign n33885 = n33537 & ~n33568 ;
  assign n33886 = n33590 & n33885 ;
  assign n33887 = ~n33884 & ~n33886 ;
  assign n33888 = n33567 & ~n33887 ;
  assign n33901 = ~n33543 & n33593 ;
  assign n33902 = n33590 & n33901 ;
  assign n33910 = ~n33888 & ~n33902 ;
  assign n33911 = ~n33900 & n33910 ;
  assign n33912 = ~n33909 & n33911 ;
  assign n33913 = ~\u1_L10_reg[1]/NET0131  & ~n33912 ;
  assign n33914 = \u1_L10_reg[1]/NET0131  & n33912 ;
  assign n33915 = ~n33913 & ~n33914 ;
  assign n33920 = ~n33807 & n33869 ;
  assign n33916 = n33807 & n33814 ;
  assign n33917 = ~n33801 & ~n33831 ;
  assign n33918 = ~n33844 & ~n33917 ;
  assign n33919 = n33916 & ~n33918 ;
  assign n33928 = ~n33842 & ~n33854 ;
  assign n33931 = ~n33919 & n33928 ;
  assign n33932 = ~n33920 & n33931 ;
  assign n33921 = n33821 & n33834 ;
  assign n33922 = ~n33869 & ~n33921 ;
  assign n33923 = n33831 & ~n33922 ;
  assign n33926 = n33801 & ~n33831 ;
  assign n33927 = n33823 & n33926 ;
  assign n33924 = n33821 & ~n33831 ;
  assign n33925 = n33850 & n33924 ;
  assign n33929 = ~n33867 & ~n33925 ;
  assign n33930 = ~n33927 & n33929 ;
  assign n33933 = ~n33923 & n33930 ;
  assign n33934 = n33932 & n33933 ;
  assign n33935 = ~n33808 & ~n33848 ;
  assign n33936 = n33814 & ~n33935 ;
  assign n33937 = ~n33831 & ~n33936 ;
  assign n33938 = n33814 & n33853 ;
  assign n33942 = n33831 & ~n33938 ;
  assign n33939 = n33807 & n33821 ;
  assign n33940 = ~n33814 & n33939 ;
  assign n33941 = n33807 & n33833 ;
  assign n33943 = ~n33940 & ~n33941 ;
  assign n33944 = n33942 & n33943 ;
  assign n33945 = ~n33937 & ~n33944 ;
  assign n33946 = ~n33851 & ~n33921 ;
  assign n33947 = n33801 & ~n33946 ;
  assign n33948 = n33842 & ~n33860 ;
  assign n33949 = ~n33947 & n33948 ;
  assign n33950 = ~n33945 & n33949 ;
  assign n33951 = ~n33934 & ~n33950 ;
  assign n33952 = n33833 & n33846 ;
  assign n33953 = ~n33831 & n33844 ;
  assign n33954 = n33916 & n33953 ;
  assign n33955 = ~n33952 & ~n33954 ;
  assign n33956 = ~n33951 & n33955 ;
  assign n33957 = ~\u1_L10_reg[21]/NET0131  & ~n33956 ;
  assign n33958 = \u1_L10_reg[21]/NET0131  & n33956 ;
  assign n33959 = ~n33957 & ~n33958 ;
  assign n33963 = ~n33679 & ~n33685 ;
  assign n33964 = ~n33693 & n33963 ;
  assign n33962 = ~n33678 & ~n33692 ;
  assign n33965 = ~n33712 & ~n33962 ;
  assign n33966 = ~n33964 & n33965 ;
  assign n33967 = n33700 & ~n33966 ;
  assign n33968 = ~n33692 & n33711 ;
  assign n33969 = ~n33694 & ~n33968 ;
  assign n33970 = ~n33700 & ~n33969 ;
  assign n33960 = ~n33672 & n33685 ;
  assign n33961 = n33692 & n33960 ;
  assign n33971 = n33672 & n33733 ;
  assign n33972 = ~n33961 & ~n33971 ;
  assign n33973 = ~n33970 & n33972 ;
  assign n33974 = ~n33967 & n33973 ;
  assign n33975 = n33730 & ~n33974 ;
  assign n33983 = ~n33678 & n33706 ;
  assign n33984 = ~n33709 & ~n33983 ;
  assign n33985 = ~n33700 & ~n33984 ;
  assign n33987 = ~n33685 & n33700 ;
  assign n33988 = n33693 & n33987 ;
  assign n33982 = n33742 & n33962 ;
  assign n33986 = n33706 & n33714 ;
  assign n33989 = ~n33982 & ~n33986 ;
  assign n33990 = ~n33988 & n33989 ;
  assign n33991 = ~n33985 & n33990 ;
  assign n33992 = ~n33730 & ~n33991 ;
  assign n33976 = ~n33755 & ~n33971 ;
  assign n33977 = ~n33672 & n33714 ;
  assign n33978 = ~n33692 & n33977 ;
  assign n33979 = n33976 & ~n33978 ;
  assign n33980 = n33700 & ~n33979 ;
  assign n33981 = n33708 & n33744 ;
  assign n33993 = ~n33713 & ~n33981 ;
  assign n33994 = ~n33980 & n33993 ;
  assign n33995 = ~n33992 & n33994 ;
  assign n33996 = ~n33975 & n33995 ;
  assign n33997 = ~\u1_L10_reg[25]/NET0131  & ~n33996 ;
  assign n33998 = \u1_L10_reg[25]/NET0131  & n33996 ;
  assign n33999 = ~n33997 & ~n33998 ;
  assign n34034 = decrypt_pad & ~\u1_uk_K_r10_reg[55]/NET0131  ;
  assign n34035 = ~decrypt_pad & ~\u1_uk_K_r10_reg[46]/NET0131  ;
  assign n34036 = ~n34034 & ~n34035 ;
  assign n34037 = \u1_R10_reg[6]/NET0131  & ~n34036 ;
  assign n34038 = ~\u1_R10_reg[6]/NET0131  & n34036 ;
  assign n34039 = ~n34037 & ~n34038 ;
  assign n34012 = decrypt_pad & ~\u1_uk_K_r10_reg[53]/NET0131  ;
  assign n34013 = ~decrypt_pad & ~\u1_uk_K_r10_reg[19]/NET0131  ;
  assign n34014 = ~n34012 & ~n34013 ;
  assign n34015 = \u1_R10_reg[4]/NET0131  & ~n34014 ;
  assign n34016 = ~\u1_R10_reg[4]/NET0131  & n34014 ;
  assign n34017 = ~n34015 & ~n34016 ;
  assign n34018 = decrypt_pad & ~\u1_uk_K_r10_reg[20]/NET0131  ;
  assign n34019 = ~decrypt_pad & ~\u1_uk_K_r10_reg[11]/NET0131  ;
  assign n34020 = ~n34018 & ~n34019 ;
  assign n34021 = \u1_R10_reg[9]/NET0131  & ~n34020 ;
  assign n34022 = ~\u1_R10_reg[9]/NET0131  & n34020 ;
  assign n34023 = ~n34021 & ~n34022 ;
  assign n34025 = decrypt_pad & ~\u1_uk_K_r10_reg[32]/NET0131  ;
  assign n34026 = ~decrypt_pad & ~\u1_uk_K_r10_reg[55]/NET0131  ;
  assign n34027 = ~n34025 & ~n34026 ;
  assign n34028 = \u1_R10_reg[5]/NET0131  & ~n34027 ;
  assign n34029 = ~\u1_R10_reg[5]/NET0131  & n34027 ;
  assign n34030 = ~n34028 & ~n34029 ;
  assign n34040 = ~n34023 & n34030 ;
  assign n34041 = ~n34017 & n34040 ;
  assign n34042 = n34039 & n34041 ;
  assign n34032 = ~n34023 & ~n34030 ;
  assign n34033 = n34017 & n34032 ;
  assign n34006 = decrypt_pad & ~\u1_uk_K_r10_reg[17]/NET0131  ;
  assign n34007 = ~decrypt_pad & ~\u1_uk_K_r10_reg[40]/NET0131  ;
  assign n34008 = ~n34006 & ~n34007 ;
  assign n34009 = \u1_R10_reg[7]/NET0131  & ~n34008 ;
  assign n34010 = ~\u1_R10_reg[7]/NET0131  & n34008 ;
  assign n34011 = ~n34009 & ~n34010 ;
  assign n34024 = n34017 & n34023 ;
  assign n34031 = n34024 & n34030 ;
  assign n34043 = n34011 & ~n34031 ;
  assign n34044 = ~n34033 & n34043 ;
  assign n34045 = ~n34042 & n34044 ;
  assign n34051 = ~n34030 & n34039 ;
  assign n34052 = ~n34011 & ~n34051 ;
  assign n34053 = ~n34011 & n34017 ;
  assign n34054 = ~n34052 & ~n34053 ;
  assign n34046 = ~n34017 & ~n34023 ;
  assign n34047 = ~n34039 & n34046 ;
  assign n34048 = ~n34017 & n34023 ;
  assign n34049 = n34030 & n34048 ;
  assign n34050 = ~n34047 & ~n34049 ;
  assign n34055 = n34017 & n34039 ;
  assign n34056 = n34040 & n34055 ;
  assign n34057 = n34050 & ~n34056 ;
  assign n34058 = ~n34054 & n34057 ;
  assign n34059 = ~n34045 & ~n34058 ;
  assign n34064 = n34039 & n34048 ;
  assign n34065 = ~n34030 & n34064 ;
  assign n34000 = decrypt_pad & ~\u1_uk_K_r10_reg[40]/NET0131  ;
  assign n34001 = ~decrypt_pad & ~\u1_uk_K_r10_reg[6]/NET0131  ;
  assign n34002 = ~n34000 & ~n34001 ;
  assign n34003 = \u1_R10_reg[8]/NET0131  & ~n34002 ;
  assign n34004 = ~\u1_R10_reg[8]/NET0131  & n34002 ;
  assign n34005 = ~n34003 & ~n34004 ;
  assign n34060 = n34017 & ~n34039 ;
  assign n34061 = n34023 & ~n34030 ;
  assign n34062 = ~n34011 & ~n34061 ;
  assign n34063 = n34060 & ~n34062 ;
  assign n34066 = n34005 & ~n34063 ;
  assign n34067 = ~n34065 & n34066 ;
  assign n34068 = ~n34059 & n34067 ;
  assign n34069 = n34011 & n34050 ;
  assign n34072 = ~n34030 & n34048 ;
  assign n34070 = ~n34023 & n34060 ;
  assign n34071 = n34017 & n34030 ;
  assign n34073 = ~n34070 & ~n34071 ;
  assign n34074 = ~n34072 & n34073 ;
  assign n34075 = ~n34054 & n34074 ;
  assign n34076 = ~n34069 & ~n34075 ;
  assign n34077 = ~n34024 & ~n34046 ;
  assign n34078 = n34051 & ~n34077 ;
  assign n34079 = ~n34005 & ~n34056 ;
  assign n34080 = ~n34078 & n34079 ;
  assign n34081 = ~n34076 & n34080 ;
  assign n34082 = ~n34068 & ~n34081 ;
  assign n34083 = ~\u1_L10_reg[28]/NET0131  & n34082 ;
  assign n34084 = \u1_L10_reg[28]/NET0131  & ~n34082 ;
  assign n34085 = ~n34083 & ~n34084 ;
  assign n34104 = ~n33426 & n33457 ;
  assign n34105 = ~n33491 & ~n34104 ;
  assign n34106 = ~n33440 & ~n33479 ;
  assign n34107 = ~n33456 & ~n34106 ;
  assign n34108 = n34105 & ~n34107 ;
  assign n34109 = n33449 & ~n34108 ;
  assign n34086 = n33426 & n33457 ;
  assign n34087 = n33439 & n34086 ;
  assign n34094 = ~n33439 & ~n33499 ;
  assign n34102 = ~n34087 & ~n34094 ;
  assign n34103 = ~n33449 & ~n34102 ;
  assign n34110 = n33462 & n33480 ;
  assign n34111 = ~n34103 & ~n34110 ;
  assign n34112 = ~n34109 & n34111 ;
  assign n34113 = ~n33420 & ~n34112 ;
  assign n34088 = n33426 & n33464 ;
  assign n34089 = ~n33497 & ~n34088 ;
  assign n34090 = ~n34087 & n34089 ;
  assign n34091 = n33449 & ~n34090 ;
  assign n34095 = ~n33466 & n33476 ;
  assign n34092 = ~n33426 & ~n33484 ;
  assign n34093 = n33449 & ~n34092 ;
  assign n34096 = ~n34093 & ~n34094 ;
  assign n34097 = ~n34095 & n34096 ;
  assign n34098 = ~n34091 & ~n34097 ;
  assign n34099 = n33420 & ~n34098 ;
  assign n34100 = n33449 & n33456 ;
  assign n34101 = n33441 & n34100 ;
  assign n34114 = ~n33490 & ~n34101 ;
  assign n34115 = ~n34099 & n34114 ;
  assign n34116 = ~n34113 & n34115 ;
  assign n34117 = \u1_L10_reg[29]/NET0131  & ~n34116 ;
  assign n34118 = ~\u1_L10_reg[29]/NET0131  & n34116 ;
  assign n34119 = ~n34117 & ~n34118 ;
  assign n34128 = ~n34011 & ~n34030 ;
  assign n34129 = n34046 & n34128 ;
  assign n34126 = n34030 & ~n34039 ;
  assign n34127 = n34024 & n34126 ;
  assign n34135 = n34005 & ~n34127 ;
  assign n34136 = ~n34129 & n34135 ;
  assign n34132 = ~n34011 & n34039 ;
  assign n34133 = ~n34071 & n34132 ;
  assign n34134 = ~n34077 & n34133 ;
  assign n34125 = ~n34030 & n34070 ;
  assign n34130 = ~n34071 & ~n34126 ;
  assign n34131 = n34011 & ~n34130 ;
  assign n34137 = ~n34125 & ~n34131 ;
  assign n34138 = ~n34134 & n34137 ;
  assign n34139 = n34136 & n34138 ;
  assign n34140 = ~n34040 & ~n34072 ;
  assign n34141 = ~n34039 & ~n34140 ;
  assign n34146 = n34055 & n34061 ;
  assign n34147 = n34011 & n34146 ;
  assign n34152 = ~n34005 & ~n34147 ;
  assign n34153 = ~n34141 & n34152 ;
  assign n34142 = ~n34055 & ~n34061 ;
  assign n34143 = n34024 & ~n34030 ;
  assign n34144 = ~n34011 & ~n34143 ;
  assign n34145 = ~n34142 & n34144 ;
  assign n34148 = n34023 & ~n34039 ;
  assign n34149 = n34128 & n34148 ;
  assign n34150 = n34030 & n34064 ;
  assign n34151 = ~n34149 & ~n34150 ;
  assign n34154 = ~n34145 & n34151 ;
  assign n34155 = n34153 & n34154 ;
  assign n34156 = ~n34139 & ~n34155 ;
  assign n34120 = ~n34023 & n34051 ;
  assign n34121 = ~n34017 & n34120 ;
  assign n34122 = n34030 & n34060 ;
  assign n34123 = ~n34121 & ~n34122 ;
  assign n34124 = n34011 & ~n34123 ;
  assign n34157 = n34048 & ~n34126 ;
  assign n34158 = n34052 & n34157 ;
  assign n34159 = ~n34124 & ~n34158 ;
  assign n34160 = ~n34156 & n34159 ;
  assign n34161 = \u1_L10_reg[2]/NET0131  & n34160 ;
  assign n34162 = ~\u1_L10_reg[2]/NET0131  & ~n34160 ;
  assign n34163 = ~n34161 & ~n34162 ;
  assign n34167 = n33456 & ~n33458 ;
  assign n34168 = n33465 & n34167 ;
  assign n34169 = n33420 & ~n34168 ;
  assign n34170 = ~n33432 & n33484 ;
  assign n34171 = n33426 & n34170 ;
  assign n34172 = n34169 & ~n34171 ;
  assign n34173 = ~n33420 & ~n33490 ;
  assign n34174 = ~n33495 & n34173 ;
  assign n34175 = ~n33439 & n33480 ;
  assign n34176 = ~n33463 & ~n34086 ;
  assign n34177 = ~n34175 & n34176 ;
  assign n34178 = n34174 & n34177 ;
  assign n34179 = ~n34172 & ~n34178 ;
  assign n34164 = ~n33488 & ~n33497 ;
  assign n34165 = ~n34086 & n34164 ;
  assign n34166 = n33439 & ~n34165 ;
  assign n34180 = n33449 & ~n34166 ;
  assign n34181 = ~n34179 & n34180 ;
  assign n34183 = ~n33464 & ~n33485 ;
  assign n34184 = n34169 & n34183 ;
  assign n34185 = ~n33474 & ~n34110 ;
  assign n34186 = n34174 & n34185 ;
  assign n34187 = ~n34184 & ~n34186 ;
  assign n34182 = n33439 & ~n34105 ;
  assign n34188 = ~n33449 & ~n34170 ;
  assign n34189 = ~n34182 & n34188 ;
  assign n34190 = ~n34187 & n34189 ;
  assign n34191 = ~n34181 & ~n34190 ;
  assign n34192 = ~\u1_L10_reg[4]/NET0131  & n34191 ;
  assign n34193 = \u1_L10_reg[4]/NET0131  & ~n34191 ;
  assign n34194 = ~n34192 & ~n34193 ;
  assign n34195 = ~n33545 & n33622 ;
  assign n34196 = ~n33543 & ~n33590 ;
  assign n34197 = ~n33569 & ~n34196 ;
  assign n34198 = ~n33537 & ~n34197 ;
  assign n34199 = ~n33524 & n33548 ;
  assign n34200 = ~n33551 & ~n34199 ;
  assign n34201 = ~n33567 & ~n34200 ;
  assign n34202 = ~n33518 & ~n34201 ;
  assign n34203 = ~n34198 & n34202 ;
  assign n34204 = ~n34195 & ~n34203 ;
  assign n34206 = ~n33573 & ~n33890 ;
  assign n34207 = n33530 & ~n34206 ;
  assign n34205 = n33518 & n33552 ;
  assign n34214 = n33567 & ~n34205 ;
  assign n34215 = ~n34207 & n34214 ;
  assign n34208 = ~n33586 & ~n33882 ;
  assign n34209 = n33537 & ~n34208 ;
  assign n34210 = ~n33530 & n33544 ;
  assign n34211 = ~n33568 & ~n34210 ;
  assign n34212 = ~n33518 & ~n33903 ;
  assign n34213 = ~n34211 & n34212 ;
  assign n34216 = ~n34209 & ~n34213 ;
  assign n34217 = n34215 & n34216 ;
  assign n34218 = n33577 & ~n33585 ;
  assign n34219 = ~n33567 & ~n33904 ;
  assign n34220 = n33588 & n34219 ;
  assign n34221 = ~n34218 & n34220 ;
  assign n34222 = ~n34217 & ~n34221 ;
  assign n34223 = ~n34204 & ~n34222 ;
  assign n34224 = ~\u1_L10_reg[26]/NET0131  & ~n34223 ;
  assign n34225 = \u1_L10_reg[26]/NET0131  & n34223 ;
  assign n34226 = ~n34224 & ~n34225 ;
  assign n34238 = n33432 & ~n33441 ;
  assign n34239 = ~n33474 & ~n34238 ;
  assign n34240 = n33449 & ~n34239 ;
  assign n34236 = n33439 & n33491 ;
  assign n34237 = ~n33449 & ~n34164 ;
  assign n34241 = ~n34236 & ~n34237 ;
  assign n34242 = ~n34240 & n34241 ;
  assign n34243 = ~n33420 & ~n34242 ;
  assign n34229 = ~n33481 & ~n33483 ;
  assign n34230 = ~n34175 & n34229 ;
  assign n34231 = ~n33426 & ~n34230 ;
  assign n34227 = n33439 & ~n34164 ;
  assign n34228 = n33442 & n33449 ;
  assign n34232 = ~n33485 & ~n34228 ;
  assign n34233 = ~n34227 & n34232 ;
  assign n34234 = ~n34231 & n34233 ;
  assign n34235 = n33420 & ~n34234 ;
  assign n34244 = n33487 & ~n33496 ;
  assign n34245 = ~n34235 & n34244 ;
  assign n34246 = ~n34243 & n34245 ;
  assign n34247 = ~\u1_L10_reg[19]/P0001  & ~n34246 ;
  assign n34248 = \u1_L10_reg[19]/P0001  & n34246 ;
  assign n34249 = ~n34247 & ~n34248 ;
  assign n34268 = n33330 & n33783 ;
  assign n34269 = ~n33784 & ~n34268 ;
  assign n34267 = n33349 & ~n33384 ;
  assign n34270 = ~n33343 & ~n34267 ;
  assign n34271 = n34269 & n34270 ;
  assign n34272 = n33343 & n33769 ;
  assign n34273 = ~n34267 & n34272 ;
  assign n34274 = ~n33352 & ~n33772 ;
  assign n34275 = ~n34273 & n34274 ;
  assign n34276 = ~n34271 & n34275 ;
  assign n34277 = n33368 & ~n34276 ;
  assign n34259 = ~n33360 & ~n33362 ;
  assign n34260 = ~n33361 & n33368 ;
  assign n34261 = ~n34259 & ~n34260 ;
  assign n34262 = n33353 & n33400 ;
  assign n34263 = n33349 & n33371 ;
  assign n34264 = ~n34262 & ~n34263 ;
  assign n34265 = ~n34261 & n34264 ;
  assign n34266 = ~n33343 & ~n34265 ;
  assign n34250 = ~n33349 & ~n33370 ;
  assign n34251 = ~n33336 & n33343 ;
  assign n34252 = ~n33362 & n34251 ;
  assign n34253 = ~n34250 & n34252 ;
  assign n34255 = n33398 & n33780 ;
  assign n34254 = n33350 & n33370 ;
  assign n34256 = ~n33377 & ~n34254 ;
  assign n34257 = ~n34255 & n34256 ;
  assign n34258 = ~n33368 & ~n34257 ;
  assign n34278 = ~n34253 & ~n34258 ;
  assign n34279 = ~n34266 & n34278 ;
  assign n34280 = ~n34277 & n34279 ;
  assign n34281 = \u1_L10_reg[23]/NET0131  & ~n34280 ;
  assign n34282 = ~\u1_L10_reg[23]/NET0131  & n34280 ;
  assign n34283 = ~n34281 & ~n34282 ;
  assign n34303 = ~n33814 & n33833 ;
  assign n34304 = ~n33921 & ~n33940 ;
  assign n34305 = ~n34303 & n34304 ;
  assign n34306 = n33842 & ~n34305 ;
  assign n34308 = n33814 & n33941 ;
  assign n34307 = n33834 & n33844 ;
  assign n34309 = ~n33855 & ~n34307 ;
  assign n34310 = ~n34308 & n34309 ;
  assign n34311 = ~n34306 & n34310 ;
  assign n34312 = ~n33831 & ~n34311 ;
  assign n34297 = n33831 & ~n33834 ;
  assign n34298 = n33822 & n34297 ;
  assign n34299 = ~n33861 & ~n33941 ;
  assign n34300 = ~n33920 & n34299 ;
  assign n34301 = ~n34298 & n34300 ;
  assign n34302 = n33842 & ~n34301 ;
  assign n34284 = ~n33807 & n33831 ;
  assign n34285 = n33823 & ~n33842 ;
  assign n34286 = ~n34284 & ~n34285 ;
  assign n34287 = n33847 & ~n34286 ;
  assign n34291 = n33831 & ~n33854 ;
  assign n34289 = ~n33807 & n33844 ;
  assign n34290 = n33807 & ~n33844 ;
  assign n34292 = ~n34289 & ~n34290 ;
  assign n34293 = n34291 & n34292 ;
  assign n34288 = n33916 & n33926 ;
  assign n34294 = ~n33925 & ~n34288 ;
  assign n34295 = ~n34293 & n34294 ;
  assign n34296 = ~n33842 & ~n34295 ;
  assign n34313 = ~n34287 & ~n34296 ;
  assign n34314 = ~n34302 & n34313 ;
  assign n34315 = ~n34312 & n34314 ;
  assign n34316 = ~\u1_L10_reg[27]/NET0131  & ~n34315 ;
  assign n34317 = \u1_L10_reg[27]/NET0131  & n34315 ;
  assign n34318 = ~n34316 & ~n34317 ;
  assign n34324 = ~n33286 & ~n33307 ;
  assign n34326 = ~n33273 & n33645 ;
  assign n34327 = n34324 & ~n34326 ;
  assign n34325 = ~n33273 & ~n34324 ;
  assign n34328 = ~n33265 & ~n34325 ;
  assign n34329 = ~n34327 & n34328 ;
  assign n34319 = n33275 & n33307 ;
  assign n34320 = n33238 & ~n33307 ;
  assign n34321 = n33296 & ~n34320 ;
  assign n34322 = ~n33258 & ~n34321 ;
  assign n34323 = n33265 & ~n34322 ;
  assign n34330 = ~n34319 & ~n34323 ;
  assign n34331 = ~n34329 & n34330 ;
  assign n34332 = n33232 & ~n34331 ;
  assign n34334 = ~n33637 & ~n33645 ;
  assign n34335 = ~n33265 & ~n34334 ;
  assign n34336 = ~n33244 & n33289 ;
  assign n34337 = n33265 & ~n33637 ;
  assign n34338 = ~n34336 & n34337 ;
  assign n34339 = ~n34335 & ~n34338 ;
  assign n34333 = n33244 & ~n33639 ;
  assign n34340 = n33306 & ~n34333 ;
  assign n34341 = ~n34339 & n34340 ;
  assign n34342 = ~n33232 & ~n34341 ;
  assign n34343 = n33265 & n33288 ;
  assign n34344 = ~n33276 & n33303 ;
  assign n34345 = n33269 & n34344 ;
  assign n34346 = ~n34343 & ~n34345 ;
  assign n34347 = ~n34342 & n34346 ;
  assign n34348 = ~n34332 & n34347 ;
  assign n34349 = \u1_L10_reg[32]/NET0131  & n34348 ;
  assign n34350 = ~\u1_L10_reg[32]/NET0131  & ~n34348 ;
  assign n34351 = ~n34349 & ~n34350 ;
  assign n34386 = decrypt_pad & ~\u1_uk_K_r10_reg[3]/NET0131  ;
  assign n34387 = ~decrypt_pad & ~\u1_uk_K_r10_reg[26]/NET0131  ;
  assign n34388 = ~n34386 & ~n34387 ;
  assign n34389 = \u1_R10_reg[11]/NET0131  & ~n34388 ;
  assign n34390 = ~\u1_R10_reg[11]/NET0131  & n34388 ;
  assign n34391 = ~n34389 & ~n34390 ;
  assign n34378 = decrypt_pad & ~\u1_uk_K_r10_reg[18]/NET0131  ;
  assign n34379 = ~decrypt_pad & ~\u1_uk_K_r10_reg[41]/P0001  ;
  assign n34380 = ~n34378 & ~n34379 ;
  assign n34381 = \u1_R10_reg[12]/NET0131  & ~n34380 ;
  assign n34382 = ~\u1_R10_reg[12]/NET0131  & n34380 ;
  assign n34383 = ~n34381 & ~n34382 ;
  assign n34352 = decrypt_pad & ~\u1_uk_K_r10_reg[6]/NET0131  ;
  assign n34353 = ~decrypt_pad & ~\u1_uk_K_r10_reg[54]/NET0131  ;
  assign n34354 = ~n34352 & ~n34353 ;
  assign n34355 = \u1_R10_reg[13]/NET0131  & ~n34354 ;
  assign n34356 = ~\u1_R10_reg[13]/NET0131  & n34354 ;
  assign n34357 = ~n34355 & ~n34356 ;
  assign n34365 = decrypt_pad & ~\u1_uk_K_r10_reg[26]/NET0131  ;
  assign n34366 = ~decrypt_pad & ~\u1_uk_K_r10_reg[17]/NET0131  ;
  assign n34367 = ~n34365 & ~n34366 ;
  assign n34368 = \u1_R10_reg[9]/NET0131  & ~n34367 ;
  assign n34369 = ~\u1_R10_reg[9]/NET0131  & n34367 ;
  assign n34370 = ~n34368 & ~n34369 ;
  assign n34392 = n34357 & ~n34370 ;
  assign n34371 = decrypt_pad & ~\u1_uk_K_r10_reg[34]/NET0131  ;
  assign n34372 = ~decrypt_pad & ~\u1_uk_K_r10_reg[25]/NET0131  ;
  assign n34373 = ~n34371 & ~n34372 ;
  assign n34374 = \u1_R10_reg[10]/NET0131  & ~n34373 ;
  assign n34375 = ~\u1_R10_reg[10]/NET0131  & n34373 ;
  assign n34376 = ~n34374 & ~n34375 ;
  assign n34358 = decrypt_pad & ~\u1_uk_K_r10_reg[54]/NET0131  ;
  assign n34359 = ~decrypt_pad & ~\u1_uk_K_r10_reg[20]/NET0131  ;
  assign n34360 = ~n34358 & ~n34359 ;
  assign n34361 = \u1_R10_reg[8]/NET0131  & ~n34360 ;
  assign n34362 = ~\u1_R10_reg[8]/NET0131  & n34360 ;
  assign n34363 = ~n34361 & ~n34362 ;
  assign n34394 = n34357 & ~n34363 ;
  assign n34395 = n34376 & n34394 ;
  assign n34396 = ~n34357 & n34363 ;
  assign n34397 = n34370 & n34396 ;
  assign n34398 = ~n34395 & ~n34397 ;
  assign n34399 = ~n34392 & n34398 ;
  assign n34400 = n34383 & ~n34399 ;
  assign n34393 = n34376 & n34392 ;
  assign n34364 = ~n34357 & ~n34363 ;
  assign n34401 = ~n34370 & ~n34376 ;
  assign n34402 = n34364 & n34401 ;
  assign n34403 = ~n34393 & ~n34402 ;
  assign n34404 = ~n34400 & n34403 ;
  assign n34405 = n34391 & ~n34404 ;
  assign n34377 = n34370 & n34376 ;
  assign n34413 = ~n34377 & ~n34401 ;
  assign n34406 = n34357 & n34363 ;
  assign n34407 = ~n34364 & ~n34406 ;
  assign n34414 = n34357 & n34391 ;
  assign n34415 = n34407 & ~n34414 ;
  assign n34416 = ~n34413 & ~n34415 ;
  assign n34408 = ~n34401 & n34407 ;
  assign n34409 = ~n34376 & n34391 ;
  assign n34410 = n34357 & n34409 ;
  assign n34411 = ~n34377 & ~n34410 ;
  assign n34412 = n34408 & n34411 ;
  assign n34417 = ~n34383 & ~n34412 ;
  assign n34418 = ~n34416 & n34417 ;
  assign n34384 = n34377 & n34383 ;
  assign n34385 = n34364 & n34384 ;
  assign n34421 = n34370 & ~n34376 ;
  assign n34422 = ~n34363 & ~n34421 ;
  assign n34419 = ~n34357 & n34370 ;
  assign n34420 = ~n34392 & ~n34419 ;
  assign n34423 = n34383 & ~n34391 ;
  assign n34424 = n34420 & n34423 ;
  assign n34425 = ~n34422 & n34424 ;
  assign n34426 = ~n34385 & ~n34425 ;
  assign n34427 = ~n34418 & n34426 ;
  assign n34428 = ~n34405 & n34427 ;
  assign n34429 = ~\u1_L10_reg[6]/NET0131  & ~n34428 ;
  assign n34430 = \u1_L10_reg[6]/NET0131  & n34428 ;
  assign n34431 = ~n34429 & ~n34430 ;
  assign n34449 = ~n33257 & ~n33643 ;
  assign n34432 = n33244 & ~n34324 ;
  assign n34450 = n33238 & n33307 ;
  assign n34451 = ~n34432 & ~n34450 ;
  assign n34452 = ~n34449 & n34451 ;
  assign n34453 = ~n33265 & ~n34452 ;
  assign n34433 = ~n34336 & ~n34432 ;
  assign n34434 = n33238 & ~n34433 ;
  assign n34443 = ~n33238 & ~n33251 ;
  assign n34444 = n34324 & n34443 ;
  assign n34454 = n33265 & n34444 ;
  assign n34455 = ~n34434 & ~n34454 ;
  assign n34456 = ~n34453 & n34455 ;
  assign n34457 = n33232 & ~n34456 ;
  assign n34435 = ~n33265 & n34434 ;
  assign n34436 = n33232 & ~n33265 ;
  assign n34437 = n33295 & ~n34324 ;
  assign n34438 = n33250 & ~n33655 ;
  assign n34439 = n33265 & n34320 ;
  assign n34440 = ~n34438 & n34439 ;
  assign n34441 = ~n34437 & ~n34440 ;
  assign n34442 = ~n33232 & ~n34441 ;
  assign n34445 = ~n33265 & n34444 ;
  assign n34446 = ~n33259 & ~n34445 ;
  assign n34447 = ~n34442 & n34446 ;
  assign n34448 = ~n34436 & ~n34447 ;
  assign n34458 = ~n34435 & ~n34448 ;
  assign n34459 = ~n34457 & n34458 ;
  assign n34460 = ~\u1_L10_reg[7]/NET0131  & ~n34459 ;
  assign n34461 = \u1_L10_reg[7]/NET0131  & n34459 ;
  assign n34462 = ~n34460 & ~n34461 ;
  assign n34475 = n33700 & ~n33710 ;
  assign n34476 = ~n33712 & n34475 ;
  assign n34477 = n33714 & ~n33747 ;
  assign n34478 = ~n33700 & ~n33968 ;
  assign n34479 = ~n34477 & n34478 ;
  assign n34480 = ~n34476 & ~n34479 ;
  assign n34481 = ~n33694 & n33976 ;
  assign n34482 = ~n34480 & n34481 ;
  assign n34483 = ~n33730 & ~n34482 ;
  assign n34463 = ~n33672 & n33702 ;
  assign n34464 = ~n33968 & ~n34463 ;
  assign n34465 = n33700 & ~n34464 ;
  assign n34466 = n33678 & n33742 ;
  assign n34467 = n33760 & ~n34466 ;
  assign n34468 = ~n34465 & n34467 ;
  assign n34469 = n33730 & ~n34468 ;
  assign n34470 = n33685 & n33694 ;
  assign n34471 = ~n33707 & ~n33758 ;
  assign n34472 = ~n34470 & n34471 ;
  assign n34473 = n33700 & ~n34472 ;
  assign n34474 = ~n33685 & n33981 ;
  assign n34484 = ~n34473 & ~n34474 ;
  assign n34485 = ~n34469 & n34484 ;
  assign n34486 = ~n34483 & n34485 ;
  assign n34487 = ~\u1_L10_reg[8]/NET0131  & ~n34486 ;
  assign n34488 = \u1_L10_reg[8]/NET0131  & n34486 ;
  assign n34489 = ~n34487 & ~n34488 ;
  assign n34501 = ~n34056 & ~n34127 ;
  assign n34502 = ~n34041 & ~n34065 ;
  assign n34503 = ~n34125 & n34502 ;
  assign n34504 = ~n34005 & ~n34503 ;
  assign n34505 = n34501 & ~n34504 ;
  assign n34506 = ~n34011 & ~n34505 ;
  assign n34495 = ~n34030 & n34077 ;
  assign n34494 = n34030 & ~n34070 ;
  assign n34496 = n34011 & ~n34494 ;
  assign n34497 = ~n34495 & n34496 ;
  assign n34490 = n34011 & ~n34040 ;
  assign n34491 = n34055 & n34490 ;
  assign n34492 = ~n34017 & ~n34128 ;
  assign n34493 = n34148 & n34492 ;
  assign n34498 = ~n34491 & ~n34493 ;
  assign n34499 = ~n34497 & n34498 ;
  assign n34500 = ~n34005 & ~n34499 ;
  assign n34507 = ~n34120 & n34144 ;
  assign n34508 = n34032 & ~n34039 ;
  assign n34509 = n34011 & ~n34064 ;
  assign n34510 = ~n34508 & n34509 ;
  assign n34511 = ~n34507 & ~n34510 ;
  assign n34512 = n34046 & n34126 ;
  assign n34513 = n34501 & ~n34512 ;
  assign n34514 = n34151 & n34513 ;
  assign n34515 = ~n34511 & n34514 ;
  assign n34516 = n34005 & ~n34515 ;
  assign n34517 = ~n34500 & ~n34516 ;
  assign n34518 = ~n34506 & n34517 ;
  assign n34519 = ~\u1_L10_reg[13]/NET0131  & n34518 ;
  assign n34520 = \u1_L10_reg[13]/NET0131  & ~n34518 ;
  assign n34521 = ~n34519 & ~n34520 ;
  assign n34522 = n34364 & n34370 ;
  assign n34523 = n34391 & n34522 ;
  assign n34524 = ~n34363 & ~n34370 ;
  assign n34525 = n34363 & n34370 ;
  assign n34526 = ~n34524 & ~n34525 ;
  assign n34527 = n34357 & n34526 ;
  assign n34528 = ~n34419 & ~n34527 ;
  assign n34529 = ~n34364 & n34528 ;
  assign n34530 = ~n34523 & ~n34529 ;
  assign n34531 = ~n34376 & ~n34530 ;
  assign n34532 = n34363 & n34376 ;
  assign n34533 = ~n34391 & ~n34532 ;
  assign n34534 = ~n34357 & n34376 ;
  assign n34535 = ~n34396 & ~n34534 ;
  assign n34536 = n34533 & ~n34535 ;
  assign n34537 = n34370 & n34395 ;
  assign n34538 = ~n34536 & ~n34537 ;
  assign n34539 = ~n34531 & n34538 ;
  assign n34540 = n34383 & ~n34539 ;
  assign n34543 = ~n34364 & n34391 ;
  assign n34544 = ~n34528 & n34543 ;
  assign n34541 = ~n34391 & n34535 ;
  assign n34542 = ~n34527 & n34541 ;
  assign n34545 = ~n34402 & ~n34542 ;
  assign n34546 = ~n34544 & n34545 ;
  assign n34547 = ~n34383 & ~n34546 ;
  assign n34548 = ~n34526 & n34534 ;
  assign n34549 = n34391 & ~n34548 ;
  assign n34550 = ~n34370 & n34532 ;
  assign n34551 = ~n34391 & ~n34550 ;
  assign n34552 = ~n34549 & ~n34551 ;
  assign n34553 = ~n34547 & ~n34552 ;
  assign n34554 = ~n34540 & n34553 ;
  assign n34555 = ~\u1_L10_reg[16]/NET0131  & ~n34554 ;
  assign n34556 = \u1_L10_reg[16]/NET0131  & n34554 ;
  assign n34557 = ~n34555 & ~n34556 ;
  assign n34562 = ~n34376 & n34394 ;
  assign n34563 = n34364 & n34376 ;
  assign n34564 = ~n34562 & ~n34563 ;
  assign n34565 = ~n34522 & ~n34550 ;
  assign n34566 = n34564 & n34565 ;
  assign n34567 = n34391 & ~n34566 ;
  assign n34558 = ~n34357 & n34550 ;
  assign n34559 = n34401 & ~n34407 ;
  assign n34560 = n34398 & ~n34559 ;
  assign n34561 = ~n34391 & ~n34560 ;
  assign n34568 = ~n34558 & ~n34561 ;
  assign n34569 = ~n34567 & n34568 ;
  assign n34570 = ~n34383 & ~n34569 ;
  assign n34571 = n34376 & ~n34394 ;
  assign n34572 = ~n34525 & n34571 ;
  assign n34573 = n34391 & ~n34421 ;
  assign n34574 = ~n34562 & n34573 ;
  assign n34575 = ~n34572 & n34574 ;
  assign n34576 = ~n34391 & ~n34408 ;
  assign n34577 = ~n34559 & n34576 ;
  assign n34578 = ~n34575 & ~n34577 ;
  assign n34579 = n34383 & ~n34578 ;
  assign n34580 = n34376 & ~n34391 ;
  assign n34581 = n34370 & n34406 ;
  assign n34582 = n34580 & n34581 ;
  assign n34583 = n34407 & n34409 ;
  assign n34584 = n34420 & n34583 ;
  assign n34585 = ~n34582 & ~n34584 ;
  assign n34586 = ~n34579 & n34585 ;
  assign n34587 = ~n34570 & n34586 ;
  assign n34588 = ~\u1_L10_reg[24]/NET0131  & ~n34587 ;
  assign n34589 = \u1_L10_reg[24]/NET0131  & n34587 ;
  assign n34590 = ~n34588 & ~n34589 ;
  assign n34592 = ~n34522 & n34533 ;
  assign n34593 = n34396 & n34401 ;
  assign n34594 = n34391 & ~n34593 ;
  assign n34595 = n34564 & n34594 ;
  assign n34596 = ~n34592 & ~n34595 ;
  assign n34597 = n34383 & ~n34596 ;
  assign n34599 = ~n34419 & n34532 ;
  assign n34600 = ~n34357 & n34421 ;
  assign n34601 = ~n34599 & ~n34600 ;
  assign n34602 = n34391 & ~n34601 ;
  assign n34605 = ~n34383 & ~n34559 ;
  assign n34598 = ~n34370 & n34395 ;
  assign n34603 = ~n34419 & ~n34524 ;
  assign n34604 = n34533 & n34603 ;
  assign n34606 = ~n34598 & ~n34604 ;
  assign n34607 = n34605 & n34606 ;
  assign n34608 = ~n34602 & n34607 ;
  assign n34609 = ~n34597 & ~n34608 ;
  assign n34610 = n34384 & ~n34406 ;
  assign n34591 = n34414 & n34550 ;
  assign n34611 = n34419 & n34580 ;
  assign n34612 = ~n34591 & ~n34611 ;
  assign n34613 = ~n34610 & n34612 ;
  assign n34614 = ~n34609 & n34613 ;
  assign n34615 = ~\u1_L10_reg[30]/NET0131  & n34614 ;
  assign n34616 = \u1_L10_reg[30]/NET0131  & ~n34614 ;
  assign n34617 = ~n34615 & ~n34616 ;
  assign n34619 = n33692 & n33701 ;
  assign n34620 = ~n33738 & ~n34619 ;
  assign n34621 = n33700 & ~n34620 ;
  assign n34618 = ~n33700 & n33740 ;
  assign n34622 = n33730 & ~n33748 ;
  assign n34623 = ~n33713 & n34622 ;
  assign n34624 = ~n34618 & n34623 ;
  assign n34625 = ~n34621 & n34624 ;
  assign n34630 = ~n33733 & ~n33977 ;
  assign n34631 = n33700 & ~n34630 ;
  assign n34627 = ~n33708 & n33960 ;
  assign n34626 = n33700 & ~n33747 ;
  assign n34628 = ~n33732 & ~n34626 ;
  assign n34629 = ~n34627 & n34628 ;
  assign n34632 = ~n33730 & ~n34629 ;
  assign n34633 = ~n34631 & n34632 ;
  assign n34634 = ~n34625 & ~n34633 ;
  assign n34635 = ~n33758 & n34475 ;
  assign n34636 = ~n33700 & ~n33746 ;
  assign n34637 = ~n33721 & n34636 ;
  assign n34638 = ~n34463 & n34637 ;
  assign n34639 = ~n34635 & ~n34638 ;
  assign n34640 = ~n34634 & ~n34639 ;
  assign n34641 = ~\u1_L10_reg[3]/NET0131  & ~n34640 ;
  assign n34642 = \u1_L10_reg[3]/NET0131  & n34640 ;
  assign n34643 = ~n34641 & ~n34642 ;
  assign n34645 = n33336 & n34269 ;
  assign n34644 = n33780 & n34252 ;
  assign n34646 = n33368 & ~n34263 ;
  assign n34647 = ~n34644 & n34646 ;
  assign n34648 = ~n34645 & n34647 ;
  assign n34652 = n33343 & ~n33401 ;
  assign n34653 = ~n33780 & n34652 ;
  assign n34651 = n33337 & ~n33783 ;
  assign n34649 = n33379 & n33780 ;
  assign n34650 = n33362 & n33397 ;
  assign n34654 = ~n33368 & ~n34650 ;
  assign n34655 = ~n34649 & n34654 ;
  assign n34656 = ~n34651 & n34655 ;
  assign n34657 = ~n34653 & n34656 ;
  assign n34658 = ~n34648 & ~n34657 ;
  assign n34659 = n33324 & n33387 ;
  assign n34660 = ~n33381 & n34659 ;
  assign n34661 = ~n34658 & ~n34660 ;
  assign n34662 = ~\u1_L10_reg[9]/NET0131  & ~n34661 ;
  assign n34663 = \u1_L10_reg[9]/NET0131  & n34661 ;
  assign n34664 = ~n34662 & ~n34663 ;
  assign n34676 = ~n34056 & ~n34146 ;
  assign n34677 = ~n34508 & n34676 ;
  assign n34672 = n34011 & n34031 ;
  assign n34673 = n34030 & ~n34132 ;
  assign n34674 = ~n34017 & ~n34051 ;
  assign n34675 = ~n34673 & n34674 ;
  assign n34678 = ~n34672 & ~n34675 ;
  assign n34679 = n34677 & n34678 ;
  assign n34680 = ~n34005 & ~n34679 ;
  assign n34668 = n34011 & ~n34140 ;
  assign n34666 = ~n34032 & ~n34148 ;
  assign n34667 = n34053 & ~n34666 ;
  assign n34669 = ~n34121 & ~n34667 ;
  assign n34670 = ~n34668 & n34669 ;
  assign n34671 = n34005 & ~n34670 ;
  assign n34665 = ~n34011 & n34049 ;
  assign n34681 = n34024 & n34039 ;
  assign n34682 = ~n34512 & ~n34681 ;
  assign n34683 = n34011 & ~n34682 ;
  assign n34684 = ~n34665 & ~n34683 ;
  assign n34685 = ~n34671 & n34684 ;
  assign n34686 = ~n34680 & n34685 ;
  assign n34687 = \u1_L10_reg[18]/P0001  & n34686 ;
  assign n34688 = ~\u1_L10_reg[18]/P0001  & ~n34686 ;
  assign n34689 = ~n34687 & ~n34688 ;
  assign n34742 = decrypt_pad & ~\u1_uk_K_r9_reg[25]/NET0131  ;
  assign n34743 = ~decrypt_pad & ~\u1_uk_K_r9_reg[19]/NET0131  ;
  assign n34744 = ~n34742 & ~n34743 ;
  assign n34745 = \u1_R9_reg[4]/NET0131  & ~n34744 ;
  assign n34746 = ~\u1_R9_reg[4]/NET0131  & n34744 ;
  assign n34747 = ~n34745 & ~n34746 ;
  assign n34690 = decrypt_pad & ~\u1_uk_K_r9_reg[47]/NET0131  ;
  assign n34691 = ~decrypt_pad & ~\u1_uk_K_r9_reg[41]/NET0131  ;
  assign n34692 = ~n34690 & ~n34691 ;
  assign n34693 = \u1_R9_reg[3]/NET0131  & ~n34692 ;
  assign n34694 = ~\u1_R9_reg[3]/NET0131  & n34692 ;
  assign n34695 = ~n34693 & ~n34694 ;
  assign n34709 = decrypt_pad & ~\u1_uk_K_r9_reg[53]/NET0131  ;
  assign n34710 = ~decrypt_pad & ~\u1_uk_K_r9_reg[47]/NET0131  ;
  assign n34711 = ~n34709 & ~n34710 ;
  assign n34712 = \u1_R9_reg[5]/NET0131  & ~n34711 ;
  assign n34713 = ~\u1_R9_reg[5]/NET0131  & n34711 ;
  assign n34714 = ~n34712 & ~n34713 ;
  assign n34722 = decrypt_pad & ~\u1_uk_K_r9_reg[55]/NET0131  ;
  assign n34723 = ~decrypt_pad & ~\u1_uk_K_r9_reg[17]/NET0131  ;
  assign n34724 = ~n34722 & ~n34723 ;
  assign n34725 = \u1_R9_reg[1]/NET0131  & ~n34724 ;
  assign n34726 = ~\u1_R9_reg[1]/NET0131  & n34724 ;
  assign n34727 = ~n34725 & ~n34726 ;
  assign n34734 = n34714 & ~n34727 ;
  assign n34696 = decrypt_pad & ~\u1_uk_K_r9_reg[13]/NET0131  ;
  assign n34697 = ~decrypt_pad & ~\u1_uk_K_r9_reg[32]/NET0131  ;
  assign n34698 = ~n34696 & ~n34697 ;
  assign n34699 = \u1_R9_reg[2]/NET0131  & ~n34698 ;
  assign n34700 = ~\u1_R9_reg[2]/NET0131  & n34698 ;
  assign n34701 = ~n34699 & ~n34700 ;
  assign n34703 = decrypt_pad & ~\u1_uk_K_r9_reg[34]/NET0131  ;
  assign n34704 = ~decrypt_pad & ~\u1_uk_K_r9_reg[53]/NET0131  ;
  assign n34705 = ~n34703 & ~n34704 ;
  assign n34706 = \u1_R9_reg[32]/NET0131  & ~n34705 ;
  assign n34707 = ~\u1_R9_reg[32]/NET0131  & n34705 ;
  assign n34708 = ~n34706 & ~n34707 ;
  assign n34733 = n34701 & ~n34708 ;
  assign n34750 = ~n34714 & n34733 ;
  assign n34751 = ~n34734 & ~n34750 ;
  assign n34752 = n34695 & ~n34751 ;
  assign n34729 = ~n34701 & n34708 ;
  assign n34757 = ~n34729 & ~n34733 ;
  assign n34716 = n34708 & n34714 ;
  assign n34758 = ~n34716 & ~n34727 ;
  assign n34759 = ~n34757 & n34758 ;
  assign n34730 = ~n34695 & n34727 ;
  assign n34749 = n34708 & n34730 ;
  assign n34753 = ~n34708 & n34714 ;
  assign n34754 = n34695 & ~n34701 ;
  assign n34755 = n34727 & ~n34754 ;
  assign n34756 = n34753 & ~n34755 ;
  assign n34760 = ~n34749 & ~n34756 ;
  assign n34761 = ~n34759 & n34760 ;
  assign n34762 = ~n34752 & n34761 ;
  assign n34763 = n34747 & ~n34762 ;
  assign n34702 = n34695 & n34701 ;
  assign n34715 = ~n34708 & ~n34714 ;
  assign n34717 = ~n34715 & ~n34716 ;
  assign n34718 = n34702 & n34717 ;
  assign n34719 = ~n34701 & ~n34714 ;
  assign n34720 = ~n34708 & n34719 ;
  assign n34721 = ~n34718 & ~n34720 ;
  assign n34728 = ~n34721 & n34727 ;
  assign n34731 = n34714 & n34729 ;
  assign n34732 = ~n34730 & n34731 ;
  assign n34735 = n34701 & ~n34727 ;
  assign n34736 = n34708 & ~n34735 ;
  assign n34737 = ~n34695 & ~n34733 ;
  assign n34738 = ~n34734 & n34737 ;
  assign n34739 = ~n34736 & n34738 ;
  assign n34740 = ~n34732 & ~n34739 ;
  assign n34741 = ~n34728 & n34740 ;
  assign n34748 = ~n34741 & ~n34747 ;
  assign n34766 = n34701 & n34716 ;
  assign n34767 = ~n34719 & ~n34766 ;
  assign n34768 = n34727 & ~n34767 ;
  assign n34769 = n34733 & n34734 ;
  assign n34770 = ~n34768 & ~n34769 ;
  assign n34771 = ~n34695 & ~n34770 ;
  assign n34764 = n34695 & n34715 ;
  assign n34765 = n34735 & n34764 ;
  assign n34772 = ~n34701 & ~n34727 ;
  assign n34773 = n34695 & n34708 ;
  assign n34774 = n34772 & n34773 ;
  assign n34775 = ~n34765 & ~n34774 ;
  assign n34776 = ~n34771 & n34775 ;
  assign n34777 = ~n34748 & n34776 ;
  assign n34778 = ~n34763 & n34777 ;
  assign n34779 = ~\u1_L9_reg[31]/NET0131  & ~n34778 ;
  assign n34780 = \u1_L9_reg[31]/NET0131  & n34778 ;
  assign n34781 = ~n34779 & ~n34780 ;
  assign n34782 = decrypt_pad & ~\u1_uk_K_r9_reg[51]/NET0131  ;
  assign n34783 = ~decrypt_pad & ~\u1_uk_K_r9_reg[43]/NET0131  ;
  assign n34784 = ~n34782 & ~n34783 ;
  assign n34785 = \u1_R9_reg[24]/NET0131  & ~n34784 ;
  assign n34786 = ~\u1_R9_reg[24]/NET0131  & n34784 ;
  assign n34787 = ~n34785 & ~n34786 ;
  assign n34788 = decrypt_pad & ~\u1_uk_K_r9_reg[49]/NET0131  ;
  assign n34789 = ~decrypt_pad & ~\u1_uk_K_r9_reg[45]/NET0131  ;
  assign n34790 = ~n34788 & ~n34789 ;
  assign n34791 = \u1_R9_reg[23]/NET0131  & ~n34790 ;
  assign n34792 = ~\u1_R9_reg[23]/NET0131  & n34790 ;
  assign n34793 = ~n34791 & ~n34792 ;
  assign n34814 = decrypt_pad & ~\u1_uk_K_r9_reg[36]/NET0131  ;
  assign n34815 = ~decrypt_pad & ~\u1_uk_K_r9_reg[28]/NET0131  ;
  assign n34816 = ~n34814 & ~n34815 ;
  assign n34817 = \u1_R9_reg[22]/NET0131  & ~n34816 ;
  assign n34818 = ~\u1_R9_reg[22]/NET0131  & n34816 ;
  assign n34819 = ~n34817 & ~n34818 ;
  assign n34794 = decrypt_pad & ~\u1_uk_K_r9_reg[30]/NET0131  ;
  assign n34795 = ~decrypt_pad & ~\u1_uk_K_r9_reg[22]/NET0131  ;
  assign n34796 = ~n34794 & ~n34795 ;
  assign n34797 = \u1_R9_reg[20]/NET0131  & ~n34796 ;
  assign n34798 = ~\u1_R9_reg[20]/NET0131  & n34796 ;
  assign n34799 = ~n34797 & ~n34798 ;
  assign n34807 = decrypt_pad & ~\u1_uk_K_r9_reg[14]/NET0131  ;
  assign n34808 = ~decrypt_pad & ~\u1_uk_K_r9_reg[37]/NET0131  ;
  assign n34809 = ~n34807 & ~n34808 ;
  assign n34810 = \u1_R9_reg[21]/NET0131  & ~n34809 ;
  assign n34811 = ~\u1_R9_reg[21]/NET0131  & n34809 ;
  assign n34812 = ~n34810 & ~n34811 ;
  assign n34830 = n34799 & ~n34812 ;
  assign n34855 = n34819 & n34830 ;
  assign n34856 = ~n34799 & ~n34819 ;
  assign n34857 = ~n34855 & ~n34856 ;
  assign n34858 = n34793 & n34857 ;
  assign n34820 = n34812 & n34819 ;
  assign n34821 = ~n34799 & n34820 ;
  assign n34828 = ~n34793 & ~n34821 ;
  assign n34846 = n34812 & ~n34819 ;
  assign n34859 = n34799 & n34846 ;
  assign n34860 = n34828 & ~n34859 ;
  assign n34861 = ~n34858 & ~n34860 ;
  assign n34800 = decrypt_pad & ~\u1_uk_K_r9_reg[15]/NET0131  ;
  assign n34801 = ~decrypt_pad & ~\u1_uk_K_r9_reg[7]/NET0131  ;
  assign n34802 = ~n34800 & ~n34801 ;
  assign n34803 = \u1_R9_reg[25]/NET0131  & ~n34802 ;
  assign n34804 = ~\u1_R9_reg[25]/NET0131  & n34802 ;
  assign n34805 = ~n34803 & ~n34804 ;
  assign n34822 = n34799 & ~n34805 ;
  assign n34840 = ~n34793 & ~n34819 ;
  assign n34862 = n34822 & n34840 ;
  assign n34831 = n34805 & n34830 ;
  assign n34863 = n34819 & n34831 ;
  assign n34864 = ~n34862 & ~n34863 ;
  assign n34832 = ~n34799 & n34805 ;
  assign n34849 = ~n34812 & n34832 ;
  assign n34854 = n34793 & n34849 ;
  assign n34847 = ~n34805 & n34846 ;
  assign n34865 = n34799 & n34847 ;
  assign n34866 = ~n34854 & ~n34865 ;
  assign n34867 = n34864 & n34866 ;
  assign n34868 = ~n34861 & n34867 ;
  assign n34869 = ~n34787 & ~n34868 ;
  assign n34823 = ~n34812 & ~n34819 ;
  assign n34824 = n34822 & n34823 ;
  assign n34806 = n34799 & n34805 ;
  assign n34813 = n34806 & n34812 ;
  assign n34825 = ~n34813 & ~n34821 ;
  assign n34826 = ~n34824 & n34825 ;
  assign n34827 = n34793 & ~n34826 ;
  assign n34833 = n34812 & n34832 ;
  assign n34834 = ~n34819 & ~n34831 ;
  assign n34835 = ~n34833 & n34834 ;
  assign n34829 = n34806 & n34819 ;
  assign n34836 = n34828 & ~n34829 ;
  assign n34837 = ~n34835 & n34836 ;
  assign n34838 = ~n34827 & ~n34837 ;
  assign n34839 = n34787 & ~n34838 ;
  assign n34841 = n34812 & n34822 ;
  assign n34842 = ~n34799 & ~n34805 ;
  assign n34843 = ~n34812 & n34842 ;
  assign n34844 = ~n34841 & ~n34843 ;
  assign n34845 = n34840 & ~n34844 ;
  assign n34850 = ~n34819 & n34849 ;
  assign n34848 = ~n34799 & n34847 ;
  assign n34851 = ~n34829 & ~n34848 ;
  assign n34852 = ~n34850 & n34851 ;
  assign n34853 = n34793 & ~n34852 ;
  assign n34870 = ~n34845 & ~n34853 ;
  assign n34871 = ~n34839 & n34870 ;
  assign n34872 = ~n34869 & n34871 ;
  assign n34873 = \u1_L9_reg[11]/NET0131  & ~n34872 ;
  assign n34874 = ~\u1_L9_reg[11]/NET0131  & n34872 ;
  assign n34875 = ~n34873 & ~n34874 ;
  assign n34876 = decrypt_pad & ~\u1_uk_K_r9_reg[31]/P0001  ;
  assign n34877 = ~decrypt_pad & ~\u1_uk_K_r9_reg[50]/NET0131  ;
  assign n34878 = ~n34876 & ~n34877 ;
  assign n34879 = \u1_R9_reg[28]/NET0131  & ~n34878 ;
  assign n34880 = ~\u1_R9_reg[28]/NET0131  & n34878 ;
  assign n34881 = ~n34879 & ~n34880 ;
  assign n34882 = decrypt_pad & ~\u1_uk_K_r9_reg[7]/NET0131  ;
  assign n34883 = ~decrypt_pad & ~\u1_uk_K_r9_reg[30]/NET0131  ;
  assign n34884 = ~n34882 & ~n34883 ;
  assign n34885 = \u1_R9_reg[26]/NET0131  & ~n34884 ;
  assign n34886 = ~\u1_R9_reg[26]/NET0131  & n34884 ;
  assign n34887 = ~n34885 & ~n34886 ;
  assign n34888 = decrypt_pad & ~\u1_uk_K_r9_reg[22]/NET0131  ;
  assign n34889 = ~decrypt_pad & ~\u1_uk_K_r9_reg[14]/NET0131  ;
  assign n34890 = ~n34888 & ~n34889 ;
  assign n34891 = \u1_R9_reg[25]/NET0131  & ~n34890 ;
  assign n34892 = ~\u1_R9_reg[25]/NET0131  & n34890 ;
  assign n34893 = ~n34891 & ~n34892 ;
  assign n34922 = ~n34887 & ~n34893 ;
  assign n34894 = decrypt_pad & ~\u1_uk_K_r9_reg[50]/NET0131  ;
  assign n34895 = ~decrypt_pad & ~\u1_uk_K_r9_reg[42]/NET0131  ;
  assign n34896 = ~n34894 & ~n34895 ;
  assign n34897 = \u1_R9_reg[29]/NET0131  & ~n34896 ;
  assign n34898 = ~\u1_R9_reg[29]/NET0131  & n34896 ;
  assign n34899 = ~n34897 & ~n34898 ;
  assign n34925 = ~n34887 & ~n34899 ;
  assign n34945 = ~n34922 & ~n34925 ;
  assign n34901 = decrypt_pad & ~\u1_uk_K_r9_reg[42]/NET0131  ;
  assign n34902 = ~decrypt_pad & ~\u1_uk_K_r9_reg[38]/NET0131  ;
  assign n34903 = ~n34901 & ~n34902 ;
  assign n34904 = \u1_R9_reg[24]/NET0131  & ~n34903 ;
  assign n34905 = ~\u1_R9_reg[24]/NET0131  & n34903 ;
  assign n34906 = ~n34904 & ~n34905 ;
  assign n34909 = decrypt_pad & ~\u1_uk_K_r9_reg[16]/NET0131  ;
  assign n34910 = ~decrypt_pad & ~\u1_uk_K_r9_reg[8]/NET0131  ;
  assign n34911 = ~n34909 & ~n34910 ;
  assign n34912 = \u1_R9_reg[27]/NET0131  & ~n34911 ;
  assign n34913 = ~\u1_R9_reg[27]/NET0131  & n34911 ;
  assign n34914 = ~n34912 & ~n34913 ;
  assign n34924 = n34887 & n34893 ;
  assign n34944 = n34914 & ~n34924 ;
  assign n34946 = n34906 & n34944 ;
  assign n34947 = n34945 & n34946 ;
  assign n34938 = n34899 & n34906 ;
  assign n34939 = n34922 & n34938 ;
  assign n34940 = n34893 & n34899 ;
  assign n34941 = ~n34906 & n34940 ;
  assign n34942 = ~n34939 & ~n34941 ;
  assign n34943 = ~n34914 & ~n34942 ;
  assign n34933 = ~n34899 & ~n34906 ;
  assign n34934 = n34922 & n34933 ;
  assign n34935 = n34899 & ~n34906 ;
  assign n34936 = n34887 & ~n34893 ;
  assign n34937 = n34935 & n34936 ;
  assign n34948 = ~n34934 & ~n34937 ;
  assign n34949 = ~n34943 & n34948 ;
  assign n34950 = ~n34947 & n34949 ;
  assign n34951 = n34881 & ~n34950 ;
  assign n34926 = ~n34914 & ~n34924 ;
  assign n34927 = ~n34925 & n34926 ;
  assign n34923 = n34914 & ~n34922 ;
  assign n34928 = n34906 & ~n34923 ;
  assign n34929 = ~n34927 & n34928 ;
  assign n34900 = ~n34893 & ~n34899 ;
  assign n34907 = n34900 & ~n34906 ;
  assign n34908 = n34887 & n34907 ;
  assign n34915 = n34908 & ~n34914 ;
  assign n34916 = ~n34887 & ~n34906 ;
  assign n34917 = n34887 & n34906 ;
  assign n34918 = ~n34916 & ~n34917 ;
  assign n34919 = ~n34893 & n34914 ;
  assign n34920 = n34899 & ~n34919 ;
  assign n34921 = ~n34918 & n34920 ;
  assign n34930 = ~n34915 & ~n34921 ;
  assign n34931 = ~n34929 & n34930 ;
  assign n34932 = ~n34881 & ~n34931 ;
  assign n34954 = n34924 & n34933 ;
  assign n34955 = ~n34937 & ~n34954 ;
  assign n34956 = ~n34899 & n34906 ;
  assign n34957 = ~n34893 & n34956 ;
  assign n34958 = n34955 & ~n34957 ;
  assign n34959 = n34914 & ~n34958 ;
  assign n34952 = n34893 & ~n34914 ;
  assign n34953 = ~n34918 & n34952 ;
  assign n34960 = n34919 & n34925 ;
  assign n34961 = ~n34953 & ~n34960 ;
  assign n34962 = ~n34959 & n34961 ;
  assign n34963 = ~n34932 & n34962 ;
  assign n34964 = ~n34951 & n34963 ;
  assign n34965 = ~\u1_L9_reg[22]/NET0131  & ~n34964 ;
  assign n34966 = \u1_L9_reg[22]/NET0131  & n34964 ;
  assign n34967 = ~n34965 & ~n34966 ;
  assign n34981 = decrypt_pad & ~\u1_uk_K_r9_reg[10]/NET0131  ;
  assign n34982 = ~decrypt_pad & ~\u1_uk_K_r9_reg[4]/NET0131  ;
  assign n34983 = ~n34981 & ~n34982 ;
  assign n34984 = \u1_R9_reg[13]/NET0131  & ~n34983 ;
  assign n34985 = ~\u1_R9_reg[13]/NET0131  & n34983 ;
  assign n34986 = ~n34984 & ~n34985 ;
  assign n34987 = decrypt_pad & ~\u1_uk_K_r9_reg[19]/NET0131  ;
  assign n34988 = ~decrypt_pad & ~\u1_uk_K_r9_reg[13]/NET0131  ;
  assign n34989 = ~n34987 & ~n34988 ;
  assign n34990 = \u1_R9_reg[15]/NET0131  & ~n34989 ;
  assign n34991 = ~\u1_R9_reg[15]/NET0131  & n34989 ;
  assign n34992 = ~n34990 & ~n34991 ;
  assign n34993 = n34986 & n34992 ;
  assign n34968 = decrypt_pad & ~\u1_uk_K_r9_reg[48]/NET0131  ;
  assign n34969 = ~decrypt_pad & ~\u1_uk_K_r9_reg[10]/NET0131  ;
  assign n34970 = ~n34968 & ~n34969 ;
  assign n34971 = \u1_R9_reg[12]/NET0131  & ~n34970 ;
  assign n34972 = ~\u1_R9_reg[12]/NET0131  & n34970 ;
  assign n34973 = ~n34971 & ~n34972 ;
  assign n34995 = decrypt_pad & ~\u1_uk_K_r9_reg[11]/NET0131  ;
  assign n34996 = ~decrypt_pad & ~\u1_uk_K_r9_reg[5]/NET0131  ;
  assign n34997 = ~n34995 & ~n34996 ;
  assign n34998 = \u1_R9_reg[14]/NET0131  & ~n34997 ;
  assign n34999 = ~\u1_R9_reg[14]/NET0131  & n34997 ;
  assign n35000 = ~n34998 & ~n34999 ;
  assign n35015 = ~n34973 & n35000 ;
  assign n35016 = n34993 & n35015 ;
  assign n35017 = decrypt_pad & ~\u1_uk_K_r9_reg[27]/P0001  ;
  assign n35018 = ~decrypt_pad & ~\u1_uk_K_r9_reg[46]/NET0131  ;
  assign n35019 = ~n35017 & ~n35018 ;
  assign n35020 = \u1_R9_reg[16]/NET0131  & ~n35019 ;
  assign n35021 = ~\u1_R9_reg[16]/NET0131  & n35019 ;
  assign n35022 = ~n35020 & ~n35021 ;
  assign n35032 = ~n35016 & ~n35022 ;
  assign n34974 = decrypt_pad & ~\u1_uk_K_r9_reg[32]/NET0131  ;
  assign n34975 = ~decrypt_pad & ~\u1_uk_K_r9_reg[26]/NET0131  ;
  assign n34976 = ~n34974 & ~n34975 ;
  assign n34977 = \u1_R9_reg[17]/NET0131  & ~n34976 ;
  assign n34978 = ~\u1_R9_reg[17]/NET0131  & n34976 ;
  assign n34979 = ~n34977 & ~n34978 ;
  assign n35030 = n34973 & n34979 ;
  assign n35031 = n34993 & n35030 ;
  assign n35003 = n34979 & ~n35000 ;
  assign n35023 = n34973 & ~n34986 ;
  assign n35024 = n35003 & n35023 ;
  assign n35006 = ~n34986 & n34992 ;
  assign n35007 = ~n34973 & ~n34979 ;
  assign n35025 = n35006 & n35007 ;
  assign n35033 = ~n35024 & ~n35025 ;
  assign n35034 = ~n35031 & n35033 ;
  assign n35035 = n35032 & n35034 ;
  assign n34980 = n34973 & ~n34979 ;
  assign n35009 = n34980 & n35000 ;
  assign n35012 = n34979 & ~n34986 ;
  assign n35013 = ~n35009 & ~n35012 ;
  assign n35014 = ~n34992 & ~n35013 ;
  assign n35008 = ~n35000 & n35007 ;
  assign n35026 = ~n34986 & n35008 ;
  assign n35002 = ~n34973 & n34986 ;
  assign n35027 = ~n34979 & n35000 ;
  assign n35028 = n35002 & n35027 ;
  assign n35029 = ~n35026 & ~n35028 ;
  assign n35036 = ~n35014 & n35029 ;
  assign n35037 = n35035 & n35036 ;
  assign n35045 = n34986 & n35030 ;
  assign n35046 = ~n34986 & ~n34992 ;
  assign n35047 = n35007 & n35046 ;
  assign n35048 = ~n35045 & ~n35047 ;
  assign n35049 = n35000 & ~n35048 ;
  assign n35042 = ~n35002 & ~n35023 ;
  assign n35043 = ~n34992 & ~n35000 ;
  assign n35044 = ~n35042 & n35043 ;
  assign n34994 = n34980 & n34993 ;
  assign n35038 = n35002 & n35003 ;
  assign n35039 = ~n34994 & ~n35038 ;
  assign n35040 = ~n34973 & n34979 ;
  assign n35041 = n35006 & n35040 ;
  assign n35050 = n35022 & ~n35041 ;
  assign n35051 = n35039 & n35050 ;
  assign n35052 = ~n35044 & n35051 ;
  assign n35053 = ~n35049 & n35052 ;
  assign n35054 = ~n35037 & ~n35053 ;
  assign n35010 = ~n35008 & ~n35009 ;
  assign n35011 = n35006 & ~n35010 ;
  assign n35001 = n34994 & ~n35000 ;
  assign n35004 = ~n34992 & n35003 ;
  assign n35005 = n35002 & n35004 ;
  assign n35055 = ~n35001 & ~n35005 ;
  assign n35056 = ~n35011 & n35055 ;
  assign n35057 = ~n35054 & n35056 ;
  assign n35058 = ~\u1_L9_reg[20]/NET0131  & ~n35057 ;
  assign n35059 = \u1_L9_reg[20]/NET0131  & n35057 ;
  assign n35060 = ~n35058 & ~n35059 ;
  assign n35073 = decrypt_pad & ~\u1_uk_K_r9_reg[41]/NET0131  ;
  assign n35074 = ~decrypt_pad & ~\u1_uk_K_r9_reg[3]/NET0131  ;
  assign n35075 = ~n35073 & ~n35074 ;
  assign n35076 = \u1_R9_reg[6]/NET0131  & ~n35075 ;
  assign n35077 = ~\u1_R9_reg[6]/NET0131  & n35075 ;
  assign n35078 = ~n35076 & ~n35077 ;
  assign n35080 = decrypt_pad & ~\u1_uk_K_r9_reg[6]/NET0131  ;
  assign n35081 = ~decrypt_pad & ~\u1_uk_K_r9_reg[25]/NET0131  ;
  assign n35082 = ~n35080 & ~n35081 ;
  assign n35083 = \u1_R9_reg[9]/NET0131  & ~n35082 ;
  assign n35084 = ~\u1_R9_reg[9]/NET0131  & n35082 ;
  assign n35085 = ~n35083 & ~n35084 ;
  assign n35086 = decrypt_pad & ~\u1_uk_K_r9_reg[18]/NET0131  ;
  assign n35087 = ~decrypt_pad & ~\u1_uk_K_r9_reg[12]/NET0131  ;
  assign n35088 = ~n35086 & ~n35087 ;
  assign n35089 = \u1_R9_reg[5]/NET0131  & ~n35088 ;
  assign n35090 = ~\u1_R9_reg[5]/NET0131  & n35088 ;
  assign n35091 = ~n35089 & ~n35090 ;
  assign n35101 = ~n35085 & n35091 ;
  assign n35067 = decrypt_pad & ~\u1_uk_K_r9_reg[39]/NET0131  ;
  assign n35068 = ~decrypt_pad & ~\u1_uk_K_r9_reg[33]/NET0131  ;
  assign n35069 = ~n35067 & ~n35068 ;
  assign n35070 = \u1_R9_reg[4]/NET0131  & ~n35069 ;
  assign n35071 = ~\u1_R9_reg[4]/NET0131  & n35069 ;
  assign n35072 = ~n35070 & ~n35071 ;
  assign n35102 = n35085 & ~n35091 ;
  assign n35103 = ~n35072 & n35102 ;
  assign n35104 = ~n35101 & ~n35103 ;
  assign n35105 = ~n35078 & ~n35104 ;
  assign n35061 = decrypt_pad & ~\u1_uk_K_r9_reg[3]/NET0131  ;
  assign n35062 = ~decrypt_pad & ~\u1_uk_K_r9_reg[54]/NET0131  ;
  assign n35063 = ~n35061 & ~n35062 ;
  assign n35064 = \u1_R9_reg[7]/NET0131  & ~n35063 ;
  assign n35065 = ~\u1_R9_reg[7]/NET0131  & n35063 ;
  assign n35066 = ~n35064 & ~n35065 ;
  assign n35098 = ~n35066 & ~n35091 ;
  assign n35099 = ~n35072 & n35085 ;
  assign n35100 = n35098 & n35099 ;
  assign n35116 = decrypt_pad & ~\u1_uk_K_r9_reg[26]/NET0131  ;
  assign n35117 = ~decrypt_pad & ~\u1_uk_K_r9_reg[20]/NET0131  ;
  assign n35118 = ~n35116 & ~n35117 ;
  assign n35119 = \u1_R9_reg[8]/NET0131  & ~n35118 ;
  assign n35120 = ~\u1_R9_reg[8]/NET0131  & n35118 ;
  assign n35121 = ~n35119 & ~n35120 ;
  assign n35122 = ~n35100 & ~n35121 ;
  assign n35123 = ~n35105 & n35122 ;
  assign n35106 = ~n35078 & n35085 ;
  assign n35107 = n35098 & n35106 ;
  assign n35108 = n35091 & n35099 ;
  assign n35109 = n35078 & n35108 ;
  assign n35110 = ~n35107 & ~n35109 ;
  assign n35111 = n35072 & n35078 ;
  assign n35112 = ~n35066 & ~n35102 ;
  assign n35113 = n35066 & n35102 ;
  assign n35114 = ~n35112 & ~n35113 ;
  assign n35115 = n35111 & ~n35114 ;
  assign n35124 = n35110 & ~n35115 ;
  assign n35125 = n35123 & n35124 ;
  assign n35079 = ~n35072 & n35078 ;
  assign n35135 = n35066 & n35091 ;
  assign n35136 = ~n35078 & ~n35085 ;
  assign n35137 = n35072 & n35136 ;
  assign n35138 = ~n35091 & n35137 ;
  assign n35139 = ~n35135 & ~n35138 ;
  assign n35140 = ~n35079 & ~n35139 ;
  assign n35127 = ~n35072 & ~n35085 ;
  assign n35131 = n35072 & n35085 ;
  assign n35132 = ~n35127 & ~n35131 ;
  assign n35129 = ~n35066 & n35078 ;
  assign n35130 = n35072 & n35091 ;
  assign n35133 = n35129 & ~n35130 ;
  assign n35134 = ~n35132 & n35133 ;
  assign n35094 = n35072 & ~n35078 ;
  assign n35095 = n35091 & n35094 ;
  assign n35126 = n35085 & n35095 ;
  assign n35128 = n35098 & n35127 ;
  assign n35141 = n35121 & ~n35128 ;
  assign n35142 = ~n35126 & n35141 ;
  assign n35143 = ~n35134 & n35142 ;
  assign n35144 = ~n35140 & n35143 ;
  assign n35145 = ~n35125 & ~n35144 ;
  assign n35092 = ~n35085 & ~n35091 ;
  assign n35093 = n35079 & n35092 ;
  assign n35096 = ~n35093 & ~n35095 ;
  assign n35097 = n35066 & ~n35096 ;
  assign n35148 = ~n35098 & ~n35129 ;
  assign n35146 = n35078 & ~n35091 ;
  assign n35147 = ~n35072 & ~n35146 ;
  assign n35149 = n35085 & n35147 ;
  assign n35150 = ~n35148 & n35149 ;
  assign n35151 = ~n35097 & ~n35150 ;
  assign n35152 = ~n35145 & n35151 ;
  assign n35153 = \u1_L9_reg[2]/NET0131  & n35152 ;
  assign n35154 = ~\u1_L9_reg[2]/NET0131  & ~n35152 ;
  assign n35155 = ~n35153 & ~n35154 ;
  assign n35156 = n34819 & n34822 ;
  assign n35157 = ~n34856 & ~n35156 ;
  assign n35158 = n34812 & ~n35157 ;
  assign n35178 = n34806 & ~n34819 ;
  assign n35179 = ~n35158 & ~n35178 ;
  assign n35180 = ~n34793 & ~n35179 ;
  assign n35172 = ~n34812 & n34822 ;
  assign n35173 = ~n34813 & ~n35172 ;
  assign n35174 = ~n34821 & ~n34823 ;
  assign n35175 = ~n34805 & ~n35174 ;
  assign n35176 = n35173 & ~n35175 ;
  assign n35177 = n34793 & ~n35176 ;
  assign n35181 = n34819 & n34849 ;
  assign n35182 = ~n35177 & ~n35181 ;
  assign n35183 = ~n35180 & n35182 ;
  assign n35184 = ~n34787 & ~n35183 ;
  assign n35159 = ~n34833 & ~n35158 ;
  assign n35160 = n34793 & ~n35159 ;
  assign n35161 = n34842 & ~n34846 ;
  assign n35162 = ~n34829 & ~n35161 ;
  assign n35163 = ~n34793 & ~n35162 ;
  assign n35164 = n34819 & n34843 ;
  assign n35165 = ~n34850 & ~n35164 ;
  assign n35166 = n34864 & n35165 ;
  assign n35167 = ~n35163 & n35166 ;
  assign n35168 = ~n35160 & n35167 ;
  assign n35169 = n34787 & ~n35168 ;
  assign n35170 = n34793 & n34805 ;
  assign n35171 = n34846 & n35170 ;
  assign n35185 = ~n34824 & ~n35171 ;
  assign n35186 = ~n35169 & n35185 ;
  assign n35187 = ~n35184 & n35186 ;
  assign n35188 = \u1_L9_reg[29]/NET0131  & ~n35187 ;
  assign n35189 = ~\u1_L9_reg[29]/NET0131  & n35187 ;
  assign n35190 = ~n35188 & ~n35189 ;
  assign n35191 = n34805 & ~n34857 ;
  assign n35192 = ~n34841 & ~n35191 ;
  assign n35193 = ~n34787 & ~n35192 ;
  assign n35194 = ~n34833 & ~n34843 ;
  assign n35195 = ~n34841 & n35194 ;
  assign n35196 = n34819 & ~n35195 ;
  assign n35197 = ~n35193 & ~n35196 ;
  assign n35198 = n34793 & ~n35197 ;
  assign n35207 = ~n34847 & ~n34856 ;
  assign n35208 = n34787 & ~n35207 ;
  assign n35205 = ~n34819 & n34842 ;
  assign n35206 = n34819 & ~n35173 ;
  assign n35209 = ~n35205 & ~n35206 ;
  assign n35210 = ~n35208 & n35209 ;
  assign n35211 = ~n34793 & ~n35210 ;
  assign n35199 = n34812 & n34842 ;
  assign n35200 = ~n35178 & ~n35199 ;
  assign n35201 = ~n35181 & n35200 ;
  assign n35202 = ~n34793 & ~n35201 ;
  assign n35203 = ~n34824 & ~n35202 ;
  assign n35204 = ~n34787 & ~n35203 ;
  assign n35213 = n34793 & n35178 ;
  assign n35212 = n34805 & n34820 ;
  assign n35214 = ~n34848 & ~n35212 ;
  assign n35215 = ~n35213 & n35214 ;
  assign n35216 = n34787 & ~n35215 ;
  assign n35217 = ~n35204 & ~n35216 ;
  assign n35218 = ~n35211 & n35217 ;
  assign n35219 = ~n35198 & n35218 ;
  assign n35220 = ~\u1_L9_reg[4]/NET0131  & ~n35219 ;
  assign n35221 = \u1_L9_reg[4]/NET0131  & n35219 ;
  assign n35222 = ~n35220 & ~n35221 ;
  assign n35273 = decrypt_pad & ~\u1_uk_K_r9_reg[23]/NET0131  ;
  assign n35274 = ~decrypt_pad & ~\u1_uk_K_r9_reg[15]/NET0131  ;
  assign n35275 = ~n35273 & ~n35274 ;
  assign n35276 = \u1_R9_reg[32]/NET0131  & ~n35275 ;
  assign n35277 = ~\u1_R9_reg[32]/NET0131  & n35275 ;
  assign n35278 = ~n35276 & ~n35277 ;
  assign n35249 = decrypt_pad & ~\u1_uk_K_r9_reg[45]/NET0131  ;
  assign n35250 = ~decrypt_pad & ~\u1_uk_K_r9_reg[9]/NET0131  ;
  assign n35251 = ~n35249 & ~n35250 ;
  assign n35252 = \u1_R9_reg[31]/NET0131  & ~n35251 ;
  assign n35253 = ~\u1_R9_reg[31]/NET0131  & n35251 ;
  assign n35254 = ~n35252 & ~n35253 ;
  assign n35229 = decrypt_pad & ~\u1_uk_K_r9_reg[28]/NET0131  ;
  assign n35230 = ~decrypt_pad & ~\u1_uk_K_r9_reg[51]/NET0131  ;
  assign n35231 = ~n35229 & ~n35230 ;
  assign n35232 = \u1_R9_reg[29]/NET0131  & ~n35231 ;
  assign n35233 = ~\u1_R9_reg[29]/NET0131  & n35231 ;
  assign n35234 = ~n35232 & ~n35233 ;
  assign n35235 = decrypt_pad & ~\u1_uk_K_r9_reg[44]/NET0131  ;
  assign n35236 = ~decrypt_pad & ~\u1_uk_K_r9_reg[36]/NET0131  ;
  assign n35237 = ~n35235 & ~n35236 ;
  assign n35238 = \u1_R9_reg[1]/NET0131  & ~n35237 ;
  assign n35239 = ~\u1_R9_reg[1]/NET0131  & n35237 ;
  assign n35240 = ~n35238 & ~n35239 ;
  assign n35242 = decrypt_pad & ~\u1_uk_K_r9_reg[29]/NET0131  ;
  assign n35243 = ~decrypt_pad & ~\u1_uk_K_r9_reg[21]/NET0131  ;
  assign n35244 = ~n35242 & ~n35243 ;
  assign n35245 = \u1_R9_reg[30]/NET0131  & ~n35244 ;
  assign n35246 = ~\u1_R9_reg[30]/NET0131  & n35244 ;
  assign n35247 = ~n35245 & ~n35246 ;
  assign n35263 = ~n35240 & n35247 ;
  assign n35223 = decrypt_pad & ~\u1_uk_K_r9_reg[1]/NET0131  ;
  assign n35224 = ~decrypt_pad & ~\u1_uk_K_r9_reg[52]/NET0131  ;
  assign n35225 = ~n35223 & ~n35224 ;
  assign n35226 = \u1_R9_reg[28]/NET0131  & ~n35225 ;
  assign n35227 = ~\u1_R9_reg[28]/NET0131  & n35225 ;
  assign n35228 = ~n35226 & ~n35227 ;
  assign n35294 = ~n35228 & ~n35240 ;
  assign n35300 = ~n35263 & ~n35294 ;
  assign n35301 = n35234 & ~n35300 ;
  assign n35289 = n35228 & n35240 ;
  assign n35290 = ~n35247 & n35289 ;
  assign n35264 = n35228 & ~n35234 ;
  assign n35302 = ~n35247 & n35264 ;
  assign n35303 = ~n35290 & ~n35302 ;
  assign n35304 = ~n35301 & n35303 ;
  assign n35305 = n35254 & ~n35304 ;
  assign n35306 = ~n35234 & ~n35247 ;
  assign n35307 = ~n35228 & n35306 ;
  assign n35308 = ~n35254 & n35307 ;
  assign n35241 = n35234 & n35240 ;
  assign n35248 = n35241 & n35247 ;
  assign n35309 = ~n35228 & n35248 ;
  assign n35310 = ~n35308 & ~n35309 ;
  assign n35311 = ~n35305 & n35310 ;
  assign n35312 = n35278 & ~n35311 ;
  assign n35256 = n35234 & ~n35247 ;
  assign n35257 = ~n35240 & n35256 ;
  assign n35255 = ~n35247 & ~n35254 ;
  assign n35258 = ~n35248 & ~n35255 ;
  assign n35259 = ~n35257 & n35258 ;
  assign n35260 = n35228 & ~n35259 ;
  assign n35265 = n35263 & n35264 ;
  assign n35261 = ~n35234 & n35240 ;
  assign n35262 = ~n35228 & n35261 ;
  assign n35266 = n35254 & ~n35262 ;
  assign n35267 = ~n35265 & n35266 ;
  assign n35268 = ~n35228 & n35263 ;
  assign n35269 = ~n35241 & ~n35254 ;
  assign n35270 = ~n35268 & n35269 ;
  assign n35271 = ~n35267 & ~n35270 ;
  assign n35272 = ~n35260 & ~n35271 ;
  assign n35279 = ~n35272 & ~n35278 ;
  assign n35286 = n35234 & n35247 ;
  assign n35287 = ~n35228 & n35286 ;
  assign n35288 = ~n35240 & n35287 ;
  assign n35291 = ~n35234 & n35290 ;
  assign n35292 = ~n35288 & ~n35291 ;
  assign n35293 = n35247 & n35262 ;
  assign n35295 = ~n35234 & n35294 ;
  assign n35296 = ~n35247 & n35295 ;
  assign n35297 = ~n35293 & ~n35296 ;
  assign n35298 = n35292 & n35297 ;
  assign n35299 = n35254 & ~n35298 ;
  assign n35280 = n35247 & ~n35254 ;
  assign n35281 = n35264 & n35278 ;
  assign n35282 = n35280 & n35281 ;
  assign n35283 = n35228 & n35234 ;
  assign n35284 = ~n35240 & n35283 ;
  assign n35285 = n35255 & n35284 ;
  assign n35313 = ~n35282 & ~n35285 ;
  assign n35314 = ~n35299 & n35313 ;
  assign n35315 = ~n35279 & n35314 ;
  assign n35316 = ~n35312 & n35315 ;
  assign n35317 = \u1_L9_reg[5]/NET0131  & ~n35316 ;
  assign n35318 = ~\u1_L9_reg[5]/NET0131  & n35316 ;
  assign n35319 = ~n35317 & ~n35318 ;
  assign n35335 = n35000 & n35042 ;
  assign n35336 = n34979 & n35335 ;
  assign n35332 = n34986 & n35007 ;
  assign n35333 = ~n35024 & ~n35332 ;
  assign n35334 = n34992 & ~n35333 ;
  assign n35322 = n34986 & ~n35000 ;
  assign n35337 = ~n34992 & ~n35322 ;
  assign n35338 = n34980 & n35337 ;
  assign n35339 = ~n35005 & ~n35338 ;
  assign n35340 = ~n35334 & n35339 ;
  assign n35341 = ~n35336 & n35340 ;
  assign n35342 = n35022 & ~n35341 ;
  assign n35325 = n34992 & n35003 ;
  assign n35326 = ~n34973 & n35325 ;
  assign n35320 = n34973 & ~n35003 ;
  assign n35321 = n35006 & n35320 ;
  assign n35327 = ~n35047 & ~n35321 ;
  assign n35328 = ~n35326 & n35327 ;
  assign n35323 = ~n35004 & ~n35322 ;
  assign n35324 = n34973 & ~n35323 ;
  assign n35329 = n35029 & ~n35324 ;
  assign n35330 = n35328 & n35329 ;
  assign n35331 = ~n35022 & ~n35330 ;
  assign n35343 = ~n35026 & ~n35336 ;
  assign n35344 = ~n34992 & ~n35343 ;
  assign n35345 = ~n35001 & ~n35016 ;
  assign n35346 = ~n35344 & n35345 ;
  assign n35347 = ~n35331 & n35346 ;
  assign n35348 = ~n35342 & n35347 ;
  assign n35349 = ~\u1_L9_reg[10]/NET0131  & ~n35348 ;
  assign n35350 = \u1_L9_reg[10]/NET0131  & n35348 ;
  assign n35351 = ~n35349 & ~n35350 ;
  assign n35358 = ~n34922 & ~n34924 ;
  assign n35359 = n34933 & n35358 ;
  assign n35356 = ~n34919 & ~n34924 ;
  assign n35357 = n34935 & ~n35356 ;
  assign n35363 = ~n34881 & ~n35357 ;
  assign n35364 = ~n35359 & n35363 ;
  assign n35352 = n34906 & n34925 ;
  assign n35353 = n34899 & n34917 ;
  assign n35354 = ~n35352 & ~n35353 ;
  assign n35355 = ~n34893 & ~n35354 ;
  assign n35360 = ~n34900 & ~n34940 ;
  assign n35361 = ~n34917 & n35360 ;
  assign n35362 = ~n34914 & ~n35361 ;
  assign n35365 = ~n35355 & ~n35362 ;
  assign n35366 = n35364 & n35365 ;
  assign n35367 = ~n34914 & n34937 ;
  assign n35373 = n34881 & ~n34939 ;
  assign n35374 = ~n34954 & n35373 ;
  assign n35375 = ~n35367 & n35374 ;
  assign n35368 = ~n34916 & ~n34957 ;
  assign n35369 = n34945 & ~n35368 ;
  assign n35370 = n34893 & n34906 ;
  assign n35371 = ~n34934 & ~n35370 ;
  assign n35372 = n34914 & ~n35371 ;
  assign n35376 = ~n35369 & ~n35372 ;
  assign n35377 = n35375 & n35376 ;
  assign n35378 = ~n35366 & ~n35377 ;
  assign n35379 = \u1_L9_reg[12]/NET0131  & n35378 ;
  assign n35380 = ~\u1_L9_reg[12]/NET0131  & ~n35378 ;
  assign n35381 = ~n35379 & ~n35380 ;
  assign n35382 = n35072 & n35092 ;
  assign n35383 = n35066 & ~n35382 ;
  assign n35384 = ~n35091 & ~n35099 ;
  assign n35385 = ~n35137 & ~n35384 ;
  assign n35386 = n35383 & ~n35385 ;
  assign n35389 = ~n35072 & ~n35098 ;
  assign n35390 = n35106 & n35389 ;
  assign n35387 = n35066 & ~n35101 ;
  assign n35388 = n35111 & n35387 ;
  assign n35391 = ~n35121 & ~n35388 ;
  assign n35392 = ~n35390 & n35391 ;
  assign n35393 = ~n35386 & n35392 ;
  assign n35394 = ~n35136 & n35384 ;
  assign n35395 = ~n35066 & ~n35394 ;
  assign n35397 = n35078 & n35099 ;
  assign n35396 = ~n35078 & n35092 ;
  assign n35398 = n35066 & ~n35396 ;
  assign n35399 = ~n35397 & n35398 ;
  assign n35400 = ~n35395 & ~n35399 ;
  assign n35401 = n35101 & n35111 ;
  assign n35402 = ~n35126 & ~n35401 ;
  assign n35403 = n35091 & n35127 ;
  assign n35404 = ~n35078 & n35403 ;
  assign n35405 = n35121 & ~n35404 ;
  assign n35406 = n35110 & n35405 ;
  assign n35407 = n35402 & n35406 ;
  assign n35408 = ~n35400 & n35407 ;
  assign n35409 = ~n35393 & ~n35408 ;
  assign n35410 = n35079 & n35102 ;
  assign n35411 = ~n35403 & ~n35410 ;
  assign n35412 = ~n35138 & n35411 ;
  assign n35413 = ~n35121 & ~n35412 ;
  assign n35414 = n35402 & ~n35413 ;
  assign n35415 = ~n35066 & ~n35414 ;
  assign n35416 = ~n35409 & ~n35415 ;
  assign n35417 = ~\u1_L9_reg[13]/NET0131  & n35416 ;
  assign n35418 = \u1_L9_reg[13]/NET0131  & ~n35416 ;
  assign n35419 = ~n35417 & ~n35418 ;
  assign n35478 = decrypt_pad & ~\u1_uk_K_r9_reg[8]/NET0131  ;
  assign n35479 = ~decrypt_pad & ~\u1_uk_K_r9_reg[0]/P0001  ;
  assign n35480 = ~n35478 & ~n35479 ;
  assign n35481 = \u1_R9_reg[20]/NET0131  & ~n35480 ;
  assign n35482 = ~\u1_R9_reg[20]/NET0131  & n35480 ;
  assign n35483 = ~n35481 & ~n35482 ;
  assign n35452 = decrypt_pad & ~\u1_uk_K_r9_reg[52]/NET0131  ;
  assign n35453 = ~decrypt_pad & ~\u1_uk_K_r9_reg[16]/NET0131  ;
  assign n35454 = ~n35452 & ~n35453 ;
  assign n35455 = \u1_R9_reg[19]/NET0131  & ~n35454 ;
  assign n35456 = ~\u1_R9_reg[19]/NET0131  & n35454 ;
  assign n35457 = ~n35455 & ~n35456 ;
  assign n35433 = decrypt_pad & ~\u1_uk_K_r9_reg[21]/NET0131  ;
  assign n35434 = ~decrypt_pad & ~\u1_uk_K_r9_reg[44]/NET0131  ;
  assign n35435 = ~n35433 & ~n35434 ;
  assign n35436 = \u1_R9_reg[16]/NET0131  & ~n35435 ;
  assign n35437 = ~\u1_R9_reg[16]/NET0131  & n35435 ;
  assign n35438 = ~n35436 & ~n35437 ;
  assign n35426 = decrypt_pad & ~\u1_uk_K_r9_reg[9]/NET0131  ;
  assign n35427 = ~decrypt_pad & ~\u1_uk_K_r9_reg[1]/NET0131  ;
  assign n35428 = ~n35426 & ~n35427 ;
  assign n35429 = \u1_R9_reg[21]/NET0131  & ~n35428 ;
  assign n35430 = ~\u1_R9_reg[21]/NET0131  & n35428 ;
  assign n35431 = ~n35429 & ~n35430 ;
  assign n35441 = decrypt_pad & ~\u1_uk_K_r9_reg[43]/NET0131  ;
  assign n35442 = ~decrypt_pad & ~\u1_uk_K_r9_reg[35]/NET0131  ;
  assign n35443 = ~n35441 & ~n35442 ;
  assign n35444 = \u1_R9_reg[17]/NET0131  & ~n35443 ;
  assign n35445 = ~\u1_R9_reg[17]/NET0131  & n35443 ;
  assign n35446 = ~n35444 & ~n35445 ;
  assign n35465 = ~n35431 & n35446 ;
  assign n35500 = n35438 & n35465 ;
  assign n35420 = decrypt_pad & ~\u1_uk_K_r9_reg[37]/NET0131  ;
  assign n35421 = ~decrypt_pad & ~\u1_uk_K_r9_reg[29]/NET0131  ;
  assign n35422 = ~n35420 & ~n35421 ;
  assign n35423 = \u1_R9_reg[18]/NET0131  & ~n35422 ;
  assign n35424 = ~\u1_R9_reg[18]/NET0131  & n35422 ;
  assign n35425 = ~n35423 & ~n35424 ;
  assign n35447 = ~n35425 & n35446 ;
  assign n35486 = n35431 & ~n35438 ;
  assign n35498 = ~n35447 & n35486 ;
  assign n35469 = n35431 & n35438 ;
  assign n35499 = ~n35425 & n35469 ;
  assign n35501 = ~n35498 & ~n35499 ;
  assign n35502 = ~n35500 & n35501 ;
  assign n35503 = n35457 & ~n35502 ;
  assign n35485 = ~n35425 & ~n35457 ;
  assign n35439 = ~n35431 & ~n35438 ;
  assign n35458 = n35439 & ~n35446 ;
  assign n35487 = n35446 & n35486 ;
  assign n35488 = ~n35458 & ~n35487 ;
  assign n35489 = n35485 & ~n35488 ;
  assign n35470 = n35446 & n35469 ;
  assign n35494 = n35425 & ~n35457 ;
  assign n35495 = n35470 & n35494 ;
  assign n35490 = ~n35446 & n35469 ;
  assign n35491 = ~n35425 & n35490 ;
  assign n35492 = ~n35431 & n35438 ;
  assign n35493 = n35447 & n35492 ;
  assign n35496 = n35425 & ~n35446 ;
  assign n35497 = n35492 & n35496 ;
  assign n35504 = ~n35493 & ~n35497 ;
  assign n35505 = ~n35491 & n35504 ;
  assign n35506 = ~n35495 & n35505 ;
  assign n35507 = ~n35489 & n35506 ;
  assign n35508 = ~n35503 & n35507 ;
  assign n35509 = n35483 & ~n35508 ;
  assign n35432 = n35425 & n35431 ;
  assign n35440 = ~n35432 & ~n35439 ;
  assign n35448 = n35438 & ~n35446 ;
  assign n35449 = ~n35447 & ~n35448 ;
  assign n35450 = ~n35440 & ~n35449 ;
  assign n35451 = n35432 & n35438 ;
  assign n35460 = ~n35451 & n35457 ;
  assign n35459 = ~n35438 & n35447 ;
  assign n35461 = ~n35458 & ~n35459 ;
  assign n35462 = n35460 & n35461 ;
  assign n35471 = ~n35425 & n35470 ;
  assign n35463 = ~n35425 & ~n35431 ;
  assign n35464 = n35448 & n35463 ;
  assign n35472 = ~n35457 & ~n35464 ;
  assign n35466 = n35425 & n35465 ;
  assign n35467 = ~n35438 & ~n35446 ;
  assign n35468 = n35431 & n35467 ;
  assign n35473 = ~n35466 & ~n35468 ;
  assign n35474 = n35472 & n35473 ;
  assign n35475 = ~n35471 & n35474 ;
  assign n35476 = ~n35462 & ~n35475 ;
  assign n35477 = ~n35450 & ~n35476 ;
  assign n35484 = ~n35477 & ~n35483 ;
  assign n35510 = n35432 & n35467 ;
  assign n35511 = ~n35466 & ~n35510 ;
  assign n35512 = ~n35438 & ~n35511 ;
  assign n35513 = ~n35457 & n35512 ;
  assign n35514 = n35425 & n35458 ;
  assign n35515 = ~n35493 & ~n35514 ;
  assign n35516 = n35457 & ~n35515 ;
  assign n35517 = ~n35513 & ~n35516 ;
  assign n35518 = ~n35484 & n35517 ;
  assign n35519 = ~n35509 & n35518 ;
  assign n35520 = ~\u1_L9_reg[14]/NET0131  & ~n35519 ;
  assign n35521 = \u1_L9_reg[14]/NET0131  & n35519 ;
  assign n35522 = ~n35520 & ~n35521 ;
  assign n35523 = ~n35257 & ~n35283 ;
  assign n35524 = ~n35262 & n35523 ;
  assign n35525 = n35254 & ~n35524 ;
  assign n35526 = n35228 & ~n35240 ;
  assign n35527 = n35306 & n35526 ;
  assign n35528 = ~n35525 & ~n35527 ;
  assign n35529 = ~n35278 & ~n35528 ;
  assign n35531 = n35247 & n35264 ;
  assign n35545 = ~n35228 & n35240 ;
  assign n35546 = n35256 & n35545 ;
  assign n35547 = ~n35531 & ~n35546 ;
  assign n35548 = ~n35288 & n35547 ;
  assign n35549 = ~n35296 & n35548 ;
  assign n35550 = ~n35254 & ~n35549 ;
  assign n35530 = n35228 & n35256 ;
  assign n35534 = n35261 & n35280 ;
  assign n35535 = ~n35530 & ~n35534 ;
  assign n35536 = ~n35288 & n35535 ;
  assign n35532 = n35240 & n35531 ;
  assign n35533 = n35254 & n35295 ;
  assign n35537 = ~n35532 & ~n35533 ;
  assign n35538 = n35536 & n35537 ;
  assign n35539 = n35278 & ~n35538 ;
  assign n35540 = n35240 & n35307 ;
  assign n35541 = ~n35309 & ~n35540 ;
  assign n35542 = n35254 & ~n35541 ;
  assign n35543 = ~n35254 & ~n35278 ;
  assign n35544 = n35264 & n35543 ;
  assign n35551 = ~n35542 & ~n35544 ;
  assign n35552 = ~n35539 & n35551 ;
  assign n35553 = ~n35550 & n35552 ;
  assign n35554 = ~n35529 & n35553 ;
  assign n35555 = ~\u1_L9_reg[15]/P0001  & ~n35554 ;
  assign n35556 = \u1_L9_reg[15]/P0001  & n35554 ;
  assign n35557 = ~n35555 & ~n35556 ;
  assign n35558 = ~n34979 & n35335 ;
  assign n35559 = ~n34992 & ~n35558 ;
  assign n35560 = ~n35000 & n35023 ;
  assign n35561 = ~n35012 & ~n35560 ;
  assign n35562 = n35022 & ~n35561 ;
  assign n35563 = n34992 & ~n35028 ;
  assign n35564 = ~n35336 & n35563 ;
  assign n35565 = ~n35562 & n35564 ;
  assign n35566 = ~n35559 & ~n35565 ;
  assign n35567 = ~n35030 & n35335 ;
  assign n35568 = n34986 & ~n34992 ;
  assign n35569 = ~n35027 & n35568 ;
  assign n35570 = ~n35320 & n35569 ;
  assign n35571 = n35022 & ~n35570 ;
  assign n35572 = ~n35567 & n35571 ;
  assign n35576 = n34986 & n35003 ;
  assign n35577 = n34973 & ~n35006 ;
  assign n35578 = ~n35027 & n35577 ;
  assign n35579 = ~n35576 & n35578 ;
  assign n35573 = n35023 & n35027 ;
  assign n35574 = ~n35008 & ~n35573 ;
  assign n35575 = n34992 & ~n35574 ;
  assign n35580 = ~n35022 & ~n35038 ;
  assign n35581 = ~n35575 & n35580 ;
  assign n35582 = ~n35579 & n35581 ;
  assign n35583 = ~n35572 & ~n35582 ;
  assign n35584 = ~n35566 & ~n35583 ;
  assign n35585 = ~\u1_L9_reg[1]/NET0131  & ~n35584 ;
  assign n35586 = \u1_L9_reg[1]/NET0131  & n35584 ;
  assign n35587 = ~n35585 & ~n35586 ;
  assign n35588 = ~n34831 & ~n34841 ;
  assign n35589 = ~n34793 & ~n35588 ;
  assign n35590 = ~n34854 & ~n35589 ;
  assign n35591 = ~n34819 & ~n35590 ;
  assign n35596 = ~n34793 & ~n35194 ;
  assign n35592 = n34799 & ~n34846 ;
  assign n35593 = ~n35199 & ~n35592 ;
  assign n35594 = n34793 & ~n35593 ;
  assign n35595 = n34813 & n34819 ;
  assign n35597 = ~n34787 & ~n35595 ;
  assign n35598 = ~n35594 & n35597 ;
  assign n35599 = ~n35596 & n35598 ;
  assign n35601 = ~n34793 & n34830 ;
  assign n35604 = n34787 & ~n34847 ;
  assign n35605 = ~n35601 & n35604 ;
  assign n35606 = ~n34850 & n35605 ;
  assign n35600 = n34819 & ~n35194 ;
  assign n35602 = ~n34849 & ~n34859 ;
  assign n35603 = n34793 & ~n35602 ;
  assign n35607 = ~n35600 & ~n35603 ;
  assign n35608 = n35606 & n35607 ;
  assign n35609 = ~n35599 & ~n35608 ;
  assign n35610 = ~n35591 & ~n35609 ;
  assign n35611 = ~\u1_L9_reg[19]/NET0131  & ~n35610 ;
  assign n35612 = \u1_L9_reg[19]/NET0131  & n35610 ;
  assign n35613 = ~n35611 & ~n35612 ;
  assign n35616 = n35228 & n35286 ;
  assign n35614 = n35240 & n35306 ;
  assign n35615 = ~n35228 & n35241 ;
  assign n35617 = ~n35614 & ~n35615 ;
  assign n35618 = ~n35616 & n35617 ;
  assign n35619 = n35254 & ~n35618 ;
  assign n35622 = ~n35526 & ~n35531 ;
  assign n35623 = ~n35254 & ~n35263 ;
  assign n35624 = ~n35622 & n35623 ;
  assign n35620 = ~n35284 & ~n35295 ;
  assign n35621 = n35247 & ~n35620 ;
  assign n35625 = ~n35540 & ~n35621 ;
  assign n35626 = ~n35624 & n35625 ;
  assign n35627 = ~n35619 & n35626 ;
  assign n35628 = n35278 & ~n35627 ;
  assign n35638 = ~n35265 & ~n35287 ;
  assign n35633 = n35280 & n35545 ;
  assign n35634 = n35234 & ~n35254 ;
  assign n35635 = n35294 & n35634 ;
  assign n35639 = ~n35633 & ~n35635 ;
  assign n35640 = n35638 & n35639 ;
  assign n35636 = ~n35234 & n35254 ;
  assign n35637 = n35290 & ~n35636 ;
  assign n35641 = ~n35296 & ~n35637 ;
  assign n35642 = n35640 & n35641 ;
  assign n35643 = ~n35278 & ~n35642 ;
  assign n35629 = ~n35284 & ~n35531 ;
  assign n35630 = ~n35278 & ~n35629 ;
  assign n35631 = ~n35307 & ~n35630 ;
  assign n35632 = n35254 & ~n35631 ;
  assign n35644 = n35228 & n35241 ;
  assign n35645 = n35255 & n35644 ;
  assign n35646 = ~n35632 & ~n35645 ;
  assign n35647 = ~n35643 & n35646 ;
  assign n35648 = ~n35628 & n35647 ;
  assign n35649 = ~\u1_L9_reg[21]/NET0131  & ~n35648 ;
  assign n35650 = \u1_L9_reg[21]/NET0131  & n35648 ;
  assign n35651 = ~n35649 & ~n35650 ;
  assign n35668 = n34708 & n34727 ;
  assign n35669 = ~n34766 & ~n35668 ;
  assign n35670 = ~n34695 & ~n35669 ;
  assign n35673 = ~n34714 & ~n34730 ;
  assign n35674 = ~n34735 & ~n35668 ;
  assign n35675 = n35673 & n35674 ;
  assign n35671 = n34701 & n34727 ;
  assign n35672 = n34714 & n35671 ;
  assign n35667 = n34702 & n34753 ;
  assign n35676 = ~n34747 & ~n35667 ;
  assign n35677 = ~n35672 & n35676 ;
  assign n35678 = ~n35675 & n35677 ;
  assign n35679 = ~n35670 & n35678 ;
  assign n35652 = n34695 & n34727 ;
  assign n35681 = ~n34719 & n35652 ;
  assign n35682 = n34717 & n35681 ;
  assign n35680 = n34729 & n34734 ;
  assign n35683 = n34747 & ~n35680 ;
  assign n35684 = ~n34765 & n35683 ;
  assign n35685 = ~n35682 & n35684 ;
  assign n35686 = ~n35679 & ~n35685 ;
  assign n35654 = ~n34714 & n34727 ;
  assign n35655 = ~n34734 & ~n35654 ;
  assign n35659 = ~n34708 & ~n35655 ;
  assign n35660 = n34708 & n35655 ;
  assign n35661 = ~n35659 & ~n35660 ;
  assign n35662 = ~n34736 & n34747 ;
  assign n35663 = ~n35661 & n35662 ;
  assign n35656 = n34717 & ~n35655 ;
  assign n35657 = ~n34701 & n35656 ;
  assign n35658 = n34727 & n34766 ;
  assign n35664 = ~n35657 & ~n35658 ;
  assign n35665 = ~n35663 & n35664 ;
  assign n35666 = ~n34695 & ~n35665 ;
  assign n35653 = n34720 & n35652 ;
  assign n35687 = ~n34774 & ~n35653 ;
  assign n35688 = ~n35666 & n35687 ;
  assign n35689 = ~n35686 & n35688 ;
  assign n35690 = \u1_L9_reg[23]/NET0131  & ~n35689 ;
  assign n35691 = ~\u1_L9_reg[23]/NET0131  & n35689 ;
  assign n35692 = ~n35690 & ~n35691 ;
  assign n35693 = ~n35439 & ~n35463 ;
  assign n35694 = ~n35467 & n35693 ;
  assign n35695 = ~n35447 & ~n35694 ;
  assign n35696 = ~n35470 & ~n35695 ;
  assign n35697 = n35457 & ~n35696 ;
  assign n35698 = ~n35459 & ~n35490 ;
  assign n35699 = ~n35457 & ~n35698 ;
  assign n35700 = n35446 & ~n35463 ;
  assign n35701 = n35440 & n35700 ;
  assign n35702 = ~n35699 & ~n35701 ;
  assign n35703 = ~n35697 & n35702 ;
  assign n35704 = n35483 & ~n35703 ;
  assign n35718 = ~n35458 & ~n35500 ;
  assign n35719 = n35425 & ~n35718 ;
  assign n35720 = ~n35425 & n35468 ;
  assign n35721 = ~n35719 & ~n35720 ;
  assign n35722 = n35457 & ~n35721 ;
  assign n35705 = ~n35431 & n35457 ;
  assign n35706 = ~n35431 & n35448 ;
  assign n35707 = n35425 & ~n35438 ;
  assign n35708 = n35446 & n35707 ;
  assign n35709 = ~n35706 & ~n35708 ;
  assign n35710 = ~n35705 & ~n35709 ;
  assign n35712 = n35457 & ~n35465 ;
  assign n35711 = ~n35457 & ~n35467 ;
  assign n35713 = ~n35425 & ~n35711 ;
  assign n35714 = ~n35712 & n35713 ;
  assign n35715 = ~n35710 & ~n35714 ;
  assign n35716 = ~n35483 & ~n35715 ;
  assign n35717 = n35448 & n35494 ;
  assign n35723 = ~n35471 & ~n35717 ;
  assign n35724 = ~n35716 & n35723 ;
  assign n35725 = ~n35722 & n35724 ;
  assign n35726 = ~n35704 & n35725 ;
  assign n35727 = ~\u1_L9_reg[25]/NET0131  & ~n35726 ;
  assign n35728 = \u1_L9_reg[25]/NET0131  & n35726 ;
  assign n35729 = ~n35727 & ~n35728 ;
  assign n35748 = ~n34979 & ~n35042 ;
  assign n35749 = ~n35045 & ~n35748 ;
  assign n35750 = ~n35000 & ~n35749 ;
  assign n35730 = n34979 & ~n35015 ;
  assign n35751 = ~n34986 & ~n35022 ;
  assign n35752 = ~n35730 & n35751 ;
  assign n35753 = ~n35750 & ~n35752 ;
  assign n35754 = ~n34992 & ~n35753 ;
  assign n35734 = n34986 & ~n35010 ;
  assign n35731 = n34973 & ~n35000 ;
  assign n35732 = n35337 & ~n35731 ;
  assign n35733 = n35730 & n35732 ;
  assign n35735 = n35000 & n35040 ;
  assign n35736 = ~n35046 & n35735 ;
  assign n35737 = n35022 & ~n35025 ;
  assign n35738 = ~n35736 & n35737 ;
  assign n35739 = ~n35733 & n35738 ;
  assign n35740 = ~n35734 & n35739 ;
  assign n35741 = n34993 & n35000 ;
  assign n35742 = ~n35040 & n35741 ;
  assign n35743 = ~n35022 & ~n35560 ;
  assign n35744 = n35039 & n35743 ;
  assign n35745 = ~n35742 & n35744 ;
  assign n35746 = ~n35740 & ~n35745 ;
  assign n35747 = ~n35042 & n35325 ;
  assign n35755 = ~n35746 & ~n35747 ;
  assign n35756 = ~n35754 & n35755 ;
  assign n35757 = ~\u1_L9_reg[26]/NET0131  & ~n35756 ;
  assign n35758 = \u1_L9_reg[26]/NET0131  & n35756 ;
  assign n35759 = ~n35757 & ~n35758 ;
  assign n35760 = ~n35078 & n35127 ;
  assign n35761 = ~n35108 & ~n35760 ;
  assign n35762 = n35066 & n35761 ;
  assign n35763 = ~n35072 & n35146 ;
  assign n35764 = ~n35066 & ~n35763 ;
  assign n35765 = ~n35103 & ~n35130 ;
  assign n35766 = ~n35137 & n35765 ;
  assign n35767 = n35764 & n35766 ;
  assign n35768 = ~n35762 & ~n35767 ;
  assign n35769 = ~n35132 & n35146 ;
  assign n35770 = ~n35121 & ~n35401 ;
  assign n35771 = ~n35769 & n35770 ;
  assign n35772 = ~n35768 & n35771 ;
  assign n35773 = n35091 & ~n35136 ;
  assign n35774 = ~n35132 & n35773 ;
  assign n35775 = n35383 & ~n35774 ;
  assign n35776 = ~n35401 & n35761 ;
  assign n35777 = n35764 & n35776 ;
  assign n35778 = ~n35775 & ~n35777 ;
  assign n35779 = n35094 & ~n35112 ;
  assign n35780 = n35121 & ~n35410 ;
  assign n35781 = ~n35779 & n35780 ;
  assign n35782 = ~n35778 & n35781 ;
  assign n35783 = ~n35772 & ~n35782 ;
  assign n35784 = ~\u1_L9_reg[28]/NET0131  & n35783 ;
  assign n35785 = \u1_L9_reg[28]/NET0131  & ~n35783 ;
  assign n35786 = ~n35784 & ~n35785 ;
  assign n35800 = ~n35425 & n35458 ;
  assign n35801 = ~n35490 & ~n35800 ;
  assign n35802 = n35457 & ~n35801 ;
  assign n35803 = n35438 & n35485 ;
  assign n35804 = ~n35512 & ~n35803 ;
  assign n35805 = ~n35802 & n35804 ;
  assign n35806 = n35483 & ~n35805 ;
  assign n35791 = n35457 & ~n35464 ;
  assign n35792 = ~n35470 & n35791 ;
  assign n35793 = n35486 & ~n35496 ;
  assign n35794 = ~n35457 & ~n35490 ;
  assign n35795 = ~n35793 & n35794 ;
  assign n35796 = ~n35792 & ~n35795 ;
  assign n35797 = ~n35459 & ~n35719 ;
  assign n35798 = ~n35796 & n35797 ;
  assign n35799 = ~n35483 & ~n35798 ;
  assign n35787 = n35447 & n35486 ;
  assign n35788 = n35511 & ~n35787 ;
  assign n35789 = n35457 & ~n35788 ;
  assign n35790 = ~n35431 & n35717 ;
  assign n35807 = ~n35789 & ~n35790 ;
  assign n35808 = ~n35799 & n35807 ;
  assign n35809 = ~n35806 & n35808 ;
  assign n35810 = ~\u1_L9_reg[8]/NET0131  & ~n35809 ;
  assign n35811 = \u1_L9_reg[8]/NET0131  & n35809 ;
  assign n35812 = ~n35810 & ~n35811 ;
  assign n35813 = ~n35284 & ~n35307 ;
  assign n35814 = ~n35615 & n35813 ;
  assign n35815 = ~n35254 & ~n35814 ;
  assign n35816 = n35254 & ~n35526 ;
  assign n35817 = ~n35523 & n35816 ;
  assign n35818 = ~n35265 & ~n35614 ;
  assign n35819 = ~n35309 & n35818 ;
  assign n35820 = ~n35817 & n35819 ;
  assign n35821 = ~n35815 & n35820 ;
  assign n35822 = n35278 & ~n35821 ;
  assign n35825 = n35254 & ~n35257 ;
  assign n35824 = n35240 & ~n35256 ;
  assign n35826 = ~n35287 & ~n35824 ;
  assign n35827 = n35825 & n35826 ;
  assign n35823 = n35280 & n35289 ;
  assign n35828 = ~n35635 & ~n35823 ;
  assign n35829 = ~n35293 & n35828 ;
  assign n35830 = ~n35827 & n35829 ;
  assign n35831 = ~n35278 & ~n35830 ;
  assign n35833 = ~n35254 & ~n35292 ;
  assign n35832 = n35263 & n35636 ;
  assign n35834 = ~n35285 & ~n35832 ;
  assign n35835 = ~n35833 & n35834 ;
  assign n35836 = ~n35831 & n35835 ;
  assign n35837 = ~n35822 & n35836 ;
  assign n35838 = ~\u1_L9_reg[27]/NET0131  & ~n35837 ;
  assign n35839 = \u1_L9_reg[27]/NET0131  & n35837 ;
  assign n35840 = ~n35838 & ~n35839 ;
  assign n35841 = ~n35510 & n35791 ;
  assign n35842 = ~n35485 & ~n35794 ;
  assign n35843 = ~n35425 & ~n35718 ;
  assign n35844 = ~n35842 & ~n35843 ;
  assign n35845 = ~n35841 & ~n35844 ;
  assign n35847 = n35440 & n35794 ;
  assign n35848 = ~n35425 & n35486 ;
  assign n35849 = n35457 & ~n35500 ;
  assign n35850 = ~n35848 & n35849 ;
  assign n35851 = ~n35847 & ~n35850 ;
  assign n35846 = ~n35492 & n35496 ;
  assign n35852 = ~n35483 & ~n35846 ;
  assign n35853 = ~n35851 & n35852 ;
  assign n35854 = n35439 & n35446 ;
  assign n35855 = ~n35499 & ~n35854 ;
  assign n35856 = n35457 & ~n35855 ;
  assign n35857 = ~n35457 & n35487 ;
  assign n35858 = n35483 & ~n35497 ;
  assign n35859 = ~n35471 & n35858 ;
  assign n35860 = ~n35857 & n35859 ;
  assign n35861 = ~n35856 & n35860 ;
  assign n35862 = ~n35853 & ~n35861 ;
  assign n35863 = ~n35845 & ~n35862 ;
  assign n35864 = ~\u1_L9_reg[3]/NET0131  & ~n35863 ;
  assign n35865 = \u1_L9_reg[3]/NET0131  & n35863 ;
  assign n35866 = ~n35864 & ~n35865 ;
  assign n35901 = decrypt_pad & ~\u1_uk_K_r9_reg[46]/NET0131  ;
  assign n35902 = ~decrypt_pad & ~\u1_uk_K_r9_reg[40]/NET0131  ;
  assign n35903 = ~n35901 & ~n35902 ;
  assign n35904 = \u1_R9_reg[11]/NET0131  & ~n35903 ;
  assign n35905 = ~\u1_R9_reg[11]/NET0131  & n35903 ;
  assign n35906 = ~n35904 & ~n35905 ;
  assign n35893 = decrypt_pad & ~\u1_uk_K_r9_reg[4]/NET0131  ;
  assign n35894 = ~decrypt_pad & ~\u1_uk_K_r9_reg[55]/NET0131  ;
  assign n35895 = ~n35893 & ~n35894 ;
  assign n35896 = \u1_R9_reg[12]/NET0131  & ~n35895 ;
  assign n35897 = ~\u1_R9_reg[12]/NET0131  & n35895 ;
  assign n35898 = ~n35896 & ~n35897 ;
  assign n35886 = decrypt_pad & ~\u1_uk_K_r9_reg[20]/NET0131  ;
  assign n35887 = ~decrypt_pad & ~\u1_uk_K_r9_reg[39]/NET0131  ;
  assign n35888 = ~n35886 & ~n35887 ;
  assign n35889 = \u1_R9_reg[10]/NET0131  & ~n35888 ;
  assign n35890 = ~\u1_R9_reg[10]/NET0131  & n35888 ;
  assign n35891 = ~n35889 & ~n35890 ;
  assign n35867 = decrypt_pad & ~\u1_uk_K_r9_reg[40]/NET0131  ;
  assign n35868 = ~decrypt_pad & ~\u1_uk_K_r9_reg[34]/NET0131  ;
  assign n35869 = ~n35867 & ~n35868 ;
  assign n35870 = \u1_R9_reg[8]/NET0131  & ~n35869 ;
  assign n35871 = ~\u1_R9_reg[8]/NET0131  & n35869 ;
  assign n35872 = ~n35870 & ~n35871 ;
  assign n35873 = decrypt_pad & ~\u1_uk_K_r9_reg[17]/NET0131  ;
  assign n35874 = ~decrypt_pad & ~\u1_uk_K_r9_reg[11]/NET0131  ;
  assign n35875 = ~n35873 & ~n35874 ;
  assign n35876 = \u1_R9_reg[13]/NET0131  & ~n35875 ;
  assign n35877 = ~\u1_R9_reg[13]/NET0131  & n35875 ;
  assign n35878 = ~n35876 & ~n35877 ;
  assign n35912 = ~n35872 & n35878 ;
  assign n35913 = n35891 & n35912 ;
  assign n35880 = decrypt_pad & ~\u1_uk_K_r9_reg[12]/NET0131  ;
  assign n35881 = ~decrypt_pad & ~\u1_uk_K_r9_reg[6]/NET0131  ;
  assign n35882 = ~n35880 & ~n35881 ;
  assign n35883 = \u1_R9_reg[9]/NET0131  & ~n35882 ;
  assign n35884 = ~\u1_R9_reg[9]/NET0131  & n35882 ;
  assign n35885 = ~n35883 & ~n35884 ;
  assign n35910 = n35872 & ~n35878 ;
  assign n35911 = n35885 & n35910 ;
  assign n35914 = n35878 & ~n35885 ;
  assign n35915 = ~n35911 & ~n35914 ;
  assign n35916 = ~n35913 & n35915 ;
  assign n35917 = n35898 & ~n35916 ;
  assign n35907 = ~n35872 & ~n35891 ;
  assign n35908 = ~n35878 & n35907 ;
  assign n35909 = ~n35885 & n35908 ;
  assign n35918 = n35891 & n35914 ;
  assign n35919 = ~n35909 & ~n35918 ;
  assign n35920 = ~n35917 & n35919 ;
  assign n35921 = n35906 & ~n35920 ;
  assign n35922 = n35878 & n35906 ;
  assign n35928 = n35885 & n35922 ;
  assign n35923 = ~n35910 & ~n35912 ;
  assign n35892 = n35885 & n35891 ;
  assign n35925 = ~n35885 & ~n35891 ;
  assign n35926 = ~n35892 & ~n35925 ;
  assign n35929 = ~n35923 & n35926 ;
  assign n35930 = ~n35928 & n35929 ;
  assign n35924 = ~n35922 & ~n35923 ;
  assign n35927 = ~n35924 & ~n35926 ;
  assign n35931 = ~n35898 & ~n35927 ;
  assign n35932 = ~n35930 & n35931 ;
  assign n35879 = ~n35872 & ~n35878 ;
  assign n35899 = n35892 & n35898 ;
  assign n35900 = n35879 & n35899 ;
  assign n35933 = n35885 & ~n35891 ;
  assign n35934 = n35872 & ~n35914 ;
  assign n35935 = ~n35933 & ~n35934 ;
  assign n35936 = ~n35878 & n35885 ;
  assign n35937 = n35898 & ~n35906 ;
  assign n35938 = ~n35936 & n35937 ;
  assign n35939 = ~n35935 & n35938 ;
  assign n35940 = ~n35900 & ~n35939 ;
  assign n35941 = ~n35932 & n35940 ;
  assign n35942 = ~n35921 & n35941 ;
  assign n35943 = ~\u1_L9_reg[6]/NET0131  & ~n35942 ;
  assign n35944 = \u1_L9_reg[6]/NET0131  & n35942 ;
  assign n35945 = ~n35943 & ~n35944 ;
  assign n35948 = n34701 & ~n35661 ;
  assign n35946 = ~n34716 & n35655 ;
  assign n35947 = n34754 & n35946 ;
  assign n35949 = n34719 & n35668 ;
  assign n35950 = n34747 & ~n35949 ;
  assign n35951 = ~n35947 & n35950 ;
  assign n35952 = ~n35948 & n35951 ;
  assign n35953 = ~n34695 & n35946 ;
  assign n35960 = ~n34747 & ~n35953 ;
  assign n35954 = ~n34717 & ~n35671 ;
  assign n35955 = ~n34701 & ~n35668 ;
  assign n35956 = n35954 & ~n35955 ;
  assign n35957 = ~n34714 & n34729 ;
  assign n35958 = n34695 & ~n35655 ;
  assign n35959 = ~n35957 & n35958 ;
  assign n35961 = ~n35956 & ~n35959 ;
  assign n35962 = n35960 & n35961 ;
  assign n35963 = ~n35952 & ~n35962 ;
  assign n35964 = n34714 & n34730 ;
  assign n35965 = ~n34757 & n35964 ;
  assign n35966 = ~n35963 & ~n35965 ;
  assign n35967 = ~\u1_L9_reg[9]/NET0131  & ~n35966 ;
  assign n35968 = \u1_L9_reg[9]/NET0131  & n35966 ;
  assign n35969 = ~n35967 & ~n35968 ;
  assign n35975 = ~n34935 & ~n34956 ;
  assign n35977 = ~n34922 & n35360 ;
  assign n35978 = n35975 & ~n35977 ;
  assign n35976 = ~n34922 & ~n35975 ;
  assign n35979 = ~n34914 & ~n35976 ;
  assign n35980 = ~n35978 & n35979 ;
  assign n35970 = n34924 & n34956 ;
  assign n35971 = n34887 & ~n34956 ;
  assign n35972 = n34945 & ~n35971 ;
  assign n35973 = ~n34907 & ~n35972 ;
  assign n35974 = n34914 & ~n35973 ;
  assign n35981 = ~n35970 & ~n35974 ;
  assign n35982 = ~n35980 & n35981 ;
  assign n35983 = n34881 & ~n35982 ;
  assign n35985 = ~n35352 & ~n35360 ;
  assign n35986 = ~n34914 & ~n35985 ;
  assign n35987 = ~n34893 & n34938 ;
  assign n35988 = n34914 & ~n35352 ;
  assign n35989 = ~n35987 & n35988 ;
  assign n35990 = ~n35986 & ~n35989 ;
  assign n35984 = n34893 & ~n35354 ;
  assign n35991 = n34955 & ~n35984 ;
  assign n35992 = ~n35990 & n35991 ;
  assign n35993 = ~n34881 & ~n35992 ;
  assign n35994 = n34914 & n34937 ;
  assign n35995 = ~n34925 & n34952 ;
  assign n35996 = n34918 & n35995 ;
  assign n35997 = ~n35994 & ~n35996 ;
  assign n35998 = ~n35993 & n35997 ;
  assign n35999 = ~n35983 & n35998 ;
  assign n36000 = \u1_L9_reg[32]/NET0131  & n35999 ;
  assign n36001 = ~\u1_L9_reg[32]/NET0131  & ~n35999 ;
  assign n36002 = ~n36000 & ~n36001 ;
  assign n36020 = ~n34906 & ~n35358 ;
  assign n36003 = n34893 & ~n35975 ;
  assign n36021 = n34887 & n34956 ;
  assign n36022 = ~n36003 & ~n36021 ;
  assign n36023 = ~n36020 & n36022 ;
  assign n36024 = ~n34914 & ~n36023 ;
  assign n36004 = ~n35987 & ~n36003 ;
  assign n36005 = n34887 & ~n36004 ;
  assign n36014 = ~n34887 & ~n34900 ;
  assign n36015 = n35975 & n36014 ;
  assign n36025 = n34914 & n36015 ;
  assign n36026 = ~n36005 & ~n36025 ;
  assign n36027 = ~n36024 & n36026 ;
  assign n36028 = n34881 & ~n36027 ;
  assign n36006 = ~n34914 & n36005 ;
  assign n36007 = n34881 & ~n34914 ;
  assign n36008 = n34944 & ~n35975 ;
  assign n36009 = n34899 & ~n35370 ;
  assign n36010 = n34914 & n35971 ;
  assign n36011 = ~n36009 & n36010 ;
  assign n36012 = ~n36008 & ~n36011 ;
  assign n36013 = ~n34881 & ~n36012 ;
  assign n36016 = ~n34914 & n36015 ;
  assign n36017 = ~n34908 & ~n36016 ;
  assign n36018 = ~n36013 & n36017 ;
  assign n36019 = ~n36007 & ~n36018 ;
  assign n36029 = ~n36006 & ~n36019 ;
  assign n36030 = ~n36028 & n36029 ;
  assign n36031 = ~\u1_L9_reg[7]/NET0131  & ~n36030 ;
  assign n36032 = \u1_L9_reg[7]/NET0131  & n36030 ;
  assign n36033 = ~n36031 & ~n36032 ;
  assign n36062 = n35879 & n35885 ;
  assign n36063 = n35906 & n36062 ;
  assign n36035 = n35872 & n35878 ;
  assign n36036 = n35885 & n36035 ;
  assign n36037 = ~n35885 & n35912 ;
  assign n36038 = ~n36036 & ~n36037 ;
  assign n36064 = ~n35885 & n35910 ;
  assign n36065 = n36038 & ~n36064 ;
  assign n36066 = ~n36063 & n36065 ;
  assign n36067 = ~n35891 & ~n36066 ;
  assign n36057 = n35885 & n35912 ;
  assign n36058 = n35891 & n36057 ;
  assign n36047 = ~n35885 & n35891 ;
  assign n36050 = n35879 & n36047 ;
  assign n36051 = n35906 & ~n36050 ;
  assign n36052 = n35872 & n35891 ;
  assign n36059 = ~n35878 & ~n35907 ;
  assign n36060 = ~n36052 & n36059 ;
  assign n36061 = ~n36051 & n36060 ;
  assign n36068 = ~n36058 & ~n36061 ;
  assign n36069 = ~n36067 & n36068 ;
  assign n36070 = n35898 & ~n36069 ;
  assign n36034 = n35906 & ~n35909 ;
  assign n36039 = ~n35908 & n36038 ;
  assign n36040 = ~n36034 & ~n36039 ;
  assign n36041 = ~n35885 & ~n36035 ;
  assign n36042 = ~n35879 & n35906 ;
  assign n36043 = ~n36036 & n36042 ;
  assign n36044 = ~n36041 & n36043 ;
  assign n36045 = ~n36040 & ~n36044 ;
  assign n36046 = ~n35898 & ~n36045 ;
  assign n36048 = n35872 & n36047 ;
  assign n36049 = ~n35906 & ~n36048 ;
  assign n36053 = n35885 & n36052 ;
  assign n36054 = ~n35878 & n36053 ;
  assign n36055 = n36051 & ~n36054 ;
  assign n36056 = ~n36049 & ~n36055 ;
  assign n36071 = ~n36046 & ~n36056 ;
  assign n36072 = ~n36070 & n36071 ;
  assign n36073 = ~\u1_L9_reg[16]/NET0131  & ~n36072 ;
  assign n36074 = \u1_L9_reg[16]/NET0131  & n36072 ;
  assign n36075 = ~n36073 & ~n36074 ;
  assign n36085 = n35066 & ~n35104 ;
  assign n36086 = ~n35092 & ~n35106 ;
  assign n36087 = ~n35066 & n35072 ;
  assign n36088 = ~n36086 & n36087 ;
  assign n36089 = ~n35093 & ~n36088 ;
  assign n36090 = ~n36085 & n36089 ;
  assign n36091 = n35121 & ~n36090 ;
  assign n36079 = n35091 & ~n35129 ;
  assign n36080 = n35147 & ~n36079 ;
  assign n36077 = ~n35135 & ~n35146 ;
  assign n36078 = n35131 & ~n36077 ;
  assign n36081 = ~n35396 & ~n35401 ;
  assign n36082 = ~n36078 & n36081 ;
  assign n36083 = ~n36080 & n36082 ;
  assign n36084 = ~n35121 & ~n36083 ;
  assign n36076 = ~n35066 & n35108 ;
  assign n36092 = n35085 & n35111 ;
  assign n36093 = ~n35404 & ~n36092 ;
  assign n36094 = n35066 & ~n36093 ;
  assign n36095 = ~n36076 & ~n36094 ;
  assign n36096 = ~n36084 & n36095 ;
  assign n36097 = ~n36091 & n36096 ;
  assign n36098 = \u1_L9_reg[18]/P0001  & n36097 ;
  assign n36099 = ~\u1_L9_reg[18]/P0001  & ~n36097 ;
  assign n36100 = ~n36098 & ~n36099 ;
  assign n36103 = ~n35891 & ~n35936 ;
  assign n36104 = ~n35923 & ~n36103 ;
  assign n36105 = ~n35912 & n35925 ;
  assign n36106 = ~n35910 & n36105 ;
  assign n36107 = ~n36104 & ~n36106 ;
  assign n36108 = ~n35898 & ~n36107 ;
  assign n36109 = ~n35906 & ~n36108 ;
  assign n36110 = ~n36057 & ~n36064 ;
  assign n36111 = ~n35891 & ~n36110 ;
  assign n36113 = ~n35891 & n35912 ;
  assign n36112 = n35879 & n35891 ;
  assign n36114 = n35906 & ~n36112 ;
  assign n36115 = ~n36113 & n36114 ;
  assign n36116 = ~n36048 & ~n36062 ;
  assign n36117 = n36115 & n36116 ;
  assign n36118 = ~n35898 & ~n36117 ;
  assign n36119 = ~n36111 & ~n36118 ;
  assign n36120 = ~n36109 & ~n36119 ;
  assign n36101 = n35891 & ~n35906 ;
  assign n36102 = n36036 & n36101 ;
  assign n36122 = ~n35913 & ~n36053 ;
  assign n36123 = ~n36105 & n36122 ;
  assign n36124 = n35906 & ~n36123 ;
  assign n36121 = n35924 & n35925 ;
  assign n36125 = ~n35906 & ~n35925 ;
  assign n36126 = n35923 & n36125 ;
  assign n36127 = ~n36121 & ~n36126 ;
  assign n36128 = ~n36124 & n36127 ;
  assign n36129 = n35898 & ~n36128 ;
  assign n36130 = ~n36102 & ~n36129 ;
  assign n36131 = ~n36120 & n36130 ;
  assign n36132 = ~\u1_L9_reg[24]/NET0131  & ~n36131 ;
  assign n36133 = \u1_L9_reg[24]/NET0131  & n36131 ;
  assign n36134 = ~n36132 & ~n36133 ;
  assign n36135 = n35910 & n35925 ;
  assign n36136 = n36115 & ~n36135 ;
  assign n36137 = ~n35906 & ~n36052 ;
  assign n36138 = ~n36062 & n36137 ;
  assign n36139 = ~n36136 & ~n36138 ;
  assign n36140 = n35898 & ~n36139 ;
  assign n36142 = n35872 & n36103 ;
  assign n36143 = ~n35906 & ~n36057 ;
  assign n36144 = ~n36142 & n36143 ;
  assign n36146 = ~n35936 & n36052 ;
  assign n36145 = ~n35878 & n35933 ;
  assign n36147 = n35906 & ~n36145 ;
  assign n36148 = ~n36146 & n36147 ;
  assign n36149 = ~n36144 & ~n36148 ;
  assign n36141 = n35912 & n36047 ;
  assign n36150 = ~n35898 & ~n36141 ;
  assign n36151 = ~n36106 & n36150 ;
  assign n36152 = ~n36149 & n36151 ;
  assign n36153 = ~n36140 & ~n36152 ;
  assign n36155 = n35922 & n36048 ;
  assign n36154 = n35899 & ~n36035 ;
  assign n36156 = n35936 & n36101 ;
  assign n36157 = ~n36154 & ~n36156 ;
  assign n36158 = ~n36155 & n36157 ;
  assign n36159 = ~n36153 & n36158 ;
  assign n36160 = \u1_L9_reg[30]/NET0131  & ~n36159 ;
  assign n36161 = ~\u1_L9_reg[30]/NET0131  & n36159 ;
  assign n36162 = ~n36160 & ~n36161 ;
  assign n36212 = decrypt_pad & ~\u1_uk_K_r8_reg[44]/NET0131  ;
  assign n36213 = ~decrypt_pad & ~\u1_uk_K_r8_reg[9]/NET0131  ;
  assign n36214 = ~n36212 & ~n36213 ;
  assign n36215 = \u1_R8_reg[28]/NET0131  & ~n36214 ;
  assign n36216 = ~\u1_R8_reg[28]/NET0131  & n36214 ;
  assign n36217 = ~n36215 & ~n36216 ;
  assign n36163 = decrypt_pad & ~\u1_uk_K_r8_reg[2]/NET0131  ;
  assign n36164 = ~decrypt_pad & ~\u1_uk_K_r8_reg[22]/NET0131  ;
  assign n36165 = ~n36163 & ~n36164 ;
  assign n36166 = \u1_R8_reg[27]/NET0131  & ~n36165 ;
  assign n36167 = ~\u1_R8_reg[27]/NET0131  & n36165 ;
  assign n36168 = ~n36166 & ~n36167 ;
  assign n36182 = decrypt_pad & ~\u1_uk_K_r8_reg[28]/NET0131  ;
  assign n36183 = ~decrypt_pad & ~\u1_uk_K_r8_reg[52]/NET0131  ;
  assign n36184 = ~n36182 & ~n36183 ;
  assign n36185 = \u1_R8_reg[24]/NET0131  & ~n36184 ;
  assign n36186 = ~\u1_R8_reg[24]/NET0131  & n36184 ;
  assign n36187 = ~n36185 & ~n36186 ;
  assign n36205 = n36168 & n36187 ;
  assign n36169 = decrypt_pad & ~\u1_uk_K_r8_reg[52]/NET0131  ;
  assign n36170 = ~decrypt_pad & ~\u1_uk_K_r8_reg[44]/NET0131  ;
  assign n36171 = ~n36169 & ~n36170 ;
  assign n36172 = \u1_R8_reg[26]/NET0131  & ~n36171 ;
  assign n36173 = ~\u1_R8_reg[26]/NET0131  & n36171 ;
  assign n36174 = ~n36172 & ~n36173 ;
  assign n36175 = decrypt_pad & ~\u1_uk_K_r8_reg[8]/NET0131  ;
  assign n36176 = ~decrypt_pad & ~\u1_uk_K_r8_reg[28]/NET0131  ;
  assign n36177 = ~n36175 & ~n36176 ;
  assign n36178 = \u1_R8_reg[25]/NET0131  & ~n36177 ;
  assign n36179 = ~\u1_R8_reg[25]/NET0131  & n36177 ;
  assign n36180 = ~n36178 & ~n36179 ;
  assign n36181 = n36174 & ~n36180 ;
  assign n36188 = decrypt_pad & ~\u1_uk_K_r8_reg[36]/NET0131  ;
  assign n36189 = ~decrypt_pad & ~\u1_uk_K_r8_reg[1]/NET0131  ;
  assign n36190 = ~n36188 & ~n36189 ;
  assign n36191 = \u1_R8_reg[29]/NET0131  & ~n36190 ;
  assign n36192 = ~\u1_R8_reg[29]/NET0131  & n36190 ;
  assign n36193 = ~n36191 & ~n36192 ;
  assign n36236 = n36180 & n36193 ;
  assign n36237 = ~n36174 & n36236 ;
  assign n36238 = ~n36181 & ~n36237 ;
  assign n36239 = n36205 & ~n36238 ;
  assign n36206 = ~n36174 & ~n36180 ;
  assign n36231 = n36187 & n36193 ;
  assign n36232 = n36206 & n36231 ;
  assign n36220 = ~n36187 & n36193 ;
  assign n36233 = n36180 & n36220 ;
  assign n36234 = ~n36232 & ~n36233 ;
  assign n36235 = ~n36168 & ~n36234 ;
  assign n36221 = n36181 & n36220 ;
  assign n36224 = ~n36187 & ~n36193 ;
  assign n36230 = n36206 & n36224 ;
  assign n36240 = ~n36221 & ~n36230 ;
  assign n36241 = ~n36235 & n36240 ;
  assign n36242 = ~n36239 & n36241 ;
  assign n36243 = n36217 & ~n36242 ;
  assign n36196 = n36174 & ~n36187 ;
  assign n36197 = ~n36174 & n36187 ;
  assign n36198 = ~n36196 & ~n36197 ;
  assign n36199 = n36193 & n36198 ;
  assign n36194 = n36187 & ~n36193 ;
  assign n36195 = ~n36181 & n36194 ;
  assign n36200 = ~n36180 & ~n36193 ;
  assign n36201 = n36196 & n36200 ;
  assign n36202 = ~n36195 & ~n36201 ;
  assign n36203 = ~n36199 & n36202 ;
  assign n36204 = ~n36168 & ~n36203 ;
  assign n36207 = n36205 & n36206 ;
  assign n36208 = n36180 & n36198 ;
  assign n36209 = n36193 & n36208 ;
  assign n36210 = ~n36207 & ~n36209 ;
  assign n36211 = ~n36204 & n36210 ;
  assign n36218 = ~n36211 & ~n36217 ;
  assign n36219 = ~n36168 & ~n36208 ;
  assign n36222 = n36168 & ~n36221 ;
  assign n36223 = ~n36196 & n36200 ;
  assign n36225 = n36174 & n36180 ;
  assign n36226 = n36224 & n36225 ;
  assign n36227 = ~n36223 & ~n36226 ;
  assign n36228 = n36222 & n36227 ;
  assign n36229 = ~n36219 & ~n36228 ;
  assign n36244 = ~n36218 & ~n36229 ;
  assign n36245 = ~n36243 & n36244 ;
  assign n36246 = ~\u1_L8_reg[22]/NET0131  & ~n36245 ;
  assign n36247 = \u1_L8_reg[22]/NET0131  & n36245 ;
  assign n36248 = ~n36246 & ~n36247 ;
  assign n36249 = decrypt_pad & ~\u1_uk_K_r8_reg[37]/P0001  ;
  assign n36250 = ~decrypt_pad & ~\u1_uk_K_r8_reg[2]/NET0131  ;
  assign n36251 = ~n36249 & ~n36250 ;
  assign n36252 = \u1_R8_reg[24]/NET0131  & ~n36251 ;
  assign n36253 = ~\u1_R8_reg[24]/NET0131  & n36251 ;
  assign n36254 = ~n36252 & ~n36253 ;
  assign n36255 = decrypt_pad & ~\u1_uk_K_r8_reg[35]/NET0131  ;
  assign n36256 = ~decrypt_pad & ~\u1_uk_K_r8_reg[0]/NET0131  ;
  assign n36257 = ~n36255 & ~n36256 ;
  assign n36258 = \u1_R8_reg[23]/NET0131  & ~n36257 ;
  assign n36259 = ~\u1_R8_reg[23]/NET0131  & n36257 ;
  assign n36260 = ~n36258 & ~n36259 ;
  assign n36280 = decrypt_pad & ~\u1_uk_K_r8_reg[0]/NET0131  ;
  assign n36281 = ~decrypt_pad & ~\u1_uk_K_r8_reg[51]/NET0131  ;
  assign n36282 = ~n36280 & ~n36281 ;
  assign n36283 = \u1_R8_reg[21]/NET0131  & ~n36282 ;
  assign n36284 = ~\u1_R8_reg[21]/NET0131  & n36282 ;
  assign n36285 = ~n36283 & ~n36284 ;
  assign n36267 = decrypt_pad & ~\u1_uk_K_r8_reg[16]/NET0131  ;
  assign n36268 = ~decrypt_pad & ~\u1_uk_K_r8_reg[36]/NET0131  ;
  assign n36269 = ~n36267 & ~n36268 ;
  assign n36270 = \u1_R8_reg[20]/NET0131  & ~n36269 ;
  assign n36271 = ~\u1_R8_reg[20]/NET0131  & n36269 ;
  assign n36272 = ~n36270 & ~n36271 ;
  assign n36274 = decrypt_pad & ~\u1_uk_K_r8_reg[22]/NET0131  ;
  assign n36275 = ~decrypt_pad & ~\u1_uk_K_r8_reg[42]/NET0131  ;
  assign n36276 = ~n36274 & ~n36275 ;
  assign n36277 = \u1_R8_reg[22]/NET0131  & ~n36276 ;
  assign n36278 = ~\u1_R8_reg[22]/NET0131  & n36276 ;
  assign n36279 = ~n36277 & ~n36278 ;
  assign n36288 = ~n36272 & n36279 ;
  assign n36289 = n36285 & n36288 ;
  assign n36298 = ~n36260 & ~n36289 ;
  assign n36307 = ~n36279 & n36285 ;
  assign n36327 = n36272 & n36307 ;
  assign n36328 = n36298 & ~n36327 ;
  assign n36261 = decrypt_pad & ~\u1_uk_K_r8_reg[1]/NET0131  ;
  assign n36262 = ~decrypt_pad & ~\u1_uk_K_r8_reg[21]/NET0131  ;
  assign n36263 = ~n36261 & ~n36262 ;
  assign n36264 = \u1_R8_reg[25]/NET0131  & ~n36263 ;
  assign n36265 = ~\u1_R8_reg[25]/NET0131  & n36263 ;
  assign n36266 = ~n36264 & ~n36265 ;
  assign n36317 = ~n36272 & ~n36285 ;
  assign n36318 = n36266 & n36317 ;
  assign n36319 = n36260 & ~n36318 ;
  assign n36322 = n36272 & ~n36285 ;
  assign n36323 = n36279 & n36322 ;
  assign n36329 = ~n36272 & ~n36279 ;
  assign n36330 = ~n36323 & ~n36329 ;
  assign n36331 = n36319 & n36330 ;
  assign n36332 = ~n36328 & ~n36331 ;
  assign n36324 = n36266 & n36323 ;
  assign n36273 = ~n36266 & n36272 ;
  assign n36295 = ~n36260 & ~n36279 ;
  assign n36325 = ~n36295 & ~n36307 ;
  assign n36326 = n36273 & ~n36325 ;
  assign n36333 = ~n36324 & ~n36326 ;
  assign n36334 = ~n36332 & n36333 ;
  assign n36335 = ~n36254 & ~n36334 ;
  assign n36290 = n36266 & n36272 ;
  assign n36291 = n36285 & n36290 ;
  assign n36286 = ~n36279 & ~n36285 ;
  assign n36287 = n36273 & n36286 ;
  assign n36292 = ~n36287 & ~n36289 ;
  assign n36293 = ~n36291 & n36292 ;
  assign n36294 = n36260 & ~n36293 ;
  assign n36296 = n36290 & n36295 ;
  assign n36297 = ~n36285 & n36296 ;
  assign n36299 = n36266 & n36285 ;
  assign n36300 = ~n36279 & ~n36299 ;
  assign n36301 = ~n36290 & ~n36300 ;
  assign n36302 = n36298 & n36301 ;
  assign n36303 = ~n36297 & ~n36302 ;
  assign n36304 = ~n36294 & n36303 ;
  assign n36305 = n36254 & ~n36304 ;
  assign n36315 = n36273 & n36285 ;
  assign n36316 = ~n36260 & ~n36315 ;
  assign n36320 = ~n36279 & ~n36316 ;
  assign n36321 = ~n36319 & n36320 ;
  assign n36306 = n36279 & n36290 ;
  assign n36308 = ~n36266 & n36307 ;
  assign n36309 = ~n36272 & n36308 ;
  assign n36310 = ~n36306 & ~n36309 ;
  assign n36311 = n36260 & ~n36310 ;
  assign n36312 = ~n36266 & ~n36272 ;
  assign n36313 = ~n36285 & n36312 ;
  assign n36314 = n36295 & n36313 ;
  assign n36336 = ~n36311 & ~n36314 ;
  assign n36337 = ~n36321 & n36336 ;
  assign n36338 = ~n36305 & n36337 ;
  assign n36339 = ~n36335 & n36338 ;
  assign n36340 = \u1_L8_reg[11]/NET0131  & ~n36339 ;
  assign n36341 = ~\u1_L8_reg[11]/NET0131  & n36339 ;
  assign n36342 = ~n36340 & ~n36341 ;
  assign n36343 = decrypt_pad & ~\u1_uk_K_r8_reg[13]/P0001  ;
  assign n36344 = ~decrypt_pad & ~\u1_uk_K_r8_reg[3]/NET0131  ;
  assign n36345 = ~n36343 & ~n36344 ;
  assign n36346 = \u1_R8_reg[16]/NET0131  & ~n36345 ;
  assign n36347 = ~\u1_R8_reg[16]/NET0131  & n36345 ;
  assign n36348 = ~n36346 & ~n36347 ;
  assign n36384 = decrypt_pad & ~\u1_uk_K_r8_reg[5]/NET0131  ;
  assign n36385 = ~decrypt_pad & ~\u1_uk_K_r8_reg[27]/NET0131  ;
  assign n36386 = ~n36384 & ~n36385 ;
  assign n36387 = \u1_R8_reg[15]/NET0131  & ~n36386 ;
  assign n36388 = ~\u1_R8_reg[15]/NET0131  & n36386 ;
  assign n36389 = ~n36387 & ~n36388 ;
  assign n36349 = decrypt_pad & ~\u1_uk_K_r8_reg[18]/NET0131  ;
  assign n36350 = ~decrypt_pad & ~\u1_uk_K_r8_reg[40]/NET0131  ;
  assign n36351 = ~n36349 & ~n36350 ;
  assign n36352 = \u1_R8_reg[17]/NET0131  & ~n36351 ;
  assign n36353 = ~\u1_R8_reg[17]/NET0131  & n36351 ;
  assign n36354 = ~n36352 & ~n36353 ;
  assign n36369 = decrypt_pad & ~\u1_uk_K_r8_reg[53]/NET0131  ;
  assign n36370 = ~decrypt_pad & ~\u1_uk_K_r8_reg[18]/NET0131  ;
  assign n36371 = ~n36369 & ~n36370 ;
  assign n36372 = \u1_R8_reg[13]/NET0131  & ~n36371 ;
  assign n36373 = ~\u1_R8_reg[13]/NET0131  & n36371 ;
  assign n36374 = ~n36372 & ~n36373 ;
  assign n36414 = n36354 & ~n36374 ;
  assign n36362 = decrypt_pad & ~\u1_uk_K_r8_reg[54]/NET0131  ;
  assign n36363 = ~decrypt_pad & ~\u1_uk_K_r8_reg[19]/NET0131  ;
  assign n36364 = ~n36362 & ~n36363 ;
  assign n36365 = \u1_R8_reg[14]/NET0131  & ~n36364 ;
  assign n36366 = ~\u1_R8_reg[14]/NET0131  & n36364 ;
  assign n36367 = ~n36365 & ~n36366 ;
  assign n36355 = decrypt_pad & ~\u1_uk_K_r8_reg[34]/NET0131  ;
  assign n36356 = ~decrypt_pad & ~\u1_uk_K_r8_reg[24]/NET0131  ;
  assign n36357 = ~n36355 & ~n36356 ;
  assign n36358 = \u1_R8_reg[12]/NET0131  & ~n36357 ;
  assign n36359 = ~\u1_R8_reg[12]/NET0131  & n36357 ;
  assign n36360 = ~n36358 & ~n36359 ;
  assign n36395 = ~n36354 & n36360 ;
  assign n36415 = n36367 & n36395 ;
  assign n36416 = ~n36414 & ~n36415 ;
  assign n36417 = ~n36389 & ~n36416 ;
  assign n36361 = n36354 & n36360 ;
  assign n36396 = n36374 & n36389 ;
  assign n36424 = n36361 & n36396 ;
  assign n36380 = ~n36360 & n36374 ;
  assign n36412 = ~n36354 & n36367 ;
  assign n36413 = n36380 & n36412 ;
  assign n36418 = n36367 & n36389 ;
  assign n36419 = n36380 & n36418 ;
  assign n36425 = ~n36413 & ~n36419 ;
  assign n36426 = ~n36424 & n36425 ;
  assign n36381 = n36360 & ~n36374 ;
  assign n36420 = ~n36367 & n36381 ;
  assign n36421 = n36354 & n36420 ;
  assign n36390 = ~n36354 & ~n36374 ;
  assign n36391 = ~n36360 & n36390 ;
  assign n36422 = n36367 & ~n36389 ;
  assign n36423 = n36391 & ~n36422 ;
  assign n36427 = ~n36421 & ~n36423 ;
  assign n36428 = n36426 & n36427 ;
  assign n36429 = ~n36417 & n36428 ;
  assign n36430 = ~n36348 & ~n36429 ;
  assign n36392 = n36367 & ~n36391 ;
  assign n36382 = ~n36380 & ~n36381 ;
  assign n36383 = ~n36367 & n36382 ;
  assign n36393 = ~n36383 & ~n36389 ;
  assign n36394 = ~n36392 & n36393 ;
  assign n36368 = n36361 & n36367 ;
  assign n36375 = n36368 & n36374 ;
  assign n36376 = n36354 & n36374 ;
  assign n36377 = ~n36360 & ~n36367 ;
  assign n36378 = n36376 & n36377 ;
  assign n36379 = ~n36375 & ~n36378 ;
  assign n36397 = n36395 & n36396 ;
  assign n36398 = n36354 & ~n36360 ;
  assign n36399 = n36389 & n36398 ;
  assign n36400 = ~n36374 & n36399 ;
  assign n36401 = ~n36397 & ~n36400 ;
  assign n36402 = n36379 & n36401 ;
  assign n36403 = ~n36394 & n36402 ;
  assign n36404 = n36348 & ~n36403 ;
  assign n36406 = n36377 & n36390 ;
  assign n36407 = n36367 & ~n36374 ;
  assign n36408 = n36395 & n36407 ;
  assign n36409 = ~n36406 & ~n36408 ;
  assign n36410 = n36389 & ~n36409 ;
  assign n36405 = n36378 & ~n36389 ;
  assign n36411 = ~n36367 & n36397 ;
  assign n36431 = ~n36405 & ~n36411 ;
  assign n36432 = ~n36410 & n36431 ;
  assign n36433 = ~n36404 & n36432 ;
  assign n36434 = ~n36430 & n36433 ;
  assign n36435 = ~\u1_L8_reg[20]/NET0131  & ~n36434 ;
  assign n36436 = \u1_L8_reg[20]/NET0131  & n36434 ;
  assign n36437 = ~n36435 & ~n36436 ;
  assign n36444 = decrypt_pad & ~\u1_uk_K_r8_reg[31]/NET0131  ;
  assign n36445 = ~decrypt_pad & ~\u1_uk_K_r8_reg[23]/NET0131  ;
  assign n36446 = ~n36444 & ~n36445 ;
  assign n36447 = \u1_R8_reg[31]/P0001  & ~n36446 ;
  assign n36448 = ~\u1_R8_reg[31]/P0001  & n36446 ;
  assign n36449 = ~n36447 & ~n36448 ;
  assign n36450 = decrypt_pad & ~\u1_uk_K_r8_reg[42]/NET0131  ;
  assign n36451 = ~decrypt_pad & ~\u1_uk_K_r8_reg[7]/NET0131  ;
  assign n36452 = ~n36450 & ~n36451 ;
  assign n36453 = \u1_R8_reg[28]/NET0131  & ~n36452 ;
  assign n36454 = ~\u1_R8_reg[28]/NET0131  & n36452 ;
  assign n36455 = ~n36453 & ~n36454 ;
  assign n36471 = decrypt_pad & ~\u1_uk_K_r8_reg[15]/NET0131  ;
  assign n36472 = ~decrypt_pad & ~\u1_uk_K_r8_reg[35]/NET0131  ;
  assign n36473 = ~n36471 & ~n36472 ;
  assign n36474 = \u1_R8_reg[30]/NET0131  & ~n36473 ;
  assign n36475 = ~\u1_R8_reg[30]/NET0131  & n36473 ;
  assign n36476 = ~n36474 & ~n36475 ;
  assign n36487 = n36455 & ~n36476 ;
  assign n36456 = decrypt_pad & ~\u1_uk_K_r8_reg[30]/NET0131  ;
  assign n36457 = ~decrypt_pad & ~\u1_uk_K_r8_reg[50]/NET0131  ;
  assign n36458 = ~n36456 & ~n36457 ;
  assign n36459 = \u1_R8_reg[1]/NET0131  & ~n36458 ;
  assign n36460 = ~\u1_R8_reg[1]/NET0131  & n36458 ;
  assign n36461 = ~n36459 & ~n36460 ;
  assign n36463 = decrypt_pad & ~\u1_uk_K_r8_reg[14]/NET0131  ;
  assign n36464 = ~decrypt_pad & ~\u1_uk_K_r8_reg[38]/NET0131  ;
  assign n36465 = ~n36463 & ~n36464 ;
  assign n36466 = \u1_R8_reg[29]/NET0131  & ~n36465 ;
  assign n36467 = ~\u1_R8_reg[29]/NET0131  & n36465 ;
  assign n36468 = ~n36466 & ~n36467 ;
  assign n36488 = ~n36461 & n36468 ;
  assign n36513 = ~n36487 & ~n36488 ;
  assign n36438 = decrypt_pad & ~\u1_uk_K_r8_reg[9]/NET0131  ;
  assign n36439 = ~decrypt_pad & ~\u1_uk_K_r8_reg[29]/NET0131  ;
  assign n36440 = ~n36438 & ~n36439 ;
  assign n36441 = \u1_R8_reg[32]/NET0131  & ~n36440 ;
  assign n36442 = ~\u1_R8_reg[32]/NET0131  & n36440 ;
  assign n36443 = ~n36441 & ~n36442 ;
  assign n36489 = n36487 & n36488 ;
  assign n36514 = n36443 & ~n36489 ;
  assign n36515 = ~n36513 & n36514 ;
  assign n36481 = ~n36455 & ~n36461 ;
  assign n36491 = n36468 & n36476 ;
  assign n36507 = n36481 & n36491 ;
  assign n36501 = ~n36468 & ~n36476 ;
  assign n36508 = n36461 & n36501 ;
  assign n36509 = n36455 & n36508 ;
  assign n36510 = ~n36507 & ~n36509 ;
  assign n36462 = ~n36455 & n36461 ;
  assign n36469 = n36462 & ~n36468 ;
  assign n36511 = n36469 & n36476 ;
  assign n36502 = ~n36455 & n36501 ;
  assign n36512 = ~n36461 & n36502 ;
  assign n36516 = ~n36511 & ~n36512 ;
  assign n36517 = n36510 & n36516 ;
  assign n36518 = ~n36515 & n36517 ;
  assign n36519 = n36449 & ~n36518 ;
  assign n36470 = n36455 & ~n36468 ;
  assign n36477 = n36470 & n36476 ;
  assign n36478 = ~n36461 & n36477 ;
  assign n36479 = n36449 & ~n36469 ;
  assign n36480 = ~n36478 & n36479 ;
  assign n36482 = n36476 & n36481 ;
  assign n36483 = n36461 & n36468 ;
  assign n36484 = ~n36449 & ~n36483 ;
  assign n36485 = ~n36482 & n36484 ;
  assign n36486 = ~n36480 & ~n36485 ;
  assign n36492 = n36455 & n36461 ;
  assign n36493 = n36491 & n36492 ;
  assign n36490 = ~n36449 & n36487 ;
  assign n36494 = ~n36489 & ~n36490 ;
  assign n36495 = ~n36493 & n36494 ;
  assign n36496 = ~n36486 & n36495 ;
  assign n36497 = ~n36443 & ~n36496 ;
  assign n36498 = ~n36449 & n36489 ;
  assign n36499 = n36462 & n36491 ;
  assign n36503 = ~n36477 & ~n36499 ;
  assign n36504 = ~n36502 & n36503 ;
  assign n36500 = n36449 & ~n36499 ;
  assign n36505 = n36443 & ~n36500 ;
  assign n36506 = ~n36504 & n36505 ;
  assign n36520 = ~n36498 & ~n36506 ;
  assign n36521 = ~n36497 & n36520 ;
  assign n36522 = ~n36519 & n36521 ;
  assign n36523 = \u1_L8_reg[5]/NET0131  & ~n36522 ;
  assign n36524 = ~\u1_L8_reg[5]/NET0131  & n36522 ;
  assign n36525 = ~n36523 & ~n36524 ;
  assign n36542 = ~n36391 & ~n36399 ;
  assign n36543 = ~n36418 & ~n36542 ;
  assign n36529 = ~n36390 & ~n36407 ;
  assign n36546 = n36360 & n36389 ;
  assign n36547 = ~n36529 & n36546 ;
  assign n36544 = ~n36367 & ~n36389 ;
  assign n36545 = n36361 & n36544 ;
  assign n36530 = n36360 & n36374 ;
  assign n36534 = ~n36367 & n36530 ;
  assign n36548 = ~n36413 & ~n36534 ;
  assign n36549 = ~n36545 & n36548 ;
  assign n36550 = ~n36547 & n36549 ;
  assign n36551 = ~n36543 & n36550 ;
  assign n36552 = ~n36348 & ~n36551 ;
  assign n36535 = ~n36367 & n36376 ;
  assign n36536 = ~n36395 & ~n36535 ;
  assign n36537 = ~n36389 & ~n36534 ;
  assign n36538 = ~n36536 & n36537 ;
  assign n36526 = n36367 & n36398 ;
  assign n36527 = ~n36374 & n36526 ;
  assign n36528 = ~n36375 & ~n36527 ;
  assign n36531 = n36389 & ~n36398 ;
  assign n36532 = ~n36530 & n36531 ;
  assign n36533 = n36529 & n36532 ;
  assign n36539 = n36528 & ~n36533 ;
  assign n36540 = ~n36538 & n36539 ;
  assign n36541 = n36348 & ~n36540 ;
  assign n36553 = ~n36406 & n36528 ;
  assign n36554 = ~n36389 & ~n36553 ;
  assign n36555 = ~n36411 & ~n36419 ;
  assign n36556 = ~n36554 & n36555 ;
  assign n36557 = ~n36541 & n36556 ;
  assign n36558 = ~n36552 & n36557 ;
  assign n36559 = ~\u1_L8_reg[10]/NET0131  & ~n36558 ;
  assign n36560 = \u1_L8_reg[10]/NET0131  & n36558 ;
  assign n36561 = ~n36559 & ~n36560 ;
  assign n36571 = ~n36180 & n36231 ;
  assign n36572 = n36174 & n36571 ;
  assign n36569 = ~n36206 & ~n36225 ;
  assign n36570 = n36224 & n36569 ;
  assign n36576 = n36220 & n36225 ;
  assign n36577 = ~n36217 & ~n36576 ;
  assign n36578 = ~n36570 & n36577 ;
  assign n36579 = ~n36572 & n36578 ;
  assign n36563 = ~n36193 & n36197 ;
  assign n36564 = ~n36168 & ~n36563 ;
  assign n36562 = ~n36224 & ~n36231 ;
  assign n36565 = n36174 & n36187 ;
  assign n36566 = ~n36180 & ~n36565 ;
  assign n36567 = n36562 & n36566 ;
  assign n36568 = ~n36564 & n36567 ;
  assign n36573 = ~n36200 & ~n36236 ;
  assign n36574 = ~n36565 & n36573 ;
  assign n36575 = ~n36168 & ~n36574 ;
  assign n36580 = ~n36568 & ~n36575 ;
  assign n36581 = n36579 & n36580 ;
  assign n36588 = ~n36174 & ~n36234 ;
  assign n36585 = n36180 & n36187 ;
  assign n36586 = ~n36230 & ~n36585 ;
  assign n36587 = n36168 & ~n36586 ;
  assign n36582 = n36168 & ~n36187 ;
  assign n36583 = n36181 & ~n36582 ;
  assign n36584 = n36562 & n36583 ;
  assign n36589 = n36217 & ~n36226 ;
  assign n36590 = ~n36584 & n36589 ;
  assign n36591 = ~n36587 & n36590 ;
  assign n36592 = ~n36588 & n36591 ;
  assign n36593 = ~n36581 & ~n36592 ;
  assign n36594 = \u1_L8_reg[12]/NET0131  & n36593 ;
  assign n36595 = ~\u1_L8_reg[12]/NET0131  & ~n36593 ;
  assign n36596 = ~n36594 & ~n36595 ;
  assign n36631 = decrypt_pad & ~\u1_uk_K_r8_reg[38]/NET0131  ;
  assign n36632 = ~decrypt_pad & ~\u1_uk_K_r8_reg[30]/NET0131  ;
  assign n36633 = ~n36631 & ~n36632 ;
  assign n36634 = \u1_R8_reg[19]/NET0131  & ~n36633 ;
  assign n36635 = ~\u1_R8_reg[19]/NET0131  & n36633 ;
  assign n36636 = ~n36634 & ~n36635 ;
  assign n36603 = decrypt_pad & ~\u1_uk_K_r8_reg[50]/NET0131  ;
  assign n36604 = ~decrypt_pad & ~\u1_uk_K_r8_reg[15]/NET0131  ;
  assign n36605 = ~n36603 & ~n36604 ;
  assign n36606 = \u1_R8_reg[21]/NET0131  & ~n36605 ;
  assign n36607 = ~\u1_R8_reg[21]/NET0131  & n36605 ;
  assign n36608 = ~n36606 & ~n36607 ;
  assign n36612 = decrypt_pad & ~\u1_uk_K_r8_reg[29]/NET0131  ;
  assign n36613 = ~decrypt_pad & ~\u1_uk_K_r8_reg[49]/NET0131  ;
  assign n36614 = ~n36612 & ~n36613 ;
  assign n36615 = \u1_R8_reg[17]/NET0131  & ~n36614 ;
  assign n36616 = ~\u1_R8_reg[17]/NET0131  & n36614 ;
  assign n36617 = ~n36615 & ~n36616 ;
  assign n36618 = ~n36608 & n36617 ;
  assign n36597 = decrypt_pad & ~\u1_uk_K_r8_reg[7]/NET0131  ;
  assign n36598 = ~decrypt_pad & ~\u1_uk_K_r8_reg[31]/NET0131  ;
  assign n36599 = ~n36597 & ~n36598 ;
  assign n36600 = \u1_R8_reg[16]/NET0131  & ~n36599 ;
  assign n36601 = ~\u1_R8_reg[16]/NET0131  & n36599 ;
  assign n36602 = ~n36600 & ~n36601 ;
  assign n36619 = decrypt_pad & ~\u1_uk_K_r8_reg[23]/NET0131  ;
  assign n36620 = ~decrypt_pad & ~\u1_uk_K_r8_reg[43]/NET0131  ;
  assign n36621 = ~n36619 & ~n36620 ;
  assign n36622 = \u1_R8_reg[18]/NET0131  & ~n36621 ;
  assign n36623 = ~\u1_R8_reg[18]/NET0131  & n36621 ;
  assign n36624 = ~n36622 & ~n36623 ;
  assign n36625 = n36602 & ~n36624 ;
  assign n36626 = ~n36618 & ~n36625 ;
  assign n36638 = n36608 & n36617 ;
  assign n36639 = ~n36608 & ~n36617 ;
  assign n36640 = ~n36638 & ~n36639 ;
  assign n36641 = ~n36624 & n36640 ;
  assign n36642 = ~n36626 & ~n36641 ;
  assign n36643 = ~n36602 & ~n36617 ;
  assign n36644 = n36608 & n36643 ;
  assign n36645 = ~n36642 & ~n36644 ;
  assign n36646 = ~n36636 & ~n36645 ;
  assign n36609 = n36602 & ~n36608 ;
  assign n36610 = ~n36602 & n36608 ;
  assign n36611 = ~n36609 & ~n36610 ;
  assign n36627 = n36611 & n36626 ;
  assign n36628 = n36617 & ~n36624 ;
  assign n36629 = ~n36602 & n36628 ;
  assign n36630 = ~n36627 & ~n36629 ;
  assign n36637 = ~n36630 & n36636 ;
  assign n36647 = ~n36602 & ~n36608 ;
  assign n36648 = n36608 & n36624 ;
  assign n36649 = ~n36647 & ~n36648 ;
  assign n36650 = n36602 & ~n36617 ;
  assign n36651 = ~n36628 & ~n36650 ;
  assign n36652 = ~n36649 & ~n36651 ;
  assign n36653 = ~n36637 & ~n36652 ;
  assign n36654 = ~n36646 & n36653 ;
  assign n36655 = decrypt_pad & ~\u1_uk_K_r8_reg[49]/NET0131  ;
  assign n36656 = ~decrypt_pad & ~\u1_uk_K_r8_reg[14]/NET0131  ;
  assign n36657 = ~n36655 & ~n36656 ;
  assign n36658 = \u1_R8_reg[20]/NET0131  & ~n36657 ;
  assign n36659 = ~\u1_R8_reg[20]/NET0131  & n36657 ;
  assign n36660 = ~n36658 & ~n36659 ;
  assign n36661 = ~n36654 & ~n36660 ;
  assign n36666 = n36624 & ~n36636 ;
  assign n36667 = n36602 & n36638 ;
  assign n36668 = n36666 & n36667 ;
  assign n36663 = ~n36602 & ~n36624 ;
  assign n36664 = ~n36636 & n36663 ;
  assign n36665 = ~n36640 & n36664 ;
  assign n36669 = ~n36617 & n36624 ;
  assign n36670 = n36609 & n36669 ;
  assign n36675 = ~n36665 & ~n36670 ;
  assign n36676 = ~n36668 & n36675 ;
  assign n36662 = n36602 & n36641 ;
  assign n36671 = n36611 & n36624 ;
  assign n36672 = n36636 & ~n36639 ;
  assign n36673 = ~n36629 & n36672 ;
  assign n36674 = ~n36671 & n36673 ;
  assign n36677 = ~n36662 & ~n36674 ;
  assign n36678 = n36676 & n36677 ;
  assign n36679 = n36660 & ~n36678 ;
  assign n36680 = n36609 & n36628 ;
  assign n36681 = n36624 & n36647 ;
  assign n36682 = ~n36617 & n36681 ;
  assign n36683 = ~n36680 & ~n36682 ;
  assign n36684 = n36636 & ~n36683 ;
  assign n36685 = n36643 & n36648 ;
  assign n36686 = n36617 & n36681 ;
  assign n36687 = ~n36685 & ~n36686 ;
  assign n36688 = ~n36636 & ~n36687 ;
  assign n36689 = ~n36684 & ~n36688 ;
  assign n36690 = ~n36679 & n36689 ;
  assign n36691 = ~n36661 & n36690 ;
  assign n36692 = ~\u1_L8_reg[14]/NET0131  & ~n36691 ;
  assign n36693 = \u1_L8_reg[14]/NET0131  & n36691 ;
  assign n36694 = ~n36692 & ~n36693 ;
  assign n36695 = n36455 & n36468 ;
  assign n36696 = ~n36476 & n36488 ;
  assign n36697 = ~n36695 & ~n36696 ;
  assign n36698 = ~n36469 & n36697 ;
  assign n36699 = n36449 & ~n36698 ;
  assign n36700 = n36455 & ~n36461 ;
  assign n36701 = ~n36476 & n36700 ;
  assign n36702 = ~n36468 & n36701 ;
  assign n36703 = ~n36699 & ~n36702 ;
  assign n36704 = ~n36443 & ~n36703 ;
  assign n36705 = n36461 & n36502 ;
  assign n36706 = n36500 & ~n36705 ;
  assign n36711 = ~n36449 & ~n36507 ;
  assign n36707 = n36468 & ~n36476 ;
  assign n36708 = n36462 & n36707 ;
  assign n36709 = n36443 & ~n36476 ;
  assign n36710 = n36470 & ~n36709 ;
  assign n36712 = ~n36708 & ~n36710 ;
  assign n36713 = n36711 & n36712 ;
  assign n36714 = ~n36512 & n36713 ;
  assign n36715 = ~n36706 & ~n36714 ;
  assign n36719 = ~n36449 & n36476 ;
  assign n36720 = ~n36481 & ~n36719 ;
  assign n36718 = ~n36449 & ~n36461 ;
  assign n36721 = ~n36468 & ~n36718 ;
  assign n36722 = ~n36720 & n36721 ;
  assign n36717 = n36461 & n36477 ;
  assign n36716 = n36455 & n36707 ;
  assign n36723 = ~n36507 & ~n36716 ;
  assign n36724 = ~n36717 & n36723 ;
  assign n36725 = ~n36722 & n36724 ;
  assign n36726 = n36443 & ~n36725 ;
  assign n36727 = ~n36715 & ~n36726 ;
  assign n36728 = ~n36704 & n36727 ;
  assign n36729 = \u1_L8_reg[15]/P0001  & n36728 ;
  assign n36730 = ~\u1_L8_reg[15]/P0001  & ~n36728 ;
  assign n36731 = ~n36729 & ~n36730 ;
  assign n36732 = n36382 & n36412 ;
  assign n36733 = ~n36389 & ~n36732 ;
  assign n36734 = ~n36414 & ~n36420 ;
  assign n36735 = n36348 & ~n36734 ;
  assign n36736 = n36389 & ~n36413 ;
  assign n36737 = n36528 & n36736 ;
  assign n36738 = ~n36735 & n36737 ;
  assign n36739 = ~n36733 & ~n36738 ;
  assign n36744 = ~n36354 & n36377 ;
  assign n36745 = ~n36408 & ~n36744 ;
  assign n36746 = n36389 & ~n36745 ;
  assign n36741 = n36360 & ~n36376 ;
  assign n36740 = ~n36374 & n36389 ;
  assign n36742 = ~n36412 & ~n36740 ;
  assign n36743 = n36741 & n36742 ;
  assign n36747 = ~n36348 & ~n36743 ;
  assign n36748 = n36379 & n36747 ;
  assign n36749 = ~n36746 & n36748 ;
  assign n36750 = n36367 & ~n36398 ;
  assign n36751 = ~n36395 & ~n36750 ;
  assign n36752 = ~n36389 & n36751 ;
  assign n36753 = ~n36415 & ~n36752 ;
  assign n36754 = n36374 & ~n36753 ;
  assign n36755 = ~n36360 & n36407 ;
  assign n36756 = n36348 & ~n36755 ;
  assign n36757 = ~n36754 & n36756 ;
  assign n36758 = ~n36749 & ~n36757 ;
  assign n36759 = ~n36739 & ~n36758 ;
  assign n36760 = ~\u1_L8_reg[1]/NET0131  & ~n36759 ;
  assign n36761 = \u1_L8_reg[1]/NET0131  & n36759 ;
  assign n36762 = ~n36760 & ~n36761 ;
  assign n36769 = decrypt_pad & ~\u1_uk_K_r8_reg[39]/NET0131  ;
  assign n36770 = ~decrypt_pad & ~\u1_uk_K_r8_reg[4]/NET0131  ;
  assign n36771 = ~n36769 & ~n36770 ;
  assign n36772 = \u1_R8_reg[5]/NET0131  & ~n36771 ;
  assign n36773 = ~\u1_R8_reg[5]/NET0131  & n36771 ;
  assign n36774 = ~n36772 & ~n36773 ;
  assign n36791 = decrypt_pad & ~\u1_uk_K_r8_reg[24]/NET0131  ;
  assign n36792 = ~decrypt_pad & ~\u1_uk_K_r8_reg[46]/NET0131  ;
  assign n36793 = ~n36791 & ~n36792 ;
  assign n36794 = \u1_R8_reg[2]/NET0131  & ~n36793 ;
  assign n36795 = ~\u1_R8_reg[2]/NET0131  & n36793 ;
  assign n36796 = ~n36794 & ~n36795 ;
  assign n36797 = n36774 & n36796 ;
  assign n36798 = ~n36774 & ~n36796 ;
  assign n36799 = ~n36797 & ~n36798 ;
  assign n36763 = decrypt_pad & ~\u1_uk_K_r8_reg[41]/NET0131  ;
  assign n36764 = ~decrypt_pad & ~\u1_uk_K_r8_reg[6]/NET0131  ;
  assign n36765 = ~n36763 & ~n36764 ;
  assign n36766 = \u1_R8_reg[1]/NET0131  & ~n36765 ;
  assign n36767 = ~\u1_R8_reg[1]/NET0131  & n36765 ;
  assign n36768 = ~n36766 & ~n36767 ;
  assign n36778 = decrypt_pad & ~\u1_uk_K_r8_reg[20]/NET0131  ;
  assign n36779 = ~decrypt_pad & ~\u1_uk_K_r8_reg[10]/NET0131  ;
  assign n36780 = ~n36778 & ~n36779 ;
  assign n36781 = \u1_R8_reg[32]/NET0131  & ~n36780 ;
  assign n36782 = ~\u1_R8_reg[32]/NET0131  & n36780 ;
  assign n36783 = ~n36781 & ~n36782 ;
  assign n36800 = n36768 & ~n36783 ;
  assign n36801 = n36799 & n36800 ;
  assign n36775 = n36768 & ~n36774 ;
  assign n36776 = ~n36768 & n36774 ;
  assign n36777 = ~n36775 & ~n36776 ;
  assign n36784 = n36777 & n36783 ;
  assign n36785 = decrypt_pad & ~\u1_uk_K_r8_reg[33]/NET0131  ;
  assign n36786 = ~decrypt_pad & ~\u1_uk_K_r8_reg[55]/NET0131  ;
  assign n36787 = ~n36785 & ~n36786 ;
  assign n36788 = \u1_R8_reg[3]/NET0131  & ~n36787 ;
  assign n36789 = ~\u1_R8_reg[3]/NET0131  & n36787 ;
  assign n36790 = ~n36788 & ~n36789 ;
  assign n36802 = ~n36784 & n36790 ;
  assign n36803 = ~n36801 & n36802 ;
  assign n36804 = n36774 & n36783 ;
  assign n36805 = ~n36774 & ~n36783 ;
  assign n36806 = ~n36804 & ~n36805 ;
  assign n36807 = ~n36768 & ~n36806 ;
  assign n36808 = ~n36783 & n36798 ;
  assign n36809 = ~n36790 & ~n36808 ;
  assign n36810 = ~n36807 & n36809 ;
  assign n36811 = ~n36803 & ~n36810 ;
  assign n36812 = ~n36777 & n36806 ;
  assign n36813 = n36796 & n36812 ;
  assign n36814 = decrypt_pad & ~\u1_uk_K_r8_reg[11]/NET0131  ;
  assign n36815 = ~decrypt_pad & ~\u1_uk_K_r8_reg[33]/NET0131  ;
  assign n36816 = ~n36814 & ~n36815 ;
  assign n36817 = \u1_R8_reg[4]/NET0131  & ~n36816 ;
  assign n36818 = ~\u1_R8_reg[4]/NET0131  & n36816 ;
  assign n36819 = ~n36817 & ~n36818 ;
  assign n36820 = ~n36813 & ~n36819 ;
  assign n36821 = ~n36811 & n36820 ;
  assign n36824 = ~n36768 & ~n36796 ;
  assign n36825 = ~n36783 & ~n36824 ;
  assign n36829 = n36804 & n36824 ;
  assign n36830 = ~n36825 & ~n36829 ;
  assign n36831 = n36790 & ~n36830 ;
  assign n36826 = n36783 & ~n36796 ;
  assign n36827 = ~n36790 & ~n36826 ;
  assign n36828 = ~n36825 & n36827 ;
  assign n36822 = n36775 & n36783 ;
  assign n36823 = ~n36796 & n36822 ;
  assign n36832 = n36768 & n36797 ;
  assign n36833 = n36819 & ~n36832 ;
  assign n36834 = ~n36823 & n36833 ;
  assign n36835 = ~n36828 & n36834 ;
  assign n36836 = ~n36831 & n36835 ;
  assign n36837 = ~n36821 & ~n36836 ;
  assign n36838 = \u1_L8_reg[17]/NET0131  & n36837 ;
  assign n36839 = ~\u1_L8_reg[17]/NET0131  & ~n36837 ;
  assign n36840 = ~n36838 & ~n36839 ;
  assign n36841 = ~n36449 & ~n36701 ;
  assign n36842 = ~n36717 & n36841 ;
  assign n36843 = n36468 & ~n36481 ;
  assign n36844 = ~n36487 & n36843 ;
  assign n36845 = n36449 & ~n36508 ;
  assign n36846 = ~n36844 & n36845 ;
  assign n36847 = ~n36842 & ~n36846 ;
  assign n36848 = ~n36461 & ~n36468 ;
  assign n36849 = ~n36700 & ~n36848 ;
  assign n36850 = ~n36470 & n36476 ;
  assign n36851 = ~n36849 & n36850 ;
  assign n36852 = n36443 & ~n36705 ;
  assign n36853 = ~n36851 & n36852 ;
  assign n36854 = ~n36847 & n36853 ;
  assign n36867 = ~n36478 & ~n36512 ;
  assign n36855 = n36461 & n36490 ;
  assign n36862 = n36449 & n36455 ;
  assign n36863 = ~n36483 & n36862 ;
  assign n36864 = ~n36501 & n36863 ;
  assign n36868 = ~n36855 & ~n36864 ;
  assign n36869 = n36867 & n36868 ;
  assign n36856 = ~n36455 & n36468 ;
  assign n36858 = ~n36449 & n36462 ;
  assign n36859 = ~n36856 & ~n36858 ;
  assign n36860 = n36476 & ~n36859 ;
  assign n36861 = n36492 & n36707 ;
  assign n36857 = n36718 & n36856 ;
  assign n36865 = ~n36443 & ~n36857 ;
  assign n36866 = ~n36861 & n36865 ;
  assign n36870 = ~n36860 & n36866 ;
  assign n36871 = n36869 & n36870 ;
  assign n36872 = ~n36854 & ~n36871 ;
  assign n36873 = n36449 & n36502 ;
  assign n36874 = ~n36449 & n36861 ;
  assign n36875 = ~n36873 & ~n36874 ;
  assign n36876 = ~n36872 & n36875 ;
  assign n36877 = ~\u1_L8_reg[21]/NET0131  & ~n36876 ;
  assign n36878 = \u1_L8_reg[21]/NET0131  & n36876 ;
  assign n36879 = ~n36877 & ~n36878 ;
  assign n36888 = n36608 & n36650 ;
  assign n36889 = ~n36636 & ~n36888 ;
  assign n36890 = ~n36629 & n36889 ;
  assign n36892 = n36636 & ~n36643 ;
  assign n36893 = ~n36667 & n36892 ;
  assign n36891 = ~n36624 & n36639 ;
  assign n36894 = ~n36681 & ~n36891 ;
  assign n36895 = n36893 & n36894 ;
  assign n36896 = ~n36890 & ~n36895 ;
  assign n36882 = n36618 & n36624 ;
  assign n36883 = n36602 & n36882 ;
  assign n36897 = n36608 & n36628 ;
  assign n36898 = n36660 & ~n36897 ;
  assign n36899 = ~n36883 & n36898 ;
  assign n36900 = ~n36896 & n36899 ;
  assign n36907 = ~n36618 & n36636 ;
  assign n36904 = ~n36636 & ~n36643 ;
  assign n36908 = ~n36624 & ~n36904 ;
  assign n36909 = ~n36907 & n36908 ;
  assign n36903 = n36602 & ~n36639 ;
  assign n36905 = ~n36663 & ~n36903 ;
  assign n36906 = n36904 & n36905 ;
  assign n36901 = ~n36602 & n36638 ;
  assign n36902 = n36624 & n36901 ;
  assign n36910 = ~n36660 & ~n36902 ;
  assign n36911 = ~n36906 & n36910 ;
  assign n36912 = ~n36909 & n36911 ;
  assign n36913 = ~n36900 & ~n36912 ;
  assign n36884 = ~n36682 & ~n36883 ;
  assign n36885 = ~n36624 & n36644 ;
  assign n36886 = n36884 & ~n36885 ;
  assign n36887 = n36636 & ~n36886 ;
  assign n36880 = n36650 & n36666 ;
  assign n36881 = n36625 & n36638 ;
  assign n36914 = ~n36880 & ~n36881 ;
  assign n36915 = ~n36887 & n36914 ;
  assign n36916 = ~n36913 & n36915 ;
  assign n36917 = ~\u1_L8_reg[25]/NET0131  & ~n36916 ;
  assign n36918 = \u1_L8_reg[25]/NET0131  & n36916 ;
  assign n36919 = ~n36917 & ~n36918 ;
  assign n36920 = ~n36415 & ~n36526 ;
  assign n36921 = ~n36744 & n36920 ;
  assign n36922 = n36374 & ~n36921 ;
  assign n36926 = ~n36391 & ~n36526 ;
  assign n36927 = n36389 & ~n36926 ;
  assign n36923 = n36377 & n36414 ;
  assign n36924 = ~n36368 & ~n36923 ;
  assign n36925 = ~n36389 & ~n36924 ;
  assign n36928 = n36348 & ~n36925 ;
  assign n36929 = ~n36927 & n36928 ;
  assign n36930 = ~n36922 & n36929 ;
  assign n36931 = n36396 & ~n36751 ;
  assign n36932 = ~n36348 & ~n36378 ;
  assign n36933 = ~n36420 & n36932 ;
  assign n36934 = ~n36931 & n36933 ;
  assign n36935 = ~n36930 & ~n36934 ;
  assign n36939 = ~n36374 & ~n36395 ;
  assign n36938 = ~n36354 & n36530 ;
  assign n36940 = ~n36367 & ~n36398 ;
  assign n36941 = ~n36938 & n36940 ;
  assign n36942 = ~n36939 & n36941 ;
  assign n36936 = ~n36390 & ~n36755 ;
  assign n36937 = ~n36348 & ~n36936 ;
  assign n36943 = ~n36389 & ~n36937 ;
  assign n36944 = ~n36942 & n36943 ;
  assign n36945 = ~n36378 & n36389 ;
  assign n36946 = ~n36421 & n36945 ;
  assign n36947 = ~n36944 & ~n36946 ;
  assign n36948 = ~n36935 & ~n36947 ;
  assign n36949 = ~\u1_L8_reg[26]/NET0131  & ~n36948 ;
  assign n36950 = \u1_L8_reg[26]/NET0131  & n36948 ;
  assign n36951 = ~n36949 & ~n36950 ;
  assign n36977 = n36273 & ~n36285 ;
  assign n36978 = ~n36291 & ~n36977 ;
  assign n36979 = ~n36286 & ~n36289 ;
  assign n36980 = ~n36266 & ~n36979 ;
  assign n36981 = n36978 & ~n36980 ;
  assign n36982 = n36260 & ~n36981 ;
  assign n36953 = n36279 & n36315 ;
  assign n36973 = ~n36273 & ~n36279 ;
  assign n36974 = ~n36317 & n36973 ;
  assign n36975 = ~n36953 & ~n36974 ;
  assign n36976 = ~n36260 & ~n36975 ;
  assign n36983 = n36279 & n36318 ;
  assign n36984 = ~n36976 & ~n36983 ;
  assign n36985 = ~n36982 & n36984 ;
  assign n36986 = ~n36254 & ~n36985 ;
  assign n36952 = ~n36272 & n36299 ;
  assign n36954 = n36285 & n36329 ;
  assign n36955 = ~n36952 & ~n36954 ;
  assign n36956 = ~n36953 & n36955 ;
  assign n36957 = n36260 & ~n36956 ;
  assign n36962 = ~n36307 & n36312 ;
  assign n36963 = ~n36306 & ~n36962 ;
  assign n36964 = ~n36260 & ~n36963 ;
  assign n36958 = n36266 & n36329 ;
  assign n36959 = n36279 & n36312 ;
  assign n36960 = ~n36958 & ~n36959 ;
  assign n36961 = ~n36285 & ~n36960 ;
  assign n36965 = n36273 & n36295 ;
  assign n36966 = ~n36324 & ~n36965 ;
  assign n36967 = ~n36961 & n36966 ;
  assign n36968 = ~n36964 & n36967 ;
  assign n36969 = ~n36957 & n36968 ;
  assign n36970 = n36254 & ~n36969 ;
  assign n36971 = n36260 & ~n36279 ;
  assign n36972 = n36299 & n36971 ;
  assign n36987 = ~n36287 & ~n36972 ;
  assign n36988 = ~n36970 & n36987 ;
  assign n36989 = ~n36986 & n36988 ;
  assign n36990 = \u1_L8_reg[29]/NET0131  & ~n36989 ;
  assign n36991 = ~\u1_L8_reg[29]/NET0131  & n36989 ;
  assign n36992 = ~n36990 & ~n36991 ;
  assign n36993 = decrypt_pad & ~\u1_uk_K_r8_reg[12]/NET0131  ;
  assign n36994 = ~decrypt_pad & ~\u1_uk_K_r8_reg[34]/NET0131  ;
  assign n36995 = ~n36993 & ~n36994 ;
  assign n36996 = \u1_R8_reg[8]/NET0131  & ~n36995 ;
  assign n36997 = ~\u1_R8_reg[8]/NET0131  & n36995 ;
  assign n36998 = ~n36996 & ~n36997 ;
  assign n36999 = decrypt_pad & ~\u1_uk_K_r8_reg[46]/NET0131  ;
  assign n37000 = ~decrypt_pad & ~\u1_uk_K_r8_reg[11]/NET0131  ;
  assign n37001 = ~n36999 & ~n37000 ;
  assign n37002 = \u1_R8_reg[7]/NET0131  & ~n37001 ;
  assign n37003 = ~\u1_R8_reg[7]/NET0131  & n37001 ;
  assign n37004 = ~n37002 & ~n37003 ;
  assign n37018 = decrypt_pad & ~\u1_uk_K_r8_reg[4]/NET0131  ;
  assign n37019 = ~decrypt_pad & ~\u1_uk_K_r8_reg[26]/NET0131  ;
  assign n37020 = ~n37018 & ~n37019 ;
  assign n37021 = \u1_R8_reg[5]/NET0131  & ~n37020 ;
  assign n37022 = ~\u1_R8_reg[5]/NET0131  & n37020 ;
  assign n37023 = ~n37021 & ~n37022 ;
  assign n37005 = decrypt_pad & ~\u1_uk_K_r8_reg[25]/NET0131  ;
  assign n37006 = ~decrypt_pad & ~\u1_uk_K_r8_reg[47]/NET0131  ;
  assign n37007 = ~n37005 & ~n37006 ;
  assign n37008 = \u1_R8_reg[4]/NET0131  & ~n37007 ;
  assign n37009 = ~\u1_R8_reg[4]/NET0131  & n37007 ;
  assign n37010 = ~n37008 & ~n37009 ;
  assign n37011 = decrypt_pad & ~\u1_uk_K_r8_reg[17]/NET0131  ;
  assign n37012 = ~decrypt_pad & ~\u1_uk_K_r8_reg[39]/NET0131  ;
  assign n37013 = ~n37011 & ~n37012 ;
  assign n37014 = \u1_R8_reg[9]/NET0131  & ~n37013 ;
  assign n37015 = ~\u1_R8_reg[9]/NET0131  & n37013 ;
  assign n37016 = ~n37014 & ~n37015 ;
  assign n37033 = ~n37010 & n37016 ;
  assign n37034 = ~n37023 & n37033 ;
  assign n37025 = decrypt_pad & ~\u1_uk_K_r8_reg[27]/NET0131  ;
  assign n37026 = ~decrypt_pad & ~\u1_uk_K_r8_reg[17]/NET0131  ;
  assign n37027 = ~n37025 & ~n37026 ;
  assign n37028 = \u1_R8_reg[6]/NET0131  & ~n37027 ;
  assign n37029 = ~\u1_R8_reg[6]/NET0131  & n37027 ;
  assign n37030 = ~n37028 & ~n37029 ;
  assign n37035 = n37010 & n37023 ;
  assign n37036 = n37010 & ~n37016 ;
  assign n37037 = ~n37035 & ~n37036 ;
  assign n37038 = n37030 & ~n37037 ;
  assign n37039 = ~n37034 & ~n37038 ;
  assign n37040 = ~n37004 & ~n37039 ;
  assign n37041 = ~n37016 & n37023 ;
  assign n37042 = ~n37034 & ~n37041 ;
  assign n37043 = ~n37030 & ~n37042 ;
  assign n37017 = n37010 & n37016 ;
  assign n37024 = n37017 & ~n37023 ;
  assign n37031 = n37024 & n37030 ;
  assign n37032 = n37004 & n37031 ;
  assign n37044 = ~n37004 & ~n37023 ;
  assign n37045 = n37016 & ~n37030 ;
  assign n37046 = n37044 & n37045 ;
  assign n37047 = n37023 & n37030 ;
  assign n37048 = n37033 & n37047 ;
  assign n37049 = ~n37046 & ~n37048 ;
  assign n37050 = ~n37032 & n37049 ;
  assign n37051 = ~n37043 & n37050 ;
  assign n37052 = ~n37040 & n37051 ;
  assign n37053 = ~n36998 & ~n37052 ;
  assign n37059 = ~n37023 & n37036 ;
  assign n37060 = ~n37030 & n37059 ;
  assign n37054 = ~n37010 & ~n37016 ;
  assign n37055 = n37044 & n37054 ;
  assign n37056 = ~n37010 & n37030 ;
  assign n37057 = n37004 & n37023 ;
  assign n37058 = ~n37056 & n37057 ;
  assign n37066 = ~n37055 & ~n37058 ;
  assign n37067 = ~n37060 & n37066 ;
  assign n37061 = n37017 & n37023 ;
  assign n37062 = ~n37030 & n37061 ;
  assign n37063 = ~n37004 & n37030 ;
  assign n37064 = ~n37033 & n37063 ;
  assign n37065 = n37037 & n37064 ;
  assign n37068 = ~n37062 & ~n37065 ;
  assign n37069 = n37067 & n37068 ;
  assign n37070 = n36998 & ~n37069 ;
  assign n37071 = ~n37023 & ~n37030 ;
  assign n37072 = ~n37047 & ~n37071 ;
  assign n37073 = n37033 & ~n37072 ;
  assign n37074 = ~n37004 & ~n37073 ;
  assign n37076 = ~n37023 & n37030 ;
  assign n37077 = ~n37016 & n37076 ;
  assign n37078 = ~n37010 & n37077 ;
  assign n37075 = ~n37030 & n37035 ;
  assign n37079 = n37004 & ~n37075 ;
  assign n37080 = ~n37078 & n37079 ;
  assign n37081 = ~n37074 & ~n37080 ;
  assign n37082 = ~n37070 & ~n37081 ;
  assign n37083 = ~n37053 & n37082 ;
  assign n37084 = \u1_L8_reg[2]/NET0131  & n37083 ;
  assign n37085 = ~\u1_L8_reg[2]/NET0131  & ~n37083 ;
  assign n37086 = ~n37084 & ~n37085 ;
  assign n37109 = n37023 & n37054 ;
  assign n37110 = n37030 & n37109 ;
  assign n37111 = ~n37059 & ~n37061 ;
  assign n37112 = ~n37110 & n37111 ;
  assign n37113 = n37004 & ~n37112 ;
  assign n37091 = n37023 & n37033 ;
  assign n37092 = ~n37030 & n37054 ;
  assign n37093 = ~n37091 & ~n37092 ;
  assign n37108 = ~n37004 & ~n37093 ;
  assign n37105 = n37004 & n37010 ;
  assign n37106 = ~n37024 & ~n37105 ;
  assign n37107 = ~n37030 & ~n37106 ;
  assign n37114 = n37033 & n37076 ;
  assign n37115 = ~n37107 & ~n37114 ;
  assign n37116 = ~n37108 & n37115 ;
  assign n37117 = ~n37113 & n37116 ;
  assign n37118 = n36998 & ~n37117 ;
  assign n37087 = n37036 & n37047 ;
  assign n37088 = ~n37023 & n37056 ;
  assign n37089 = ~n37087 & ~n37088 ;
  assign n37090 = ~n37004 & ~n37089 ;
  assign n37094 = n37004 & n37093 ;
  assign n37095 = ~n37030 & n37036 ;
  assign n37096 = ~n37004 & ~n37035 ;
  assign n37097 = ~n37034 & n37096 ;
  assign n37098 = ~n37095 & n37097 ;
  assign n37099 = ~n37094 & ~n37098 ;
  assign n37100 = ~n37033 & ~n37036 ;
  assign n37101 = n37076 & n37100 ;
  assign n37102 = ~n37087 & ~n37101 ;
  assign n37103 = ~n37099 & n37102 ;
  assign n37104 = ~n36998 & ~n37103 ;
  assign n37119 = ~n37090 & ~n37104 ;
  assign n37120 = ~n37118 & n37119 ;
  assign n37121 = ~\u1_L8_reg[28]/NET0131  & ~n37120 ;
  assign n37122 = \u1_L8_reg[28]/NET0131  & n37120 ;
  assign n37123 = ~n37121 & ~n37122 ;
  assign n37133 = ~n36315 & ~n36958 ;
  assign n37134 = ~n36324 & n37133 ;
  assign n37135 = n36260 & ~n37134 ;
  assign n37136 = ~n36254 & ~n36287 ;
  assign n37137 = ~n36296 & n37136 ;
  assign n37138 = ~n37135 & n37137 ;
  assign n37140 = n36279 & n36299 ;
  assign n37139 = n36290 & n36971 ;
  assign n37141 = n36254 & ~n37139 ;
  assign n37142 = ~n37140 & n37141 ;
  assign n37143 = ~n36309 & n37142 ;
  assign n37144 = ~n37138 & ~n37143 ;
  assign n37125 = n36285 & n36312 ;
  assign n37126 = ~n36983 & ~n37125 ;
  assign n37127 = ~n36254 & ~n37126 ;
  assign n37124 = ~n36279 & n36312 ;
  assign n37128 = ~n36308 & ~n36329 ;
  assign n37129 = n36254 & ~n37128 ;
  assign n37130 = ~n37124 & ~n37129 ;
  assign n37131 = ~n37127 & n37130 ;
  assign n37132 = ~n36260 & ~n37131 ;
  assign n37148 = ~n36260 & n36978 ;
  assign n37145 = ~n36313 & ~n36952 ;
  assign n37146 = n36260 & ~n36315 ;
  assign n37147 = n37145 & n37146 ;
  assign n37149 = n36279 & ~n37147 ;
  assign n37150 = ~n37148 & n37149 ;
  assign n37151 = ~n37132 & ~n37150 ;
  assign n37152 = ~n37144 & n37151 ;
  assign n37153 = ~\u1_L8_reg[4]/NET0131  & ~n37152 ;
  assign n37154 = \u1_L8_reg[4]/NET0131  & n37152 ;
  assign n37155 = ~n37153 & ~n37154 ;
  assign n37160 = ~n37062 & ~n37087 ;
  assign n37161 = ~n37109 & ~n37114 ;
  assign n37162 = ~n37060 & n37161 ;
  assign n37163 = n37160 & n37162 ;
  assign n37164 = ~n37004 & ~n37163 ;
  assign n37165 = n37023 & ~n37095 ;
  assign n37166 = n37004 & ~n37034 ;
  assign n37167 = ~n37059 & n37166 ;
  assign n37168 = ~n37165 & n37167 ;
  assign n37158 = n37030 & ~n37041 ;
  assign n37159 = n37105 & n37158 ;
  assign n37156 = ~n37010 & ~n37044 ;
  assign n37157 = n37045 & n37156 ;
  assign n37169 = ~n36998 & ~n37157 ;
  assign n37170 = ~n37159 & n37169 ;
  assign n37171 = ~n37168 & n37170 ;
  assign n37172 = ~n37164 & n37171 ;
  assign n37175 = ~n37016 & n37071 ;
  assign n37174 = n37016 & n37056 ;
  assign n37176 = n37004 & ~n37174 ;
  assign n37177 = ~n37175 & n37176 ;
  assign n37178 = ~n37004 & ~n37024 ;
  assign n37179 = ~n37077 & n37178 ;
  assign n37180 = ~n37177 & ~n37179 ;
  assign n37173 = n37023 & n37092 ;
  assign n37181 = n36998 & n37049 ;
  assign n37182 = ~n37173 & n37181 ;
  assign n37183 = n37160 & n37182 ;
  assign n37184 = ~n37180 & n37183 ;
  assign n37185 = ~n37172 & ~n37184 ;
  assign n37186 = ~\u1_L8_reg[13]/NET0131  & ~n37185 ;
  assign n37187 = \u1_L8_reg[13]/NET0131  & n37185 ;
  assign n37188 = ~n37186 & ~n37187 ;
  assign n37193 = ~n36260 & ~n37145 ;
  assign n37189 = n36272 & ~n36307 ;
  assign n37190 = ~n37125 & ~n37189 ;
  assign n37191 = n36260 & ~n37190 ;
  assign n37192 = n36285 & n36306 ;
  assign n37194 = ~n36254 & ~n37192 ;
  assign n37195 = ~n37191 & n37194 ;
  assign n37196 = ~n37193 & n37195 ;
  assign n37200 = n36260 & n36327 ;
  assign n37197 = n36279 & n36952 ;
  assign n37201 = n36254 & ~n36308 ;
  assign n37202 = ~n37197 & n37201 ;
  assign n37203 = ~n37200 & n37202 ;
  assign n37198 = ~n36260 & ~n36322 ;
  assign n37199 = ~n36319 & ~n37198 ;
  assign n37204 = ~n36961 & ~n37199 ;
  assign n37205 = n37203 & n37204 ;
  assign n37206 = ~n37196 & ~n37205 ;
  assign n37207 = ~n36297 & ~n36321 ;
  assign n37208 = ~n37206 & n37207 ;
  assign n37209 = ~\u1_L8_reg[19]/P0001  & ~n37208 ;
  assign n37210 = \u1_L8_reg[19]/P0001  & n37208 ;
  assign n37211 = ~n37209 & ~n37210 ;
  assign n37212 = ~n36777 & ~n36783 ;
  assign n37213 = ~n36768 & n36783 ;
  assign n37214 = n36796 & n37213 ;
  assign n37215 = ~n36774 & n37214 ;
  assign n37216 = ~n37212 & ~n37215 ;
  assign n37217 = n36819 & ~n37216 ;
  assign n37218 = n36783 & n36832 ;
  assign n37219 = ~n37217 & ~n37218 ;
  assign n37220 = ~n36790 & ~n37219 ;
  assign n37221 = n36768 & n36790 ;
  assign n37222 = n36774 & ~n36783 ;
  assign n37223 = n37221 & n37222 ;
  assign n37229 = n36819 & ~n36829 ;
  assign n37230 = ~n37223 & n37229 ;
  assign n37224 = n36790 & n36796 ;
  assign n37225 = n36822 & n37224 ;
  assign n37226 = n36796 & n36805 ;
  assign n37227 = ~n36768 & n36790 ;
  assign n37228 = n37226 & n37227 ;
  assign n37231 = ~n37225 & ~n37228 ;
  assign n37232 = n37230 & n37231 ;
  assign n37235 = n37222 & n37224 ;
  assign n37234 = n36805 & n37221 ;
  assign n37239 = ~n36819 & ~n37234 ;
  assign n37240 = ~n37235 & n37239 ;
  assign n37233 = n36777 & ~n36799 ;
  assign n37236 = ~n36768 & ~n36797 ;
  assign n37237 = n36783 & ~n36790 ;
  assign n37238 = ~n37236 & n37237 ;
  assign n37241 = ~n37233 & ~n37238 ;
  assign n37242 = n37240 & n37241 ;
  assign n37243 = ~n37232 & ~n37242 ;
  assign n37244 = ~n36790 & n36812 ;
  assign n37245 = n36790 & n37213 ;
  assign n37246 = ~n37234 & ~n37245 ;
  assign n37247 = ~n37244 & n37246 ;
  assign n37248 = ~n36796 & ~n37247 ;
  assign n37249 = ~n37243 & ~n37248 ;
  assign n37250 = ~n37220 & n37249 ;
  assign n37251 = \u1_L8_reg[23]/NET0131  & ~n37250 ;
  assign n37252 = ~\u1_L8_reg[23]/NET0131  & n37250 ;
  assign n37253 = ~n37251 & ~n37252 ;
  assign n37265 = ~n36697 & ~n36700 ;
  assign n37266 = n36449 & ~n37265 ;
  assign n37267 = ~n36492 & n36843 ;
  assign n37268 = ~n36449 & ~n36502 ;
  assign n37269 = ~n37267 & n37268 ;
  assign n37270 = ~n37266 & ~n37269 ;
  assign n37271 = ~n36499 & ~n36508 ;
  assign n37272 = ~n36478 & n37271 ;
  assign n37273 = ~n37270 & n37272 ;
  assign n37274 = n36443 & ~n37273 ;
  assign n37254 = ~n36707 & n36849 ;
  assign n37255 = n36449 & ~n36696 ;
  assign n37256 = ~n37254 & n37255 ;
  assign n37257 = ~n36511 & ~n37256 ;
  assign n37258 = ~n36443 & ~n37257 ;
  assign n37261 = ~n36449 & ~n36510 ;
  assign n37262 = n36492 & n36719 ;
  assign n37263 = ~n36857 & ~n37262 ;
  assign n37264 = ~n36443 & ~n37263 ;
  assign n37259 = n36449 & n36476 ;
  assign n37260 = n36848 & n37259 ;
  assign n37275 = ~n36498 & ~n37260 ;
  assign n37276 = ~n37264 & n37275 ;
  assign n37277 = ~n37261 & n37276 ;
  assign n37278 = ~n37258 & n37277 ;
  assign n37279 = ~n37274 & n37278 ;
  assign n37280 = ~\u1_L8_reg[27]/NET0131  & ~n37279 ;
  assign n37281 = \u1_L8_reg[27]/NET0131  & n37279 ;
  assign n37282 = ~n37280 & ~n37281 ;
  assign n37299 = n36174 & ~n36562 ;
  assign n37300 = ~n36563 & ~n37299 ;
  assign n37301 = n36180 & ~n37300 ;
  assign n37302 = ~n36563 & ~n36571 ;
  assign n37303 = n36168 & ~n37302 ;
  assign n37298 = n36564 & ~n36573 ;
  assign n37304 = ~n36221 & ~n37298 ;
  assign n37305 = ~n37303 & n37304 ;
  assign n37306 = ~n37301 & n37305 ;
  assign n37307 = ~n36217 & ~n37306 ;
  assign n37285 = ~n36174 & ~n36562 ;
  assign n37286 = ~n36180 & n37285 ;
  assign n37283 = ~n36562 & n36573 ;
  assign n37284 = ~n36206 & ~n37283 ;
  assign n37287 = ~n36168 & ~n37284 ;
  assign n37288 = ~n37286 & n37287 ;
  assign n37289 = ~n36180 & n36224 ;
  assign n37290 = ~n36237 & ~n37289 ;
  assign n37291 = n36168 & ~n37290 ;
  assign n37292 = ~n36168 & ~n36180 ;
  assign n37293 = n36174 & n36194 ;
  assign n37294 = ~n37292 & n37293 ;
  assign n37295 = ~n37291 & ~n37294 ;
  assign n37296 = ~n37288 & n37295 ;
  assign n37297 = n36217 & ~n37296 ;
  assign n37308 = ~n36194 & ~n36198 ;
  assign n37309 = ~n36168 & ~n37308 ;
  assign n37310 = ~n36222 & ~n37292 ;
  assign n37311 = ~n37309 & n37310 ;
  assign n37312 = ~n37297 & ~n37311 ;
  assign n37313 = ~n37307 & n37312 ;
  assign n37314 = \u1_L8_reg[32]/NET0131  & n37313 ;
  assign n37315 = ~\u1_L8_reg[32]/NET0131  & ~n37313 ;
  assign n37316 = ~n37314 & ~n37315 ;
  assign n37317 = decrypt_pad & ~\u1_uk_K_r8_reg[32]/NET0131  ;
  assign n37318 = ~decrypt_pad & ~\u1_uk_K_r8_reg[54]/NET0131  ;
  assign n37319 = ~n37317 & ~n37318 ;
  assign n37320 = \u1_R8_reg[11]/NET0131  & ~n37319 ;
  assign n37321 = ~\u1_R8_reg[11]/NET0131  & n37319 ;
  assign n37322 = ~n37320 & ~n37321 ;
  assign n37323 = decrypt_pad & ~\u1_uk_K_r8_reg[3]/NET0131  ;
  assign n37324 = ~decrypt_pad & ~\u1_uk_K_r8_reg[25]/NET0131  ;
  assign n37325 = ~n37323 & ~n37324 ;
  assign n37326 = \u1_R8_reg[13]/NET0131  & ~n37325 ;
  assign n37327 = ~\u1_R8_reg[13]/NET0131  & n37325 ;
  assign n37328 = ~n37326 & ~n37327 ;
  assign n37343 = decrypt_pad & ~\u1_uk_K_r8_reg[55]/NET0131  ;
  assign n37344 = ~decrypt_pad & ~\u1_uk_K_r8_reg[20]/NET0131  ;
  assign n37345 = ~n37343 & ~n37344 ;
  assign n37346 = \u1_R8_reg[9]/NET0131  & ~n37345 ;
  assign n37347 = ~\u1_R8_reg[9]/NET0131  & n37345 ;
  assign n37348 = ~n37346 & ~n37347 ;
  assign n37350 = n37328 & ~n37348 ;
  assign n37336 = decrypt_pad & ~\u1_uk_K_r8_reg[6]/NET0131  ;
  assign n37337 = ~decrypt_pad & ~\u1_uk_K_r8_reg[53]/NET0131  ;
  assign n37338 = ~n37336 & ~n37337 ;
  assign n37339 = \u1_R8_reg[10]/NET0131  & ~n37338 ;
  assign n37340 = ~\u1_R8_reg[10]/NET0131  & n37338 ;
  assign n37341 = ~n37339 & ~n37340 ;
  assign n37329 = decrypt_pad & ~\u1_uk_K_r8_reg[26]/NET0131  ;
  assign n37330 = ~decrypt_pad & ~\u1_uk_K_r8_reg[48]/NET0131  ;
  assign n37331 = ~n37329 & ~n37330 ;
  assign n37332 = \u1_R8_reg[8]/NET0131  & ~n37331 ;
  assign n37333 = ~\u1_R8_reg[8]/NET0131  & n37331 ;
  assign n37334 = ~n37332 & ~n37333 ;
  assign n37351 = n37328 & ~n37334 ;
  assign n37352 = n37341 & n37351 ;
  assign n37353 = ~n37328 & n37348 ;
  assign n37354 = n37334 & n37353 ;
  assign n37355 = ~n37352 & ~n37354 ;
  assign n37356 = ~n37350 & n37355 ;
  assign n37357 = decrypt_pad & ~\u1_uk_K_r8_reg[47]/NET0131  ;
  assign n37358 = ~decrypt_pad & ~\u1_uk_K_r8_reg[12]/NET0131  ;
  assign n37359 = ~n37357 & ~n37358 ;
  assign n37360 = \u1_R8_reg[12]/NET0131  & ~n37359 ;
  assign n37361 = ~\u1_R8_reg[12]/NET0131  & n37359 ;
  assign n37362 = ~n37360 & ~n37361 ;
  assign n37363 = ~n37356 & n37362 ;
  assign n37335 = ~n37328 & ~n37334 ;
  assign n37342 = n37335 & ~n37341 ;
  assign n37349 = n37342 & ~n37348 ;
  assign n37364 = n37341 & n37350 ;
  assign n37365 = ~n37349 & ~n37364 ;
  assign n37366 = ~n37363 & n37365 ;
  assign n37367 = n37322 & ~n37366 ;
  assign n37368 = ~n37322 & ~n37353 ;
  assign n37369 = ~n37341 & n37348 ;
  assign n37370 = n37334 & ~n37350 ;
  assign n37371 = ~n37369 & ~n37370 ;
  assign n37372 = n37368 & ~n37371 ;
  assign n37373 = n37335 & n37341 ;
  assign n37374 = n37348 & n37373 ;
  assign n37375 = n37362 & ~n37374 ;
  assign n37376 = ~n37372 & n37375 ;
  assign n37386 = ~n37348 & n37351 ;
  assign n37387 = ~n37322 & n37386 ;
  assign n37381 = ~n37328 & n37334 ;
  assign n37388 = ~n37348 & n37381 ;
  assign n37389 = ~n37387 & ~n37388 ;
  assign n37390 = ~n37341 & ~n37389 ;
  assign n37377 = n37348 & n37352 ;
  assign n37378 = ~n37322 & n37377 ;
  assign n37380 = ~n37341 & ~n37348 ;
  assign n37382 = ~n37380 & ~n37381 ;
  assign n37383 = n37341 & n37348 ;
  assign n37384 = ~n37351 & ~n37383 ;
  assign n37385 = n37382 & n37384 ;
  assign n37379 = n37341 & n37354 ;
  assign n37391 = n37322 & ~n37341 ;
  assign n37392 = ~n37334 & n37348 ;
  assign n37393 = n37391 & n37392 ;
  assign n37394 = ~n37362 & ~n37393 ;
  assign n37395 = ~n37379 & n37394 ;
  assign n37396 = ~n37385 & n37395 ;
  assign n37397 = ~n37378 & n37396 ;
  assign n37398 = ~n37390 & n37397 ;
  assign n37399 = ~n37376 & ~n37398 ;
  assign n37400 = ~n37367 & ~n37399 ;
  assign n37401 = ~\u1_L8_reg[6]/NET0131  & ~n37400 ;
  assign n37402 = \u1_L8_reg[6]/NET0131  & n37400 ;
  assign n37403 = ~n37401 & ~n37402 ;
  assign n37420 = n36639 & n36663 ;
  assign n37421 = ~n36888 & ~n37420 ;
  assign n37422 = n36636 & ~n37421 ;
  assign n37423 = n36625 & ~n36636 ;
  assign n37424 = n36687 & ~n37423 ;
  assign n37425 = ~n37422 & n37424 ;
  assign n37426 = n36660 & ~n37425 ;
  assign n37404 = n36610 & ~n36669 ;
  assign n37405 = n36889 & ~n37404 ;
  assign n37406 = n36625 & n36639 ;
  assign n37407 = n36636 & ~n37406 ;
  assign n37408 = ~n37405 & ~n37407 ;
  assign n37409 = n36636 & n36667 ;
  assign n37410 = ~n36629 & ~n37409 ;
  assign n37411 = n36884 & n37410 ;
  assign n37412 = ~n37408 & n37411 ;
  assign n37413 = ~n36660 & ~n37412 ;
  assign n37414 = ~n36636 & ~n36670 ;
  assign n37415 = ~n36628 & ~n36669 ;
  assign n37416 = ~n36610 & n36636 ;
  assign n37417 = ~n37415 & ~n37416 ;
  assign n37418 = ~n36882 & ~n37417 ;
  assign n37419 = ~n37414 & ~n37418 ;
  assign n37427 = ~n37413 & ~n37419 ;
  assign n37428 = ~n37426 & n37427 ;
  assign n37429 = ~\u1_L8_reg[8]/NET0131  & ~n37428 ;
  assign n37430 = \u1_L8_reg[8]/NET0131  & n37428 ;
  assign n37431 = ~n37429 & ~n37430 ;
  assign n37432 = n36168 & ~n36217 ;
  assign n37433 = n36225 & n36562 ;
  assign n37434 = ~n36571 & ~n37285 ;
  assign n37435 = ~n37433 & n37434 ;
  assign n37436 = n37432 & ~n37435 ;
  assign n37439 = ~n36200 & n37285 ;
  assign n37437 = ~n36572 & ~n37433 ;
  assign n37438 = ~n36168 & n36217 ;
  assign n37440 = ~n37432 & ~n37438 ;
  assign n37441 = n37437 & n37440 ;
  assign n37442 = ~n37439 & n37441 ;
  assign n37443 = ~n37436 & ~n37442 ;
  assign n37444 = ~n36201 & ~n37443 ;
  assign n37446 = ~n36187 & ~n36569 ;
  assign n37445 = n36562 & ~n36566 ;
  assign n37447 = n37438 & ~n37445 ;
  assign n37448 = ~n37446 & n37447 ;
  assign n37449 = n37437 & n37448 ;
  assign n37450 = ~n37444 & ~n37449 ;
  assign n37451 = ~\u1_L8_reg[7]/NET0131  & n37450 ;
  assign n37452 = \u1_L8_reg[7]/NET0131  & ~n37450 ;
  assign n37453 = ~n37451 & ~n37452 ;
  assign n37454 = ~n37322 & n37382 ;
  assign n37455 = ~n37348 & n37391 ;
  assign n37456 = ~n37454 & ~n37455 ;
  assign n37457 = ~n37351 & ~n37456 ;
  assign n37458 = n37334 & n37383 ;
  assign n37459 = ~n37352 & ~n37458 ;
  assign n37460 = n37322 & ~n37459 ;
  assign n37461 = n37362 & ~n37460 ;
  assign n37462 = ~n37390 & n37461 ;
  assign n37463 = ~n37457 & n37462 ;
  assign n37468 = ~n37341 & n37351 ;
  assign n37469 = n37322 & ~n37373 ;
  assign n37470 = ~n37468 & n37469 ;
  assign n37466 = ~n37328 & n37392 ;
  assign n37464 = n37341 & ~n37348 ;
  assign n37467 = n37334 & n37464 ;
  assign n37471 = ~n37466 & ~n37467 ;
  assign n37472 = n37470 & n37471 ;
  assign n37473 = ~n37351 & n37380 ;
  assign n37474 = ~n37381 & n37473 ;
  assign n37475 = ~n37322 & n37355 ;
  assign n37476 = ~n37474 & n37475 ;
  assign n37477 = ~n37472 & ~n37476 ;
  assign n37465 = n37381 & n37464 ;
  assign n37478 = ~n37362 & ~n37465 ;
  assign n37479 = ~n37477 & n37478 ;
  assign n37480 = ~n37463 & ~n37479 ;
  assign n37483 = ~n37322 & n37341 ;
  assign n37484 = n37328 & n37334 ;
  assign n37485 = n37348 & n37484 ;
  assign n37486 = n37483 & n37485 ;
  assign n37481 = n37381 & n37455 ;
  assign n37482 = n37328 & n37393 ;
  assign n37487 = ~n37481 & ~n37482 ;
  assign n37488 = ~n37486 & n37487 ;
  assign n37489 = ~n37480 & n37488 ;
  assign n37490 = ~\u1_L8_reg[24]/NET0131  & ~n37489 ;
  assign n37491 = \u1_L8_reg[24]/NET0131  & n37489 ;
  assign n37492 = ~n37490 & ~n37491 ;
  assign n37496 = n37334 & n37341 ;
  assign n37497 = ~n37322 & ~n37496 ;
  assign n37498 = ~n37466 & n37497 ;
  assign n37499 = ~n37470 & ~n37498 ;
  assign n37500 = n37383 & ~n37484 ;
  assign n37501 = n37362 & ~n37500 ;
  assign n37502 = ~n37481 & n37501 ;
  assign n37503 = ~n37499 & n37502 ;
  assign n37505 = ~n37353 & n37496 ;
  assign n37506 = ~n37328 & n37369 ;
  assign n37507 = ~n37505 & ~n37506 ;
  assign n37508 = n37322 & ~n37507 ;
  assign n37509 = ~n37334 & ~n37348 ;
  assign n37510 = ~n37496 & ~n37509 ;
  assign n37511 = n37368 & n37510 ;
  assign n37504 = n37351 & n37464 ;
  assign n37512 = ~n37362 & ~n37504 ;
  assign n37513 = ~n37474 & n37512 ;
  assign n37514 = ~n37511 & n37513 ;
  assign n37515 = ~n37508 & n37514 ;
  assign n37516 = ~n37503 & ~n37515 ;
  assign n37493 = n37322 & n37464 ;
  assign n37494 = n37484 & n37493 ;
  assign n37495 = n37353 & n37483 ;
  assign n37517 = ~n37494 & ~n37495 ;
  assign n37518 = ~n37516 & n37517 ;
  assign n37519 = \u1_L8_reg[30]/NET0131  & ~n37518 ;
  assign n37520 = ~\u1_L8_reg[30]/NET0131  & n37518 ;
  assign n37521 = ~n37519 & ~n37520 ;
  assign n37523 = n36660 & ~n36670 ;
  assign n37524 = ~n36881 & n37523 ;
  assign n37525 = ~n36901 & n37524 ;
  assign n37526 = ~n36609 & n36669 ;
  assign n37527 = ~n36660 & ~n37526 ;
  assign n37528 = n36649 & ~n36888 ;
  assign n37529 = n37527 & n37528 ;
  assign n37530 = ~n37525 & ~n37529 ;
  assign n37531 = ~n36636 & ~n36680 ;
  assign n37522 = n36648 & n36650 ;
  assign n37532 = ~n37420 & ~n37522 ;
  assign n37533 = n37531 & n37532 ;
  assign n37534 = ~n37530 & n37533 ;
  assign n37535 = ~n36609 & ~n36626 ;
  assign n37536 = n37524 & ~n37535 ;
  assign n37537 = ~n36618 & ~n36663 ;
  assign n37538 = ~n36647 & ~n37537 ;
  assign n37539 = n37527 & ~n37538 ;
  assign n37540 = ~n37536 & ~n37539 ;
  assign n37541 = ~n36685 & n37407 ;
  assign n37542 = ~n37540 & n37541 ;
  assign n37543 = ~n37534 & ~n37542 ;
  assign n37544 = ~\u1_L8_reg[3]/NET0131  & n37543 ;
  assign n37545 = \u1_L8_reg[3]/NET0131  & ~n37543 ;
  assign n37546 = ~n37544 & ~n37545 ;
  assign n37563 = ~n36784 & ~n37212 ;
  assign n37564 = n36796 & ~n37563 ;
  assign n37547 = n36777 & ~n36804 ;
  assign n37561 = n36790 & ~n36796 ;
  assign n37562 = n37547 & n37561 ;
  assign n37565 = ~n36823 & ~n37562 ;
  assign n37566 = ~n37564 & n37565 ;
  assign n37567 = n36819 & ~n37566 ;
  assign n37548 = ~n36790 & n37547 ;
  assign n37550 = n36768 & n36826 ;
  assign n37551 = n36774 & n37550 ;
  assign n37554 = ~n37548 & ~n37551 ;
  assign n37549 = n36796 & n36807 ;
  assign n37552 = ~n36777 & n36790 ;
  assign n37553 = ~n37550 & n37552 ;
  assign n37555 = ~n37549 & ~n37553 ;
  assign n37556 = n37554 & n37555 ;
  assign n37557 = ~n36819 & ~n37556 ;
  assign n37558 = ~n36783 & n36832 ;
  assign n37559 = ~n37551 & ~n37558 ;
  assign n37560 = ~n36790 & ~n37559 ;
  assign n37568 = ~n37557 & ~n37560 ;
  assign n37569 = ~n37567 & n37568 ;
  assign n37570 = ~\u1_L8_reg[9]/NET0131  & ~n37569 ;
  assign n37571 = \u1_L8_reg[9]/NET0131  & n37569 ;
  assign n37572 = ~n37570 & ~n37571 ;
  assign n37577 = n37004 & ~n37042 ;
  assign n37574 = n37010 & n37045 ;
  assign n37575 = ~n37059 & ~n37574 ;
  assign n37576 = ~n37004 & ~n37575 ;
  assign n37578 = ~n37078 & ~n37576 ;
  assign n37579 = ~n37577 & n37578 ;
  assign n37580 = n36998 & ~n37579 ;
  assign n37581 = n37017 & n37057 ;
  assign n37584 = ~n37087 & ~n37175 ;
  assign n37585 = ~n37581 & n37584 ;
  assign n37582 = ~n37010 & ~n37057 ;
  assign n37583 = ~n37072 & n37582 ;
  assign n37586 = ~n37031 & ~n37583 ;
  assign n37587 = n37585 & n37586 ;
  assign n37588 = ~n36998 & ~n37587 ;
  assign n37573 = ~n37004 & n37091 ;
  assign n37589 = n37017 & n37030 ;
  assign n37590 = ~n37173 & ~n37589 ;
  assign n37591 = n37004 & ~n37590 ;
  assign n37592 = ~n37573 & ~n37591 ;
  assign n37593 = ~n37588 & n37592 ;
  assign n37594 = ~n37580 & n37593 ;
  assign n37595 = \u1_L8_reg[18]/NET0131  & n37594 ;
  assign n37596 = ~\u1_L8_reg[18]/NET0131  & ~n37594 ;
  assign n37597 = ~n37595 & ~n37596 ;
  assign n37647 = decrypt_pad & ~\u1_uk_K_r7_reg[54]/NET0131  ;
  assign n37648 = ~decrypt_pad & ~\u1_uk_K_r7_reg[47]/NET0131  ;
  assign n37649 = ~n37647 & ~n37648 ;
  assign n37650 = \u1_R7_reg[4]/NET0131  & ~n37649 ;
  assign n37651 = ~\u1_R7_reg[4]/NET0131  & n37649 ;
  assign n37652 = ~n37650 & ~n37651 ;
  assign n37598 = decrypt_pad & ~\u1_uk_K_r7_reg[6]/NET0131  ;
  assign n37599 = ~decrypt_pad & ~\u1_uk_K_r7_reg[24]/NET0131  ;
  assign n37600 = ~n37598 & ~n37599 ;
  assign n37601 = \u1_R7_reg[32]/NET0131  & ~n37600 ;
  assign n37602 = ~\u1_R7_reg[32]/NET0131  & n37600 ;
  assign n37603 = ~n37601 & ~n37602 ;
  assign n37618 = decrypt_pad & ~\u1_uk_K_r7_reg[25]/NET0131  ;
  assign n37619 = ~decrypt_pad & ~\u1_uk_K_r7_reg[18]/NET0131  ;
  assign n37620 = ~n37618 & ~n37619 ;
  assign n37621 = \u1_R7_reg[5]/NET0131  & ~n37620 ;
  assign n37622 = ~\u1_R7_reg[5]/NET0131  & n37620 ;
  assign n37623 = ~n37621 & ~n37622 ;
  assign n37628 = decrypt_pad & ~\u1_uk_K_r7_reg[27]/NET0131  ;
  assign n37629 = ~decrypt_pad & ~\u1_uk_K_r7_reg[20]/NET0131  ;
  assign n37630 = ~n37628 & ~n37629 ;
  assign n37631 = \u1_R7_reg[1]/NET0131  & ~n37630 ;
  assign n37632 = ~\u1_R7_reg[1]/NET0131  & n37630 ;
  assign n37633 = ~n37631 & ~n37632 ;
  assign n37635 = n37623 & ~n37633 ;
  assign n37611 = decrypt_pad & ~\u1_uk_K_r7_reg[19]/NET0131  ;
  assign n37612 = ~decrypt_pad & ~\u1_uk_K_r7_reg[12]/NET0131  ;
  assign n37613 = ~n37611 & ~n37612 ;
  assign n37614 = \u1_R7_reg[3]/NET0131  & ~n37613 ;
  assign n37615 = ~\u1_R7_reg[3]/NET0131  & n37613 ;
  assign n37616 = ~n37614 & ~n37615 ;
  assign n37655 = ~n37616 & n37633 ;
  assign n37604 = decrypt_pad & ~\u1_uk_K_r7_reg[10]/NET0131  ;
  assign n37605 = ~decrypt_pad & ~\u1_uk_K_r7_reg[3]/NET0131  ;
  assign n37606 = ~n37604 & ~n37605 ;
  assign n37607 = \u1_R7_reg[2]/NET0131  & ~n37606 ;
  assign n37608 = ~\u1_R7_reg[2]/NET0131  & n37606 ;
  assign n37609 = ~n37607 & ~n37608 ;
  assign n37639 = n37609 & ~n37623 ;
  assign n37642 = ~n37609 & n37623 ;
  assign n37660 = ~n37639 & ~n37642 ;
  assign n37661 = ~n37655 & ~n37660 ;
  assign n37662 = ~n37635 & ~n37661 ;
  assign n37663 = ~n37603 & ~n37662 ;
  assign n37654 = n37616 & n37635 ;
  assign n37656 = ~n37623 & ~n37633 ;
  assign n37657 = ~n37609 & n37656 ;
  assign n37658 = ~n37655 & ~n37657 ;
  assign n37659 = n37603 & ~n37658 ;
  assign n37664 = ~n37654 & ~n37659 ;
  assign n37665 = ~n37663 & n37664 ;
  assign n37666 = n37652 & ~n37665 ;
  assign n37610 = ~n37603 & n37609 ;
  assign n37617 = n37610 & n37616 ;
  assign n37624 = n37617 & n37623 ;
  assign n37625 = ~n37603 & ~n37623 ;
  assign n37626 = ~n37609 & n37625 ;
  assign n37627 = ~n37624 & ~n37626 ;
  assign n37634 = ~n37627 & n37633 ;
  assign n37636 = n37603 & ~n37609 ;
  assign n37637 = n37635 & n37636 ;
  assign n37638 = ~n37616 & ~n37637 ;
  assign n37640 = n37603 & n37633 ;
  assign n37641 = n37639 & n37640 ;
  assign n37643 = n37603 & n37642 ;
  assign n37644 = ~n37641 & ~n37643 ;
  assign n37645 = ~n37638 & ~n37644 ;
  assign n37646 = ~n37634 & ~n37645 ;
  assign n37653 = ~n37646 & ~n37652 ;
  assign n37667 = n37610 & n37635 ;
  assign n37668 = ~n37603 & n37623 ;
  assign n37669 = n37633 & ~n37668 ;
  assign n37670 = n37660 & n37669 ;
  assign n37671 = ~n37667 & ~n37670 ;
  assign n37672 = ~n37616 & ~n37671 ;
  assign n37678 = ~n37616 & ~n37640 ;
  assign n37677 = ~n37610 & ~n37636 ;
  assign n37679 = ~n37635 & ~n37652 ;
  assign n37680 = n37677 & n37679 ;
  assign n37681 = n37678 & n37680 ;
  assign n37673 = n37603 & ~n37633 ;
  assign n37674 = ~n37609 & n37616 ;
  assign n37675 = n37673 & n37674 ;
  assign n37676 = n37617 & n37656 ;
  assign n37682 = ~n37675 & ~n37676 ;
  assign n37683 = ~n37681 & n37682 ;
  assign n37684 = ~n37672 & n37683 ;
  assign n37685 = ~n37653 & n37684 ;
  assign n37686 = ~n37666 & n37685 ;
  assign n37687 = ~\u1_L7_reg[31]/NET0131  & ~n37686 ;
  assign n37688 = \u1_L7_reg[31]/NET0131  & n37686 ;
  assign n37689 = ~n37687 & ~n37688 ;
  assign n37724 = decrypt_pad & ~\u1_uk_K_r7_reg[23]/P0001  ;
  assign n37725 = ~decrypt_pad & ~\u1_uk_K_r7_reg[16]/NET0131  ;
  assign n37726 = ~n37724 & ~n37725 ;
  assign n37727 = \u1_R7_reg[24]/NET0131  & ~n37726 ;
  assign n37728 = ~\u1_R7_reg[24]/NET0131  & n37726 ;
  assign n37729 = ~n37727 & ~n37728 ;
  assign n37690 = decrypt_pad & ~\u1_uk_K_r7_reg[8]/NET0131  ;
  assign n37691 = ~decrypt_pad & ~\u1_uk_K_r7_reg[1]/NET0131  ;
  assign n37692 = ~n37690 & ~n37691 ;
  assign n37693 = \u1_R7_reg[22]/NET0131  & ~n37692 ;
  assign n37694 = ~\u1_R7_reg[22]/NET0131  & n37692 ;
  assign n37695 = ~n37693 & ~n37694 ;
  assign n37703 = decrypt_pad & ~\u1_uk_K_r7_reg[2]/NET0131  ;
  assign n37704 = ~decrypt_pad & ~\u1_uk_K_r7_reg[50]/NET0131  ;
  assign n37705 = ~n37703 & ~n37704 ;
  assign n37706 = \u1_R7_reg[20]/NET0131  & ~n37705 ;
  assign n37707 = ~\u1_R7_reg[20]/NET0131  & n37705 ;
  assign n37708 = ~n37706 & ~n37707 ;
  assign n37716 = decrypt_pad & ~\u1_uk_K_r7_reg[45]/NET0131  ;
  assign n37717 = ~decrypt_pad & ~\u1_uk_K_r7_reg[38]/NET0131  ;
  assign n37718 = ~n37716 & ~n37717 ;
  assign n37719 = \u1_R7_reg[21]/NET0131  & ~n37718 ;
  assign n37720 = ~\u1_R7_reg[21]/NET0131  & n37718 ;
  assign n37721 = ~n37719 & ~n37720 ;
  assign n37732 = ~n37708 & n37721 ;
  assign n37709 = decrypt_pad & ~\u1_uk_K_r7_reg[42]/NET0131  ;
  assign n37710 = ~decrypt_pad & ~\u1_uk_K_r7_reg[35]/NET0131  ;
  assign n37711 = ~n37709 & ~n37710 ;
  assign n37712 = \u1_R7_reg[25]/NET0131  & ~n37711 ;
  assign n37713 = ~\u1_R7_reg[25]/NET0131  & n37711 ;
  assign n37714 = ~n37712 & ~n37713 ;
  assign n37740 = n37708 & n37714 ;
  assign n37745 = ~n37732 & ~n37740 ;
  assign n37746 = n37695 & ~n37745 ;
  assign n37696 = decrypt_pad & ~\u1_uk_K_r7_reg[21]/NET0131  ;
  assign n37697 = ~decrypt_pad & ~\u1_uk_K_r7_reg[14]/NET0131  ;
  assign n37698 = ~n37696 & ~n37697 ;
  assign n37699 = \u1_R7_reg[23]/NET0131  & ~n37698 ;
  assign n37700 = ~\u1_R7_reg[23]/NET0131  & n37698 ;
  assign n37701 = ~n37699 & ~n37700 ;
  assign n37730 = n37714 & n37721 ;
  assign n37743 = ~n37708 & n37730 ;
  assign n37744 = ~n37695 & ~n37743 ;
  assign n37747 = ~n37701 & ~n37744 ;
  assign n37748 = ~n37746 & n37747 ;
  assign n37734 = n37708 & ~n37714 ;
  assign n37735 = ~n37695 & ~n37721 ;
  assign n37736 = n37734 & n37735 ;
  assign n37731 = n37708 & n37730 ;
  assign n37733 = n37695 & n37732 ;
  assign n37737 = ~n37731 & ~n37733 ;
  assign n37738 = ~n37736 & n37737 ;
  assign n37739 = n37701 & ~n37738 ;
  assign n37702 = ~n37695 & ~n37701 ;
  assign n37741 = n37702 & n37740 ;
  assign n37742 = ~n37721 & n37741 ;
  assign n37749 = ~n37739 & ~n37742 ;
  assign n37750 = ~n37748 & n37749 ;
  assign n37751 = n37729 & ~n37750 ;
  assign n37758 = ~n37714 & n37721 ;
  assign n37759 = n37708 & ~n37758 ;
  assign n37760 = ~n37701 & ~n37708 ;
  assign n37761 = ~n37695 & ~n37760 ;
  assign n37762 = ~n37759 & n37761 ;
  assign n37752 = ~n37708 & n37714 ;
  assign n37753 = ~n37721 & n37752 ;
  assign n37754 = n37701 & n37753 ;
  assign n37755 = n37708 & ~n37721 ;
  assign n37756 = n37695 & n37701 ;
  assign n37757 = n37755 & n37756 ;
  assign n37771 = ~n37754 & ~n37757 ;
  assign n37772 = ~n37762 & n37771 ;
  assign n37763 = n37695 & n37740 ;
  assign n37764 = ~n37721 & n37763 ;
  assign n37765 = n37702 & n37734 ;
  assign n37766 = ~n37764 & ~n37765 ;
  assign n37767 = ~n37695 & n37721 ;
  assign n37768 = n37708 & n37767 ;
  assign n37769 = ~n37733 & ~n37768 ;
  assign n37770 = ~n37701 & ~n37769 ;
  assign n37773 = n37766 & ~n37770 ;
  assign n37774 = n37772 & n37773 ;
  assign n37775 = ~n37729 & ~n37774 ;
  assign n37776 = n37721 & n37734 ;
  assign n37777 = ~n37701 & n37776 ;
  assign n37778 = ~n37754 & ~n37777 ;
  assign n37779 = ~n37695 & ~n37778 ;
  assign n37715 = ~n37708 & ~n37714 ;
  assign n37722 = n37715 & ~n37721 ;
  assign n37723 = n37702 & n37722 ;
  assign n37780 = n37715 & n37767 ;
  assign n37781 = ~n37763 & ~n37780 ;
  assign n37782 = n37701 & ~n37781 ;
  assign n37783 = ~n37723 & ~n37782 ;
  assign n37784 = ~n37779 & n37783 ;
  assign n37785 = ~n37775 & n37784 ;
  assign n37786 = ~n37751 & n37785 ;
  assign n37787 = \u1_L7_reg[11]/NET0131  & ~n37786 ;
  assign n37788 = ~\u1_L7_reg[11]/NET0131  & n37786 ;
  assign n37789 = ~n37787 & ~n37788 ;
  assign n37790 = decrypt_pad & ~\u1_uk_K_r7_reg[30]/P0001  ;
  assign n37791 = ~decrypt_pad & ~\u1_uk_K_r7_reg[23]/P0001  ;
  assign n37792 = ~n37790 & ~n37791 ;
  assign n37793 = \u1_R7_reg[28]/NET0131  & ~n37792 ;
  assign n37794 = ~\u1_R7_reg[28]/NET0131  & n37792 ;
  assign n37795 = ~n37793 & ~n37794 ;
  assign n37796 = decrypt_pad & ~\u1_uk_K_r7_reg[38]/NET0131  ;
  assign n37797 = ~decrypt_pad & ~\u1_uk_K_r7_reg[31]/NET0131  ;
  assign n37798 = ~n37796 & ~n37797 ;
  assign n37799 = \u1_R7_reg[26]/NET0131  & ~n37798 ;
  assign n37800 = ~\u1_R7_reg[26]/NET0131  & n37798 ;
  assign n37801 = ~n37799 & ~n37800 ;
  assign n37802 = decrypt_pad & ~\u1_uk_K_r7_reg[49]/NET0131  ;
  assign n37803 = ~decrypt_pad & ~\u1_uk_K_r7_reg[42]/NET0131  ;
  assign n37804 = ~n37802 & ~n37803 ;
  assign n37805 = \u1_R7_reg[25]/NET0131  & ~n37804 ;
  assign n37806 = ~\u1_R7_reg[25]/NET0131  & n37804 ;
  assign n37807 = ~n37805 & ~n37806 ;
  assign n37836 = ~n37801 & ~n37807 ;
  assign n37808 = decrypt_pad & ~\u1_uk_K_r7_reg[22]/NET0131  ;
  assign n37809 = ~decrypt_pad & ~\u1_uk_K_r7_reg[15]/NET0131  ;
  assign n37810 = ~n37808 & ~n37809 ;
  assign n37811 = \u1_R7_reg[29]/NET0131  & ~n37810 ;
  assign n37812 = ~\u1_R7_reg[29]/NET0131  & n37810 ;
  assign n37813 = ~n37811 & ~n37812 ;
  assign n37839 = ~n37801 & ~n37813 ;
  assign n37859 = ~n37836 & ~n37839 ;
  assign n37815 = decrypt_pad & ~\u1_uk_K_r7_reg[14]/NET0131  ;
  assign n37816 = ~decrypt_pad & ~\u1_uk_K_r7_reg[7]/NET0131  ;
  assign n37817 = ~n37815 & ~n37816 ;
  assign n37818 = \u1_R7_reg[24]/NET0131  & ~n37817 ;
  assign n37819 = ~\u1_R7_reg[24]/NET0131  & n37817 ;
  assign n37820 = ~n37818 & ~n37819 ;
  assign n37823 = decrypt_pad & ~\u1_uk_K_r7_reg[43]/NET0131  ;
  assign n37824 = ~decrypt_pad & ~\u1_uk_K_r7_reg[36]/NET0131  ;
  assign n37825 = ~n37823 & ~n37824 ;
  assign n37826 = \u1_R7_reg[27]/NET0131  & ~n37825 ;
  assign n37827 = ~\u1_R7_reg[27]/NET0131  & n37825 ;
  assign n37828 = ~n37826 & ~n37827 ;
  assign n37838 = n37801 & n37807 ;
  assign n37858 = n37828 & ~n37838 ;
  assign n37860 = n37820 & n37858 ;
  assign n37861 = n37859 & n37860 ;
  assign n37852 = n37813 & n37820 ;
  assign n37853 = n37836 & n37852 ;
  assign n37854 = n37807 & n37813 ;
  assign n37855 = ~n37820 & n37854 ;
  assign n37856 = ~n37853 & ~n37855 ;
  assign n37857 = ~n37828 & ~n37856 ;
  assign n37847 = ~n37813 & ~n37820 ;
  assign n37848 = n37836 & n37847 ;
  assign n37849 = n37813 & ~n37820 ;
  assign n37850 = n37801 & ~n37807 ;
  assign n37851 = n37849 & n37850 ;
  assign n37862 = ~n37848 & ~n37851 ;
  assign n37863 = ~n37857 & n37862 ;
  assign n37864 = ~n37861 & n37863 ;
  assign n37865 = n37795 & ~n37864 ;
  assign n37840 = ~n37828 & ~n37838 ;
  assign n37841 = ~n37839 & n37840 ;
  assign n37837 = n37828 & ~n37836 ;
  assign n37842 = n37820 & ~n37837 ;
  assign n37843 = ~n37841 & n37842 ;
  assign n37814 = ~n37807 & ~n37813 ;
  assign n37821 = n37814 & ~n37820 ;
  assign n37822 = n37801 & n37821 ;
  assign n37829 = n37822 & ~n37828 ;
  assign n37830 = ~n37801 & ~n37820 ;
  assign n37831 = n37801 & n37820 ;
  assign n37832 = ~n37830 & ~n37831 ;
  assign n37833 = ~n37807 & n37828 ;
  assign n37834 = n37813 & ~n37833 ;
  assign n37835 = ~n37832 & n37834 ;
  assign n37844 = ~n37829 & ~n37835 ;
  assign n37845 = ~n37843 & n37844 ;
  assign n37846 = ~n37795 & ~n37845 ;
  assign n37868 = n37838 & n37847 ;
  assign n37869 = ~n37851 & ~n37868 ;
  assign n37870 = ~n37813 & n37820 ;
  assign n37871 = ~n37807 & n37870 ;
  assign n37872 = n37869 & ~n37871 ;
  assign n37873 = n37828 & ~n37872 ;
  assign n37866 = n37807 & ~n37828 ;
  assign n37867 = ~n37832 & n37866 ;
  assign n37874 = n37833 & n37839 ;
  assign n37875 = ~n37867 & ~n37874 ;
  assign n37876 = ~n37873 & n37875 ;
  assign n37877 = ~n37846 & n37876 ;
  assign n37878 = ~n37865 & n37877 ;
  assign n37879 = ~\u1_L7_reg[22]/NET0131  & ~n37878 ;
  assign n37880 = \u1_L7_reg[22]/NET0131  & n37878 ;
  assign n37881 = ~n37879 & ~n37880 ;
  assign n37888 = ~n37609 & ~n37633 ;
  assign n37889 = ~n37603 & ~n37888 ;
  assign n37890 = ~n37637 & ~n37889 ;
  assign n37891 = n37616 & ~n37890 ;
  assign n37882 = ~n37623 & n37636 ;
  assign n37883 = n37633 & n37882 ;
  assign n37884 = n37652 & ~n37883 ;
  assign n37885 = ~n37603 & n37633 ;
  assign n37886 = ~n37616 & ~n37885 ;
  assign n37887 = n37677 & n37886 ;
  assign n37892 = n37623 & n37633 ;
  assign n37893 = n37609 & n37892 ;
  assign n37894 = ~n37887 & ~n37893 ;
  assign n37895 = n37884 & n37894 ;
  assign n37896 = ~n37891 & n37895 ;
  assign n37897 = n37603 & n37623 ;
  assign n37898 = ~n37625 & ~n37897 ;
  assign n37899 = ~n37633 & ~n37898 ;
  assign n37900 = ~n37616 & ~n37626 ;
  assign n37901 = ~n37899 & n37900 ;
  assign n37903 = ~n37656 & ~n37892 ;
  assign n37904 = n37603 & ~n37903 ;
  assign n37902 = ~n37660 & n37885 ;
  assign n37905 = n37616 & ~n37902 ;
  assign n37906 = ~n37904 & n37905 ;
  assign n37907 = ~n37901 & ~n37906 ;
  assign n37908 = ~n37641 & ~n37652 ;
  assign n37909 = ~n37667 & n37908 ;
  assign n37910 = ~n37907 & n37909 ;
  assign n37911 = ~n37896 & ~n37910 ;
  assign n37912 = ~\u1_L7_reg[17]/NET0131  & n37911 ;
  assign n37913 = \u1_L7_reg[17]/NET0131  & ~n37911 ;
  assign n37914 = ~n37912 & ~n37913 ;
  assign n37927 = decrypt_pad & ~\u1_uk_K_r7_reg[20]/NET0131  ;
  assign n37928 = ~decrypt_pad & ~\u1_uk_K_r7_reg[13]/NET0131  ;
  assign n37929 = ~n37927 & ~n37928 ;
  assign n37930 = \u1_R7_reg[12]/NET0131  & ~n37929 ;
  assign n37931 = ~\u1_R7_reg[12]/NET0131  & n37929 ;
  assign n37932 = ~n37930 & ~n37931 ;
  assign n37940 = decrypt_pad & ~\u1_uk_K_r7_reg[39]/NET0131  ;
  assign n37941 = ~decrypt_pad & ~\u1_uk_K_r7_reg[32]/NET0131  ;
  assign n37942 = ~n37940 & ~n37941 ;
  assign n37943 = \u1_R7_reg[13]/NET0131  & ~n37942 ;
  assign n37944 = ~\u1_R7_reg[13]/NET0131  & n37942 ;
  assign n37945 = ~n37943 & ~n37944 ;
  assign n37915 = decrypt_pad & ~\u1_uk_K_r7_reg[48]/NET0131  ;
  assign n37916 = ~decrypt_pad & ~\u1_uk_K_r7_reg[41]/NET0131  ;
  assign n37917 = ~n37915 & ~n37916 ;
  assign n37918 = \u1_R7_reg[15]/NET0131  & ~n37917 ;
  assign n37919 = ~\u1_R7_reg[15]/NET0131  & n37917 ;
  assign n37920 = ~n37918 & ~n37919 ;
  assign n37934 = decrypt_pad & ~\u1_uk_K_r7_reg[40]/NET0131  ;
  assign n37935 = ~decrypt_pad & ~\u1_uk_K_r7_reg[33]/NET0131  ;
  assign n37936 = ~n37934 & ~n37935 ;
  assign n37937 = \u1_R7_reg[14]/NET0131  & ~n37936 ;
  assign n37938 = ~\u1_R7_reg[14]/NET0131  & n37936 ;
  assign n37939 = ~n37937 & ~n37938 ;
  assign n37968 = n37920 & n37939 ;
  assign n37969 = n37945 & n37968 ;
  assign n37970 = ~n37932 & n37969 ;
  assign n37921 = decrypt_pad & ~\u1_uk_K_r7_reg[4]/NET0131  ;
  assign n37922 = ~decrypt_pad & ~\u1_uk_K_r7_reg[54]/NET0131  ;
  assign n37923 = ~n37921 & ~n37922 ;
  assign n37924 = \u1_R7_reg[17]/NET0131  & ~n37923 ;
  assign n37925 = ~\u1_R7_reg[17]/NET0131  & n37923 ;
  assign n37926 = ~n37924 & ~n37925 ;
  assign n37965 = ~n37939 & ~n37945 ;
  assign n37966 = n37932 & n37965 ;
  assign n37967 = n37926 & n37966 ;
  assign n37971 = decrypt_pad & ~\u1_uk_K_r7_reg[24]/NET0131  ;
  assign n37972 = ~decrypt_pad & ~\u1_uk_K_r7_reg[17]/NET0131  ;
  assign n37973 = ~n37971 & ~n37972 ;
  assign n37974 = \u1_R7_reg[16]/NET0131  & ~n37973 ;
  assign n37975 = ~\u1_R7_reg[16]/NET0131  & n37973 ;
  assign n37976 = ~n37974 & ~n37975 ;
  assign n37987 = ~n37967 & ~n37976 ;
  assign n37988 = ~n37970 & n37987 ;
  assign n37982 = ~n37932 & ~n37945 ;
  assign n37983 = n37932 & n37945 ;
  assign n37984 = ~n37982 & ~n37983 ;
  assign n37933 = n37926 & ~n37932 ;
  assign n37952 = ~n37926 & n37932 ;
  assign n37981 = ~n37933 & ~n37952 ;
  assign n37985 = n37920 & n37981 ;
  assign n37986 = ~n37984 & n37985 ;
  assign n37949 = ~n37926 & ~n37939 ;
  assign n37950 = ~n37932 & n37949 ;
  assign n37951 = ~n37945 & n37950 ;
  assign n37958 = ~n37926 & n37945 ;
  assign n37962 = ~n37932 & n37958 ;
  assign n37963 = n37939 & n37962 ;
  assign n37964 = ~n37951 & ~n37963 ;
  assign n37977 = n37926 & ~n37945 ;
  assign n37978 = n37939 & n37952 ;
  assign n37979 = ~n37977 & ~n37978 ;
  assign n37980 = ~n37920 & ~n37979 ;
  assign n37989 = n37964 & ~n37980 ;
  assign n37990 = ~n37986 & n37989 ;
  assign n37991 = n37988 & n37990 ;
  assign n37992 = ~n37926 & n37982 ;
  assign n37993 = ~n37920 & n37992 ;
  assign n37994 = n37939 & n37993 ;
  assign n37997 = ~n37920 & ~n37939 ;
  assign n37998 = n37984 & n37997 ;
  assign n37995 = n37926 & n37939 ;
  assign n37996 = n37983 & n37995 ;
  assign n38002 = n37976 & ~n37996 ;
  assign n38003 = ~n37998 & n38002 ;
  assign n37946 = ~n37939 & n37945 ;
  assign n37947 = n37933 & n37946 ;
  assign n37959 = n37920 & n37932 ;
  assign n37960 = n37958 & n37959 ;
  assign n37999 = ~n37947 & ~n37960 ;
  assign n38000 = n37920 & n37933 ;
  assign n38001 = ~n37945 & n38000 ;
  assign n38004 = n37999 & ~n38001 ;
  assign n38005 = n38003 & n38004 ;
  assign n38006 = ~n37994 & n38005 ;
  assign n38007 = ~n37991 & ~n38006 ;
  assign n37948 = ~n37920 & ~n37947 ;
  assign n37953 = n37939 & ~n37945 ;
  assign n37954 = n37952 & n37953 ;
  assign n37955 = n37920 & ~n37954 ;
  assign n37956 = ~n37951 & n37955 ;
  assign n37957 = ~n37948 & ~n37956 ;
  assign n37961 = ~n37939 & n37960 ;
  assign n38008 = ~n37957 & ~n37961 ;
  assign n38009 = ~n38007 & n38008 ;
  assign n38010 = ~\u1_L7_reg[20]/NET0131  & ~n38009 ;
  assign n38011 = \u1_L7_reg[20]/NET0131  & n38009 ;
  assign n38012 = ~n38010 & ~n38011 ;
  assign n38037 = n37695 & ~n37734 ;
  assign n38038 = ~n37752 & n38037 ;
  assign n38039 = ~n37722 & ~n38038 ;
  assign n38040 = ~n37701 & ~n38039 ;
  assign n38019 = n37695 & n37776 ;
  assign n38030 = n37695 & ~n37714 ;
  assign n38034 = n37732 & ~n38030 ;
  assign n38035 = ~n38019 & ~n38034 ;
  assign n38036 = n37701 & ~n38035 ;
  assign n38029 = ~n37695 & n37752 ;
  assign n38031 = ~n37708 & n38030 ;
  assign n38032 = ~n38029 & ~n38031 ;
  assign n38033 = ~n37721 & ~n38032 ;
  assign n38041 = n37766 & ~n38033 ;
  assign n38042 = ~n38036 & n38041 ;
  assign n38043 = ~n38040 & n38042 ;
  assign n38044 = n37729 & ~n38043 ;
  assign n38013 = ~n37721 & n37734 ;
  assign n38014 = ~n37731 & ~n38013 ;
  assign n38015 = ~n37733 & ~n37735 ;
  assign n38016 = ~n37714 & ~n38015 ;
  assign n38017 = n38014 & ~n38016 ;
  assign n38018 = n37701 & ~n38017 ;
  assign n38020 = ~n37695 & ~n37745 ;
  assign n38021 = ~n38019 & ~n38020 ;
  assign n38022 = ~n37701 & ~n38021 ;
  assign n38023 = n37695 & n37753 ;
  assign n38024 = ~n38022 & ~n38023 ;
  assign n38025 = ~n38018 & n38024 ;
  assign n38026 = ~n37729 & ~n38025 ;
  assign n38027 = ~n37695 & n37701 ;
  assign n38028 = n37730 & n38027 ;
  assign n38045 = ~n37736 & ~n38028 ;
  assign n38046 = ~n38026 & n38045 ;
  assign n38047 = ~n38044 & n38046 ;
  assign n38048 = \u1_L7_reg[29]/NET0131  & ~n38047 ;
  assign n38049 = ~\u1_L7_reg[29]/NET0131  & n38047 ;
  assign n38050 = ~n38048 & ~n38049 ;
  assign n38051 = decrypt_pad & ~\u1_uk_K_r7_reg[55]/P0001  ;
  assign n38052 = ~decrypt_pad & ~\u1_uk_K_r7_reg[48]/NET0131  ;
  assign n38053 = ~n38051 & ~n38052 ;
  assign n38054 = \u1_R7_reg[8]/NET0131  & ~n38053 ;
  assign n38055 = ~\u1_R7_reg[8]/NET0131  & n38053 ;
  assign n38056 = ~n38054 & ~n38055 ;
  assign n38057 = decrypt_pad & ~\u1_uk_K_r7_reg[32]/NET0131  ;
  assign n38058 = ~decrypt_pad & ~\u1_uk_K_r7_reg[25]/NET0131  ;
  assign n38059 = ~n38057 & ~n38058 ;
  assign n38060 = \u1_R7_reg[7]/NET0131  & ~n38059 ;
  assign n38061 = ~\u1_R7_reg[7]/NET0131  & n38059 ;
  assign n38062 = ~n38060 & ~n38061 ;
  assign n38076 = decrypt_pad & ~\u1_uk_K_r7_reg[47]/NET0131  ;
  assign n38077 = ~decrypt_pad & ~\u1_uk_K_r7_reg[40]/NET0131  ;
  assign n38078 = ~n38076 & ~n38077 ;
  assign n38079 = \u1_R7_reg[5]/NET0131  & ~n38078 ;
  assign n38080 = ~\u1_R7_reg[5]/NET0131  & n38078 ;
  assign n38081 = ~n38079 & ~n38080 ;
  assign n38063 = decrypt_pad & ~\u1_uk_K_r7_reg[11]/NET0131  ;
  assign n38064 = ~decrypt_pad & ~\u1_uk_K_r7_reg[4]/NET0131  ;
  assign n38065 = ~n38063 & ~n38064 ;
  assign n38066 = \u1_R7_reg[4]/NET0131  & ~n38065 ;
  assign n38067 = ~\u1_R7_reg[4]/NET0131  & n38065 ;
  assign n38068 = ~n38066 & ~n38067 ;
  assign n38069 = decrypt_pad & ~\u1_uk_K_r7_reg[3]/NET0131  ;
  assign n38070 = ~decrypt_pad & ~\u1_uk_K_r7_reg[53]/NET0131  ;
  assign n38071 = ~n38069 & ~n38070 ;
  assign n38072 = \u1_R7_reg[9]/NET0131  & ~n38071 ;
  assign n38073 = ~\u1_R7_reg[9]/NET0131  & n38071 ;
  assign n38074 = ~n38072 & ~n38073 ;
  assign n38091 = ~n38068 & n38074 ;
  assign n38092 = ~n38081 & n38091 ;
  assign n38083 = decrypt_pad & ~\u1_uk_K_r7_reg[13]/NET0131  ;
  assign n38084 = ~decrypt_pad & ~\u1_uk_K_r7_reg[6]/NET0131  ;
  assign n38085 = ~n38083 & ~n38084 ;
  assign n38086 = \u1_R7_reg[6]/NET0131  & ~n38085 ;
  assign n38087 = ~\u1_R7_reg[6]/NET0131  & n38085 ;
  assign n38088 = ~n38086 & ~n38087 ;
  assign n38093 = n38068 & n38081 ;
  assign n38094 = n38068 & ~n38074 ;
  assign n38095 = ~n38093 & ~n38094 ;
  assign n38096 = n38088 & ~n38095 ;
  assign n38097 = ~n38092 & ~n38096 ;
  assign n38098 = ~n38062 & ~n38097 ;
  assign n38099 = ~n38074 & n38081 ;
  assign n38100 = ~n38092 & ~n38099 ;
  assign n38101 = ~n38088 & ~n38100 ;
  assign n38075 = n38068 & n38074 ;
  assign n38082 = n38075 & ~n38081 ;
  assign n38089 = n38082 & n38088 ;
  assign n38090 = n38062 & n38089 ;
  assign n38102 = ~n38062 & ~n38081 ;
  assign n38103 = n38074 & ~n38088 ;
  assign n38104 = n38102 & n38103 ;
  assign n38105 = n38081 & n38088 ;
  assign n38106 = n38091 & n38105 ;
  assign n38107 = ~n38104 & ~n38106 ;
  assign n38108 = ~n38090 & n38107 ;
  assign n38109 = ~n38101 & n38108 ;
  assign n38110 = ~n38098 & n38109 ;
  assign n38111 = ~n38056 & ~n38110 ;
  assign n38128 = ~n38068 & ~n38074 ;
  assign n38129 = ~n38089 & ~n38128 ;
  assign n38130 = n38056 & ~n38129 ;
  assign n38112 = ~n38081 & n38088 ;
  assign n38131 = n38091 & ~n38112 ;
  assign n38132 = ~n38130 & ~n38131 ;
  assign n38127 = n38081 & ~n38088 ;
  assign n38133 = ~n38062 & ~n38127 ;
  assign n38134 = ~n38132 & n38133 ;
  assign n38113 = ~n38074 & n38112 ;
  assign n38114 = ~n38068 & n38113 ;
  assign n38115 = ~n38088 & n38093 ;
  assign n38116 = ~n38114 & ~n38115 ;
  assign n38117 = n38062 & ~n38116 ;
  assign n38118 = ~n38081 & n38094 ;
  assign n38119 = n38075 & n38081 ;
  assign n38120 = ~n38118 & ~n38119 ;
  assign n38121 = ~n38088 & ~n38120 ;
  assign n38122 = ~n38068 & n38088 ;
  assign n38123 = n38062 & n38081 ;
  assign n38124 = ~n38122 & n38123 ;
  assign n38125 = ~n38121 & ~n38124 ;
  assign n38126 = n38056 & ~n38125 ;
  assign n38135 = ~n38117 & ~n38126 ;
  assign n38136 = ~n38134 & n38135 ;
  assign n38137 = ~n38111 & n38136 ;
  assign n38138 = \u1_L7_reg[2]/NET0131  & n38137 ;
  assign n38139 = ~\u1_L7_reg[2]/NET0131  & ~n38137 ;
  assign n38140 = ~n38138 & ~n38139 ;
  assign n38158 = ~n37708 & n37758 ;
  assign n38159 = ~n38023 & ~n38158 ;
  assign n38160 = ~n37701 & ~n38159 ;
  assign n38155 = ~n37776 & ~n38029 ;
  assign n38156 = ~n37764 & n38155 ;
  assign n38157 = n37701 & ~n38156 ;
  assign n38161 = ~n37736 & ~n37741 ;
  assign n38162 = ~n38157 & n38161 ;
  assign n38163 = ~n38160 & n38162 ;
  assign n38164 = ~n37729 & ~n38163 ;
  assign n38142 = n37702 & ~n37759 ;
  assign n38143 = n37740 & n38027 ;
  assign n38141 = n37695 & n37730 ;
  assign n38144 = ~n37780 & ~n38141 ;
  assign n38145 = ~n38143 & n38144 ;
  assign n38146 = ~n38142 & n38145 ;
  assign n38147 = n37729 & ~n38146 ;
  assign n38148 = ~n37722 & ~n37743 ;
  assign n38149 = ~n37776 & n38148 ;
  assign n38150 = n37756 & ~n38149 ;
  assign n38151 = n37695 & n38014 ;
  assign n38152 = ~n37695 & ~n37715 ;
  assign n38153 = ~n37701 & ~n38152 ;
  assign n38154 = ~n38151 & n38153 ;
  assign n38165 = ~n38150 & ~n38154 ;
  assign n38166 = ~n38147 & n38165 ;
  assign n38167 = ~n38164 & n38166 ;
  assign n38168 = ~\u1_L7_reg[4]/NET0131  & ~n38167 ;
  assign n38169 = \u1_L7_reg[4]/NET0131  & n38167 ;
  assign n38170 = ~n38168 & ~n38169 ;
  assign n38217 = decrypt_pad & ~\u1_uk_K_r7_reg[50]/NET0131  ;
  assign n38218 = ~decrypt_pad & ~\u1_uk_K_r7_reg[43]/NET0131  ;
  assign n38219 = ~n38217 & ~n38218 ;
  assign n38220 = \u1_R7_reg[32]/NET0131  & ~n38219 ;
  assign n38221 = ~\u1_R7_reg[32]/NET0131  & n38219 ;
  assign n38222 = ~n38220 & ~n38221 ;
  assign n38191 = decrypt_pad & ~\u1_uk_K_r7_reg[44]/NET0131  ;
  assign n38192 = ~decrypt_pad & ~\u1_uk_K_r7_reg[37]/NET0131  ;
  assign n38193 = ~n38191 & ~n38192 ;
  assign n38194 = \u1_R7_reg[31]/P0001  & ~n38193 ;
  assign n38195 = ~\u1_R7_reg[31]/P0001  & n38193 ;
  assign n38196 = ~n38194 & ~n38195 ;
  assign n38184 = decrypt_pad & ~\u1_uk_K_r7_reg[28]/NET0131  ;
  assign n38185 = ~decrypt_pad & ~\u1_uk_K_r7_reg[21]/NET0131  ;
  assign n38186 = ~n38184 & ~n38185 ;
  assign n38187 = \u1_R7_reg[28]/NET0131  & ~n38186 ;
  assign n38188 = ~\u1_R7_reg[28]/NET0131  & n38186 ;
  assign n38189 = ~n38187 & ~n38188 ;
  assign n38177 = decrypt_pad & ~\u1_uk_K_r7_reg[0]/NET0131  ;
  assign n38178 = ~decrypt_pad & ~\u1_uk_K_r7_reg[52]/NET0131  ;
  assign n38179 = ~n38177 & ~n38178 ;
  assign n38180 = \u1_R7_reg[29]/NET0131  & ~n38179 ;
  assign n38181 = ~\u1_R7_reg[29]/NET0131  & n38179 ;
  assign n38182 = ~n38180 & ~n38181 ;
  assign n38199 = decrypt_pad & ~\u1_uk_K_r7_reg[16]/NET0131  ;
  assign n38200 = ~decrypt_pad & ~\u1_uk_K_r7_reg[9]/NET0131  ;
  assign n38201 = ~n38199 & ~n38200 ;
  assign n38202 = \u1_R7_reg[1]/NET0131  & ~n38201 ;
  assign n38203 = ~\u1_R7_reg[1]/NET0131  & n38201 ;
  assign n38204 = ~n38202 & ~n38203 ;
  assign n38224 = ~n38182 & n38204 ;
  assign n38225 = ~n38189 & n38224 ;
  assign n38171 = decrypt_pad & ~\u1_uk_K_r7_reg[1]/NET0131  ;
  assign n38172 = ~decrypt_pad & ~\u1_uk_K_r7_reg[49]/NET0131  ;
  assign n38173 = ~n38171 & ~n38172 ;
  assign n38174 = \u1_R7_reg[30]/NET0131  & ~n38173 ;
  assign n38175 = ~\u1_R7_reg[30]/NET0131  & n38173 ;
  assign n38176 = ~n38174 & ~n38175 ;
  assign n38235 = ~n38182 & n38189 ;
  assign n38236 = n38176 & n38235 ;
  assign n38247 = ~n38204 & n38236 ;
  assign n38248 = ~n38225 & ~n38247 ;
  assign n38249 = n38196 & ~n38248 ;
  assign n38198 = ~n38176 & n38189 ;
  assign n38241 = ~n38176 & ~n38204 ;
  assign n38207 = n38189 & ~n38204 ;
  assign n38242 = ~n38207 & ~n38224 ;
  assign n38243 = ~n38241 & n38242 ;
  assign n38244 = ~n38198 & ~n38243 ;
  assign n38245 = ~n38196 & ~n38244 ;
  assign n38208 = ~n38176 & n38182 ;
  assign n38209 = n38207 & n38208 ;
  assign n38213 = n38176 & n38182 ;
  assign n38230 = n38189 & n38204 ;
  assign n38246 = n38213 & n38230 ;
  assign n38250 = ~n38209 & ~n38246 ;
  assign n38251 = ~n38245 & n38250 ;
  assign n38252 = ~n38249 & n38251 ;
  assign n38253 = ~n38222 & ~n38252 ;
  assign n38183 = ~n38176 & ~n38182 ;
  assign n38190 = n38183 & ~n38189 ;
  assign n38197 = ~n38190 & ~n38196 ;
  assign n38205 = n38182 & ~n38204 ;
  assign n38206 = ~n38198 & ~n38205 ;
  assign n38210 = ~n38206 & ~n38209 ;
  assign n38211 = n38196 & ~n38210 ;
  assign n38212 = ~n38197 & ~n38211 ;
  assign n38214 = ~n38189 & n38213 ;
  assign n38215 = n38204 & n38214 ;
  assign n38216 = ~n38212 & ~n38215 ;
  assign n38223 = ~n38216 & n38222 ;
  assign n38227 = ~n38204 & n38214 ;
  assign n38228 = n38190 & ~n38204 ;
  assign n38229 = ~n38227 & ~n38228 ;
  assign n38226 = n38176 & n38225 ;
  assign n38231 = n38183 & n38230 ;
  assign n38232 = n38196 & ~n38231 ;
  assign n38233 = ~n38226 & n38232 ;
  assign n38234 = n38229 & n38233 ;
  assign n38237 = n38222 & n38236 ;
  assign n38238 = ~n38196 & ~n38209 ;
  assign n38239 = ~n38237 & n38238 ;
  assign n38240 = ~n38234 & ~n38239 ;
  assign n38254 = ~n38223 & ~n38240 ;
  assign n38255 = ~n38253 & n38254 ;
  assign n38256 = \u1_L7_reg[5]/NET0131  & ~n38255 ;
  assign n38257 = ~\u1_L7_reg[5]/NET0131  & n38255 ;
  assign n38258 = ~n38256 & ~n38257 ;
  assign n38265 = ~n37836 & ~n37838 ;
  assign n38266 = n37847 & n38265 ;
  assign n38263 = ~n37833 & ~n37838 ;
  assign n38264 = n37849 & ~n38263 ;
  assign n38270 = ~n37795 & ~n38264 ;
  assign n38271 = ~n38266 & n38270 ;
  assign n38259 = n37820 & n37839 ;
  assign n38260 = n37813 & n37831 ;
  assign n38261 = ~n38259 & ~n38260 ;
  assign n38262 = ~n37807 & ~n38261 ;
  assign n38267 = ~n37814 & ~n37854 ;
  assign n38268 = ~n37831 & n38267 ;
  assign n38269 = ~n37828 & ~n38268 ;
  assign n38272 = ~n38262 & ~n38269 ;
  assign n38273 = n38271 & n38272 ;
  assign n38274 = ~n37828 & n37851 ;
  assign n38280 = n37795 & ~n37853 ;
  assign n38281 = ~n37868 & n38280 ;
  assign n38282 = ~n38274 & n38281 ;
  assign n38275 = ~n37830 & ~n37871 ;
  assign n38276 = n37859 & ~n38275 ;
  assign n38277 = n37807 & n37820 ;
  assign n38278 = ~n37848 & ~n38277 ;
  assign n38279 = n37828 & ~n38278 ;
  assign n38283 = ~n38276 & ~n38279 ;
  assign n38284 = n38282 & n38283 ;
  assign n38285 = ~n38273 & ~n38284 ;
  assign n38286 = \u1_L7_reg[12]/NET0131  & n38285 ;
  assign n38287 = ~\u1_L7_reg[12]/NET0131  & ~n38285 ;
  assign n38288 = ~n38286 & ~n38287 ;
  assign n38293 = ~n38062 & ~n38082 ;
  assign n38294 = ~n38113 & n38293 ;
  assign n38297 = n38074 & n38122 ;
  assign n38295 = ~n38081 & ~n38088 ;
  assign n38296 = ~n38074 & n38295 ;
  assign n38298 = n38062 & ~n38296 ;
  assign n38299 = ~n38297 & n38298 ;
  assign n38300 = ~n38294 & ~n38299 ;
  assign n38291 = n38081 & n38128 ;
  assign n38292 = ~n38088 & n38291 ;
  assign n38301 = n38056 & n38107 ;
  assign n38302 = ~n38292 & n38301 ;
  assign n38303 = ~n38300 & n38302 ;
  assign n38307 = ~n38068 & ~n38102 ;
  assign n38308 = n38103 & n38307 ;
  assign n38304 = n38062 & n38068 ;
  assign n38305 = n38088 & ~n38099 ;
  assign n38306 = n38304 & n38305 ;
  assign n38309 = ~n38056 & ~n38306 ;
  assign n38310 = ~n38308 & n38309 ;
  assign n38313 = ~n38062 & ~n38291 ;
  assign n38311 = n38091 & n38112 ;
  assign n38312 = n38094 & n38295 ;
  assign n38314 = ~n38311 & ~n38312 ;
  assign n38315 = n38313 & n38314 ;
  assign n38316 = n38310 & n38315 ;
  assign n38317 = ~n38303 & ~n38316 ;
  assign n38289 = n38094 & n38105 ;
  assign n38290 = n38074 & n38115 ;
  assign n38318 = ~n38289 & ~n38290 ;
  assign n38319 = ~n38317 & n38318 ;
  assign n38322 = ~n38075 & ~n38128 ;
  assign n38323 = ~n38081 & ~n38322 ;
  assign n38320 = ~n38088 & n38094 ;
  assign n38321 = n38081 & n38320 ;
  assign n38324 = n38062 & ~n38321 ;
  assign n38325 = ~n38323 & n38324 ;
  assign n38326 = n38310 & n38325 ;
  assign n38327 = ~n38319 & ~n38326 ;
  assign n38328 = ~\u1_L7_reg[13]/NET0131  & ~n38327 ;
  assign n38329 = \u1_L7_reg[13]/NET0131  & n38327 ;
  assign n38330 = ~n38328 & ~n38329 ;
  assign n38331 = decrypt_pad & ~\u1_uk_K_r7_reg[51]/NET0131  ;
  assign n38332 = ~decrypt_pad & ~\u1_uk_K_r7_reg[44]/NET0131  ;
  assign n38333 = ~n38331 & ~n38332 ;
  assign n38334 = \u1_R7_reg[19]/NET0131  & ~n38333 ;
  assign n38335 = ~\u1_R7_reg[19]/NET0131  & n38333 ;
  assign n38336 = ~n38334 & ~n38335 ;
  assign n38337 = decrypt_pad & ~\u1_uk_K_r7_reg[9]/NET0131  ;
  assign n38338 = ~decrypt_pad & ~\u1_uk_K_r7_reg[2]/NET0131  ;
  assign n38339 = ~n38337 & ~n38338 ;
  assign n38340 = \u1_R7_reg[18]/NET0131  & ~n38339 ;
  assign n38341 = ~\u1_R7_reg[18]/NET0131  & n38339 ;
  assign n38342 = ~n38340 & ~n38341 ;
  assign n38343 = decrypt_pad & ~\u1_uk_K_r7_reg[15]/NET0131  ;
  assign n38344 = ~decrypt_pad & ~\u1_uk_K_r7_reg[8]/NET0131  ;
  assign n38345 = ~n38343 & ~n38344 ;
  assign n38346 = \u1_R7_reg[17]/NET0131  & ~n38345 ;
  assign n38347 = ~\u1_R7_reg[17]/NET0131  & n38345 ;
  assign n38348 = ~n38346 & ~n38347 ;
  assign n38349 = ~n38342 & n38348 ;
  assign n38350 = decrypt_pad & ~\u1_uk_K_r7_reg[36]/NET0131  ;
  assign n38351 = ~decrypt_pad & ~\u1_uk_K_r7_reg[29]/NET0131  ;
  assign n38352 = ~n38350 & ~n38351 ;
  assign n38353 = \u1_R7_reg[21]/NET0131  & ~n38352 ;
  assign n38354 = ~\u1_R7_reg[21]/NET0131  & n38352 ;
  assign n38355 = ~n38353 & ~n38354 ;
  assign n38356 = n38349 & n38355 ;
  assign n38357 = decrypt_pad & ~\u1_uk_K_r7_reg[52]/NET0131  ;
  assign n38358 = ~decrypt_pad & ~\u1_uk_K_r7_reg[45]/NET0131  ;
  assign n38359 = ~n38357 & ~n38358 ;
  assign n38360 = \u1_R7_reg[16]/NET0131  & ~n38359 ;
  assign n38361 = ~\u1_R7_reg[16]/NET0131  & n38359 ;
  assign n38362 = ~n38360 & ~n38361 ;
  assign n38363 = n38356 & n38362 ;
  assign n38369 = n38355 & ~n38362 ;
  assign n38370 = ~n38348 & n38369 ;
  assign n38364 = n38348 & ~n38355 ;
  assign n38365 = n38342 & n38364 ;
  assign n38366 = ~n38355 & n38362 ;
  assign n38367 = ~n38342 & ~n38348 ;
  assign n38368 = n38366 & n38367 ;
  assign n38371 = ~n38365 & ~n38368 ;
  assign n38372 = ~n38370 & n38371 ;
  assign n38373 = ~n38363 & n38372 ;
  assign n38374 = ~n38336 & ~n38373 ;
  assign n38382 = n38342 & n38355 ;
  assign n38383 = n38362 & n38382 ;
  assign n38378 = n38349 & ~n38362 ;
  assign n38380 = ~n38355 & ~n38362 ;
  assign n38381 = ~n38348 & n38380 ;
  assign n38384 = ~n38378 & ~n38381 ;
  assign n38385 = ~n38383 & n38384 ;
  assign n38386 = n38336 & ~n38385 ;
  assign n38375 = n38355 & n38362 ;
  assign n38376 = n38342 & ~n38348 ;
  assign n38377 = n38375 & n38376 ;
  assign n38379 = ~n38355 & n38378 ;
  assign n38387 = ~n38377 & ~n38379 ;
  assign n38388 = ~n38386 & n38387 ;
  assign n38389 = ~n38374 & n38388 ;
  assign n38390 = decrypt_pad & ~\u1_uk_K_r7_reg[35]/NET0131  ;
  assign n38391 = ~decrypt_pad & ~\u1_uk_K_r7_reg[28]/NET0131  ;
  assign n38392 = ~n38390 & ~n38391 ;
  assign n38393 = \u1_R7_reg[20]/NET0131  & ~n38392 ;
  assign n38394 = ~\u1_R7_reg[20]/NET0131  & n38392 ;
  assign n38395 = ~n38393 & ~n38394 ;
  assign n38396 = ~n38389 & ~n38395 ;
  assign n38399 = ~n38342 & n38375 ;
  assign n38402 = ~n38370 & ~n38399 ;
  assign n38400 = n38362 & n38364 ;
  assign n38401 = n38342 & n38369 ;
  assign n38403 = ~n38400 & ~n38401 ;
  assign n38404 = n38402 & n38403 ;
  assign n38405 = n38336 & ~n38404 ;
  assign n38406 = ~n38336 & ~n38342 ;
  assign n38407 = n38348 & n38369 ;
  assign n38408 = ~n38381 & ~n38407 ;
  assign n38409 = n38406 & ~n38408 ;
  assign n38397 = ~n38349 & ~n38376 ;
  assign n38398 = n38366 & ~n38397 ;
  assign n38410 = ~n38336 & n38348 ;
  assign n38411 = n38342 & ~n38410 ;
  assign n38412 = ~n38349 & n38375 ;
  assign n38413 = ~n38411 & n38412 ;
  assign n38414 = ~n38398 & ~n38413 ;
  assign n38415 = ~n38409 & n38414 ;
  assign n38416 = ~n38405 & n38415 ;
  assign n38417 = n38395 & ~n38416 ;
  assign n38418 = ~n38342 & n38400 ;
  assign n38419 = n38342 & n38381 ;
  assign n38420 = ~n38418 & ~n38419 ;
  assign n38421 = n38336 & ~n38420 ;
  assign n38422 = ~n38348 & n38401 ;
  assign n38423 = n38342 & ~n38362 ;
  assign n38424 = n38364 & n38423 ;
  assign n38425 = ~n38422 & ~n38424 ;
  assign n38426 = ~n38336 & ~n38425 ;
  assign n38427 = ~n38421 & ~n38426 ;
  assign n38428 = ~n38417 & n38427 ;
  assign n38429 = ~n38396 & n38428 ;
  assign n38430 = ~\u1_L7_reg[14]/NET0131  & ~n38429 ;
  assign n38431 = \u1_L7_reg[14]/NET0131  & n38429 ;
  assign n38432 = ~n38430 & ~n38431 ;
  assign n38433 = ~n38189 & ~n38241 ;
  assign n38434 = n38182 & ~n38433 ;
  assign n38435 = ~n38225 & ~n38434 ;
  assign n38436 = n38196 & ~n38435 ;
  assign n38437 = n38235 & n38241 ;
  assign n38438 = ~n38436 & ~n38437 ;
  assign n38439 = ~n38222 & ~n38438 ;
  assign n38453 = ~n38189 & n38204 ;
  assign n38454 = n38208 & n38453 ;
  assign n38455 = ~n38236 & ~n38454 ;
  assign n38456 = n38229 & n38455 ;
  assign n38457 = ~n38196 & ~n38456 ;
  assign n38446 = n38176 & ~n38196 ;
  assign n38447 = n38224 & n38446 ;
  assign n38440 = n38189 & n38208 ;
  assign n38441 = n38176 & ~n38182 ;
  assign n38442 = n38230 & n38441 ;
  assign n38448 = ~n38440 & ~n38442 ;
  assign n38449 = ~n38447 & n38448 ;
  assign n38443 = ~n38189 & ~n38204 ;
  assign n38444 = ~n38182 & n38443 ;
  assign n38445 = n38196 & n38444 ;
  assign n38450 = ~n38227 & ~n38445 ;
  assign n38451 = n38449 & n38450 ;
  assign n38452 = n38222 & ~n38451 ;
  assign n38458 = n38190 & n38204 ;
  assign n38459 = ~n38215 & ~n38458 ;
  assign n38460 = n38196 & ~n38459 ;
  assign n38461 = ~n38196 & ~n38222 ;
  assign n38462 = n38235 & n38461 ;
  assign n38463 = ~n38460 & ~n38462 ;
  assign n38464 = ~n38452 & n38463 ;
  assign n38465 = ~n38457 & n38464 ;
  assign n38466 = ~n38439 & n38465 ;
  assign n38467 = \u1_L7_reg[15]/P0001  & n38466 ;
  assign n38468 = ~\u1_L7_reg[15]/P0001  & ~n38466 ;
  assign n38469 = ~n38467 & ~n38468 ;
  assign n38473 = ~n37701 & ~n38148 ;
  assign n38474 = n37701 & n38158 ;
  assign n38470 = ~n37701 & ~n37730 ;
  assign n38471 = n37708 & ~n37767 ;
  assign n38472 = ~n38470 & n38471 ;
  assign n38475 = ~n37729 & ~n38472 ;
  assign n38476 = ~n38474 & n38475 ;
  assign n38477 = ~n38473 & n38476 ;
  assign n38482 = ~n37708 & n38141 ;
  assign n38481 = ~n37701 & n37755 ;
  assign n38478 = ~n37695 & n37758 ;
  assign n38483 = n37729 & ~n38478 ;
  assign n38484 = ~n38481 & n38483 ;
  assign n38485 = ~n38482 & n38484 ;
  assign n38479 = ~n37753 & ~n37768 ;
  assign n38480 = n37701 & ~n38479 ;
  assign n38486 = ~n38033 & ~n38480 ;
  assign n38487 = n38485 & n38486 ;
  assign n38488 = ~n38477 & ~n38487 ;
  assign n38489 = ~n37742 & ~n37779 ;
  assign n38490 = ~n38488 & n38489 ;
  assign n38491 = ~\u1_L7_reg[19]/P0001  & ~n38490 ;
  assign n38492 = \u1_L7_reg[19]/P0001  & n38490 ;
  assign n38493 = ~n38491 & ~n38492 ;
  assign n38510 = ~n37949 & ~n37977 ;
  assign n38511 = n37932 & ~n38510 ;
  assign n38512 = ~n37920 & ~n38511 ;
  assign n38513 = ~n37950 & n37955 ;
  assign n38514 = ~n38512 & ~n38513 ;
  assign n38515 = n37946 & ~n37981 ;
  assign n38516 = ~n37996 & ~n38515 ;
  assign n38517 = ~n38514 & n38516 ;
  assign n38518 = ~n37976 & ~n38517 ;
  assign n38499 = ~n37966 & ~n37977 ;
  assign n38500 = n37920 & ~n38499 ;
  assign n38495 = n37933 & n37945 ;
  assign n38496 = n37946 & ~n37952 ;
  assign n38497 = ~n38495 & ~n38496 ;
  assign n38498 = ~n37920 & ~n38497 ;
  assign n38494 = ~n37932 & n37953 ;
  assign n38501 = n37945 & n37978 ;
  assign n38502 = ~n38494 & ~n38501 ;
  assign n38503 = ~n38498 & n38502 ;
  assign n38504 = ~n38500 & n38503 ;
  assign n38505 = n37976 & ~n38504 ;
  assign n38507 = ~n37984 & n37995 ;
  assign n38508 = ~n37963 & ~n38507 ;
  assign n38509 = n37920 & ~n38508 ;
  assign n38506 = ~n37920 & n38501 ;
  assign n38519 = ~n37994 & ~n38506 ;
  assign n38520 = ~n38509 & n38519 ;
  assign n38521 = ~n38505 & n38520 ;
  assign n38522 = ~n38518 & n38521 ;
  assign n38523 = ~\u1_L7_reg[1]/NET0131  & ~n38522 ;
  assign n38524 = \u1_L7_reg[1]/NET0131  & n38522 ;
  assign n38525 = ~n38523 & ~n38524 ;
  assign n38526 = ~n38190 & n38196 ;
  assign n38527 = n38198 & ~n38224 ;
  assign n38528 = ~n38441 & ~n38443 ;
  assign n38529 = ~n38527 & n38528 ;
  assign n38530 = n38526 & ~n38529 ;
  assign n38531 = ~n38196 & ~n38442 ;
  assign n38532 = ~n38527 & n38531 ;
  assign n38533 = ~n38530 & ~n38532 ;
  assign n38534 = n38189 & n38205 ;
  assign n38535 = ~n38444 & ~n38534 ;
  assign n38536 = n38176 & ~n38535 ;
  assign n38537 = n38222 & ~n38458 ;
  assign n38538 = ~n38536 & n38537 ;
  assign n38539 = ~n38533 & n38538 ;
  assign n38544 = ~n38189 & n38205 ;
  assign n38545 = ~n38196 & ~n38544 ;
  assign n38546 = ~n38236 & ~n38534 ;
  assign n38547 = n38526 & n38546 ;
  assign n38548 = ~n38545 & ~n38547 ;
  assign n38540 = n38446 & n38453 ;
  assign n38549 = ~n38214 & ~n38222 ;
  assign n38550 = ~n38540 & n38549 ;
  assign n38541 = ~n38182 & n38196 ;
  assign n38542 = n38198 & n38204 ;
  assign n38543 = ~n38541 & n38542 ;
  assign n38551 = ~n38228 & ~n38247 ;
  assign n38552 = ~n38543 & n38551 ;
  assign n38553 = n38550 & n38552 ;
  assign n38554 = ~n38548 & n38553 ;
  assign n38555 = ~n38539 & ~n38554 ;
  assign n38556 = ~\u1_L7_reg[21]/NET0131  & n38555 ;
  assign n38557 = \u1_L7_reg[21]/NET0131  & ~n38555 ;
  assign n38558 = ~n38556 & ~n38557 ;
  assign n38561 = n37625 & n37633 ;
  assign n38564 = n37616 & ~n38561 ;
  assign n38565 = n37668 & n37888 ;
  assign n38566 = ~n37883 & ~n38565 ;
  assign n38559 = n37609 & n37897 ;
  assign n38567 = n37678 & ~n38559 ;
  assign n38568 = n38566 & n38567 ;
  assign n38569 = ~n38564 & ~n38568 ;
  assign n38570 = ~n37652 & ~n37657 ;
  assign n38571 = ~n37893 & n38570 ;
  assign n38572 = ~n37624 & n38571 ;
  assign n38573 = ~n38569 & n38572 ;
  assign n38574 = ~n37603 & n37903 ;
  assign n38575 = n37639 & n37673 ;
  assign n38576 = ~n37616 & ~n38575 ;
  assign n38577 = ~n38574 & n38576 ;
  assign n38578 = n38566 & n38577 ;
  assign n38579 = n37623 & n37885 ;
  assign n38580 = n37616 & ~n37641 ;
  assign n38581 = ~n38579 & n38580 ;
  assign n38582 = ~n38578 & ~n38581 ;
  assign n38583 = ~n37637 & n37652 ;
  assign n38584 = ~n37676 & n38583 ;
  assign n38585 = ~n38582 & n38584 ;
  assign n38586 = ~n38573 & ~n38585 ;
  assign n38560 = n37655 & n38559 ;
  assign n38562 = ~n37673 & ~n38561 ;
  assign n38563 = n37674 & ~n38562 ;
  assign n38587 = ~n38560 & ~n38563 ;
  assign n38588 = ~n38586 & n38587 ;
  assign n38589 = \u1_L7_reg[23]/NET0131  & ~n38588 ;
  assign n38590 = ~\u1_L7_reg[23]/NET0131  & n38588 ;
  assign n38591 = ~n38589 & ~n38590 ;
  assign n38600 = ~n38336 & ~n38348 ;
  assign n38602 = ~n38362 & n38600 ;
  assign n38603 = n38336 & n38364 ;
  assign n38604 = ~n38602 & ~n38603 ;
  assign n38605 = ~n38342 & ~n38604 ;
  assign n38606 = n38336 & ~n38355 ;
  assign n38607 = n38348 & n38423 ;
  assign n38608 = ~n38606 & n38607 ;
  assign n38601 = n38366 & n38600 ;
  assign n38609 = ~n38395 & ~n38601 ;
  assign n38610 = ~n38608 & n38609 ;
  assign n38611 = ~n38605 & n38610 ;
  assign n38612 = ~n38348 & n38375 ;
  assign n38613 = ~n38336 & ~n38612 ;
  assign n38614 = ~n38378 & n38613 ;
  assign n38617 = ~n38367 & ~n38423 ;
  assign n38618 = ~n38355 & ~n38617 ;
  assign n38615 = n38348 & n38375 ;
  assign n38616 = ~n38348 & ~n38362 ;
  assign n38619 = n38336 & ~n38616 ;
  assign n38620 = ~n38615 & n38619 ;
  assign n38621 = ~n38618 & n38620 ;
  assign n38622 = ~n38614 & ~n38621 ;
  assign n38595 = n38362 & n38365 ;
  assign n38623 = ~n38356 & n38395 ;
  assign n38624 = ~n38595 & n38623 ;
  assign n38625 = ~n38622 & n38624 ;
  assign n38626 = ~n38611 & ~n38625 ;
  assign n38592 = ~n38336 & n38376 ;
  assign n38593 = ~n38356 & ~n38592 ;
  assign n38594 = n38362 & ~n38593 ;
  assign n38596 = ~n38419 & ~n38595 ;
  assign n38597 = n38367 & n38369 ;
  assign n38598 = n38596 & ~n38597 ;
  assign n38599 = n38336 & ~n38598 ;
  assign n38627 = ~n38594 & ~n38599 ;
  assign n38628 = ~n38626 & n38627 ;
  assign n38629 = ~\u1_L7_reg[25]/NET0131  & ~n38628 ;
  assign n38630 = \u1_L7_reg[25]/NET0131  & n38628 ;
  assign n38631 = ~n38629 & ~n38630 ;
  assign n38632 = n37920 & ~n37967 ;
  assign n38633 = ~n37947 & n38632 ;
  assign n38635 = ~n37926 & ~n37945 ;
  assign n38636 = ~n38494 & ~n38635 ;
  assign n38637 = ~n37976 & ~n38636 ;
  assign n38634 = n37946 & n37981 ;
  assign n38638 = n37932 & ~n37939 ;
  assign n38639 = n38635 & n38638 ;
  assign n38640 = ~n37920 & ~n38639 ;
  assign n38641 = ~n38634 & n38640 ;
  assign n38642 = ~n38637 & n38641 ;
  assign n38643 = ~n38633 & ~n38642 ;
  assign n38648 = ~n37932 & ~n37965 ;
  assign n38649 = ~n37920 & n37926 ;
  assign n38650 = ~n38638 & n38649 ;
  assign n38651 = ~n38648 & n38650 ;
  assign n38646 = n37920 & n37992 ;
  assign n38647 = ~n37939 & n37962 ;
  assign n38653 = ~n38646 & ~n38647 ;
  assign n38654 = ~n38651 & n38653 ;
  assign n38644 = ~n38000 & ~n38495 ;
  assign n38645 = n37939 & ~n38644 ;
  assign n38652 = n37976 & ~n38501 ;
  assign n38655 = ~n38645 & n38652 ;
  assign n38656 = n38654 & n38655 ;
  assign n38657 = ~n37933 & n37969 ;
  assign n38658 = ~n37966 & ~n37976 ;
  assign n38659 = n37999 & n38658 ;
  assign n38660 = ~n38657 & n38659 ;
  assign n38661 = ~n38656 & ~n38660 ;
  assign n38662 = ~n38643 & ~n38661 ;
  assign n38663 = ~\u1_L7_reg[26]/NET0131  & ~n38662 ;
  assign n38664 = \u1_L7_reg[26]/NET0131  & n38662 ;
  assign n38665 = ~n38663 & ~n38664 ;
  assign n38684 = n38088 & n38291 ;
  assign n38685 = n38120 & ~n38684 ;
  assign n38686 = n38062 & ~n38685 ;
  assign n38669 = ~n38088 & n38128 ;
  assign n38670 = n38081 & n38091 ;
  assign n38671 = ~n38669 & ~n38670 ;
  assign n38683 = ~n38062 & ~n38671 ;
  assign n38681 = ~n38082 & ~n38304 ;
  assign n38682 = ~n38088 & ~n38681 ;
  assign n38687 = ~n38311 & ~n38682 ;
  assign n38688 = ~n38683 & n38687 ;
  assign n38689 = ~n38686 & n38688 ;
  assign n38690 = n38056 & ~n38689 ;
  assign n38666 = ~n38081 & n38122 ;
  assign n38667 = ~n38289 & ~n38666 ;
  assign n38668 = ~n38062 & ~n38667 ;
  assign n38672 = n38062 & n38671 ;
  assign n38673 = ~n38062 & ~n38093 ;
  assign n38674 = ~n38092 & n38673 ;
  assign n38675 = ~n38320 & n38674 ;
  assign n38676 = ~n38672 & ~n38675 ;
  assign n38677 = n38112 & ~n38322 ;
  assign n38678 = ~n38289 & ~n38677 ;
  assign n38679 = ~n38676 & n38678 ;
  assign n38680 = ~n38056 & ~n38679 ;
  assign n38691 = ~n38668 & ~n38680 ;
  assign n38692 = ~n38690 & n38691 ;
  assign n38693 = ~\u1_L7_reg[28]/NET0131  & ~n38692 ;
  assign n38694 = \u1_L7_reg[28]/NET0131  & n38692 ;
  assign n38695 = ~n38693 & ~n38694 ;
  assign n38697 = n38367 & n38380 ;
  assign n38698 = ~n38612 & ~n38697 ;
  assign n38699 = n38336 & ~n38698 ;
  assign n38696 = n38362 & n38406 ;
  assign n38700 = n38395 & ~n38696 ;
  assign n38701 = n38425 & n38700 ;
  assign n38702 = ~n38699 & n38701 ;
  assign n38703 = n38369 & ~n38376 ;
  assign n38704 = n38613 & ~n38703 ;
  assign n38705 = n38336 & ~n38368 ;
  assign n38706 = ~n38615 & n38705 ;
  assign n38707 = ~n38704 & ~n38706 ;
  assign n38708 = ~n38378 & ~n38395 ;
  assign n38709 = n38596 & n38708 ;
  assign n38710 = ~n38707 & n38709 ;
  assign n38711 = ~n38702 & ~n38710 ;
  assign n38712 = n38369 & ~n38397 ;
  assign n38713 = ~n38365 & ~n38712 ;
  assign n38714 = n38336 & ~n38713 ;
  assign n38715 = n38366 & n38592 ;
  assign n38716 = ~n38714 & ~n38715 ;
  assign n38717 = ~n38711 & n38716 ;
  assign n38718 = ~\u1_L7_reg[8]/NET0131  & ~n38717 ;
  assign n38719 = \u1_L7_reg[8]/NET0131  & n38717 ;
  assign n38720 = ~n38718 & ~n38719 ;
  assign n38721 = ~n38207 & n38434 ;
  assign n38722 = n38196 & ~n38721 ;
  assign n38723 = n38182 & ~n38230 ;
  assign n38724 = ~n38443 & n38723 ;
  assign n38725 = n38197 & ~n38724 ;
  assign n38726 = ~n38722 & ~n38725 ;
  assign n38727 = n38183 & n38204 ;
  assign n38728 = ~n38215 & ~n38727 ;
  assign n38729 = ~n38247 & n38728 ;
  assign n38730 = ~n38726 & n38729 ;
  assign n38731 = n38222 & ~n38730 ;
  assign n38739 = n38196 & ~n38214 ;
  assign n38737 = ~n38204 & n38208 ;
  assign n38738 = n38204 & ~n38208 ;
  assign n38740 = ~n38737 & ~n38738 ;
  assign n38741 = n38739 & n38740 ;
  assign n38742 = n38230 & n38446 ;
  assign n38743 = ~n38226 & ~n38742 ;
  assign n38744 = ~n38741 & n38743 ;
  assign n38745 = ~n38222 & ~n38744 ;
  assign n38732 = ~n38222 & n38544 ;
  assign n38733 = ~n38209 & ~n38231 ;
  assign n38734 = ~n38227 & n38733 ;
  assign n38735 = ~n38732 & n38734 ;
  assign n38736 = ~n38196 & ~n38735 ;
  assign n38746 = n38196 & ~n38204 ;
  assign n38747 = n38441 & n38746 ;
  assign n38748 = ~n38736 & ~n38747 ;
  assign n38749 = ~n38745 & n38748 ;
  assign n38750 = ~n38731 & n38749 ;
  assign n38751 = ~\u1_L7_reg[27]/NET0131  & ~n38750 ;
  assign n38752 = \u1_L7_reg[27]/NET0131  & n38750 ;
  assign n38753 = ~n38751 & ~n38752 ;
  assign n38759 = ~n37849 & ~n37870 ;
  assign n38761 = ~n37836 & n38267 ;
  assign n38762 = n38759 & ~n38761 ;
  assign n38760 = ~n37836 & ~n38759 ;
  assign n38763 = ~n37828 & ~n38760 ;
  assign n38764 = ~n38762 & n38763 ;
  assign n38754 = n37838 & n37870 ;
  assign n38755 = n37801 & ~n37870 ;
  assign n38756 = n37859 & ~n38755 ;
  assign n38757 = ~n37821 & ~n38756 ;
  assign n38758 = n37828 & ~n38757 ;
  assign n38765 = ~n38754 & ~n38758 ;
  assign n38766 = ~n38764 & n38765 ;
  assign n38767 = n37795 & ~n38766 ;
  assign n38769 = ~n38259 & ~n38267 ;
  assign n38770 = ~n37828 & ~n38769 ;
  assign n38771 = ~n37807 & n37852 ;
  assign n38772 = n37828 & ~n38259 ;
  assign n38773 = ~n38771 & n38772 ;
  assign n38774 = ~n38770 & ~n38773 ;
  assign n38768 = n37807 & ~n38261 ;
  assign n38775 = n37869 & ~n38768 ;
  assign n38776 = ~n38774 & n38775 ;
  assign n38777 = ~n37795 & ~n38776 ;
  assign n38778 = n37828 & n37851 ;
  assign n38779 = ~n37839 & n37866 ;
  assign n38780 = n37832 & n38779 ;
  assign n38781 = ~n38778 & ~n38780 ;
  assign n38782 = ~n38777 & n38781 ;
  assign n38783 = ~n38767 & n38782 ;
  assign n38784 = \u1_L7_reg[32]/NET0131  & n38783 ;
  assign n38785 = ~\u1_L7_reg[32]/NET0131  & ~n38783 ;
  assign n38786 = ~n38784 & ~n38785 ;
  assign n38788 = n38366 & n38376 ;
  assign n38787 = n38369 & n38410 ;
  assign n38789 = n38395 & ~n38787 ;
  assign n38790 = ~n38788 & n38789 ;
  assign n38791 = ~n38363 & n38790 ;
  assign n38792 = ~n38362 & n38364 ;
  assign n38793 = ~n38399 & ~n38792 ;
  assign n38794 = n38791 & n38793 ;
  assign n38795 = ~n38366 & n38376 ;
  assign n38796 = ~n38395 & ~n38795 ;
  assign n38797 = ~n38342 & n38369 ;
  assign n38798 = ~n38400 & ~n38797 ;
  assign n38799 = n38796 & n38798 ;
  assign n38800 = ~n38794 & ~n38799 ;
  assign n38801 = ~n38422 & n38705 ;
  assign n38802 = ~n38800 & n38801 ;
  assign n38803 = ~n38380 & ~n38382 ;
  assign n38804 = ~n38612 & n38803 ;
  assign n38805 = n38796 & n38804 ;
  assign n38806 = ~n38791 & ~n38805 ;
  assign n38807 = ~n38336 & ~n38377 ;
  assign n38808 = ~n38697 & n38807 ;
  assign n38809 = ~n38418 & n38808 ;
  assign n38810 = ~n38806 & n38809 ;
  assign n38811 = ~n38802 & ~n38810 ;
  assign n38812 = ~\u1_L7_reg[3]/NET0131  & n38811 ;
  assign n38813 = \u1_L7_reg[3]/NET0131  & ~n38811 ;
  assign n38814 = ~n38812 & ~n38813 ;
  assign n38849 = decrypt_pad & ~\u1_uk_K_r7_reg[18]/NET0131  ;
  assign n38850 = ~decrypt_pad & ~\u1_uk_K_r7_reg[11]/NET0131  ;
  assign n38851 = ~n38849 & ~n38850 ;
  assign n38852 = \u1_R7_reg[11]/NET0131  & ~n38851 ;
  assign n38853 = ~\u1_R7_reg[11]/NET0131  & n38851 ;
  assign n38854 = ~n38852 & ~n38853 ;
  assign n38841 = decrypt_pad & ~\u1_uk_K_r7_reg[33]/NET0131  ;
  assign n38842 = ~decrypt_pad & ~\u1_uk_K_r7_reg[26]/P0001  ;
  assign n38843 = ~n38841 & ~n38842 ;
  assign n38844 = \u1_R7_reg[12]/NET0131  & ~n38843 ;
  assign n38845 = ~\u1_R7_reg[12]/NET0131  & n38843 ;
  assign n38846 = ~n38844 & ~n38845 ;
  assign n38815 = decrypt_pad & ~\u1_uk_K_r7_reg[46]/NET0131  ;
  assign n38816 = ~decrypt_pad & ~\u1_uk_K_r7_reg[39]/NET0131  ;
  assign n38817 = ~n38815 & ~n38816 ;
  assign n38818 = \u1_R7_reg[13]/NET0131  & ~n38817 ;
  assign n38819 = ~\u1_R7_reg[13]/NET0131  & n38817 ;
  assign n38820 = ~n38818 & ~n38819 ;
  assign n38828 = decrypt_pad & ~\u1_uk_K_r7_reg[41]/NET0131  ;
  assign n38829 = ~decrypt_pad & ~\u1_uk_K_r7_reg[34]/NET0131  ;
  assign n38830 = ~n38828 & ~n38829 ;
  assign n38831 = \u1_R7_reg[9]/NET0131  & ~n38830 ;
  assign n38832 = ~\u1_R7_reg[9]/NET0131  & n38830 ;
  assign n38833 = ~n38831 & ~n38832 ;
  assign n38855 = n38820 & ~n38833 ;
  assign n38834 = decrypt_pad & ~\u1_uk_K_r7_reg[17]/NET0131  ;
  assign n38835 = ~decrypt_pad & ~\u1_uk_K_r7_reg[10]/NET0131  ;
  assign n38836 = ~n38834 & ~n38835 ;
  assign n38837 = \u1_R7_reg[10]/NET0131  & ~n38836 ;
  assign n38838 = ~\u1_R7_reg[10]/NET0131  & n38836 ;
  assign n38839 = ~n38837 & ~n38838 ;
  assign n38821 = decrypt_pad & ~\u1_uk_K_r7_reg[12]/NET0131  ;
  assign n38822 = ~decrypt_pad & ~\u1_uk_K_r7_reg[5]/NET0131  ;
  assign n38823 = ~n38821 & ~n38822 ;
  assign n38824 = \u1_R7_reg[8]/NET0131  & ~n38823 ;
  assign n38825 = ~\u1_R7_reg[8]/NET0131  & n38823 ;
  assign n38826 = ~n38824 & ~n38825 ;
  assign n38857 = n38820 & ~n38826 ;
  assign n38858 = n38839 & n38857 ;
  assign n38859 = ~n38820 & n38833 ;
  assign n38860 = n38826 & n38859 ;
  assign n38861 = ~n38858 & ~n38860 ;
  assign n38862 = ~n38855 & n38861 ;
  assign n38863 = n38846 & ~n38862 ;
  assign n38856 = n38839 & n38855 ;
  assign n38864 = ~n38826 & ~n38833 ;
  assign n38865 = ~n38820 & n38864 ;
  assign n38866 = ~n38839 & n38865 ;
  assign n38867 = ~n38856 & ~n38866 ;
  assign n38868 = ~n38863 & n38867 ;
  assign n38869 = n38854 & ~n38868 ;
  assign n38840 = n38833 & n38839 ;
  assign n38878 = ~n38833 & ~n38839 ;
  assign n38879 = ~n38840 & ~n38878 ;
  assign n38827 = ~n38820 & ~n38826 ;
  assign n38876 = n38820 & n38826 ;
  assign n38877 = ~n38827 & ~n38876 ;
  assign n38880 = n38820 & n38854 ;
  assign n38884 = n38877 & ~n38880 ;
  assign n38885 = ~n38879 & ~n38884 ;
  assign n38881 = n38833 & n38880 ;
  assign n38882 = n38877 & n38879 ;
  assign n38883 = ~n38881 & n38882 ;
  assign n38886 = ~n38846 & ~n38883 ;
  assign n38887 = ~n38885 & n38886 ;
  assign n38847 = n38840 & n38846 ;
  assign n38848 = n38827 & n38847 ;
  assign n38870 = n38833 & ~n38839 ;
  assign n38871 = ~n38826 & ~n38870 ;
  assign n38872 = n38846 & ~n38854 ;
  assign n38873 = ~n38855 & n38872 ;
  assign n38874 = ~n38859 & n38873 ;
  assign n38875 = ~n38871 & n38874 ;
  assign n38888 = ~n38848 & ~n38875 ;
  assign n38889 = ~n38887 & n38888 ;
  assign n38890 = ~n38869 & n38889 ;
  assign n38891 = ~\u1_L7_reg[6]/NET0131  & ~n38890 ;
  assign n38892 = \u1_L7_reg[6]/NET0131  & n38890 ;
  assign n38893 = ~n38891 & ~n38892 ;
  assign n38911 = ~n37820 & ~n38265 ;
  assign n38894 = n37807 & ~n38759 ;
  assign n38912 = n37801 & n37870 ;
  assign n38913 = ~n38894 & ~n38912 ;
  assign n38914 = ~n38911 & n38913 ;
  assign n38915 = ~n37828 & ~n38914 ;
  assign n38895 = ~n38771 & ~n38894 ;
  assign n38896 = n37801 & ~n38895 ;
  assign n38905 = ~n37801 & ~n37814 ;
  assign n38906 = n38759 & n38905 ;
  assign n38916 = n37828 & n38906 ;
  assign n38917 = ~n38896 & ~n38916 ;
  assign n38918 = ~n38915 & n38917 ;
  assign n38919 = n37795 & ~n38918 ;
  assign n38897 = ~n37828 & n38896 ;
  assign n38898 = n37795 & ~n37828 ;
  assign n38899 = n37858 & ~n38759 ;
  assign n38900 = n37813 & ~n38277 ;
  assign n38901 = n37828 & n38755 ;
  assign n38902 = ~n38900 & n38901 ;
  assign n38903 = ~n38899 & ~n38902 ;
  assign n38904 = ~n37795 & ~n38903 ;
  assign n38907 = ~n37828 & n38906 ;
  assign n38908 = ~n37822 & ~n38907 ;
  assign n38909 = ~n38904 & n38908 ;
  assign n38910 = ~n38898 & ~n38909 ;
  assign n38920 = ~n38897 & ~n38910 ;
  assign n38921 = ~n38919 & n38920 ;
  assign n38922 = ~\u1_L7_reg[7]/NET0131  & ~n38921 ;
  assign n38923 = \u1_L7_reg[7]/NET0131  & n38921 ;
  assign n38924 = ~n38922 & ~n38923 ;
  assign n38927 = ~n37882 & n37903 ;
  assign n38928 = ~n37678 & ~n38927 ;
  assign n38929 = ~n37616 & n37903 ;
  assign n38930 = ~n38928 & ~n38929 ;
  assign n38925 = ~n37643 & ~n37899 ;
  assign n38926 = ~n37888 & ~n38925 ;
  assign n38931 = ~n37652 & ~n38926 ;
  assign n38932 = ~n38930 & n38931 ;
  assign n38935 = ~n37904 & ~n38574 ;
  assign n38936 = n37609 & ~n38935 ;
  assign n38933 = ~n37640 & n37674 ;
  assign n38934 = ~n37903 & n38933 ;
  assign n38937 = n37884 & ~n38934 ;
  assign n38938 = ~n38936 & n38937 ;
  assign n38939 = ~n38932 & ~n38938 ;
  assign n38940 = ~n37616 & n37892 ;
  assign n38941 = ~n37677 & n38940 ;
  assign n38942 = ~n38939 & ~n38941 ;
  assign n38943 = ~\u1_L7_reg[9]/NET0131  & ~n38942 ;
  assign n38944 = \u1_L7_reg[9]/NET0131  & n38942 ;
  assign n38945 = ~n38943 & ~n38944 ;
  assign n38959 = ~n38833 & ~n38876 ;
  assign n38947 = n38833 & n38876 ;
  assign n38960 = ~n38827 & ~n38947 ;
  assign n38961 = ~n38959 & n38960 ;
  assign n38971 = ~n38846 & n38961 ;
  assign n38969 = ~n38860 & ~n38865 ;
  assign n38970 = n38839 & ~n38969 ;
  assign n38972 = n38854 & ~n38970 ;
  assign n38973 = ~n38971 & n38972 ;
  assign n38948 = n38827 & ~n38839 ;
  assign n38946 = ~n38833 & n38857 ;
  assign n38949 = ~n38946 & ~n38947 ;
  assign n38950 = ~n38948 & n38949 ;
  assign n38951 = ~n38846 & ~n38950 ;
  assign n38974 = n38826 & n38839 ;
  assign n38975 = ~n38833 & n38974 ;
  assign n38976 = ~n38854 & ~n38975 ;
  assign n38977 = ~n38951 & n38976 ;
  assign n38978 = ~n38973 & ~n38977 ;
  assign n38952 = n38866 & n38951 ;
  assign n38962 = n38833 & n38854 ;
  assign n38963 = n38827 & ~n38962 ;
  assign n38964 = ~n38839 & ~n38963 ;
  assign n38965 = ~n38961 & n38964 ;
  assign n38953 = n38827 & n38839 ;
  assign n38954 = ~n38820 & n38826 ;
  assign n38955 = ~n38839 & n38954 ;
  assign n38956 = ~n38953 & ~n38955 ;
  assign n38957 = ~n38854 & ~n38956 ;
  assign n38958 = n38833 & n38858 ;
  assign n38966 = ~n38957 & ~n38958 ;
  assign n38967 = ~n38965 & n38966 ;
  assign n38968 = n38846 & ~n38967 ;
  assign n38979 = ~n38952 & ~n38968 ;
  assign n38980 = ~n38978 & n38979 ;
  assign n38981 = ~\u1_L7_reg[16]/NET0131  & ~n38980 ;
  assign n38982 = \u1_L7_reg[16]/NET0131  & n38980 ;
  assign n38983 = ~n38981 & ~n38982 ;
  assign n38985 = n38068 & n38103 ;
  assign n38986 = ~n38118 & ~n38985 ;
  assign n38987 = ~n38062 & ~n38986 ;
  assign n38984 = n38062 & ~n38100 ;
  assign n38988 = n38056 & ~n38114 ;
  assign n38989 = ~n38984 & n38988 ;
  assign n38990 = ~n38987 & n38989 ;
  assign n38992 = ~n38062 & n38105 ;
  assign n38993 = ~n38295 & ~n38992 ;
  assign n38994 = ~n38068 & ~n38993 ;
  assign n38995 = ~n38056 & ~n38289 ;
  assign n38996 = ~n38296 & n38995 ;
  assign n38991 = n38062 & n38119 ;
  assign n38997 = ~n38089 & ~n38991 ;
  assign n38998 = n38996 & n38997 ;
  assign n38999 = ~n38994 & n38998 ;
  assign n39000 = ~n38990 & ~n38999 ;
  assign n39001 = ~n38062 & n38670 ;
  assign n39002 = n38075 & n38088 ;
  assign n39003 = ~n38292 & ~n39002 ;
  assign n39004 = n38062 & ~n39003 ;
  assign n39005 = ~n39001 & ~n39004 ;
  assign n39006 = ~n39000 & n39005 ;
  assign n39007 = \u1_L7_reg[18]/NET0131  & n39006 ;
  assign n39008 = ~\u1_L7_reg[18]/NET0131  & ~n39006 ;
  assign n39009 = ~n39007 & ~n39008 ;
  assign n39010 = ~n38820 & n38975 ;
  assign n39011 = ~n38839 & n38857 ;
  assign n39012 = ~n38953 & ~n39011 ;
  assign n39013 = n38827 & n38833 ;
  assign n39014 = ~n38975 & ~n39013 ;
  assign n39015 = n39012 & n39014 ;
  assign n39016 = n38854 & ~n39015 ;
  assign n39017 = ~n39010 & ~n39016 ;
  assign n39018 = ~n38846 & ~n39017 ;
  assign n39027 = n38878 & n38884 ;
  assign n39029 = ~n38878 & ~n38954 ;
  assign n39030 = ~n38854 & ~n39029 ;
  assign n39028 = n38854 & ~n38878 ;
  assign n39031 = ~n38857 & ~n39028 ;
  assign n39032 = ~n39030 & n39031 ;
  assign n39033 = ~n39027 & ~n39032 ;
  assign n39034 = n38846 & ~n39033 ;
  assign n39019 = n38826 & n38840 ;
  assign n39020 = ~n38858 & ~n39019 ;
  assign n39021 = n38846 & ~n39020 ;
  assign n39022 = ~n38859 & ~n38864 ;
  assign n39023 = ~n38839 & ~n38876 ;
  assign n39024 = n39022 & n39023 ;
  assign n39025 = ~n39021 & ~n39024 ;
  assign n39026 = n38854 & ~n39025 ;
  assign n39035 = n38839 & ~n38854 ;
  assign n39036 = n38947 & n39035 ;
  assign n39037 = ~n38877 & n38878 ;
  assign n39038 = n38861 & ~n39037 ;
  assign n39039 = ~n38846 & ~n38854 ;
  assign n39040 = ~n39038 & n39039 ;
  assign n39041 = ~n39036 & ~n39040 ;
  assign n39042 = ~n39026 & n39041 ;
  assign n39043 = ~n39034 & n39042 ;
  assign n39044 = ~n39018 & n39043 ;
  assign n39045 = ~\u1_L7_reg[24]/NET0131  & ~n39044 ;
  assign n39046 = \u1_L7_reg[24]/NET0131  & n39044 ;
  assign n39047 = ~n39045 & ~n39046 ;
  assign n39048 = n38878 & n38954 ;
  assign n39049 = n38854 & ~n39048 ;
  assign n39050 = n39012 & n39049 ;
  assign n39051 = ~n38854 & ~n38974 ;
  assign n39052 = ~n39013 & n39051 ;
  assign n39053 = ~n39050 & ~n39052 ;
  assign n39054 = n38846 & ~n39053 ;
  assign n39056 = ~n38974 & n39022 ;
  assign n39057 = ~n38854 & ~n39056 ;
  assign n39059 = ~n38859 & n38974 ;
  assign n39058 = ~n38820 & n38870 ;
  assign n39060 = n38854 & ~n39058 ;
  assign n39061 = ~n39059 & n39060 ;
  assign n39062 = ~n39057 & ~n39061 ;
  assign n39055 = n38839 & n38946 ;
  assign n39063 = ~n38846 & ~n39037 ;
  assign n39064 = ~n39055 & n39063 ;
  assign n39065 = ~n39062 & n39064 ;
  assign n39066 = ~n39054 & ~n39065 ;
  assign n39068 = n38880 & n38975 ;
  assign n39067 = n38847 & ~n38876 ;
  assign n39069 = n38859 & n39035 ;
  assign n39070 = ~n39067 & ~n39069 ;
  assign n39071 = ~n39068 & n39070 ;
  assign n39072 = ~n39066 & n39071 ;
  assign n39073 = \u1_L7_reg[30]/NET0131  & ~n39072 ;
  assign n39074 = ~\u1_L7_reg[30]/NET0131  & n39072 ;
  assign n39075 = ~n39073 & ~n39074 ;
  assign n39076 = decrypt_pad & ~\u1_uk_K_r6_reg[23]/P0001  ;
  assign n39077 = ~decrypt_pad & ~\u1_uk_K_r6_reg[30]/P0001  ;
  assign n39078 = ~n39076 & ~n39077 ;
  assign n39079 = \u1_R6_reg[28]/NET0131  & ~n39078 ;
  assign n39080 = ~\u1_R6_reg[28]/NET0131  & n39078 ;
  assign n39081 = ~n39079 & ~n39080 ;
  assign n39082 = decrypt_pad & ~\u1_uk_K_r6_reg[31]/NET0131  ;
  assign n39083 = ~decrypt_pad & ~\u1_uk_K_r6_reg[38]/NET0131  ;
  assign n39084 = ~n39082 & ~n39083 ;
  assign n39085 = \u1_R6_reg[26]/NET0131  & ~n39084 ;
  assign n39086 = ~\u1_R6_reg[26]/NET0131  & n39084 ;
  assign n39087 = ~n39085 & ~n39086 ;
  assign n39088 = decrypt_pad & ~\u1_uk_K_r6_reg[42]/NET0131  ;
  assign n39089 = ~decrypt_pad & ~\u1_uk_K_r6_reg[49]/NET0131  ;
  assign n39090 = ~n39088 & ~n39089 ;
  assign n39091 = \u1_R6_reg[25]/NET0131  & ~n39090 ;
  assign n39092 = ~\u1_R6_reg[25]/NET0131  & n39090 ;
  assign n39093 = ~n39091 & ~n39092 ;
  assign n39122 = ~n39087 & ~n39093 ;
  assign n39094 = decrypt_pad & ~\u1_uk_K_r6_reg[15]/NET0131  ;
  assign n39095 = ~decrypt_pad & ~\u1_uk_K_r6_reg[22]/NET0131  ;
  assign n39096 = ~n39094 & ~n39095 ;
  assign n39097 = \u1_R6_reg[29]/NET0131  & ~n39096 ;
  assign n39098 = ~\u1_R6_reg[29]/NET0131  & n39096 ;
  assign n39099 = ~n39097 & ~n39098 ;
  assign n39125 = ~n39087 & ~n39099 ;
  assign n39145 = ~n39122 & ~n39125 ;
  assign n39101 = decrypt_pad & ~\u1_uk_K_r6_reg[7]/NET0131  ;
  assign n39102 = ~decrypt_pad & ~\u1_uk_K_r6_reg[14]/NET0131  ;
  assign n39103 = ~n39101 & ~n39102 ;
  assign n39104 = \u1_R6_reg[24]/NET0131  & ~n39103 ;
  assign n39105 = ~\u1_R6_reg[24]/NET0131  & n39103 ;
  assign n39106 = ~n39104 & ~n39105 ;
  assign n39109 = decrypt_pad & ~\u1_uk_K_r6_reg[36]/NET0131  ;
  assign n39110 = ~decrypt_pad & ~\u1_uk_K_r6_reg[43]/NET0131  ;
  assign n39111 = ~n39109 & ~n39110 ;
  assign n39112 = \u1_R6_reg[27]/NET0131  & ~n39111 ;
  assign n39113 = ~\u1_R6_reg[27]/NET0131  & n39111 ;
  assign n39114 = ~n39112 & ~n39113 ;
  assign n39124 = n39087 & n39093 ;
  assign n39144 = n39114 & ~n39124 ;
  assign n39146 = n39106 & n39144 ;
  assign n39147 = n39145 & n39146 ;
  assign n39138 = n39099 & n39106 ;
  assign n39139 = n39122 & n39138 ;
  assign n39140 = n39093 & n39099 ;
  assign n39141 = ~n39106 & n39140 ;
  assign n39142 = ~n39139 & ~n39141 ;
  assign n39143 = ~n39114 & ~n39142 ;
  assign n39133 = ~n39099 & ~n39106 ;
  assign n39134 = n39122 & n39133 ;
  assign n39135 = n39099 & ~n39106 ;
  assign n39136 = n39087 & ~n39093 ;
  assign n39137 = n39135 & n39136 ;
  assign n39148 = ~n39134 & ~n39137 ;
  assign n39149 = ~n39143 & n39148 ;
  assign n39150 = ~n39147 & n39149 ;
  assign n39151 = n39081 & ~n39150 ;
  assign n39126 = ~n39114 & ~n39124 ;
  assign n39127 = ~n39125 & n39126 ;
  assign n39123 = n39114 & ~n39122 ;
  assign n39128 = n39106 & ~n39123 ;
  assign n39129 = ~n39127 & n39128 ;
  assign n39100 = ~n39093 & ~n39099 ;
  assign n39107 = n39100 & ~n39106 ;
  assign n39108 = n39087 & n39107 ;
  assign n39115 = n39108 & ~n39114 ;
  assign n39116 = ~n39087 & ~n39106 ;
  assign n39117 = n39087 & n39106 ;
  assign n39118 = ~n39116 & ~n39117 ;
  assign n39119 = ~n39093 & n39114 ;
  assign n39120 = n39099 & ~n39119 ;
  assign n39121 = ~n39118 & n39120 ;
  assign n39130 = ~n39115 & ~n39121 ;
  assign n39131 = ~n39129 & n39130 ;
  assign n39132 = ~n39081 & ~n39131 ;
  assign n39154 = n39124 & n39133 ;
  assign n39155 = ~n39137 & ~n39154 ;
  assign n39156 = ~n39099 & n39106 ;
  assign n39157 = ~n39093 & n39156 ;
  assign n39158 = n39155 & ~n39157 ;
  assign n39159 = n39114 & ~n39158 ;
  assign n39152 = n39093 & ~n39114 ;
  assign n39153 = ~n39118 & n39152 ;
  assign n39160 = n39119 & n39125 ;
  assign n39161 = ~n39153 & ~n39160 ;
  assign n39162 = ~n39159 & n39161 ;
  assign n39163 = ~n39132 & n39162 ;
  assign n39164 = ~n39151 & n39163 ;
  assign n39165 = ~\u1_L6_reg[22]/NET0131  & ~n39164 ;
  assign n39166 = \u1_L6_reg[22]/NET0131  & n39164 ;
  assign n39167 = ~n39165 & ~n39166 ;
  assign n39205 = decrypt_pad & ~\u1_uk_K_r6_reg[12]/NET0131  ;
  assign n39206 = ~decrypt_pad & ~\u1_uk_K_r6_reg[19]/NET0131  ;
  assign n39207 = ~n39205 & ~n39206 ;
  assign n39208 = \u1_R6_reg[3]/NET0131  & ~n39207 ;
  assign n39209 = ~\u1_R6_reg[3]/NET0131  & n39207 ;
  assign n39210 = ~n39208 & ~n39209 ;
  assign n39168 = decrypt_pad & ~\u1_uk_K_r6_reg[47]/NET0131  ;
  assign n39169 = ~decrypt_pad & ~\u1_uk_K_r6_reg[54]/NET0131  ;
  assign n39170 = ~n39168 & ~n39169 ;
  assign n39171 = \u1_R6_reg[4]/NET0131  & ~n39170 ;
  assign n39172 = ~\u1_R6_reg[4]/NET0131  & n39170 ;
  assign n39173 = ~n39171 & ~n39172 ;
  assign n39187 = decrypt_pad & ~\u1_uk_K_r6_reg[3]/NET0131  ;
  assign n39188 = ~decrypt_pad & ~\u1_uk_K_r6_reg[10]/NET0131  ;
  assign n39189 = ~n39187 & ~n39188 ;
  assign n39190 = \u1_R6_reg[2]/NET0131  & ~n39189 ;
  assign n39191 = ~\u1_R6_reg[2]/NET0131  & n39189 ;
  assign n39192 = ~n39190 & ~n39191 ;
  assign n39174 = decrypt_pad & ~\u1_uk_K_r6_reg[20]/NET0131  ;
  assign n39175 = ~decrypt_pad & ~\u1_uk_K_r6_reg[27]/NET0131  ;
  assign n39176 = ~n39174 & ~n39175 ;
  assign n39177 = \u1_R6_reg[1]/NET0131  & ~n39176 ;
  assign n39178 = ~\u1_R6_reg[1]/NET0131  & n39176 ;
  assign n39179 = ~n39177 & ~n39178 ;
  assign n39180 = decrypt_pad & ~\u1_uk_K_r6_reg[18]/NET0131  ;
  assign n39181 = ~decrypt_pad & ~\u1_uk_K_r6_reg[25]/NET0131  ;
  assign n39182 = ~n39180 & ~n39181 ;
  assign n39183 = \u1_R6_reg[5]/NET0131  & ~n39182 ;
  assign n39184 = ~\u1_R6_reg[5]/NET0131  & n39182 ;
  assign n39185 = ~n39183 & ~n39184 ;
  assign n39186 = ~n39179 & ~n39185 ;
  assign n39194 = decrypt_pad & ~\u1_uk_K_r6_reg[24]/NET0131  ;
  assign n39195 = ~decrypt_pad & ~\u1_uk_K_r6_reg[6]/NET0131  ;
  assign n39196 = ~n39194 & ~n39195 ;
  assign n39197 = \u1_R6_reg[32]/NET0131  & ~n39196 ;
  assign n39198 = ~\u1_R6_reg[32]/NET0131  & n39196 ;
  assign n39199 = ~n39197 & ~n39198 ;
  assign n39243 = n39186 & n39199 ;
  assign n39244 = n39192 & n39243 ;
  assign n39201 = ~n39179 & n39185 ;
  assign n39245 = ~n39192 & ~n39199 ;
  assign n39246 = ~n39201 & n39245 ;
  assign n39247 = ~n39244 & ~n39246 ;
  assign n39248 = ~n39173 & ~n39247 ;
  assign n39230 = n39185 & n39199 ;
  assign n39241 = n39179 & n39230 ;
  assign n39242 = n39192 & n39241 ;
  assign n39202 = n39192 & ~n39199 ;
  assign n39249 = n39201 & n39202 ;
  assign n39228 = n39179 & ~n39185 ;
  assign n39250 = ~n39192 & n39228 ;
  assign n39251 = ~n39249 & ~n39250 ;
  assign n39252 = ~n39242 & n39251 ;
  assign n39253 = ~n39248 & n39252 ;
  assign n39254 = ~n39210 & ~n39253 ;
  assign n39203 = ~n39185 & n39202 ;
  assign n39204 = ~n39201 & ~n39203 ;
  assign n39211 = ~n39204 & n39210 ;
  assign n39216 = ~n39192 & n39210 ;
  assign n39217 = n39179 & ~n39216 ;
  assign n39218 = n39185 & ~n39199 ;
  assign n39219 = ~n39217 & n39218 ;
  assign n39193 = n39186 & ~n39192 ;
  assign n39200 = n39193 & n39199 ;
  assign n39212 = n39179 & ~n39199 ;
  assign n39213 = n39179 & ~n39210 ;
  assign n39214 = ~n39202 & ~n39213 ;
  assign n39215 = ~n39212 & ~n39214 ;
  assign n39220 = ~n39200 & ~n39215 ;
  assign n39221 = ~n39219 & n39220 ;
  assign n39222 = ~n39211 & n39221 ;
  assign n39223 = n39173 & ~n39222 ;
  assign n39234 = ~n39185 & ~n39199 ;
  assign n39235 = ~n39230 & ~n39234 ;
  assign n39236 = n39179 & n39235 ;
  assign n39237 = n39210 & n39236 ;
  assign n39238 = n39192 & ~n39237 ;
  assign n39231 = ~n39213 & n39230 ;
  assign n39229 = ~n39199 & n39228 ;
  assign n39232 = ~n39192 & ~n39229 ;
  assign n39233 = ~n39231 & n39232 ;
  assign n39239 = ~n39173 & ~n39233 ;
  assign n39240 = ~n39238 & n39239 ;
  assign n39224 = ~n39179 & n39210 ;
  assign n39225 = n39203 & n39224 ;
  assign n39226 = ~n39192 & n39199 ;
  assign n39227 = n39224 & n39226 ;
  assign n39255 = ~n39225 & ~n39227 ;
  assign n39256 = ~n39240 & n39255 ;
  assign n39257 = ~n39223 & n39256 ;
  assign n39258 = ~n39254 & n39257 ;
  assign n39259 = ~\u1_L6_reg[31]/NET0131  & ~n39258 ;
  assign n39260 = \u1_L6_reg[31]/NET0131  & n39258 ;
  assign n39261 = ~n39259 & ~n39260 ;
  assign n39316 = decrypt_pad & ~\u1_uk_K_r6_reg[16]/NET0131  ;
  assign n39317 = ~decrypt_pad & ~\u1_uk_K_r6_reg[23]/P0001  ;
  assign n39318 = ~n39316 & ~n39317 ;
  assign n39319 = \u1_R6_reg[24]/NET0131  & ~n39318 ;
  assign n39320 = ~\u1_R6_reg[24]/NET0131  & n39318 ;
  assign n39321 = ~n39319 & ~n39320 ;
  assign n39285 = decrypt_pad & ~\u1_uk_K_r6_reg[14]/NET0131  ;
  assign n39286 = ~decrypt_pad & ~\u1_uk_K_r6_reg[21]/NET0131  ;
  assign n39287 = ~n39285 & ~n39286 ;
  assign n39288 = \u1_R6_reg[23]/NET0131  & ~n39287 ;
  assign n39289 = ~\u1_R6_reg[23]/NET0131  & n39287 ;
  assign n39290 = ~n39288 & ~n39289 ;
  assign n39262 = decrypt_pad & ~\u1_uk_K_r6_reg[38]/NET0131  ;
  assign n39263 = ~decrypt_pad & ~\u1_uk_K_r6_reg[45]/NET0131  ;
  assign n39264 = ~n39262 & ~n39263 ;
  assign n39265 = \u1_R6_reg[21]/NET0131  & ~n39264 ;
  assign n39266 = ~\u1_R6_reg[21]/NET0131  & n39264 ;
  assign n39267 = ~n39265 & ~n39266 ;
  assign n39268 = decrypt_pad & ~\u1_uk_K_r6_reg[50]/NET0131  ;
  assign n39269 = ~decrypt_pad & ~\u1_uk_K_r6_reg[2]/NET0131  ;
  assign n39270 = ~n39268 & ~n39269 ;
  assign n39271 = \u1_R6_reg[20]/NET0131  & ~n39270 ;
  assign n39272 = ~\u1_R6_reg[20]/NET0131  & n39270 ;
  assign n39273 = ~n39271 & ~n39272 ;
  assign n39274 = n39267 & ~n39273 ;
  assign n39275 = decrypt_pad & ~\u1_uk_K_r6_reg[1]/NET0131  ;
  assign n39276 = ~decrypt_pad & ~\u1_uk_K_r6_reg[8]/NET0131  ;
  assign n39277 = ~n39275 & ~n39276 ;
  assign n39278 = \u1_R6_reg[22]/NET0131  & ~n39277 ;
  assign n39279 = ~\u1_R6_reg[22]/NET0131  & n39277 ;
  assign n39280 = ~n39278 & ~n39279 ;
  assign n39281 = n39274 & n39280 ;
  assign n39293 = decrypt_pad & ~\u1_uk_K_r6_reg[35]/NET0131  ;
  assign n39294 = ~decrypt_pad & ~\u1_uk_K_r6_reg[42]/NET0131  ;
  assign n39295 = ~n39293 & ~n39294 ;
  assign n39296 = \u1_R6_reg[25]/NET0131  & ~n39295 ;
  assign n39297 = ~\u1_R6_reg[25]/NET0131  & n39295 ;
  assign n39298 = ~n39296 & ~n39297 ;
  assign n39341 = n39267 & ~n39298 ;
  assign n39342 = n39273 & ~n39341 ;
  assign n39299 = ~n39280 & ~n39298 ;
  assign n39343 = ~n39267 & ~n39299 ;
  assign n39344 = n39342 & ~n39343 ;
  assign n39345 = ~n39281 & ~n39344 ;
  assign n39346 = n39290 & ~n39345 ;
  assign n39304 = n39273 & n39298 ;
  assign n39337 = ~n39274 & ~n39304 ;
  assign n39338 = n39280 & ~n39337 ;
  assign n39309 = ~n39273 & n39298 ;
  assign n39335 = n39267 & n39309 ;
  assign n39336 = ~n39280 & ~n39335 ;
  assign n39339 = ~n39290 & ~n39336 ;
  assign n39340 = ~n39338 & n39339 ;
  assign n39331 = ~n39280 & ~n39290 ;
  assign n39347 = n39304 & n39331 ;
  assign n39348 = ~n39267 & n39347 ;
  assign n39349 = ~n39340 & ~n39348 ;
  assign n39350 = ~n39346 & n39349 ;
  assign n39351 = n39321 & ~n39350 ;
  assign n39282 = n39267 & n39273 ;
  assign n39283 = ~n39280 & n39282 ;
  assign n39284 = ~n39281 & ~n39283 ;
  assign n39291 = ~n39284 & ~n39290 ;
  assign n39300 = ~n39267 & n39290 ;
  assign n39310 = n39300 & n39309 ;
  assign n39307 = n39282 & n39299 ;
  assign n39292 = ~n39280 & n39290 ;
  assign n39308 = ~n39273 & n39292 ;
  assign n39311 = ~n39307 & ~n39308 ;
  assign n39312 = ~n39310 & n39311 ;
  assign n39301 = ~n39299 & ~n39300 ;
  assign n39302 = n39273 & ~n39292 ;
  assign n39303 = ~n39301 & n39302 ;
  assign n39305 = n39280 & n39304 ;
  assign n39306 = ~n39267 & n39305 ;
  assign n39313 = ~n39303 & ~n39306 ;
  assign n39314 = n39312 & n39313 ;
  assign n39315 = ~n39291 & n39314 ;
  assign n39322 = ~n39315 & ~n39321 ;
  assign n39327 = n39282 & ~n39298 ;
  assign n39328 = ~n39290 & n39327 ;
  assign n39329 = ~n39310 & ~n39328 ;
  assign n39330 = ~n39280 & ~n39329 ;
  assign n39323 = n39274 & ~n39298 ;
  assign n39324 = ~n39280 & n39323 ;
  assign n39325 = ~n39305 & ~n39324 ;
  assign n39326 = n39290 & ~n39325 ;
  assign n39332 = ~n39273 & ~n39298 ;
  assign n39333 = n39331 & n39332 ;
  assign n39334 = ~n39267 & n39333 ;
  assign n39352 = ~n39326 & ~n39334 ;
  assign n39353 = ~n39330 & n39352 ;
  assign n39354 = ~n39322 & n39353 ;
  assign n39355 = ~n39351 & n39354 ;
  assign n39356 = \u1_L6_reg[11]/NET0131  & ~n39355 ;
  assign n39357 = ~\u1_L6_reg[11]/NET0131  & n39355 ;
  assign n39358 = ~n39356 & ~n39357 ;
  assign n39372 = decrypt_pad & ~\u1_uk_K_r6_reg[32]/NET0131  ;
  assign n39373 = ~decrypt_pad & ~\u1_uk_K_r6_reg[39]/NET0131  ;
  assign n39374 = ~n39372 & ~n39373 ;
  assign n39375 = \u1_R6_reg[13]/NET0131  & ~n39374 ;
  assign n39376 = ~\u1_R6_reg[13]/NET0131  & n39374 ;
  assign n39377 = ~n39375 & ~n39376 ;
  assign n39378 = decrypt_pad & ~\u1_uk_K_r6_reg[41]/NET0131  ;
  assign n39379 = ~decrypt_pad & ~\u1_uk_K_r6_reg[48]/NET0131  ;
  assign n39380 = ~n39378 & ~n39379 ;
  assign n39381 = \u1_R6_reg[15]/NET0131  & ~n39380 ;
  assign n39382 = ~\u1_R6_reg[15]/NET0131  & n39380 ;
  assign n39383 = ~n39381 & ~n39382 ;
  assign n39384 = n39377 & n39383 ;
  assign n39359 = decrypt_pad & ~\u1_uk_K_r6_reg[13]/NET0131  ;
  assign n39360 = ~decrypt_pad & ~\u1_uk_K_r6_reg[20]/NET0131  ;
  assign n39361 = ~n39359 & ~n39360 ;
  assign n39362 = \u1_R6_reg[12]/NET0131  & ~n39361 ;
  assign n39363 = ~\u1_R6_reg[12]/NET0131  & n39361 ;
  assign n39364 = ~n39362 & ~n39363 ;
  assign n39386 = decrypt_pad & ~\u1_uk_K_r6_reg[33]/NET0131  ;
  assign n39387 = ~decrypt_pad & ~\u1_uk_K_r6_reg[40]/NET0131  ;
  assign n39388 = ~n39386 & ~n39387 ;
  assign n39389 = \u1_R6_reg[14]/NET0131  & ~n39388 ;
  assign n39390 = ~\u1_R6_reg[14]/NET0131  & n39388 ;
  assign n39391 = ~n39389 & ~n39390 ;
  assign n39406 = ~n39364 & n39391 ;
  assign n39407 = n39384 & n39406 ;
  assign n39408 = decrypt_pad & ~\u1_uk_K_r6_reg[17]/NET0131  ;
  assign n39409 = ~decrypt_pad & ~\u1_uk_K_r6_reg[24]/NET0131  ;
  assign n39410 = ~n39408 & ~n39409 ;
  assign n39411 = \u1_R6_reg[16]/NET0131  & ~n39410 ;
  assign n39412 = ~\u1_R6_reg[16]/NET0131  & n39410 ;
  assign n39413 = ~n39411 & ~n39412 ;
  assign n39423 = ~n39407 & ~n39413 ;
  assign n39365 = decrypt_pad & ~\u1_uk_K_r6_reg[54]/NET0131  ;
  assign n39366 = ~decrypt_pad & ~\u1_uk_K_r6_reg[4]/NET0131  ;
  assign n39367 = ~n39365 & ~n39366 ;
  assign n39368 = \u1_R6_reg[17]/NET0131  & ~n39367 ;
  assign n39369 = ~\u1_R6_reg[17]/NET0131  & n39367 ;
  assign n39370 = ~n39368 & ~n39369 ;
  assign n39421 = n39364 & n39370 ;
  assign n39422 = n39384 & n39421 ;
  assign n39394 = n39370 & ~n39391 ;
  assign n39414 = n39364 & ~n39377 ;
  assign n39415 = n39394 & n39414 ;
  assign n39397 = ~n39377 & n39383 ;
  assign n39398 = ~n39364 & ~n39370 ;
  assign n39416 = n39397 & n39398 ;
  assign n39424 = ~n39415 & ~n39416 ;
  assign n39425 = ~n39422 & n39424 ;
  assign n39426 = n39423 & n39425 ;
  assign n39371 = n39364 & ~n39370 ;
  assign n39400 = n39371 & n39391 ;
  assign n39403 = n39370 & ~n39377 ;
  assign n39404 = ~n39400 & ~n39403 ;
  assign n39405 = ~n39383 & ~n39404 ;
  assign n39399 = ~n39391 & n39398 ;
  assign n39417 = ~n39377 & n39399 ;
  assign n39393 = ~n39364 & n39377 ;
  assign n39418 = ~n39370 & n39391 ;
  assign n39419 = n39393 & n39418 ;
  assign n39420 = ~n39417 & ~n39419 ;
  assign n39427 = ~n39405 & n39420 ;
  assign n39428 = n39426 & n39427 ;
  assign n39436 = n39377 & n39421 ;
  assign n39437 = ~n39377 & ~n39383 ;
  assign n39438 = n39398 & n39437 ;
  assign n39439 = ~n39436 & ~n39438 ;
  assign n39440 = n39391 & ~n39439 ;
  assign n39433 = ~n39393 & ~n39414 ;
  assign n39434 = ~n39383 & ~n39391 ;
  assign n39435 = ~n39433 & n39434 ;
  assign n39385 = n39371 & n39384 ;
  assign n39429 = n39393 & n39394 ;
  assign n39430 = ~n39385 & ~n39429 ;
  assign n39431 = ~n39364 & n39370 ;
  assign n39432 = n39397 & n39431 ;
  assign n39441 = n39413 & ~n39432 ;
  assign n39442 = n39430 & n39441 ;
  assign n39443 = ~n39435 & n39442 ;
  assign n39444 = ~n39440 & n39443 ;
  assign n39445 = ~n39428 & ~n39444 ;
  assign n39401 = ~n39399 & ~n39400 ;
  assign n39402 = n39397 & ~n39401 ;
  assign n39392 = n39385 & ~n39391 ;
  assign n39395 = ~n39383 & n39394 ;
  assign n39396 = n39393 & n39395 ;
  assign n39446 = ~n39392 & ~n39396 ;
  assign n39447 = ~n39402 & n39446 ;
  assign n39448 = ~n39445 & n39447 ;
  assign n39449 = ~\u1_L6_reg[20]/NET0131  & ~n39448 ;
  assign n39450 = \u1_L6_reg[20]/NET0131  & n39448 ;
  assign n39451 = ~n39449 & ~n39450 ;
  assign n39452 = decrypt_pad & ~\u1_uk_K_r6_reg[21]/NET0131  ;
  assign n39453 = ~decrypt_pad & ~\u1_uk_K_r6_reg[28]/NET0131  ;
  assign n39454 = ~n39452 & ~n39453 ;
  assign n39455 = \u1_R6_reg[28]/NET0131  & ~n39454 ;
  assign n39456 = ~\u1_R6_reg[28]/NET0131  & n39454 ;
  assign n39457 = ~n39455 & ~n39456 ;
  assign n39458 = decrypt_pad & ~\u1_uk_K_r6_reg[9]/NET0131  ;
  assign n39459 = ~decrypt_pad & ~\u1_uk_K_r6_reg[16]/NET0131  ;
  assign n39460 = ~n39458 & ~n39459 ;
  assign n39461 = \u1_R6_reg[1]/NET0131  & ~n39460 ;
  assign n39462 = ~\u1_R6_reg[1]/NET0131  & n39460 ;
  assign n39463 = ~n39461 & ~n39462 ;
  assign n39465 = decrypt_pad & ~\u1_uk_K_r6_reg[52]/NET0131  ;
  assign n39466 = ~decrypt_pad & ~\u1_uk_K_r6_reg[0]/NET0131  ;
  assign n39467 = ~n39465 & ~n39466 ;
  assign n39468 = \u1_R6_reg[29]/NET0131  & ~n39467 ;
  assign n39469 = ~\u1_R6_reg[29]/NET0131  & n39467 ;
  assign n39470 = ~n39468 & ~n39469 ;
  assign n39473 = decrypt_pad & ~\u1_uk_K_r6_reg[49]/NET0131  ;
  assign n39474 = ~decrypt_pad & ~\u1_uk_K_r6_reg[1]/NET0131  ;
  assign n39475 = ~n39473 & ~n39474 ;
  assign n39476 = \u1_R6_reg[30]/NET0131  & ~n39475 ;
  assign n39477 = ~\u1_R6_reg[30]/NET0131  & n39475 ;
  assign n39478 = ~n39476 & ~n39477 ;
  assign n39497 = n39470 & n39478 ;
  assign n39498 = n39463 & n39497 ;
  assign n39495 = n39470 & ~n39478 ;
  assign n39496 = ~n39463 & n39495 ;
  assign n39482 = decrypt_pad & ~\u1_uk_K_r6_reg[37]/NET0131  ;
  assign n39483 = ~decrypt_pad & ~\u1_uk_K_r6_reg[44]/NET0131  ;
  assign n39484 = ~n39482 & ~n39483 ;
  assign n39485 = \u1_R6_reg[31]/P0001  & ~n39484 ;
  assign n39486 = ~\u1_R6_reg[31]/P0001  & n39484 ;
  assign n39487 = ~n39485 & ~n39486 ;
  assign n39499 = ~n39478 & ~n39487 ;
  assign n39500 = ~n39496 & ~n39499 ;
  assign n39501 = ~n39498 & n39500 ;
  assign n39502 = n39457 & ~n39501 ;
  assign n39464 = ~n39457 & n39463 ;
  assign n39471 = n39464 & ~n39470 ;
  assign n39472 = n39457 & ~n39470 ;
  assign n39479 = ~n39463 & n39478 ;
  assign n39480 = n39472 & n39479 ;
  assign n39481 = ~n39471 & ~n39480 ;
  assign n39488 = ~n39481 & n39487 ;
  assign n39489 = n39457 & ~n39463 ;
  assign n39490 = ~n39487 & ~n39489 ;
  assign n39491 = n39463 & ~n39470 ;
  assign n39492 = ~n39463 & ~n39478 ;
  assign n39493 = ~n39491 & ~n39492 ;
  assign n39494 = n39490 & n39493 ;
  assign n39503 = decrypt_pad & ~\u1_uk_K_r6_reg[43]/NET0131  ;
  assign n39504 = ~decrypt_pad & ~\u1_uk_K_r6_reg[50]/NET0131  ;
  assign n39505 = ~n39503 & ~n39504 ;
  assign n39506 = \u1_R6_reg[32]/NET0131  & ~n39505 ;
  assign n39507 = ~\u1_R6_reg[32]/NET0131  & n39505 ;
  assign n39508 = ~n39506 & ~n39507 ;
  assign n39509 = ~n39494 & ~n39508 ;
  assign n39510 = ~n39488 & n39509 ;
  assign n39511 = ~n39502 & n39510 ;
  assign n39522 = n39457 & n39470 ;
  assign n39523 = ~n39463 & n39522 ;
  assign n39524 = ~n39478 & n39523 ;
  assign n39519 = ~n39463 & n39470 ;
  assign n39520 = n39457 & ~n39478 ;
  assign n39521 = ~n39519 & ~n39520 ;
  assign n39525 = n39487 & ~n39521 ;
  assign n39526 = ~n39524 & n39525 ;
  assign n39514 = n39472 & n39478 ;
  assign n39515 = ~n39470 & ~n39478 ;
  assign n39516 = ~n39457 & n39515 ;
  assign n39517 = ~n39514 & ~n39516 ;
  assign n39518 = ~n39487 & ~n39517 ;
  assign n39512 = ~n39457 & n39497 ;
  assign n39513 = n39463 & n39512 ;
  assign n39527 = n39508 & ~n39513 ;
  assign n39528 = ~n39518 & n39527 ;
  assign n39529 = ~n39526 & n39528 ;
  assign n39530 = ~n39511 & ~n39529 ;
  assign n39531 = ~n39487 & n39524 ;
  assign n39535 = ~n39463 & n39516 ;
  assign n39532 = ~n39489 & ~n39495 ;
  assign n39533 = ~n39521 & n39532 ;
  assign n39534 = n39471 & n39478 ;
  assign n39536 = ~n39533 & ~n39534 ;
  assign n39537 = ~n39535 & n39536 ;
  assign n39538 = n39487 & ~n39537 ;
  assign n39539 = ~n39531 & ~n39538 ;
  assign n39540 = ~n39530 & n39539 ;
  assign n39541 = \u1_L6_reg[5]/NET0131  & ~n39540 ;
  assign n39542 = ~\u1_L6_reg[5]/NET0131  & n39540 ;
  assign n39543 = ~n39541 & ~n39542 ;
  assign n39559 = n39391 & n39433 ;
  assign n39560 = n39370 & n39559 ;
  assign n39556 = n39377 & n39398 ;
  assign n39557 = ~n39415 & ~n39556 ;
  assign n39558 = n39383 & ~n39557 ;
  assign n39546 = n39377 & ~n39391 ;
  assign n39561 = ~n39383 & ~n39546 ;
  assign n39562 = n39371 & n39561 ;
  assign n39563 = ~n39396 & ~n39562 ;
  assign n39564 = ~n39558 & n39563 ;
  assign n39565 = ~n39560 & n39564 ;
  assign n39566 = n39413 & ~n39565 ;
  assign n39549 = n39383 & n39394 ;
  assign n39550 = ~n39364 & n39549 ;
  assign n39544 = n39364 & ~n39394 ;
  assign n39545 = n39397 & n39544 ;
  assign n39551 = ~n39438 & ~n39545 ;
  assign n39552 = ~n39550 & n39551 ;
  assign n39547 = ~n39395 & ~n39546 ;
  assign n39548 = n39364 & ~n39547 ;
  assign n39553 = n39420 & ~n39548 ;
  assign n39554 = n39552 & n39553 ;
  assign n39555 = ~n39413 & ~n39554 ;
  assign n39567 = ~n39417 & ~n39560 ;
  assign n39568 = ~n39383 & ~n39567 ;
  assign n39569 = ~n39392 & ~n39407 ;
  assign n39570 = ~n39568 & n39569 ;
  assign n39571 = ~n39555 & n39570 ;
  assign n39572 = ~n39566 & n39571 ;
  assign n39573 = ~\u1_L6_reg[10]/NET0131  & ~n39572 ;
  assign n39574 = \u1_L6_reg[10]/NET0131  & n39572 ;
  assign n39575 = ~n39573 & ~n39574 ;
  assign n39582 = ~n39122 & ~n39124 ;
  assign n39583 = n39133 & n39582 ;
  assign n39580 = ~n39119 & ~n39124 ;
  assign n39581 = n39135 & ~n39580 ;
  assign n39587 = ~n39081 & ~n39581 ;
  assign n39588 = ~n39583 & n39587 ;
  assign n39576 = n39106 & n39125 ;
  assign n39577 = n39099 & n39117 ;
  assign n39578 = ~n39576 & ~n39577 ;
  assign n39579 = ~n39093 & ~n39578 ;
  assign n39584 = ~n39100 & ~n39140 ;
  assign n39585 = ~n39117 & n39584 ;
  assign n39586 = ~n39114 & ~n39585 ;
  assign n39589 = ~n39579 & ~n39586 ;
  assign n39590 = n39588 & n39589 ;
  assign n39591 = ~n39114 & n39137 ;
  assign n39597 = n39081 & ~n39139 ;
  assign n39598 = ~n39154 & n39597 ;
  assign n39599 = ~n39591 & n39598 ;
  assign n39592 = ~n39116 & ~n39157 ;
  assign n39593 = n39145 & ~n39592 ;
  assign n39594 = n39093 & n39106 ;
  assign n39595 = ~n39134 & ~n39594 ;
  assign n39596 = n39114 & ~n39595 ;
  assign n39600 = ~n39593 & ~n39596 ;
  assign n39601 = n39599 & n39600 ;
  assign n39602 = ~n39590 & ~n39601 ;
  assign n39603 = \u1_L6_reg[12]/NET0131  & n39602 ;
  assign n39604 = ~\u1_L6_reg[12]/NET0131  & ~n39602 ;
  assign n39605 = ~n39603 & ~n39604 ;
  assign n39642 = decrypt_pad & ~\u1_uk_K_r6_reg[28]/NET0131  ;
  assign n39643 = ~decrypt_pad & ~\u1_uk_K_r6_reg[35]/NET0131  ;
  assign n39644 = ~n39642 & ~n39643 ;
  assign n39645 = \u1_R6_reg[20]/NET0131  & ~n39644 ;
  assign n39646 = ~\u1_R6_reg[20]/NET0131  & n39644 ;
  assign n39647 = ~n39645 & ~n39646 ;
  assign n39606 = decrypt_pad & ~\u1_uk_K_r6_reg[8]/NET0131  ;
  assign n39607 = ~decrypt_pad & ~\u1_uk_K_r6_reg[15]/NET0131  ;
  assign n39608 = ~n39606 & ~n39607 ;
  assign n39609 = \u1_R6_reg[17]/NET0131  & ~n39608 ;
  assign n39610 = ~\u1_R6_reg[17]/NET0131  & n39608 ;
  assign n39611 = ~n39609 & ~n39610 ;
  assign n39612 = decrypt_pad & ~\u1_uk_K_r6_reg[29]/NET0131  ;
  assign n39613 = ~decrypt_pad & ~\u1_uk_K_r6_reg[36]/NET0131  ;
  assign n39614 = ~n39612 & ~n39613 ;
  assign n39615 = \u1_R6_reg[21]/NET0131  & ~n39614 ;
  assign n39616 = ~\u1_R6_reg[21]/NET0131  & n39614 ;
  assign n39617 = ~n39615 & ~n39616 ;
  assign n39618 = ~n39611 & ~n39617 ;
  assign n39619 = n39611 & n39617 ;
  assign n39620 = ~n39618 & ~n39619 ;
  assign n39621 = decrypt_pad & ~\u1_uk_K_r6_reg[2]/NET0131  ;
  assign n39622 = ~decrypt_pad & ~\u1_uk_K_r6_reg[9]/NET0131  ;
  assign n39623 = ~n39621 & ~n39622 ;
  assign n39624 = \u1_R6_reg[18]/NET0131  & ~n39623 ;
  assign n39625 = ~\u1_R6_reg[18]/NET0131  & n39623 ;
  assign n39626 = ~n39624 & ~n39625 ;
  assign n39627 = decrypt_pad & ~\u1_uk_K_r6_reg[45]/NET0131  ;
  assign n39628 = ~decrypt_pad & ~\u1_uk_K_r6_reg[52]/NET0131  ;
  assign n39629 = ~n39627 & ~n39628 ;
  assign n39630 = \u1_R6_reg[16]/NET0131  & ~n39629 ;
  assign n39631 = ~\u1_R6_reg[16]/NET0131  & n39629 ;
  assign n39632 = ~n39630 & ~n39631 ;
  assign n39652 = ~n39626 & n39632 ;
  assign n39653 = ~n39620 & n39652 ;
  assign n39635 = decrypt_pad & ~\u1_uk_K_r6_reg[44]/NET0131  ;
  assign n39636 = ~decrypt_pad & ~\u1_uk_K_r6_reg[51]/NET0131  ;
  assign n39637 = ~n39635 & ~n39636 ;
  assign n39638 = \u1_R6_reg[19]/NET0131  & ~n39637 ;
  assign n39639 = ~\u1_R6_reg[19]/NET0131  & n39637 ;
  assign n39640 = ~n39638 & ~n39639 ;
  assign n39648 = n39611 & ~n39626 ;
  assign n39649 = n39617 & n39632 ;
  assign n39650 = ~n39648 & ~n39649 ;
  assign n39651 = n39620 & n39650 ;
  assign n39654 = ~n39640 & ~n39651 ;
  assign n39655 = ~n39653 & n39654 ;
  assign n39656 = ~n39650 & ~n39652 ;
  assign n39657 = ~n39611 & ~n39632 ;
  assign n39658 = ~n39617 & n39657 ;
  assign n39659 = n39640 & ~n39658 ;
  assign n39660 = ~n39656 & n39659 ;
  assign n39661 = ~n39655 & ~n39660 ;
  assign n39662 = n39626 & n39632 ;
  assign n39663 = ~n39648 & ~n39662 ;
  assign n39664 = ~n39617 & n39632 ;
  assign n39665 = ~n39619 & ~n39664 ;
  assign n39666 = ~n39663 & n39665 ;
  assign n39667 = ~n39661 & ~n39666 ;
  assign n39668 = ~n39647 & ~n39667 ;
  assign n39669 = n39611 & n39664 ;
  assign n39670 = ~n39632 & n39648 ;
  assign n39671 = n39617 & ~n39662 ;
  assign n39672 = ~n39670 & n39671 ;
  assign n39673 = ~n39669 & ~n39672 ;
  assign n39674 = n39640 & ~n39673 ;
  assign n39676 = n39626 & ~n39649 ;
  assign n39675 = ~n39640 & ~n39652 ;
  assign n39677 = ~n39620 & n39675 ;
  assign n39678 = ~n39676 & n39677 ;
  assign n39679 = n39620 & n39652 ;
  assign n39680 = n39618 & n39662 ;
  assign n39681 = ~n39679 & ~n39680 ;
  assign n39682 = ~n39678 & n39681 ;
  assign n39683 = ~n39674 & n39682 ;
  assign n39684 = n39647 & ~n39683 ;
  assign n39633 = n39626 & ~n39632 ;
  assign n39634 = n39620 & n39633 ;
  assign n39641 = n39634 & ~n39640 ;
  assign n39685 = n39648 & n39664 ;
  assign n39686 = n39618 & n39633 ;
  assign n39687 = ~n39685 & ~n39686 ;
  assign n39688 = n39640 & ~n39687 ;
  assign n39689 = ~n39641 & ~n39688 ;
  assign n39690 = ~n39684 & n39689 ;
  assign n39691 = ~n39668 & n39690 ;
  assign n39692 = ~\u1_L6_reg[14]/NET0131  & ~n39691 ;
  assign n39693 = \u1_L6_reg[14]/NET0131  & n39691 ;
  assign n39694 = ~n39692 & ~n39693 ;
  assign n39695 = ~n39496 & ~n39522 ;
  assign n39696 = ~n39471 & n39695 ;
  assign n39697 = n39487 & ~n39696 ;
  assign n39698 = n39489 & n39515 ;
  assign n39699 = ~n39697 & ~n39698 ;
  assign n39700 = ~n39508 & ~n39699 ;
  assign n39701 = ~n39463 & n39512 ;
  assign n39712 = n39470 & n39520 ;
  assign n39713 = n39478 & ~n39487 ;
  assign n39714 = n39491 & n39713 ;
  assign n39719 = ~n39712 & ~n39714 ;
  assign n39720 = ~n39701 & n39719 ;
  assign n39715 = n39463 & n39514 ;
  assign n39716 = ~n39457 & ~n39463 ;
  assign n39717 = ~n39470 & n39716 ;
  assign n39718 = n39487 & n39717 ;
  assign n39721 = ~n39715 & ~n39718 ;
  assign n39722 = n39720 & n39721 ;
  assign n39723 = n39508 & ~n39722 ;
  assign n39702 = n39464 & n39495 ;
  assign n39703 = ~n39514 & ~n39702 ;
  assign n39704 = ~n39535 & n39703 ;
  assign n39705 = ~n39701 & n39704 ;
  assign n39706 = ~n39487 & ~n39705 ;
  assign n39707 = n39471 & ~n39478 ;
  assign n39708 = ~n39513 & ~n39707 ;
  assign n39709 = n39487 & ~n39708 ;
  assign n39710 = ~n39487 & ~n39508 ;
  assign n39711 = n39472 & n39710 ;
  assign n39724 = ~n39709 & ~n39711 ;
  assign n39725 = ~n39706 & n39724 ;
  assign n39726 = ~n39723 & n39725 ;
  assign n39727 = ~n39700 & n39726 ;
  assign n39728 = \u1_L6_reg[15]/P0001  & n39727 ;
  assign n39729 = ~\u1_L6_reg[15]/P0001  & ~n39727 ;
  assign n39730 = ~n39728 & ~n39729 ;
  assign n39749 = ~n39202 & ~n39212 ;
  assign n39750 = n39201 & n39226 ;
  assign n39751 = n39749 & ~n39750 ;
  assign n39752 = n39210 & ~n39751 ;
  assign n39755 = ~n39210 & ~n39226 ;
  assign n39756 = n39749 & n39755 ;
  assign n39748 = n39199 & n39250 ;
  assign n39753 = n39185 & n39192 ;
  assign n39754 = n39179 & n39753 ;
  assign n39757 = ~n39748 & ~n39754 ;
  assign n39758 = ~n39756 & n39757 ;
  assign n39759 = ~n39752 & n39758 ;
  assign n39760 = n39173 & ~n39759 ;
  assign n39733 = ~n39179 & ~n39235 ;
  assign n39734 = ~n39192 & n39234 ;
  assign n39735 = ~n39733 & ~n39734 ;
  assign n39736 = ~n39210 & ~n39735 ;
  assign n39737 = ~n39241 & ~n39243 ;
  assign n39738 = n39210 & ~n39737 ;
  assign n39731 = n39192 & n39228 ;
  assign n39732 = n39199 & n39731 ;
  assign n39739 = ~n39249 & ~n39732 ;
  assign n39740 = ~n39738 & n39739 ;
  assign n39741 = ~n39736 & n39740 ;
  assign n39742 = ~n39173 & ~n39741 ;
  assign n39745 = n39192 & ~n39229 ;
  assign n39743 = n39185 & n39212 ;
  assign n39744 = ~n39192 & ~n39743 ;
  assign n39746 = n39210 & ~n39744 ;
  assign n39747 = ~n39745 & n39746 ;
  assign n39761 = ~n39742 & ~n39747 ;
  assign n39762 = ~n39760 & n39761 ;
  assign n39763 = ~\u1_L6_reg[17]/NET0131  & ~n39762 ;
  assign n39764 = \u1_L6_reg[17]/NET0131  & n39762 ;
  assign n39765 = ~n39763 & ~n39764 ;
  assign n39766 = ~n39370 & n39559 ;
  assign n39767 = ~n39383 & ~n39766 ;
  assign n39768 = ~n39391 & n39414 ;
  assign n39769 = ~n39403 & ~n39768 ;
  assign n39770 = n39413 & ~n39769 ;
  assign n39771 = n39383 & ~n39419 ;
  assign n39772 = ~n39560 & n39771 ;
  assign n39773 = ~n39770 & n39772 ;
  assign n39774 = ~n39767 & ~n39773 ;
  assign n39775 = ~n39421 & n39559 ;
  assign n39776 = n39377 & ~n39383 ;
  assign n39777 = ~n39418 & n39776 ;
  assign n39778 = ~n39544 & n39777 ;
  assign n39779 = n39413 & ~n39778 ;
  assign n39780 = ~n39775 & n39779 ;
  assign n39784 = n39377 & n39394 ;
  assign n39785 = n39364 & ~n39397 ;
  assign n39786 = ~n39418 & n39785 ;
  assign n39787 = ~n39784 & n39786 ;
  assign n39781 = n39414 & n39418 ;
  assign n39782 = ~n39399 & ~n39781 ;
  assign n39783 = n39383 & ~n39782 ;
  assign n39788 = ~n39413 & ~n39429 ;
  assign n39789 = ~n39783 & n39788 ;
  assign n39790 = ~n39787 & n39789 ;
  assign n39791 = ~n39780 & ~n39790 ;
  assign n39792 = ~n39774 & ~n39791 ;
  assign n39793 = ~\u1_L6_reg[1]/NET0131  & ~n39792 ;
  assign n39794 = \u1_L6_reg[1]/NET0131  & n39792 ;
  assign n39795 = ~n39793 & ~n39794 ;
  assign n39797 = n39463 & n39520 ;
  assign n39804 = ~n39470 & n39487 ;
  assign n39805 = n39797 & ~n39804 ;
  assign n39807 = ~n39508 & ~n39512 ;
  assign n39800 = n39464 & n39713 ;
  assign n39796 = n39470 & ~n39487 ;
  assign n39806 = n39716 & n39796 ;
  assign n39808 = ~n39800 & ~n39806 ;
  assign n39809 = n39807 & n39808 ;
  assign n39810 = ~n39805 & n39809 ;
  assign n39801 = ~n39463 & ~n39517 ;
  assign n39802 = ~n39514 & ~n39523 ;
  assign n39803 = n39487 & ~n39802 ;
  assign n39811 = ~n39801 & ~n39803 ;
  assign n39812 = n39810 & n39811 ;
  assign n39815 = ~n39490 & ~n39713 ;
  assign n39816 = ~n39715 & ~n39815 ;
  assign n39817 = n39463 & n39515 ;
  assign n39820 = n39487 & ~n39817 ;
  assign n39818 = n39464 & n39470 ;
  assign n39819 = n39478 & n39522 ;
  assign n39821 = ~n39818 & ~n39819 ;
  assign n39822 = n39820 & n39821 ;
  assign n39823 = ~n39816 & ~n39822 ;
  assign n39813 = ~n39523 & ~n39717 ;
  assign n39814 = n39478 & ~n39813 ;
  assign n39824 = n39508 & ~n39707 ;
  assign n39825 = ~n39814 & n39824 ;
  assign n39826 = ~n39823 & n39825 ;
  assign n39827 = ~n39812 & ~n39826 ;
  assign n39798 = n39796 & n39797 ;
  assign n39799 = n39487 & n39516 ;
  assign n39828 = ~n39798 & ~n39799 ;
  assign n39829 = ~n39827 & n39828 ;
  assign n39830 = ~\u1_L6_reg[21]/NET0131  & ~n39829 ;
  assign n39831 = \u1_L6_reg[21]/NET0131  & n39829 ;
  assign n39832 = ~n39830 & ~n39831 ;
  assign n39839 = n39611 & ~n39617 ;
  assign n39840 = n39640 & ~n39839 ;
  assign n39838 = ~n39640 & ~n39657 ;
  assign n39841 = ~n39626 & ~n39838 ;
  assign n39842 = ~n39840 & n39841 ;
  assign n39833 = ~n39617 & n39640 ;
  assign n39834 = n39611 & n39633 ;
  assign n39835 = ~n39833 & n39834 ;
  assign n39836 = n39632 & ~n39640 ;
  assign n39837 = n39618 & n39836 ;
  assign n39843 = ~n39647 & ~n39837 ;
  assign n39844 = ~n39835 & n39843 ;
  assign n39845 = ~n39842 & n39844 ;
  assign n39846 = ~n39611 & n39649 ;
  assign n39847 = ~n39640 & ~n39846 ;
  assign n39848 = ~n39670 & n39847 ;
  assign n39850 = ~n39617 & n39663 ;
  assign n39849 = n39611 & n39649 ;
  assign n39851 = n39640 & ~n39657 ;
  assign n39852 = ~n39849 & n39851 ;
  assign n39853 = ~n39850 & n39852 ;
  assign n39854 = ~n39848 & ~n39853 ;
  assign n39856 = n39662 & n39839 ;
  assign n39855 = n39617 & n39648 ;
  assign n39857 = n39647 & ~n39855 ;
  assign n39858 = ~n39856 & n39857 ;
  assign n39859 = ~n39854 & n39858 ;
  assign n39860 = ~n39845 & ~n39859 ;
  assign n39863 = ~n39686 & ~n39856 ;
  assign n39864 = n39617 & ~n39626 ;
  assign n39865 = n39657 & n39864 ;
  assign n39866 = n39863 & ~n39865 ;
  assign n39867 = n39640 & ~n39866 ;
  assign n39861 = ~n39611 & n39626 ;
  assign n39862 = n39836 & n39861 ;
  assign n39868 = ~n39626 & n39849 ;
  assign n39869 = ~n39862 & ~n39868 ;
  assign n39870 = ~n39867 & n39869 ;
  assign n39871 = ~n39860 & n39870 ;
  assign n39872 = ~\u1_L6_reg[25]/NET0131  & ~n39871 ;
  assign n39873 = \u1_L6_reg[25]/NET0131  & n39871 ;
  assign n39874 = ~n39872 & ~n39873 ;
  assign n39893 = ~n39370 & ~n39433 ;
  assign n39894 = ~n39436 & ~n39893 ;
  assign n39895 = ~n39391 & ~n39894 ;
  assign n39875 = n39370 & ~n39406 ;
  assign n39896 = ~n39377 & ~n39413 ;
  assign n39897 = ~n39875 & n39896 ;
  assign n39898 = ~n39895 & ~n39897 ;
  assign n39899 = ~n39383 & ~n39898 ;
  assign n39879 = n39377 & ~n39401 ;
  assign n39876 = n39364 & ~n39391 ;
  assign n39877 = n39561 & ~n39876 ;
  assign n39878 = n39875 & n39877 ;
  assign n39880 = n39391 & n39431 ;
  assign n39881 = ~n39437 & n39880 ;
  assign n39882 = n39413 & ~n39416 ;
  assign n39883 = ~n39881 & n39882 ;
  assign n39884 = ~n39878 & n39883 ;
  assign n39885 = ~n39879 & n39884 ;
  assign n39886 = n39384 & n39391 ;
  assign n39887 = ~n39431 & n39886 ;
  assign n39888 = ~n39413 & ~n39768 ;
  assign n39889 = n39430 & n39888 ;
  assign n39890 = ~n39887 & n39889 ;
  assign n39891 = ~n39885 & ~n39890 ;
  assign n39892 = ~n39433 & n39549 ;
  assign n39900 = ~n39891 & ~n39892 ;
  assign n39901 = ~n39899 & n39900 ;
  assign n39902 = ~\u1_L6_reg[26]/NET0131  & ~n39901 ;
  assign n39903 = \u1_L6_reg[26]/NET0131  & n39901 ;
  assign n39904 = ~n39902 & ~n39903 ;
  assign n39942 = decrypt_pad & ~\u1_uk_K_r6_reg[48]/NET0131  ;
  assign n39943 = ~decrypt_pad & ~\u1_uk_K_r6_reg[55]/P0001  ;
  assign n39944 = ~n39942 & ~n39943 ;
  assign n39945 = \u1_R6_reg[8]/NET0131  & ~n39944 ;
  assign n39946 = ~\u1_R6_reg[8]/NET0131  & n39944 ;
  assign n39947 = ~n39945 & ~n39946 ;
  assign n39935 = decrypt_pad & ~\u1_uk_K_r6_reg[25]/NET0131  ;
  assign n39936 = ~decrypt_pad & ~\u1_uk_K_r6_reg[32]/NET0131  ;
  assign n39937 = ~n39935 & ~n39936 ;
  assign n39938 = \u1_R6_reg[7]/NET0131  & ~n39937 ;
  assign n39939 = ~\u1_R6_reg[7]/NET0131  & n39937 ;
  assign n39940 = ~n39938 & ~n39939 ;
  assign n39905 = decrypt_pad & ~\u1_uk_K_r6_reg[40]/NET0131  ;
  assign n39906 = ~decrypt_pad & ~\u1_uk_K_r6_reg[47]/NET0131  ;
  assign n39907 = ~n39905 & ~n39906 ;
  assign n39908 = \u1_R6_reg[5]/NET0131  & ~n39907 ;
  assign n39909 = ~\u1_R6_reg[5]/NET0131  & n39907 ;
  assign n39910 = ~n39908 & ~n39909 ;
  assign n39918 = decrypt_pad & ~\u1_uk_K_r6_reg[4]/NET0131  ;
  assign n39919 = ~decrypt_pad & ~\u1_uk_K_r6_reg[11]/NET0131  ;
  assign n39920 = ~n39918 & ~n39919 ;
  assign n39921 = \u1_R6_reg[4]/NET0131  & ~n39920 ;
  assign n39922 = ~\u1_R6_reg[4]/NET0131  & n39920 ;
  assign n39923 = ~n39921 & ~n39922 ;
  assign n39926 = decrypt_pad & ~\u1_uk_K_r6_reg[53]/NET0131  ;
  assign n39927 = ~decrypt_pad & ~\u1_uk_K_r6_reg[3]/NET0131  ;
  assign n39928 = ~n39926 & ~n39927 ;
  assign n39929 = \u1_R6_reg[9]/NET0131  & ~n39928 ;
  assign n39930 = ~\u1_R6_reg[9]/NET0131  & n39928 ;
  assign n39931 = ~n39929 & ~n39930 ;
  assign n39948 = n39923 & ~n39931 ;
  assign n39949 = ~n39910 & n39948 ;
  assign n39961 = n39910 & n39923 ;
  assign n39975 = n39931 & n39961 ;
  assign n39976 = ~n39949 & ~n39975 ;
  assign n39955 = ~n39923 & ~n39931 ;
  assign n39911 = decrypt_pad & ~\u1_uk_K_r6_reg[6]/NET0131  ;
  assign n39912 = ~decrypt_pad & ~\u1_uk_K_r6_reg[13]/NET0131  ;
  assign n39913 = ~n39911 & ~n39912 ;
  assign n39914 = \u1_R6_reg[6]/NET0131  & ~n39913 ;
  assign n39915 = ~\u1_R6_reg[6]/NET0131  & n39913 ;
  assign n39916 = ~n39914 & ~n39915 ;
  assign n39977 = n39910 & n39916 ;
  assign n39978 = n39955 & n39977 ;
  assign n39979 = n39976 & ~n39978 ;
  assign n39980 = n39940 & ~n39979 ;
  assign n39956 = ~n39916 & n39955 ;
  assign n39952 = ~n39923 & n39931 ;
  assign n39957 = n39910 & n39952 ;
  assign n39958 = ~n39956 & ~n39957 ;
  assign n39974 = ~n39940 & ~n39958 ;
  assign n39962 = ~n39916 & n39923 ;
  assign n39970 = ~n39910 & n39931 ;
  assign n39971 = n39923 & n39970 ;
  assign n39972 = ~n39940 & ~n39971 ;
  assign n39973 = n39962 & ~n39972 ;
  assign n39981 = n39916 & n39952 ;
  assign n39982 = ~n39910 & n39981 ;
  assign n39983 = ~n39973 & ~n39982 ;
  assign n39984 = ~n39974 & n39983 ;
  assign n39985 = ~n39980 & n39984 ;
  assign n39986 = n39947 & ~n39985 ;
  assign n39917 = ~n39910 & n39916 ;
  assign n39924 = n39917 & ~n39923 ;
  assign n39925 = n39916 & n39923 ;
  assign n39932 = n39910 & ~n39931 ;
  assign n39933 = n39925 & n39932 ;
  assign n39934 = ~n39924 & ~n39933 ;
  assign n39941 = ~n39934 & ~n39940 ;
  assign n39963 = ~n39931 & n39962 ;
  assign n39960 = ~n39910 & n39952 ;
  assign n39964 = ~n39960 & ~n39961 ;
  assign n39965 = ~n39963 & n39964 ;
  assign n39966 = ~n39940 & ~n39965 ;
  assign n39950 = n39910 & ~n39948 ;
  assign n39951 = ~n39949 & ~n39950 ;
  assign n39953 = n39916 & ~n39952 ;
  assign n39954 = n39951 & n39953 ;
  assign n39959 = n39940 & ~n39958 ;
  assign n39967 = ~n39954 & ~n39959 ;
  assign n39968 = ~n39966 & n39967 ;
  assign n39969 = ~n39947 & ~n39968 ;
  assign n39987 = ~n39941 & ~n39969 ;
  assign n39988 = ~n39986 & n39987 ;
  assign n39989 = ~\u1_L6_reg[28]/NET0131  & ~n39988 ;
  assign n39990 = \u1_L6_reg[28]/NET0131  & n39988 ;
  assign n39991 = ~n39989 & ~n39990 ;
  assign n39997 = ~n39267 & n39298 ;
  assign n39998 = n39342 & ~n39997 ;
  assign n39999 = ~n39267 & ~n39280 ;
  assign n40000 = ~n39281 & ~n39999 ;
  assign n40001 = ~n39298 & ~n40000 ;
  assign n40002 = ~n39998 & ~n40001 ;
  assign n40003 = n39290 & ~n40002 ;
  assign n39992 = ~n39280 & ~n39337 ;
  assign n39993 = n39280 & ~n39298 ;
  assign n39994 = n39282 & n39993 ;
  assign n39995 = ~n39992 & ~n39994 ;
  assign n39996 = ~n39290 & ~n39995 ;
  assign n40004 = ~n39273 & n39997 ;
  assign n40005 = n39280 & n40004 ;
  assign n40006 = ~n39996 & ~n40005 ;
  assign n40007 = ~n40003 & n40006 ;
  assign n40008 = ~n39321 & ~n40007 ;
  assign n40013 = n39274 & ~n39993 ;
  assign n40014 = ~n39994 & ~n40013 ;
  assign n40015 = n39290 & ~n40014 ;
  assign n40017 = n39280 & ~n39304 ;
  assign n40018 = ~n39332 & n40017 ;
  assign n40016 = n39290 & ~n39343 ;
  assign n40019 = ~n39992 & ~n40016 ;
  assign n40020 = ~n40018 & n40019 ;
  assign n40021 = ~n40015 & ~n40020 ;
  assign n40022 = n39321 & ~n40021 ;
  assign n40009 = ~n39267 & n39273 ;
  assign n40010 = n39299 & n40009 ;
  assign n40011 = n39267 & n39298 ;
  assign n40012 = n39292 & n40011 ;
  assign n40023 = ~n40010 & ~n40012 ;
  assign n40024 = ~n40022 & n40023 ;
  assign n40025 = ~n40008 & n40024 ;
  assign n40026 = \u1_L6_reg[29]/NET0131  & ~n40025 ;
  assign n40027 = ~\u1_L6_reg[29]/NET0131  & n40025 ;
  assign n40028 = ~n40026 & ~n40027 ;
  assign n40029 = ~n39932 & ~n39960 ;
  assign n40030 = ~n39916 & ~n40029 ;
  assign n40031 = ~n39940 & ~n39947 ;
  assign n40032 = n39925 & n39970 ;
  assign n40033 = ~n39947 & ~n40032 ;
  assign n40034 = ~n40031 & ~n40033 ;
  assign n40041 = ~n40030 & ~n40034 ;
  assign n40035 = ~n39925 & ~n39970 ;
  assign n40036 = n39972 & ~n40035 ;
  assign n40037 = n39916 & n39957 ;
  assign n40038 = ~n39916 & ~n39940 ;
  assign n40039 = n39970 & n40038 ;
  assign n40040 = ~n40037 & ~n40039 ;
  assign n40042 = ~n40036 & n40040 ;
  assign n40043 = n40041 & n40042 ;
  assign n40047 = ~n39916 & ~n39976 ;
  assign n40044 = n39910 & ~n39916 ;
  assign n40045 = ~n39961 & ~n40044 ;
  assign n40046 = n39940 & ~n40045 ;
  assign n40048 = n39947 & ~n40046 ;
  assign n40049 = ~n40047 & n40048 ;
  assign n40050 = ~n40043 & ~n40049 ;
  assign n40051 = ~n39955 & ~n40032 ;
  assign n40052 = n39947 & ~n40051 ;
  assign n40053 = ~n39917 & n39952 ;
  assign n40054 = ~n40052 & ~n40053 ;
  assign n40055 = ~n40044 & ~n40054 ;
  assign n40056 = ~n39940 & ~n40055 ;
  assign n40058 = n39924 & ~n39931 ;
  assign n40057 = ~n39916 & n39961 ;
  assign n40059 = n39940 & ~n40057 ;
  assign n40060 = ~n40058 & n40059 ;
  assign n40061 = ~n40056 & ~n40060 ;
  assign n40062 = ~n40050 & ~n40061 ;
  assign n40063 = \u1_L6_reg[2]/NET0131  & n40062 ;
  assign n40064 = ~\u1_L6_reg[2]/NET0131  & ~n40062 ;
  assign n40065 = ~n40063 & ~n40064 ;
  assign n40068 = n39292 & n39304 ;
  assign n40066 = n39280 & n40011 ;
  assign n40069 = n39321 & ~n40066 ;
  assign n40070 = ~n40068 & n40069 ;
  assign n40067 = n39331 & ~n39342 ;
  assign n40071 = ~n39324 & ~n40067 ;
  assign n40072 = n40070 & n40071 ;
  assign n40074 = n39290 & ~n39327 ;
  assign n40073 = ~n39280 & n39309 ;
  assign n40075 = ~n39306 & ~n40073 ;
  assign n40076 = n40074 & n40075 ;
  assign n40077 = ~n39290 & ~n39323 ;
  assign n40078 = ~n40005 & n40077 ;
  assign n40079 = ~n40076 & ~n40078 ;
  assign n40080 = ~n39321 & ~n39347 ;
  assign n40081 = ~n40010 & n40080 ;
  assign n40082 = ~n40079 & n40081 ;
  assign n40083 = ~n40072 & ~n40082 ;
  assign n40085 = ~n39273 & ~n39341 ;
  assign n40086 = ~n39997 & n40085 ;
  assign n40087 = n40074 & ~n40086 ;
  assign n40084 = ~n39290 & ~n39998 ;
  assign n40088 = n39280 & ~n40084 ;
  assign n40089 = ~n40087 & n40088 ;
  assign n40090 = ~n39333 & ~n40089 ;
  assign n40091 = ~n40083 & n40090 ;
  assign n40092 = ~\u1_L6_reg[4]/NET0131  & ~n40091 ;
  assign n40093 = \u1_L6_reg[4]/NET0131  & n40091 ;
  assign n40094 = ~n40092 & ~n40093 ;
  assign n40097 = ~n39290 & n40086 ;
  assign n40095 = ~n39283 & n39290 ;
  assign n40096 = ~n40085 & n40095 ;
  assign n40098 = n39273 & n40066 ;
  assign n40099 = ~n39321 & ~n40098 ;
  assign n40100 = ~n40096 & n40099 ;
  assign n40101 = ~n40097 & n40100 ;
  assign n40102 = n39280 & n40086 ;
  assign n40107 = ~n39310 & n39321 ;
  assign n40108 = ~n40102 & n40107 ;
  assign n40103 = ~n39341 & ~n40004 ;
  assign n40104 = ~n39280 & ~n40103 ;
  assign n40105 = ~n39290 & ~n40009 ;
  assign n40106 = ~n40095 & ~n40105 ;
  assign n40109 = ~n40104 & ~n40106 ;
  assign n40110 = n40108 & n40109 ;
  assign n40111 = ~n40101 & ~n40110 ;
  assign n40112 = ~n39330 & ~n39348 ;
  assign n40113 = ~n40111 & n40112 ;
  assign n40114 = ~\u1_L6_reg[19]/NET0131  & ~n40113 ;
  assign n40115 = \u1_L6_reg[19]/NET0131  & n40113 ;
  assign n40116 = ~n40114 & ~n40115 ;
  assign n40133 = ~n39201 & ~n39229 ;
  assign n40134 = ~n39199 & ~n40133 ;
  assign n40135 = ~n39244 & ~n40134 ;
  assign n40136 = n39173 & ~n40135 ;
  assign n40137 = n39201 & n39245 ;
  assign n40138 = ~n39242 & ~n40137 ;
  assign n40139 = ~n39748 & n40138 ;
  assign n40140 = ~n40136 & n40139 ;
  assign n40141 = ~n39210 & ~n40140 ;
  assign n40123 = ~n39173 & ~n39193 ;
  assign n40124 = ~n39754 & n40123 ;
  assign n40117 = ~n39179 & ~n39753 ;
  assign n40118 = n39199 & ~n39210 ;
  assign n40119 = ~n40117 & n40118 ;
  assign n40120 = ~n39228 & ~n39753 ;
  assign n40121 = ~n39199 & n39210 ;
  assign n40122 = ~n40120 & n40121 ;
  assign n40125 = ~n40119 & ~n40122 ;
  assign n40126 = n40124 & n40125 ;
  assign n40127 = ~n39226 & n39237 ;
  assign n40128 = n39173 & ~n39750 ;
  assign n40129 = ~n39225 & n40128 ;
  assign n40130 = ~n40127 & n40129 ;
  assign n40131 = ~n40126 & ~n40130 ;
  assign n40132 = n39216 & n39229 ;
  assign n40142 = ~n39227 & ~n40132 ;
  assign n40143 = ~n40131 & n40142 ;
  assign n40144 = ~n40141 & n40143 ;
  assign n40145 = \u1_L6_reg[23]/NET0131  & ~n40144 ;
  assign n40146 = ~\u1_L6_reg[23]/NET0131  & n40144 ;
  assign n40147 = ~n40145 & ~n40146 ;
  assign n40148 = ~n39516 & ~n39523 ;
  assign n40149 = ~n39818 & n40148 ;
  assign n40150 = ~n39487 & ~n40149 ;
  assign n40151 = n39487 & ~n39489 ;
  assign n40152 = ~n39695 & n40151 ;
  assign n40153 = ~n39480 & ~n39817 ;
  assign n40154 = ~n39513 & n40153 ;
  assign n40155 = ~n40152 & n40154 ;
  assign n40156 = ~n40150 & n40155 ;
  assign n40157 = n39508 & ~n40156 ;
  assign n40163 = n39487 & ~n39496 ;
  assign n40162 = n39463 & ~n39495 ;
  assign n40164 = ~n39512 & ~n40162 ;
  assign n40165 = n40163 & n40164 ;
  assign n40160 = n39457 & n39463 ;
  assign n40161 = n39713 & n40160 ;
  assign n40166 = ~n39806 & ~n40161 ;
  assign n40167 = ~n39534 & n40166 ;
  assign n40168 = ~n40165 & n40167 ;
  assign n40169 = ~n39508 & ~n40168 ;
  assign n40158 = ~n39487 & n39533 ;
  assign n40159 = n39479 & n39804 ;
  assign n40170 = ~n39531 & ~n40159 ;
  assign n40171 = ~n40158 & n40170 ;
  assign n40172 = ~n40169 & n40171 ;
  assign n40173 = ~n40157 & n40172 ;
  assign n40174 = ~\u1_L6_reg[27]/NET0131  & ~n40173 ;
  assign n40175 = \u1_L6_reg[27]/NET0131  & n40173 ;
  assign n40176 = ~n40174 & ~n40175 ;
  assign n40182 = ~n39135 & ~n39156 ;
  assign n40184 = ~n39122 & n39584 ;
  assign n40185 = n40182 & ~n40184 ;
  assign n40183 = ~n39122 & ~n40182 ;
  assign n40186 = ~n39114 & ~n40183 ;
  assign n40187 = ~n40185 & n40186 ;
  assign n40177 = n39124 & n39156 ;
  assign n40178 = n39087 & ~n39156 ;
  assign n40179 = n39145 & ~n40178 ;
  assign n40180 = ~n39107 & ~n40179 ;
  assign n40181 = n39114 & ~n40180 ;
  assign n40188 = ~n40177 & ~n40181 ;
  assign n40189 = ~n40187 & n40188 ;
  assign n40190 = n39081 & ~n40189 ;
  assign n40192 = ~n39576 & ~n39584 ;
  assign n40193 = ~n39114 & ~n40192 ;
  assign n40194 = ~n39093 & n39138 ;
  assign n40195 = n39114 & ~n39576 ;
  assign n40196 = ~n40194 & n40195 ;
  assign n40197 = ~n40193 & ~n40196 ;
  assign n40191 = n39093 & ~n39578 ;
  assign n40198 = n39155 & ~n40191 ;
  assign n40199 = ~n40197 & n40198 ;
  assign n40200 = ~n39081 & ~n40199 ;
  assign n40201 = n39114 & n39137 ;
  assign n40202 = ~n39125 & n39152 ;
  assign n40203 = n39118 & n40202 ;
  assign n40204 = ~n40201 & ~n40203 ;
  assign n40205 = ~n40200 & n40204 ;
  assign n40206 = ~n40190 & n40205 ;
  assign n40207 = \u1_L6_reg[32]/NET0131  & n40206 ;
  assign n40208 = ~\u1_L6_reg[32]/NET0131  & ~n40206 ;
  assign n40209 = ~n40207 & ~n40208 ;
  assign n40210 = decrypt_pad & ~\u1_uk_K_r6_reg[39]/NET0131  ;
  assign n40211 = ~decrypt_pad & ~\u1_uk_K_r6_reg[46]/NET0131  ;
  assign n40212 = ~n40210 & ~n40211 ;
  assign n40213 = \u1_R6_reg[13]/NET0131  & ~n40212 ;
  assign n40214 = ~\u1_R6_reg[13]/NET0131  & n40212 ;
  assign n40215 = ~n40213 & ~n40214 ;
  assign n40230 = decrypt_pad & ~\u1_uk_K_r6_reg[34]/NET0131  ;
  assign n40231 = ~decrypt_pad & ~\u1_uk_K_r6_reg[41]/NET0131  ;
  assign n40232 = ~n40230 & ~n40231 ;
  assign n40233 = \u1_R6_reg[9]/NET0131  & ~n40232 ;
  assign n40234 = ~\u1_R6_reg[9]/NET0131  & n40232 ;
  assign n40235 = ~n40233 & ~n40234 ;
  assign n40237 = ~n40215 & n40235 ;
  assign n40238 = decrypt_pad & ~\u1_uk_K_r6_reg[11]/NET0131  ;
  assign n40239 = ~decrypt_pad & ~\u1_uk_K_r6_reg[18]/NET0131  ;
  assign n40240 = ~n40238 & ~n40239 ;
  assign n40241 = \u1_R6_reg[11]/NET0131  & ~n40240 ;
  assign n40242 = ~\u1_R6_reg[11]/NET0131  & n40240 ;
  assign n40243 = ~n40241 & ~n40242 ;
  assign n40244 = ~n40237 & ~n40243 ;
  assign n40223 = decrypt_pad & ~\u1_uk_K_r6_reg[10]/NET0131  ;
  assign n40224 = ~decrypt_pad & ~\u1_uk_K_r6_reg[17]/NET0131  ;
  assign n40225 = ~n40223 & ~n40224 ;
  assign n40226 = \u1_R6_reg[10]/NET0131  & ~n40225 ;
  assign n40227 = ~\u1_R6_reg[10]/NET0131  & n40225 ;
  assign n40228 = ~n40226 & ~n40227 ;
  assign n40245 = ~n40228 & n40235 ;
  assign n40216 = decrypt_pad & ~\u1_uk_K_r6_reg[5]/NET0131  ;
  assign n40217 = ~decrypt_pad & ~\u1_uk_K_r6_reg[12]/NET0131  ;
  assign n40218 = ~n40216 & ~n40217 ;
  assign n40219 = \u1_R6_reg[8]/NET0131  & ~n40218 ;
  assign n40220 = ~\u1_R6_reg[8]/NET0131  & n40218 ;
  assign n40221 = ~n40219 & ~n40220 ;
  assign n40246 = n40215 & ~n40235 ;
  assign n40247 = n40221 & ~n40246 ;
  assign n40248 = ~n40245 & ~n40247 ;
  assign n40249 = n40244 & ~n40248 ;
  assign n40222 = ~n40215 & ~n40221 ;
  assign n40229 = n40222 & n40228 ;
  assign n40236 = n40229 & n40235 ;
  assign n40250 = decrypt_pad & ~\u1_uk_K_r6_reg[26]/NET0131  ;
  assign n40251 = ~decrypt_pad & ~\u1_uk_K_r6_reg[33]/NET0131  ;
  assign n40252 = ~n40250 & ~n40251 ;
  assign n40253 = \u1_R6_reg[12]/NET0131  & ~n40252 ;
  assign n40254 = ~\u1_R6_reg[12]/NET0131  & n40252 ;
  assign n40255 = ~n40253 & ~n40254 ;
  assign n40256 = ~n40236 & n40255 ;
  assign n40257 = ~n40249 & n40256 ;
  assign n40260 = n40228 & ~n40235 ;
  assign n40261 = ~n40245 & ~n40260 ;
  assign n40258 = ~n40221 & n40243 ;
  assign n40262 = n40215 & n40221 ;
  assign n40263 = ~n40222 & ~n40262 ;
  assign n40264 = ~n40258 & n40263 ;
  assign n40265 = n40261 & n40264 ;
  assign n40266 = ~n40261 & ~n40263 ;
  assign n40259 = n40245 & n40258 ;
  assign n40267 = ~n40255 & ~n40259 ;
  assign n40268 = ~n40266 & n40267 ;
  assign n40269 = ~n40265 & n40268 ;
  assign n40270 = ~n40257 & ~n40269 ;
  assign n40274 = n40215 & ~n40221 ;
  assign n40275 = n40228 & n40274 ;
  assign n40276 = n40221 & n40237 ;
  assign n40277 = ~n40275 & ~n40276 ;
  assign n40278 = ~n40246 & n40277 ;
  assign n40279 = n40255 & ~n40278 ;
  assign n40271 = ~n40221 & ~n40228 ;
  assign n40272 = ~n40215 & n40271 ;
  assign n40273 = ~n40235 & n40272 ;
  assign n40280 = n40215 & n40260 ;
  assign n40281 = ~n40273 & ~n40280 ;
  assign n40282 = ~n40279 & n40281 ;
  assign n40283 = n40243 & ~n40282 ;
  assign n40284 = ~n40270 & ~n40283 ;
  assign n40285 = ~\u1_L6_reg[6]/NET0131  & ~n40284 ;
  assign n40286 = \u1_L6_reg[6]/NET0131  & n40284 ;
  assign n40287 = ~n40285 & ~n40286 ;
  assign n40305 = ~n39106 & ~n39582 ;
  assign n40288 = n39093 & ~n40182 ;
  assign n40306 = n39087 & n39156 ;
  assign n40307 = ~n40288 & ~n40306 ;
  assign n40308 = ~n40305 & n40307 ;
  assign n40309 = ~n39114 & ~n40308 ;
  assign n40289 = ~n40194 & ~n40288 ;
  assign n40290 = n39087 & ~n40289 ;
  assign n40299 = ~n39087 & ~n39100 ;
  assign n40300 = n40182 & n40299 ;
  assign n40310 = n39114 & n40300 ;
  assign n40311 = ~n40290 & ~n40310 ;
  assign n40312 = ~n40309 & n40311 ;
  assign n40313 = n39081 & ~n40312 ;
  assign n40291 = ~n39114 & n40290 ;
  assign n40292 = n39081 & ~n39114 ;
  assign n40293 = n39144 & ~n40182 ;
  assign n40294 = n39099 & ~n39594 ;
  assign n40295 = n39114 & n40178 ;
  assign n40296 = ~n40294 & n40295 ;
  assign n40297 = ~n40293 & ~n40296 ;
  assign n40298 = ~n39081 & ~n40297 ;
  assign n40301 = ~n39114 & n40300 ;
  assign n40302 = ~n39108 & ~n40301 ;
  assign n40303 = ~n40298 & n40302 ;
  assign n40304 = ~n40292 & ~n40303 ;
  assign n40314 = ~n40291 & ~n40304 ;
  assign n40315 = ~n40313 & n40314 ;
  assign n40316 = ~\u1_L6_reg[7]/NET0131  & ~n40315 ;
  assign n40317 = \u1_L6_reg[7]/NET0131  & n40315 ;
  assign n40318 = ~n40316 & ~n40317 ;
  assign n40330 = n39617 & ~n39632 ;
  assign n40331 = ~n39861 & n40330 ;
  assign n40332 = n39847 & ~n40331 ;
  assign n40333 = n39618 & n39652 ;
  assign n40334 = n39640 & ~n40333 ;
  assign n40335 = ~n39849 & n40334 ;
  assign n40336 = ~n40332 & ~n40335 ;
  assign n40337 = ~n39670 & n39863 ;
  assign n40338 = ~n40336 & n40337 ;
  assign n40339 = ~n39647 & ~n40338 ;
  assign n40319 = ~n39626 & n39658 ;
  assign n40320 = n39640 & ~n39846 ;
  assign n40321 = ~n40319 & n40320 ;
  assign n40322 = ~n39675 & ~n40321 ;
  assign n40323 = ~n39634 & ~n40322 ;
  assign n40324 = n39647 & ~n40323 ;
  assign n40325 = n39620 & n39676 ;
  assign n40326 = n39617 & n39670 ;
  assign n40327 = ~n40325 & ~n40326 ;
  assign n40328 = n39640 & ~n40327 ;
  assign n40329 = n39626 & n39837 ;
  assign n40340 = ~n40328 & ~n40329 ;
  assign n40341 = ~n40324 & n40340 ;
  assign n40342 = ~n40339 & n40341 ;
  assign n40343 = ~\u1_L6_reg[8]/NET0131  & ~n40342 ;
  assign n40344 = \u1_L6_reg[8]/NET0131  & n40342 ;
  assign n40345 = ~n40343 & ~n40344 ;
  assign n40347 = n40235 & n40262 ;
  assign n40348 = ~n40235 & ~n40262 ;
  assign n40349 = ~n40347 & ~n40348 ;
  assign n40350 = ~n40222 & ~n40349 ;
  assign n40351 = n40237 & n40258 ;
  assign n40352 = ~n40350 & ~n40351 ;
  assign n40353 = ~n40228 & ~n40352 ;
  assign n40346 = n40235 & n40275 ;
  assign n40355 = ~n40215 & ~n40243 ;
  assign n40354 = n40221 & n40228 ;
  assign n40356 = ~n40271 & ~n40354 ;
  assign n40357 = n40355 & n40356 ;
  assign n40358 = ~n40346 & ~n40357 ;
  assign n40359 = ~n40353 & n40358 ;
  assign n40360 = n40255 & ~n40359 ;
  assign n40363 = n40243 & ~n40273 ;
  assign n40364 = ~n40221 & ~n40235 ;
  assign n40365 = n40215 & n40364 ;
  assign n40366 = ~n40272 & ~n40347 ;
  assign n40367 = ~n40365 & n40366 ;
  assign n40368 = ~n40363 & ~n40367 ;
  assign n40369 = ~n40222 & n40243 ;
  assign n40370 = n40349 & n40369 ;
  assign n40371 = ~n40368 & ~n40370 ;
  assign n40372 = ~n40255 & ~n40371 ;
  assign n40361 = n40221 & n40260 ;
  assign n40362 = ~n40243 & n40361 ;
  assign n40373 = n40222 & ~n40235 ;
  assign n40374 = ~n40276 & ~n40373 ;
  assign n40375 = n40228 & n40243 ;
  assign n40376 = ~n40374 & n40375 ;
  assign n40377 = ~n40362 & ~n40376 ;
  assign n40378 = ~n40372 & n40377 ;
  assign n40379 = ~n40360 & n40378 ;
  assign n40380 = ~\u1_L6_reg[16]/NET0131  & ~n40379 ;
  assign n40381 = \u1_L6_reg[16]/NET0131  & n40379 ;
  assign n40382 = ~n40380 & ~n40381 ;
  assign n40383 = ~n40215 & n40221 ;
  assign n40384 = ~n40228 & ~n40235 ;
  assign n40396 = ~n40383 & ~n40384 ;
  assign n40397 = ~n40243 & ~n40396 ;
  assign n40395 = n40243 & ~n40384 ;
  assign n40398 = ~n40274 & ~n40395 ;
  assign n40399 = ~n40397 & n40398 ;
  assign n40403 = n40255 & ~n40399 ;
  assign n40400 = n40264 & n40384 ;
  assign n40390 = n40235 & n40354 ;
  assign n40401 = ~n40275 & ~n40390 ;
  assign n40402 = n40243 & ~n40401 ;
  assign n40404 = ~n40400 & ~n40402 ;
  assign n40405 = n40403 & n40404 ;
  assign n40406 = ~n40228 & n40274 ;
  assign n40407 = ~n40229 & ~n40406 ;
  assign n40408 = ~n40221 & n40237 ;
  assign n40409 = ~n40361 & ~n40408 ;
  assign n40410 = n40407 & n40409 ;
  assign n40411 = n40243 & ~n40410 ;
  assign n40412 = n40260 & n40383 ;
  assign n40413 = ~n40255 & ~n40412 ;
  assign n40414 = ~n40411 & n40413 ;
  assign n40415 = ~n40405 & ~n40414 ;
  assign n40387 = ~n40263 & n40384 ;
  assign n40388 = n40277 & ~n40387 ;
  assign n40389 = ~n40255 & ~n40388 ;
  assign n40391 = n40215 & n40390 ;
  assign n40392 = ~n40389 & ~n40391 ;
  assign n40393 = ~n40243 & ~n40392 ;
  assign n40385 = n40383 & n40384 ;
  assign n40386 = n40243 & n40385 ;
  assign n40394 = n40215 & n40259 ;
  assign n40416 = ~n40386 & ~n40394 ;
  assign n40417 = ~n40393 & n40416 ;
  assign n40418 = ~n40415 & n40417 ;
  assign n40419 = ~\u1_L6_reg[24]/NET0131  & ~n40418 ;
  assign n40420 = \u1_L6_reg[24]/NET0131  & n40418 ;
  assign n40421 = ~n40419 & ~n40420 ;
  assign n40441 = n40255 & ~n40385 ;
  assign n40442 = n40407 & n40441 ;
  assign n40438 = ~n40215 & n40245 ;
  assign n40437 = ~n40237 & n40354 ;
  assign n40439 = ~n40255 & ~n40437 ;
  assign n40440 = ~n40438 & n40439 ;
  assign n40443 = n40243 & ~n40440 ;
  assign n40444 = ~n40442 & n40443 ;
  assign n40422 = ~n40354 & ~n40364 ;
  assign n40423 = n40244 & n40422 ;
  assign n40424 = n40260 & n40274 ;
  assign n40425 = ~n40387 & ~n40424 ;
  assign n40426 = ~n40423 & n40425 ;
  assign n40427 = ~n40255 & ~n40426 ;
  assign n40428 = ~n40255 & ~n40262 ;
  assign n40429 = ~n40355 & n40428 ;
  assign n40430 = ~n40243 & n40262 ;
  assign n40431 = n40228 & ~n40430 ;
  assign n40432 = n40349 & n40431 ;
  assign n40433 = ~n40429 & n40432 ;
  assign n40434 = ~n40354 & ~n40408 ;
  assign n40435 = ~n40243 & n40255 ;
  assign n40436 = ~n40434 & n40435 ;
  assign n40445 = ~n40433 & ~n40436 ;
  assign n40446 = ~n40427 & n40445 ;
  assign n40447 = ~n40444 & n40446 ;
  assign n40448 = \u1_L6_reg[30]/NET0131  & ~n40447 ;
  assign n40449 = ~\u1_L6_reg[30]/NET0131  & n40447 ;
  assign n40450 = ~n40448 & ~n40449 ;
  assign n40451 = n39647 & ~n39680 ;
  assign n40452 = ~n39868 & n40451 ;
  assign n40453 = n39619 & ~n39632 ;
  assign n40454 = n40452 & ~n40453 ;
  assign n40455 = ~n39664 & n39861 ;
  assign n40456 = ~n39647 & ~n40455 ;
  assign n40457 = ~n39664 & ~n39864 ;
  assign n40458 = ~n39846 & ~n40457 ;
  assign n40459 = n40456 & n40458 ;
  assign n40460 = ~n40454 & ~n40459 ;
  assign n40461 = n39649 & n39861 ;
  assign n40462 = ~n39640 & ~n39685 ;
  assign n40463 = ~n40461 & n40462 ;
  assign n40464 = ~n40319 & n40463 ;
  assign n40465 = ~n40460 & n40464 ;
  assign n40467 = ~n39652 & ~n39839 ;
  assign n40468 = ~n39664 & ~n40467 ;
  assign n40469 = n40452 & ~n40468 ;
  assign n40470 = ~n39632 & n39864 ;
  assign n40471 = ~n39669 & ~n40470 ;
  assign n40472 = n40456 & n40471 ;
  assign n40473 = ~n40469 & ~n40472 ;
  assign n40466 = n39861 & n40330 ;
  assign n40474 = n40334 & ~n40466 ;
  assign n40475 = ~n40473 & n40474 ;
  assign n40476 = ~n40465 & ~n40475 ;
  assign n40477 = ~\u1_L6_reg[3]/NET0131  & n40476 ;
  assign n40478 = \u1_L6_reg[3]/NET0131  & ~n40476 ;
  assign n40479 = ~n40477 & ~n40478 ;
  assign n40482 = ~n39731 & n40133 ;
  assign n40483 = n39210 & ~n40482 ;
  assign n40484 = n39192 & n39733 ;
  assign n40480 = ~n39186 & ~n39743 ;
  assign n40481 = ~n39210 & ~n40480 ;
  assign n40485 = ~n39192 & n39241 ;
  assign n40486 = ~n40481 & ~n40485 ;
  assign n40487 = ~n40484 & n40486 ;
  assign n40488 = ~n40483 & n40487 ;
  assign n40489 = ~n39173 & ~n40488 ;
  assign n40490 = n39192 & n39743 ;
  assign n40491 = ~n40485 & ~n40490 ;
  assign n40492 = ~n39210 & ~n40491 ;
  assign n40494 = n39192 & ~n39236 ;
  assign n40495 = ~n39733 & n40494 ;
  assign n40493 = n39216 & ~n40480 ;
  assign n40496 = ~n39748 & ~n40493 ;
  assign n40497 = ~n40495 & n40496 ;
  assign n40498 = n39173 & ~n40497 ;
  assign n40499 = ~n40492 & ~n40498 ;
  assign n40500 = ~n40489 & n40499 ;
  assign n40501 = ~\u1_L6_reg[9]/NET0131  & ~n40500 ;
  assign n40502 = \u1_L6_reg[9]/NET0131  & n40500 ;
  assign n40503 = ~n40501 & ~n40502 ;
  assign n40505 = ~n39910 & ~n39916 ;
  assign n40507 = ~n39940 & n39977 ;
  assign n40508 = ~n40505 & ~n40507 ;
  assign n40509 = ~n39923 & ~n40508 ;
  assign n40504 = n39940 & n39975 ;
  assign n40506 = ~n39931 & n40505 ;
  assign n40510 = ~n39933 & ~n40506 ;
  assign n40511 = n40033 & n40510 ;
  assign n40512 = ~n40504 & n40511 ;
  assign n40513 = ~n40509 & n40512 ;
  assign n40517 = n39940 & ~n40029 ;
  assign n40514 = n39931 & n39962 ;
  assign n40515 = ~n39949 & ~n40514 ;
  assign n40516 = ~n39940 & ~n40515 ;
  assign n40518 = n39947 & ~n40058 ;
  assign n40519 = ~n40516 & n40518 ;
  assign n40520 = ~n40517 & n40519 ;
  assign n40521 = ~n40513 & ~n40520 ;
  assign n40522 = n39925 & n39931 ;
  assign n40523 = n39910 & n39956 ;
  assign n40524 = ~n40522 & ~n40523 ;
  assign n40525 = n39940 & ~n40524 ;
  assign n40526 = ~n39940 & n39957 ;
  assign n40527 = ~n40525 & ~n40526 ;
  assign n40528 = ~n40521 & n40527 ;
  assign n40529 = \u1_L6_reg[18]/NET0131  & n40528 ;
  assign n40530 = ~\u1_L6_reg[18]/NET0131  & ~n40528 ;
  assign n40531 = ~n40529 & ~n40530 ;
  assign n40579 = decrypt_pad & ~\u1_uk_K_r5_reg[33]/NET0131  ;
  assign n40580 = ~decrypt_pad & ~\u1_uk_K_r5_reg[11]/NET0131  ;
  assign n40581 = ~n40579 & ~n40580 ;
  assign n40582 = \u1_R5_reg[4]/NET0131  & ~n40581 ;
  assign n40583 = ~\u1_R5_reg[4]/NET0131  & n40581 ;
  assign n40584 = ~n40582 & ~n40583 ;
  assign n40532 = decrypt_pad & ~\u1_uk_K_r5_reg[55]/NET0131  ;
  assign n40533 = ~decrypt_pad & ~\u1_uk_K_r5_reg[33]/NET0131  ;
  assign n40534 = ~n40532 & ~n40533 ;
  assign n40535 = \u1_R5_reg[3]/NET0131  & ~n40534 ;
  assign n40536 = ~\u1_R5_reg[3]/NET0131  & n40534 ;
  assign n40537 = ~n40535 & ~n40536 ;
  assign n40552 = decrypt_pad & ~\u1_uk_K_r5_reg[46]/NET0131  ;
  assign n40553 = ~decrypt_pad & ~\u1_uk_K_r5_reg[24]/NET0131  ;
  assign n40554 = ~n40552 & ~n40553 ;
  assign n40555 = \u1_R5_reg[2]/NET0131  & ~n40554 ;
  assign n40556 = ~\u1_R5_reg[2]/NET0131  & n40554 ;
  assign n40557 = ~n40555 & ~n40556 ;
  assign n40538 = decrypt_pad & ~\u1_uk_K_r5_reg[6]/NET0131  ;
  assign n40539 = ~decrypt_pad & ~\u1_uk_K_r5_reg[41]/NET0131  ;
  assign n40540 = ~n40538 & ~n40539 ;
  assign n40541 = \u1_R5_reg[1]/NET0131  & ~n40540 ;
  assign n40542 = ~\u1_R5_reg[1]/NET0131  & n40540 ;
  assign n40543 = ~n40541 & ~n40542 ;
  assign n40545 = decrypt_pad & ~\u1_uk_K_r5_reg[4]/NET0131  ;
  assign n40546 = ~decrypt_pad & ~\u1_uk_K_r5_reg[39]/NET0131  ;
  assign n40547 = ~n40545 & ~n40546 ;
  assign n40548 = \u1_R5_reg[5]/NET0131  & ~n40547 ;
  assign n40549 = ~\u1_R5_reg[5]/NET0131  & n40547 ;
  assign n40550 = ~n40548 & ~n40549 ;
  assign n40551 = ~n40543 & ~n40550 ;
  assign n40560 = decrypt_pad & ~\u1_uk_K_r5_reg[10]/NET0131  ;
  assign n40561 = ~decrypt_pad & ~\u1_uk_K_r5_reg[20]/NET0131  ;
  assign n40562 = ~n40560 & ~n40561 ;
  assign n40563 = \u1_R5_reg[32]/NET0131  & ~n40562 ;
  assign n40564 = ~\u1_R5_reg[32]/NET0131  & n40562 ;
  assign n40565 = ~n40563 & ~n40564 ;
  assign n40592 = n40551 & n40565 ;
  assign n40593 = n40557 & n40592 ;
  assign n40567 = ~n40543 & n40550 ;
  assign n40594 = ~n40557 & ~n40565 ;
  assign n40595 = ~n40567 & n40594 ;
  assign n40596 = ~n40593 & ~n40595 ;
  assign n40597 = ~n40537 & ~n40596 ;
  assign n40586 = n40537 & n40557 ;
  assign n40587 = ~n40550 & ~n40565 ;
  assign n40588 = n40550 & n40565 ;
  assign n40589 = ~n40587 & ~n40588 ;
  assign n40590 = n40543 & n40589 ;
  assign n40591 = n40586 & n40590 ;
  assign n40544 = ~n40537 & n40543 ;
  assign n40598 = ~n40544 & n40588 ;
  assign n40599 = n40543 & n40587 ;
  assign n40600 = ~n40598 & ~n40599 ;
  assign n40601 = ~n40557 & ~n40600 ;
  assign n40602 = ~n40591 & ~n40601 ;
  assign n40603 = ~n40597 & n40602 ;
  assign n40604 = ~n40584 & ~n40603 ;
  assign n40568 = n40557 & ~n40565 ;
  assign n40569 = ~n40550 & n40568 ;
  assign n40570 = ~n40567 & ~n40569 ;
  assign n40571 = n40537 & ~n40570 ;
  assign n40558 = n40551 & ~n40557 ;
  assign n40559 = ~n40544 & ~n40558 ;
  assign n40566 = ~n40559 & n40565 ;
  assign n40572 = n40537 & ~n40557 ;
  assign n40573 = n40543 & ~n40572 ;
  assign n40574 = ~n40550 & ~n40557 ;
  assign n40575 = ~n40565 & ~n40574 ;
  assign n40576 = ~n40573 & n40575 ;
  assign n40577 = ~n40566 & ~n40576 ;
  assign n40578 = ~n40571 & n40577 ;
  assign n40585 = ~n40578 & n40584 ;
  assign n40609 = n40543 & n40588 ;
  assign n40610 = n40557 & n40609 ;
  assign n40611 = n40567 & n40568 ;
  assign n40612 = n40543 & n40574 ;
  assign n40613 = ~n40611 & ~n40612 ;
  assign n40614 = ~n40610 & n40613 ;
  assign n40615 = ~n40537 & ~n40614 ;
  assign n40605 = ~n40543 & n40586 ;
  assign n40606 = n40587 & n40605 ;
  assign n40607 = ~n40543 & n40565 ;
  assign n40608 = n40572 & n40607 ;
  assign n40616 = ~n40606 & ~n40608 ;
  assign n40617 = ~n40615 & n40616 ;
  assign n40618 = ~n40585 & n40617 ;
  assign n40619 = ~n40604 & n40618 ;
  assign n40620 = ~\u1_L5_reg[31]/NET0131  & ~n40619 ;
  assign n40621 = \u1_L5_reg[31]/NET0131  & n40619 ;
  assign n40622 = ~n40620 & ~n40621 ;
  assign n40670 = decrypt_pad & ~\u1_uk_K_r5_reg[2]/NET0131  ;
  assign n40671 = ~decrypt_pad & ~\u1_uk_K_r5_reg[37]/P0001  ;
  assign n40672 = ~n40670 & ~n40671 ;
  assign n40673 = \u1_R5_reg[24]/NET0131  & ~n40672 ;
  assign n40674 = ~\u1_R5_reg[24]/NET0131  & n40672 ;
  assign n40675 = ~n40673 & ~n40674 ;
  assign n40629 = decrypt_pad & ~\u1_uk_K_r5_reg[0]/NET0131  ;
  assign n40630 = ~decrypt_pad & ~\u1_uk_K_r5_reg[35]/NET0131  ;
  assign n40631 = ~n40629 & ~n40630 ;
  assign n40632 = \u1_R5_reg[23]/NET0131  & ~n40631 ;
  assign n40633 = ~\u1_R5_reg[23]/NET0131  & n40631 ;
  assign n40634 = ~n40632 & ~n40633 ;
  assign n40623 = decrypt_pad & ~\u1_uk_K_r5_reg[42]/NET0131  ;
  assign n40624 = ~decrypt_pad & ~\u1_uk_K_r5_reg[22]/NET0131  ;
  assign n40625 = ~n40623 & ~n40624 ;
  assign n40626 = \u1_R5_reg[22]/NET0131  & ~n40625 ;
  assign n40627 = ~\u1_R5_reg[22]/NET0131  & n40625 ;
  assign n40628 = ~n40626 & ~n40627 ;
  assign n40636 = decrypt_pad & ~\u1_uk_K_r5_reg[36]/NET0131  ;
  assign n40637 = ~decrypt_pad & ~\u1_uk_K_r5_reg[16]/NET0131  ;
  assign n40638 = ~n40636 & ~n40637 ;
  assign n40639 = \u1_R5_reg[20]/NET0131  & ~n40638 ;
  assign n40640 = ~\u1_R5_reg[20]/NET0131  & n40638 ;
  assign n40641 = ~n40639 & ~n40640 ;
  assign n40649 = decrypt_pad & ~\u1_uk_K_r5_reg[51]/NET0131  ;
  assign n40650 = ~decrypt_pad & ~\u1_uk_K_r5_reg[0]/NET0131  ;
  assign n40651 = ~n40649 & ~n40650 ;
  assign n40652 = \u1_R5_reg[21]/NET0131  & ~n40651 ;
  assign n40653 = ~\u1_R5_reg[21]/NET0131  & n40651 ;
  assign n40654 = ~n40652 & ~n40653 ;
  assign n40676 = ~n40641 & n40654 ;
  assign n40677 = n40628 & n40676 ;
  assign n40642 = decrypt_pad & ~\u1_uk_K_r5_reg[21]/NET0131  ;
  assign n40643 = ~decrypt_pad & ~\u1_uk_K_r5_reg[1]/NET0131  ;
  assign n40644 = ~n40642 & ~n40643 ;
  assign n40645 = \u1_R5_reg[25]/NET0131  & ~n40644 ;
  assign n40646 = ~\u1_R5_reg[25]/NET0131  & n40644 ;
  assign n40647 = ~n40645 & ~n40646 ;
  assign n40656 = ~n40647 & n40654 ;
  assign n40681 = n40641 & ~n40656 ;
  assign n40703 = ~n40628 & ~n40647 ;
  assign n40704 = ~n40654 & ~n40703 ;
  assign n40705 = n40681 & ~n40704 ;
  assign n40706 = ~n40677 & ~n40705 ;
  assign n40707 = n40634 & ~n40706 ;
  assign n40660 = ~n40641 & n40647 ;
  assign n40699 = n40654 & n40660 ;
  assign n40700 = ~n40628 & ~n40699 ;
  assign n40665 = n40641 & n40647 ;
  assign n40697 = ~n40665 & ~n40676 ;
  assign n40698 = n40628 & ~n40697 ;
  assign n40701 = ~n40634 & ~n40698 ;
  assign n40702 = ~n40700 & n40701 ;
  assign n40635 = ~n40628 & ~n40634 ;
  assign n40708 = n40635 & n40665 ;
  assign n40709 = ~n40654 & n40708 ;
  assign n40710 = ~n40702 & ~n40709 ;
  assign n40711 = ~n40707 & n40710 ;
  assign n40712 = n40675 & ~n40711 ;
  assign n40687 = n40641 & ~n40654 ;
  assign n40688 = n40628 & n40687 ;
  assign n40691 = n40647 & n40688 ;
  assign n40682 = ~n40634 & ~n40641 ;
  assign n40683 = ~n40628 & ~n40682 ;
  assign n40684 = ~n40681 & n40683 ;
  assign n40685 = n40641 & ~n40647 ;
  assign n40686 = n40635 & n40685 ;
  assign n40692 = ~n40684 & ~n40686 ;
  assign n40693 = ~n40691 & n40692 ;
  assign n40666 = ~n40628 & n40654 ;
  assign n40678 = n40641 & n40666 ;
  assign n40679 = ~n40677 & ~n40678 ;
  assign n40680 = ~n40634 & ~n40679 ;
  assign n40661 = ~n40654 & n40660 ;
  assign n40689 = ~n40661 & ~n40688 ;
  assign n40690 = n40634 & ~n40689 ;
  assign n40694 = ~n40680 & ~n40690 ;
  assign n40695 = n40693 & n40694 ;
  assign n40696 = ~n40675 & ~n40695 ;
  assign n40667 = ~n40665 & ~n40666 ;
  assign n40648 = ~n40641 & ~n40647 ;
  assign n40664 = ~n40628 & ~n40648 ;
  assign n40668 = n40634 & ~n40664 ;
  assign n40669 = ~n40667 & n40668 ;
  assign n40655 = n40648 & ~n40654 ;
  assign n40657 = n40641 & n40656 ;
  assign n40658 = ~n40655 & ~n40657 ;
  assign n40659 = n40635 & ~n40658 ;
  assign n40662 = ~n40628 & n40634 ;
  assign n40663 = n40661 & n40662 ;
  assign n40713 = ~n40659 & ~n40663 ;
  assign n40714 = ~n40669 & n40713 ;
  assign n40715 = ~n40696 & n40714 ;
  assign n40716 = ~n40712 & n40715 ;
  assign n40717 = ~\u1_L5_reg[11]/NET0131  & n40716 ;
  assign n40718 = \u1_L5_reg[11]/NET0131  & ~n40716 ;
  assign n40719 = ~n40717 & ~n40718 ;
  assign n40720 = decrypt_pad & ~\u1_uk_K_r5_reg[9]/NET0131  ;
  assign n40721 = ~decrypt_pad & ~\u1_uk_K_r5_reg[44]/NET0131  ;
  assign n40722 = ~n40720 & ~n40721 ;
  assign n40723 = \u1_R5_reg[28]/NET0131  & ~n40722 ;
  assign n40724 = ~\u1_R5_reg[28]/NET0131  & n40722 ;
  assign n40725 = ~n40723 & ~n40724 ;
  assign n40726 = decrypt_pad & ~\u1_uk_K_r5_reg[44]/NET0131  ;
  assign n40727 = ~decrypt_pad & ~\u1_uk_K_r5_reg[52]/NET0131  ;
  assign n40728 = ~n40726 & ~n40727 ;
  assign n40729 = \u1_R5_reg[26]/NET0131  & ~n40728 ;
  assign n40730 = ~\u1_R5_reg[26]/NET0131  & n40728 ;
  assign n40731 = ~n40729 & ~n40730 ;
  assign n40732 = decrypt_pad & ~\u1_uk_K_r5_reg[28]/NET0131  ;
  assign n40733 = ~decrypt_pad & ~\u1_uk_K_r5_reg[8]/NET0131  ;
  assign n40734 = ~n40732 & ~n40733 ;
  assign n40735 = \u1_R5_reg[25]/NET0131  & ~n40734 ;
  assign n40736 = ~\u1_R5_reg[25]/NET0131  & n40734 ;
  assign n40737 = ~n40735 & ~n40736 ;
  assign n40766 = ~n40731 & ~n40737 ;
  assign n40738 = decrypt_pad & ~\u1_uk_K_r5_reg[1]/NET0131  ;
  assign n40739 = ~decrypt_pad & ~\u1_uk_K_r5_reg[36]/NET0131  ;
  assign n40740 = ~n40738 & ~n40739 ;
  assign n40741 = \u1_R5_reg[29]/NET0131  & ~n40740 ;
  assign n40742 = ~\u1_R5_reg[29]/NET0131  & n40740 ;
  assign n40743 = ~n40741 & ~n40742 ;
  assign n40769 = ~n40731 & ~n40743 ;
  assign n40789 = ~n40766 & ~n40769 ;
  assign n40745 = decrypt_pad & ~\u1_uk_K_r5_reg[52]/NET0131  ;
  assign n40746 = ~decrypt_pad & ~\u1_uk_K_r5_reg[28]/NET0131  ;
  assign n40747 = ~n40745 & ~n40746 ;
  assign n40748 = \u1_R5_reg[24]/NET0131  & ~n40747 ;
  assign n40749 = ~\u1_R5_reg[24]/NET0131  & n40747 ;
  assign n40750 = ~n40748 & ~n40749 ;
  assign n40753 = decrypt_pad & ~\u1_uk_K_r5_reg[22]/NET0131  ;
  assign n40754 = ~decrypt_pad & ~\u1_uk_K_r5_reg[2]/NET0131  ;
  assign n40755 = ~n40753 & ~n40754 ;
  assign n40756 = \u1_R5_reg[27]/NET0131  & ~n40755 ;
  assign n40757 = ~\u1_R5_reg[27]/NET0131  & n40755 ;
  assign n40758 = ~n40756 & ~n40757 ;
  assign n40768 = n40731 & n40737 ;
  assign n40788 = n40758 & ~n40768 ;
  assign n40790 = n40750 & n40788 ;
  assign n40791 = n40789 & n40790 ;
  assign n40782 = n40743 & n40750 ;
  assign n40783 = n40766 & n40782 ;
  assign n40784 = n40737 & n40743 ;
  assign n40785 = ~n40750 & n40784 ;
  assign n40786 = ~n40783 & ~n40785 ;
  assign n40787 = ~n40758 & ~n40786 ;
  assign n40777 = ~n40743 & ~n40750 ;
  assign n40778 = n40766 & n40777 ;
  assign n40779 = n40743 & ~n40750 ;
  assign n40780 = n40731 & ~n40737 ;
  assign n40781 = n40779 & n40780 ;
  assign n40792 = ~n40778 & ~n40781 ;
  assign n40793 = ~n40787 & n40792 ;
  assign n40794 = ~n40791 & n40793 ;
  assign n40795 = n40725 & ~n40794 ;
  assign n40770 = ~n40758 & ~n40768 ;
  assign n40771 = ~n40769 & n40770 ;
  assign n40767 = n40758 & ~n40766 ;
  assign n40772 = n40750 & ~n40767 ;
  assign n40773 = ~n40771 & n40772 ;
  assign n40744 = ~n40737 & ~n40743 ;
  assign n40751 = n40744 & ~n40750 ;
  assign n40752 = n40731 & n40751 ;
  assign n40759 = n40752 & ~n40758 ;
  assign n40760 = ~n40731 & ~n40750 ;
  assign n40761 = n40731 & n40750 ;
  assign n40762 = ~n40760 & ~n40761 ;
  assign n40763 = ~n40737 & n40758 ;
  assign n40764 = n40743 & ~n40763 ;
  assign n40765 = ~n40762 & n40764 ;
  assign n40774 = ~n40759 & ~n40765 ;
  assign n40775 = ~n40773 & n40774 ;
  assign n40776 = ~n40725 & ~n40775 ;
  assign n40798 = n40768 & n40777 ;
  assign n40799 = ~n40781 & ~n40798 ;
  assign n40800 = ~n40743 & n40750 ;
  assign n40801 = ~n40737 & n40800 ;
  assign n40802 = n40799 & ~n40801 ;
  assign n40803 = n40758 & ~n40802 ;
  assign n40796 = n40737 & ~n40758 ;
  assign n40797 = ~n40762 & n40796 ;
  assign n40804 = n40763 & n40769 ;
  assign n40805 = ~n40797 & ~n40804 ;
  assign n40806 = ~n40803 & n40805 ;
  assign n40807 = ~n40776 & n40806 ;
  assign n40808 = ~n40795 & n40807 ;
  assign n40809 = ~\u1_L5_reg[22]/NET0131  & ~n40808 ;
  assign n40810 = \u1_L5_reg[22]/NET0131  & n40808 ;
  assign n40811 = ~n40809 & ~n40810 ;
  assign n40833 = ~n40543 & ~n40557 ;
  assign n40834 = ~n40565 & ~n40833 ;
  assign n40835 = n40588 & n40833 ;
  assign n40836 = ~n40834 & ~n40835 ;
  assign n40837 = n40537 & ~n40836 ;
  assign n40838 = ~n40557 & n40565 ;
  assign n40839 = ~n40537 & ~n40838 ;
  assign n40840 = ~n40834 & n40839 ;
  assign n40812 = n40543 & n40557 ;
  assign n40831 = n40550 & n40812 ;
  assign n40832 = n40565 & n40612 ;
  assign n40841 = ~n40831 & ~n40832 ;
  assign n40842 = ~n40840 & n40841 ;
  assign n40843 = ~n40837 & n40842 ;
  assign n40844 = n40584 & ~n40843 ;
  assign n40815 = ~n40543 & ~n40589 ;
  assign n40816 = ~n40550 & n40594 ;
  assign n40817 = ~n40815 & ~n40816 ;
  assign n40818 = ~n40537 & ~n40817 ;
  assign n40819 = ~n40592 & ~n40609 ;
  assign n40820 = n40537 & ~n40819 ;
  assign n40813 = ~n40550 & n40812 ;
  assign n40814 = n40565 & n40813 ;
  assign n40821 = ~n40611 & ~n40814 ;
  assign n40822 = ~n40820 & n40821 ;
  assign n40823 = ~n40818 & n40822 ;
  assign n40824 = ~n40584 & ~n40823 ;
  assign n40828 = n40557 & ~n40599 ;
  assign n40825 = n40550 & ~n40565 ;
  assign n40826 = n40543 & n40825 ;
  assign n40827 = ~n40557 & ~n40826 ;
  assign n40829 = n40537 & ~n40827 ;
  assign n40830 = ~n40828 & n40829 ;
  assign n40845 = ~n40824 & ~n40830 ;
  assign n40846 = ~n40844 & n40845 ;
  assign n40847 = ~\u1_L5_reg[17]/NET0131  & ~n40846 ;
  assign n40848 = \u1_L5_reg[17]/NET0131  & n40846 ;
  assign n40849 = ~n40847 & ~n40848 ;
  assign n40850 = decrypt_pad & ~\u1_uk_K_r5_reg[3]/NET0131  ;
  assign n40851 = ~decrypt_pad & ~\u1_uk_K_r5_reg[13]/P0001  ;
  assign n40852 = ~n40850 & ~n40851 ;
  assign n40853 = \u1_R5_reg[16]/NET0131  & ~n40852 ;
  assign n40854 = ~\u1_R5_reg[16]/NET0131  & n40852 ;
  assign n40855 = ~n40853 & ~n40854 ;
  assign n40862 = decrypt_pad & ~\u1_uk_K_r5_reg[18]/NET0131  ;
  assign n40863 = ~decrypt_pad & ~\u1_uk_K_r5_reg[53]/NET0131  ;
  assign n40864 = ~n40862 & ~n40863 ;
  assign n40865 = \u1_R5_reg[13]/NET0131  & ~n40864 ;
  assign n40866 = ~\u1_R5_reg[13]/NET0131  & n40864 ;
  assign n40867 = ~n40865 & ~n40866 ;
  assign n40856 = decrypt_pad & ~\u1_uk_K_r5_reg[27]/NET0131  ;
  assign n40857 = ~decrypt_pad & ~\u1_uk_K_r5_reg[5]/NET0131  ;
  assign n40858 = ~n40856 & ~n40857 ;
  assign n40859 = \u1_R5_reg[15]/NET0131  & ~n40858 ;
  assign n40860 = ~\u1_R5_reg[15]/NET0131  & n40858 ;
  assign n40861 = ~n40859 & ~n40860 ;
  assign n40869 = decrypt_pad & ~\u1_uk_K_r5_reg[24]/NET0131  ;
  assign n40870 = ~decrypt_pad & ~\u1_uk_K_r5_reg[34]/NET0131  ;
  assign n40871 = ~n40869 & ~n40870 ;
  assign n40872 = \u1_R5_reg[12]/NET0131  & ~n40871 ;
  assign n40873 = ~\u1_R5_reg[12]/NET0131  & n40871 ;
  assign n40874 = ~n40872 & ~n40873 ;
  assign n40875 = decrypt_pad & ~\u1_uk_K_r5_reg[40]/NET0131  ;
  assign n40876 = ~decrypt_pad & ~\u1_uk_K_r5_reg[18]/NET0131  ;
  assign n40877 = ~n40875 & ~n40876 ;
  assign n40878 = \u1_R5_reg[17]/NET0131  & ~n40877 ;
  assign n40879 = ~\u1_R5_reg[17]/NET0131  & n40877 ;
  assign n40880 = ~n40878 & ~n40879 ;
  assign n40918 = ~n40874 & n40880 ;
  assign n40923 = n40861 & n40918 ;
  assign n40924 = ~n40867 & n40923 ;
  assign n40882 = decrypt_pad & ~\u1_uk_K_r5_reg[19]/NET0131  ;
  assign n40883 = ~decrypt_pad & ~\u1_uk_K_r5_reg[54]/NET0131  ;
  assign n40884 = ~n40882 & ~n40883 ;
  assign n40885 = \u1_R5_reg[14]/NET0131  & ~n40884 ;
  assign n40886 = ~\u1_R5_reg[14]/NET0131  & n40884 ;
  assign n40887 = ~n40885 & ~n40886 ;
  assign n40917 = ~n40861 & ~n40887 ;
  assign n40897 = ~n40867 & n40874 ;
  assign n40902 = n40867 & ~n40874 ;
  assign n40921 = ~n40897 & ~n40902 ;
  assign n40922 = n40917 & ~n40921 ;
  assign n40868 = n40861 & n40867 ;
  assign n40881 = n40874 & ~n40880 ;
  assign n40935 = n40868 & n40881 ;
  assign n40936 = ~n40922 & ~n40935 ;
  assign n40937 = ~n40924 & n40936 ;
  assign n40925 = n40874 & n40880 ;
  assign n40926 = n40887 & n40925 ;
  assign n40927 = n40867 & n40926 ;
  assign n40928 = n40867 & ~n40887 ;
  assign n40929 = n40880 & n40928 ;
  assign n40930 = ~n40874 & n40929 ;
  assign n40931 = ~n40927 & ~n40930 ;
  assign n40913 = ~n40867 & n40887 ;
  assign n40932 = ~n40874 & n40913 ;
  assign n40933 = ~n40880 & n40932 ;
  assign n40934 = ~n40861 & n40933 ;
  assign n40938 = n40931 & ~n40934 ;
  assign n40939 = n40937 & n40938 ;
  assign n40940 = n40855 & ~n40939 ;
  assign n40903 = ~n40880 & n40902 ;
  assign n40904 = n40887 & n40903 ;
  assign n40898 = ~n40887 & n40897 ;
  assign n40899 = n40880 & n40898 ;
  assign n40895 = ~n40867 & ~n40880 ;
  assign n40900 = ~n40874 & n40895 ;
  assign n40901 = n40861 & n40900 ;
  assign n40906 = ~n40899 & ~n40901 ;
  assign n40907 = ~n40904 & n40906 ;
  assign n40891 = ~n40867 & n40880 ;
  assign n40892 = n40881 & n40887 ;
  assign n40893 = ~n40891 & ~n40892 ;
  assign n40894 = ~n40861 & ~n40893 ;
  assign n40888 = ~n40874 & ~n40887 ;
  assign n40889 = n40868 & ~n40881 ;
  assign n40890 = ~n40888 & n40889 ;
  assign n40896 = n40888 & n40895 ;
  assign n40905 = ~n40890 & ~n40896 ;
  assign n40908 = ~n40894 & n40905 ;
  assign n40909 = n40907 & n40908 ;
  assign n40910 = ~n40855 & ~n40909 ;
  assign n40914 = n40881 & n40913 ;
  assign n40915 = ~n40896 & ~n40914 ;
  assign n40916 = n40861 & ~n40915 ;
  assign n40911 = n40881 & ~n40887 ;
  assign n40912 = n40868 & n40911 ;
  assign n40919 = n40867 & n40918 ;
  assign n40920 = n40917 & n40919 ;
  assign n40941 = ~n40912 & ~n40920 ;
  assign n40942 = ~n40916 & n40941 ;
  assign n40943 = ~n40910 & n40942 ;
  assign n40944 = ~n40940 & n40943 ;
  assign n40945 = ~\u1_L5_reg[20]/NET0131  & ~n40944 ;
  assign n40946 = \u1_L5_reg[20]/NET0131  & n40944 ;
  assign n40947 = ~n40945 & ~n40946 ;
  assign n40966 = decrypt_pad & ~\u1_uk_K_r5_reg[17]/NET0131  ;
  assign n40967 = ~decrypt_pad & ~\u1_uk_K_r5_reg[27]/NET0131  ;
  assign n40968 = ~n40966 & ~n40967 ;
  assign n40969 = \u1_R5_reg[6]/NET0131  & ~n40968 ;
  assign n40970 = ~\u1_R5_reg[6]/NET0131  & n40968 ;
  assign n40971 = ~n40969 & ~n40970 ;
  assign n40954 = decrypt_pad & ~\u1_uk_K_r5_reg[39]/NET0131  ;
  assign n40955 = ~decrypt_pad & ~\u1_uk_K_r5_reg[17]/NET0131  ;
  assign n40956 = ~n40954 & ~n40955 ;
  assign n40957 = \u1_R5_reg[9]/NET0131  & ~n40956 ;
  assign n40958 = ~\u1_R5_reg[9]/NET0131  & n40956 ;
  assign n40959 = ~n40957 & ~n40958 ;
  assign n40960 = decrypt_pad & ~\u1_uk_K_r5_reg[26]/NET0131  ;
  assign n40961 = ~decrypt_pad & ~\u1_uk_K_r5_reg[4]/NET0131  ;
  assign n40962 = ~n40960 & ~n40961 ;
  assign n40963 = \u1_R5_reg[5]/NET0131  & ~n40962 ;
  assign n40964 = ~\u1_R5_reg[5]/NET0131  & n40962 ;
  assign n40965 = ~n40963 & ~n40964 ;
  assign n40985 = ~n40959 & n40965 ;
  assign n40973 = decrypt_pad & ~\u1_uk_K_r5_reg[47]/NET0131  ;
  assign n40974 = ~decrypt_pad & ~\u1_uk_K_r5_reg[25]/NET0131  ;
  assign n40975 = ~n40973 & ~n40974 ;
  assign n40976 = \u1_R5_reg[4]/NET0131  & ~n40975 ;
  assign n40977 = ~\u1_R5_reg[4]/NET0131  & n40975 ;
  assign n40978 = ~n40976 & ~n40977 ;
  assign n40986 = n40959 & ~n40965 ;
  assign n40987 = ~n40978 & n40986 ;
  assign n40988 = ~n40985 & ~n40987 ;
  assign n40989 = ~n40971 & ~n40988 ;
  assign n40948 = decrypt_pad & ~\u1_uk_K_r5_reg[11]/NET0131  ;
  assign n40949 = ~decrypt_pad & ~\u1_uk_K_r5_reg[46]/NET0131  ;
  assign n40950 = ~n40948 & ~n40949 ;
  assign n40951 = \u1_R5_reg[7]/NET0131  & ~n40950 ;
  assign n40952 = ~\u1_R5_reg[7]/NET0131  & n40950 ;
  assign n40953 = ~n40951 & ~n40952 ;
  assign n40998 = n40971 & n40978 ;
  assign n40999 = n40953 & n40998 ;
  assign n41000 = n40986 & n40999 ;
  assign n41004 = decrypt_pad & ~\u1_uk_K_r5_reg[34]/NET0131  ;
  assign n41005 = ~decrypt_pad & ~\u1_uk_K_r5_reg[12]/P0001  ;
  assign n41006 = ~n41004 & ~n41005 ;
  assign n41007 = \u1_R5_reg[8]/NET0131  & ~n41006 ;
  assign n41008 = ~\u1_R5_reg[8]/NET0131  & n41006 ;
  assign n41009 = ~n41007 & ~n41008 ;
  assign n41010 = ~n41000 & ~n41009 ;
  assign n41011 = ~n40989 & n41010 ;
  assign n40992 = n40959 & ~n40978 ;
  assign n40993 = n40965 & n40992 ;
  assign n40994 = n40971 & ~n40993 ;
  assign n40990 = ~n40953 & ~n40965 ;
  assign n40991 = ~n40971 & ~n40990 ;
  assign n40995 = ~n40959 & ~n40971 ;
  assign n40996 = ~n40991 & ~n40995 ;
  assign n40997 = ~n40994 & n40996 ;
  assign n41001 = ~n40986 & n40998 ;
  assign n41002 = ~n40987 & ~n41001 ;
  assign n41003 = ~n40953 & ~n41002 ;
  assign n41012 = ~n40997 & ~n41003 ;
  assign n41013 = n41011 & n41012 ;
  assign n41021 = ~n40971 & n40978 ;
  assign n41022 = n40959 & n41021 ;
  assign n41023 = n40971 & ~n40978 ;
  assign n41024 = n40953 & ~n41023 ;
  assign n41025 = ~n41022 & ~n41024 ;
  assign n41026 = n40965 & ~n41025 ;
  assign n40972 = ~n40965 & n40971 ;
  assign n41017 = n40959 & ~n40972 ;
  assign n41015 = ~n40953 & n40971 ;
  assign n41016 = ~n40990 & ~n41015 ;
  assign n41014 = ~n40959 & n40978 ;
  assign n41018 = ~n40992 & ~n41014 ;
  assign n41019 = ~n41016 & n41018 ;
  assign n41020 = ~n41017 & n41019 ;
  assign n41027 = ~n40965 & n40995 ;
  assign n41028 = n40978 & n41027 ;
  assign n41029 = n41009 & ~n41028 ;
  assign n41030 = ~n41020 & n41029 ;
  assign n41031 = ~n41026 & n41030 ;
  assign n41032 = ~n41013 & ~n41031 ;
  assign n40979 = n40972 & ~n40978 ;
  assign n40980 = ~n40959 & n40979 ;
  assign n40981 = n40965 & n40978 ;
  assign n40982 = ~n40971 & n40981 ;
  assign n40983 = ~n40980 & ~n40982 ;
  assign n40984 = n40953 & ~n40983 ;
  assign n41033 = ~n40972 & ~n40978 ;
  assign n41034 = n40959 & ~n41016 ;
  assign n41035 = n41033 & n41034 ;
  assign n41036 = ~n40984 & ~n41035 ;
  assign n41037 = ~n41032 & n41036 ;
  assign n41038 = \u1_L5_reg[2]/NET0131  & n41037 ;
  assign n41039 = ~\u1_L5_reg[2]/NET0131  & ~n41037 ;
  assign n41040 = ~n41038 & ~n41039 ;
  assign n41045 = n40654 & n40665 ;
  assign n41046 = ~n40654 & n40685 ;
  assign n41047 = ~n41045 & ~n41046 ;
  assign n41048 = n40628 & ~n40676 ;
  assign n41049 = ~n40647 & ~n40666 ;
  assign n41050 = ~n41048 & n41049 ;
  assign n41051 = n41047 & ~n41050 ;
  assign n41052 = n40634 & ~n41051 ;
  assign n41041 = n40628 & n40657 ;
  assign n41042 = ~n40628 & ~n40697 ;
  assign n41043 = ~n41041 & ~n41042 ;
  assign n41044 = ~n40634 & ~n41043 ;
  assign n41053 = n40628 & n40661 ;
  assign n41054 = ~n41044 & ~n41053 ;
  assign n41055 = ~n41052 & n41054 ;
  assign n41056 = ~n40675 & ~n41055 ;
  assign n41059 = n40628 & ~n40647 ;
  assign n41060 = n40676 & ~n41059 ;
  assign n41061 = ~n41041 & ~n41060 ;
  assign n41062 = n40634 & ~n41061 ;
  assign n41064 = n40628 & ~n40648 ;
  assign n41065 = ~n40665 & n41064 ;
  assign n41063 = n40634 & ~n40704 ;
  assign n41066 = ~n41042 & ~n41063 ;
  assign n41067 = ~n41065 & n41066 ;
  assign n41068 = ~n41062 & ~n41067 ;
  assign n41069 = n40675 & ~n41068 ;
  assign n41057 = n40634 & n40647 ;
  assign n41058 = n40666 & n41057 ;
  assign n41070 = ~n40628 & n41046 ;
  assign n41071 = ~n41058 & ~n41070 ;
  assign n41072 = ~n41069 & n41071 ;
  assign n41073 = ~n41056 & n41072 ;
  assign n41074 = \u1_L5_reg[29]/NET0131  & ~n41073 ;
  assign n41075 = ~\u1_L5_reg[29]/NET0131  & n41073 ;
  assign n41076 = ~n41074 & ~n41075 ;
  assign n41077 = decrypt_pad & ~\u1_uk_K_r5_reg[35]/NET0131  ;
  assign n41078 = ~decrypt_pad & ~\u1_uk_K_r5_reg[15]/NET0131  ;
  assign n41079 = ~n41077 & ~n41078 ;
  assign n41080 = \u1_R5_reg[30]/NET0131  & ~n41079 ;
  assign n41081 = ~\u1_R5_reg[30]/NET0131  & n41079 ;
  assign n41082 = ~n41080 & ~n41081 ;
  assign n41083 = decrypt_pad & ~\u1_uk_K_r5_reg[38]/NET0131  ;
  assign n41084 = ~decrypt_pad & ~\u1_uk_K_r5_reg[14]/NET0131  ;
  assign n41085 = ~n41083 & ~n41084 ;
  assign n41086 = \u1_R5_reg[29]/NET0131  & ~n41085 ;
  assign n41087 = ~\u1_R5_reg[29]/NET0131  & n41085 ;
  assign n41088 = ~n41086 & ~n41087 ;
  assign n41089 = decrypt_pad & ~\u1_uk_K_r5_reg[50]/NET0131  ;
  assign n41090 = ~decrypt_pad & ~\u1_uk_K_r5_reg[30]/NET0131  ;
  assign n41091 = ~n41089 & ~n41090 ;
  assign n41092 = \u1_R5_reg[1]/NET0131  & ~n41091 ;
  assign n41093 = ~\u1_R5_reg[1]/NET0131  & n41091 ;
  assign n41094 = ~n41092 & ~n41093 ;
  assign n41095 = n41088 & n41094 ;
  assign n41096 = decrypt_pad & ~\u1_uk_K_r5_reg[7]/NET0131  ;
  assign n41097 = ~decrypt_pad & ~\u1_uk_K_r5_reg[42]/NET0131  ;
  assign n41098 = ~n41096 & ~n41097 ;
  assign n41099 = \u1_R5_reg[28]/NET0131  & ~n41098 ;
  assign n41100 = ~\u1_R5_reg[28]/NET0131  & n41098 ;
  assign n41101 = ~n41099 & ~n41100 ;
  assign n41102 = n41095 & ~n41101 ;
  assign n41103 = n41082 & n41102 ;
  assign n41104 = ~n41082 & n41101 ;
  assign n41105 = n41088 & ~n41094 ;
  assign n41106 = ~n41104 & ~n41105 ;
  assign n41107 = ~n41094 & n41104 ;
  assign n41108 = n41088 & n41107 ;
  assign n41109 = ~n41106 & ~n41108 ;
  assign n41110 = decrypt_pad & ~\u1_uk_K_r5_reg[23]/NET0131  ;
  assign n41111 = ~decrypt_pad & ~\u1_uk_K_r5_reg[31]/NET0131  ;
  assign n41112 = ~n41110 & ~n41111 ;
  assign n41113 = \u1_R5_reg[31]/P0001  & ~n41112 ;
  assign n41114 = ~\u1_R5_reg[31]/P0001  & n41112 ;
  assign n41115 = ~n41113 & ~n41114 ;
  assign n41116 = ~n41109 & n41115 ;
  assign n41117 = ~n41082 & ~n41088 ;
  assign n41118 = ~n41101 & n41117 ;
  assign n41119 = ~n41088 & n41101 ;
  assign n41120 = n41082 & n41119 ;
  assign n41121 = ~n41115 & ~n41120 ;
  assign n41122 = ~n41118 & n41121 ;
  assign n41123 = ~n41116 & ~n41122 ;
  assign n41124 = ~n41103 & ~n41123 ;
  assign n41125 = decrypt_pad & ~\u1_uk_K_r5_reg[29]/NET0131  ;
  assign n41126 = ~decrypt_pad & ~\u1_uk_K_r5_reg[9]/NET0131  ;
  assign n41127 = ~n41125 & ~n41126 ;
  assign n41128 = \u1_R5_reg[32]/NET0131  & ~n41127 ;
  assign n41129 = ~\u1_R5_reg[32]/NET0131  & n41127 ;
  assign n41130 = ~n41128 & ~n41129 ;
  assign n41131 = ~n41124 & n41130 ;
  assign n41147 = ~n41094 & n41120 ;
  assign n41139 = n41094 & ~n41101 ;
  assign n41140 = ~n41088 & n41139 ;
  assign n41148 = n41115 & ~n41140 ;
  assign n41149 = ~n41147 & n41148 ;
  assign n41134 = n41082 & ~n41094 ;
  assign n41135 = ~n41101 & n41134 ;
  assign n41150 = ~n41095 & ~n41115 ;
  assign n41151 = ~n41135 & n41150 ;
  assign n41152 = ~n41149 & ~n41151 ;
  assign n41153 = n41088 & n41101 ;
  assign n41154 = n41082 & n41153 ;
  assign n41155 = n41094 & n41154 ;
  assign n41132 = n41104 & ~n41115 ;
  assign n41156 = ~n41108 & ~n41132 ;
  assign n41157 = ~n41155 & n41156 ;
  assign n41158 = ~n41152 & n41157 ;
  assign n41159 = ~n41130 & ~n41158 ;
  assign n41133 = n41105 & n41132 ;
  assign n41136 = n41088 & n41135 ;
  assign n41137 = ~n41094 & n41118 ;
  assign n41138 = ~n41136 & ~n41137 ;
  assign n41141 = n41082 & n41140 ;
  assign n41142 = ~n41088 & n41094 ;
  assign n41143 = n41104 & n41142 ;
  assign n41144 = ~n41141 & ~n41143 ;
  assign n41145 = n41138 & n41144 ;
  assign n41146 = n41115 & ~n41145 ;
  assign n41160 = ~n41133 & ~n41146 ;
  assign n41161 = ~n41159 & n41160 ;
  assign n41162 = ~n41131 & n41161 ;
  assign n41163 = \u1_L5_reg[5]/NET0131  & ~n41162 ;
  assign n41164 = ~\u1_L5_reg[5]/NET0131  & n41162 ;
  assign n41165 = ~n41163 & ~n41164 ;
  assign n41182 = n40648 & n40654 ;
  assign n41183 = ~n41053 & ~n41182 ;
  assign n41184 = ~n40634 & ~n41183 ;
  assign n41185 = ~n40708 & ~n41070 ;
  assign n41186 = ~n41184 & n41185 ;
  assign n41187 = ~n40675 & ~n41186 ;
  assign n41173 = ~n40655 & ~n40699 ;
  assign n41174 = ~n40657 & n41173 ;
  assign n41175 = n40628 & ~n41174 ;
  assign n41176 = ~n40628 & n40660 ;
  assign n41177 = ~n40657 & ~n41176 ;
  assign n41178 = ~n40691 & n41177 ;
  assign n41179 = ~n40675 & ~n41178 ;
  assign n41180 = ~n41175 & ~n41179 ;
  assign n41181 = n40634 & ~n41180 ;
  assign n41168 = n40654 & ~n41059 ;
  assign n41169 = ~n40664 & n41168 ;
  assign n41166 = n40635 & ~n40681 ;
  assign n41167 = n40662 & n40665 ;
  assign n41170 = ~n41166 & ~n41167 ;
  assign n41171 = ~n41169 & n41170 ;
  assign n41172 = n40675 & ~n41171 ;
  assign n41188 = n40628 & n41047 ;
  assign n41189 = ~n40634 & ~n40664 ;
  assign n41190 = ~n41188 & n41189 ;
  assign n41191 = ~n41172 & ~n41190 ;
  assign n41192 = ~n41181 & n41191 ;
  assign n41193 = ~n41187 & n41192 ;
  assign n41194 = ~\u1_L5_reg[4]/NET0131  & ~n41193 ;
  assign n41195 = \u1_L5_reg[4]/NET0131  & n41193 ;
  assign n41196 = ~n41194 & ~n41195 ;
  assign n41215 = ~n40899 & ~n40903 ;
  assign n41216 = n40861 & ~n41215 ;
  assign n41210 = n40880 & n40932 ;
  assign n41211 = ~n40927 & ~n41210 ;
  assign n41217 = ~n40881 & ~n40929 ;
  assign n41203 = n40874 & n40928 ;
  assign n41218 = ~n40861 & ~n41203 ;
  assign n41219 = ~n41217 & n41218 ;
  assign n41220 = n41211 & ~n41219 ;
  assign n41221 = ~n41216 & n41220 ;
  assign n41222 = n40855 & ~n41221 ;
  assign n41197 = n40861 & n40887 ;
  assign n41198 = ~n40900 & ~n40923 ;
  assign n41199 = ~n41197 & ~n41198 ;
  assign n41200 = ~n40895 & ~n40913 ;
  assign n41201 = n40861 & n40874 ;
  assign n41202 = ~n41200 & n41201 ;
  assign n41204 = n40917 & n40925 ;
  assign n41205 = ~n41203 & ~n41204 ;
  assign n41206 = ~n40904 & n41205 ;
  assign n41207 = ~n41202 & n41206 ;
  assign n41208 = ~n41199 & n41207 ;
  assign n41209 = ~n40855 & ~n41208 ;
  assign n41212 = ~n40896 & n41211 ;
  assign n41213 = ~n40861 & ~n41212 ;
  assign n41214 = n40902 & n41197 ;
  assign n41223 = ~n40912 & ~n41214 ;
  assign n41224 = ~n41213 & n41223 ;
  assign n41225 = ~n41209 & n41224 ;
  assign n41226 = ~n41222 & n41225 ;
  assign n41227 = ~\u1_L5_reg[10]/NET0131  & ~n41226 ;
  assign n41228 = \u1_L5_reg[10]/NET0131  & n41226 ;
  assign n41229 = ~n41227 & ~n41228 ;
  assign n41236 = ~n40766 & ~n40768 ;
  assign n41237 = n40777 & n41236 ;
  assign n41234 = ~n40763 & ~n40768 ;
  assign n41235 = n40779 & ~n41234 ;
  assign n41241 = ~n40725 & ~n41235 ;
  assign n41242 = ~n41237 & n41241 ;
  assign n41230 = n40750 & n40769 ;
  assign n41231 = n40743 & n40761 ;
  assign n41232 = ~n41230 & ~n41231 ;
  assign n41233 = ~n40737 & ~n41232 ;
  assign n41238 = ~n40744 & ~n40784 ;
  assign n41239 = ~n40761 & n41238 ;
  assign n41240 = ~n40758 & ~n41239 ;
  assign n41243 = ~n41233 & ~n41240 ;
  assign n41244 = n41242 & n41243 ;
  assign n41245 = ~n40758 & n40781 ;
  assign n41251 = n40725 & ~n40783 ;
  assign n41252 = ~n40798 & n41251 ;
  assign n41253 = ~n41245 & n41252 ;
  assign n41246 = ~n40760 & ~n40801 ;
  assign n41247 = n40789 & ~n41246 ;
  assign n41248 = n40737 & n40750 ;
  assign n41249 = ~n40778 & ~n41248 ;
  assign n41250 = n40758 & ~n41249 ;
  assign n41254 = ~n41247 & ~n41250 ;
  assign n41255 = n41253 & n41254 ;
  assign n41256 = ~n41244 & ~n41255 ;
  assign n41257 = \u1_L5_reg[12]/NET0131  & n41256 ;
  assign n41258 = ~\u1_L5_reg[12]/NET0131  & ~n41256 ;
  assign n41259 = ~n41257 & ~n41258 ;
  assign n41260 = ~n40959 & n41021 ;
  assign n41261 = ~n40985 & ~n41260 ;
  assign n41262 = ~n40981 & ~n41261 ;
  assign n41263 = n40959 & n40979 ;
  assign n41264 = ~n41262 & ~n41263 ;
  assign n41265 = ~n41009 & ~n41264 ;
  assign n41266 = n40985 & n40998 ;
  assign n41267 = n40959 & n40982 ;
  assign n41268 = ~n41266 & ~n41267 ;
  assign n41269 = ~n41265 & n41268 ;
  assign n41270 = ~n40953 & ~n41269 ;
  assign n41271 = ~n40965 & ~n40992 ;
  assign n41272 = ~n41014 & n41271 ;
  assign n41273 = n40965 & n41260 ;
  assign n41274 = ~n41272 & ~n41273 ;
  assign n41275 = n40953 & ~n41274 ;
  assign n41277 = n40991 & n40992 ;
  assign n41276 = ~n40985 & n40999 ;
  assign n41278 = ~n41009 & ~n41276 ;
  assign n41279 = ~n41277 & n41278 ;
  assign n41280 = ~n41275 & n41279 ;
  assign n41281 = ~n40995 & n41271 ;
  assign n41282 = ~n40953 & ~n41281 ;
  assign n41283 = n40959 & n41023 ;
  assign n41284 = n40953 & ~n41027 ;
  assign n41285 = ~n41283 & n41284 ;
  assign n41286 = ~n41282 & ~n41285 ;
  assign n41287 = ~n40978 & n40995 ;
  assign n41288 = n40965 & n41287 ;
  assign n41289 = n41009 & ~n41288 ;
  assign n41290 = ~n40997 & n41289 ;
  assign n41291 = n41268 & n41290 ;
  assign n41292 = ~n41286 & n41291 ;
  assign n41293 = ~n41280 & ~n41292 ;
  assign n41294 = ~n41270 & ~n41293 ;
  assign n41295 = ~\u1_L5_reg[13]/NET0131  & n41294 ;
  assign n41296 = \u1_L5_reg[13]/NET0131  & ~n41294 ;
  assign n41297 = ~n41295 & ~n41296 ;
  assign n41298 = decrypt_pad & ~\u1_uk_K_r5_reg[30]/NET0131  ;
  assign n41299 = ~decrypt_pad & ~\u1_uk_K_r5_reg[38]/NET0131  ;
  assign n41300 = ~n41298 & ~n41299 ;
  assign n41301 = \u1_R5_reg[19]/NET0131  & ~n41300 ;
  assign n41302 = ~\u1_R5_reg[19]/NET0131  & n41300 ;
  assign n41303 = ~n41301 & ~n41302 ;
  assign n41304 = decrypt_pad & ~\u1_uk_K_r5_reg[43]/NET0131  ;
  assign n41305 = ~decrypt_pad & ~\u1_uk_K_r5_reg[23]/NET0131  ;
  assign n41306 = ~n41304 & ~n41305 ;
  assign n41307 = \u1_R5_reg[18]/NET0131  & ~n41306 ;
  assign n41308 = ~\u1_R5_reg[18]/NET0131  & n41306 ;
  assign n41309 = ~n41307 & ~n41308 ;
  assign n41310 = decrypt_pad & ~\u1_uk_K_r5_reg[49]/NET0131  ;
  assign n41311 = ~decrypt_pad & ~\u1_uk_K_r5_reg[29]/NET0131  ;
  assign n41312 = ~n41310 & ~n41311 ;
  assign n41313 = \u1_R5_reg[17]/NET0131  & ~n41312 ;
  assign n41314 = ~\u1_R5_reg[17]/NET0131  & n41312 ;
  assign n41315 = ~n41313 & ~n41314 ;
  assign n41316 = ~n41309 & n41315 ;
  assign n41317 = decrypt_pad & ~\u1_uk_K_r5_reg[15]/NET0131  ;
  assign n41318 = ~decrypt_pad & ~\u1_uk_K_r5_reg[50]/NET0131  ;
  assign n41319 = ~n41317 & ~n41318 ;
  assign n41320 = \u1_R5_reg[21]/NET0131  & ~n41319 ;
  assign n41321 = ~\u1_R5_reg[21]/NET0131  & n41319 ;
  assign n41322 = ~n41320 & ~n41321 ;
  assign n41323 = n41316 & n41322 ;
  assign n41324 = decrypt_pad & ~\u1_uk_K_r5_reg[31]/NET0131  ;
  assign n41325 = ~decrypt_pad & ~\u1_uk_K_r5_reg[7]/NET0131  ;
  assign n41326 = ~n41324 & ~n41325 ;
  assign n41327 = \u1_R5_reg[16]/NET0131  & ~n41326 ;
  assign n41328 = ~\u1_R5_reg[16]/NET0131  & n41326 ;
  assign n41329 = ~n41327 & ~n41328 ;
  assign n41330 = n41323 & n41329 ;
  assign n41336 = n41322 & ~n41329 ;
  assign n41337 = ~n41315 & n41336 ;
  assign n41331 = n41315 & ~n41322 ;
  assign n41332 = n41309 & n41331 ;
  assign n41333 = ~n41322 & n41329 ;
  assign n41334 = ~n41309 & ~n41315 ;
  assign n41335 = n41333 & n41334 ;
  assign n41338 = ~n41332 & ~n41335 ;
  assign n41339 = ~n41337 & n41338 ;
  assign n41340 = ~n41330 & n41339 ;
  assign n41341 = ~n41303 & ~n41340 ;
  assign n41349 = n41309 & n41322 ;
  assign n41350 = n41329 & n41349 ;
  assign n41345 = n41316 & ~n41329 ;
  assign n41347 = ~n41322 & ~n41329 ;
  assign n41348 = ~n41315 & n41347 ;
  assign n41351 = ~n41345 & ~n41348 ;
  assign n41352 = ~n41350 & n41351 ;
  assign n41353 = n41303 & ~n41352 ;
  assign n41342 = n41322 & n41329 ;
  assign n41343 = n41309 & ~n41315 ;
  assign n41344 = n41342 & n41343 ;
  assign n41346 = ~n41322 & n41345 ;
  assign n41354 = ~n41344 & ~n41346 ;
  assign n41355 = ~n41353 & n41354 ;
  assign n41356 = ~n41341 & n41355 ;
  assign n41357 = decrypt_pad & ~\u1_uk_K_r5_reg[14]/NET0131  ;
  assign n41358 = ~decrypt_pad & ~\u1_uk_K_r5_reg[49]/NET0131  ;
  assign n41359 = ~n41357 & ~n41358 ;
  assign n41360 = \u1_R5_reg[20]/NET0131  & ~n41359 ;
  assign n41361 = ~\u1_R5_reg[20]/NET0131  & n41359 ;
  assign n41362 = ~n41360 & ~n41361 ;
  assign n41363 = ~n41356 & ~n41362 ;
  assign n41366 = ~n41309 & n41342 ;
  assign n41369 = ~n41337 & ~n41366 ;
  assign n41367 = n41329 & n41331 ;
  assign n41368 = n41309 & n41336 ;
  assign n41370 = ~n41367 & ~n41368 ;
  assign n41371 = n41369 & n41370 ;
  assign n41372 = n41303 & ~n41371 ;
  assign n41373 = ~n41303 & ~n41309 ;
  assign n41374 = n41315 & n41336 ;
  assign n41375 = ~n41348 & ~n41374 ;
  assign n41376 = n41373 & ~n41375 ;
  assign n41364 = ~n41316 & ~n41343 ;
  assign n41365 = n41333 & ~n41364 ;
  assign n41377 = n41303 & n41309 ;
  assign n41378 = n41342 & ~n41377 ;
  assign n41379 = n41364 & n41378 ;
  assign n41380 = ~n41365 & ~n41379 ;
  assign n41381 = ~n41376 & n41380 ;
  assign n41382 = ~n41372 & n41381 ;
  assign n41383 = n41362 & ~n41382 ;
  assign n41384 = ~n41309 & n41367 ;
  assign n41385 = n41309 & n41348 ;
  assign n41386 = ~n41384 & ~n41385 ;
  assign n41387 = n41303 & ~n41386 ;
  assign n41388 = ~n41315 & n41368 ;
  assign n41389 = n41309 & ~n41329 ;
  assign n41390 = n41331 & n41389 ;
  assign n41391 = ~n41388 & ~n41390 ;
  assign n41392 = ~n41303 & ~n41391 ;
  assign n41393 = ~n41387 & ~n41392 ;
  assign n41394 = ~n41383 & n41393 ;
  assign n41395 = ~n41363 & n41394 ;
  assign n41396 = ~\u1_L5_reg[14]/NET0131  & ~n41395 ;
  assign n41397 = \u1_L5_reg[14]/NET0131  & n41395 ;
  assign n41398 = ~n41396 & ~n41397 ;
  assign n41399 = ~n41082 & n41105 ;
  assign n41400 = ~n41140 & ~n41153 ;
  assign n41401 = ~n41399 & n41400 ;
  assign n41402 = n41115 & ~n41401 ;
  assign n41403 = ~n41088 & n41107 ;
  assign n41404 = ~n41130 & ~n41403 ;
  assign n41405 = ~n41402 & n41404 ;
  assign n41406 = ~n41082 & n41088 ;
  assign n41407 = n41101 & n41406 ;
  assign n41414 = n41130 & ~n41407 ;
  assign n41408 = ~n41094 & ~n41101 ;
  assign n41409 = ~n41088 & n41115 ;
  assign n41410 = n41408 & n41409 ;
  assign n41411 = n41082 & ~n41115 ;
  assign n41412 = n41142 & n41411 ;
  assign n41415 = ~n41410 & ~n41412 ;
  assign n41416 = n41414 & n41415 ;
  assign n41413 = n41094 & n41120 ;
  assign n41417 = ~n41136 & ~n41413 ;
  assign n41418 = n41416 & n41417 ;
  assign n41419 = ~n41405 & ~n41418 ;
  assign n41420 = n41139 & n41406 ;
  assign n41421 = n41121 & ~n41420 ;
  assign n41422 = n41138 & n41421 ;
  assign n41423 = ~n41082 & n41140 ;
  assign n41424 = ~n41103 & n41115 ;
  assign n41425 = ~n41423 & n41424 ;
  assign n41426 = ~n41422 & ~n41425 ;
  assign n41427 = ~n41115 & ~n41130 ;
  assign n41428 = n41119 & n41427 ;
  assign n41429 = ~n41426 & ~n41428 ;
  assign n41430 = ~n41419 & n41429 ;
  assign n41431 = \u1_L5_reg[15]/P0001  & n41430 ;
  assign n41432 = ~\u1_L5_reg[15]/P0001  & ~n41430 ;
  assign n41433 = ~n41431 & ~n41432 ;
  assign n41434 = ~n40634 & ~n40687 ;
  assign n41435 = n40634 & ~n40678 ;
  assign n41436 = ~n40661 & n41435 ;
  assign n41437 = ~n41434 & ~n41436 ;
  assign n41439 = ~n40656 & ~n40661 ;
  assign n41440 = ~n40628 & ~n41439 ;
  assign n41438 = n40628 & ~n41173 ;
  assign n41441 = n40675 & ~n41438 ;
  assign n41442 = ~n41440 & n41441 ;
  assign n41443 = ~n41437 & n41442 ;
  assign n41445 = ~n40641 & ~n40656 ;
  assign n41446 = n41435 & ~n41445 ;
  assign n41444 = ~n40634 & ~n41173 ;
  assign n41447 = n40628 & n41045 ;
  assign n41448 = ~n40675 & ~n41447 ;
  assign n41449 = ~n41444 & n41448 ;
  assign n41450 = ~n41446 & n41449 ;
  assign n41451 = ~n41443 & ~n41450 ;
  assign n41452 = n40635 & n40657 ;
  assign n41453 = ~n40663 & ~n40709 ;
  assign n41454 = ~n41452 & n41453 ;
  assign n41455 = ~n41451 & n41454 ;
  assign n41456 = ~\u1_L5_reg[19]/NET0131  & ~n41455 ;
  assign n41457 = \u1_L5_reg[19]/NET0131  & n41455 ;
  assign n41458 = ~n41456 & ~n41457 ;
  assign n41459 = ~n40891 & ~n40898 ;
  assign n41460 = n40855 & ~n41459 ;
  assign n41461 = n40861 & ~n40904 ;
  assign n41462 = n41211 & n41461 ;
  assign n41463 = ~n41460 & n41462 ;
  assign n41464 = n40867 & n40892 ;
  assign n41465 = ~n40861 & ~n40933 ;
  assign n41466 = ~n41464 & n41465 ;
  assign n41467 = ~n41463 & ~n41466 ;
  assign n41469 = n40874 & n40891 ;
  assign n41470 = ~n40861 & ~n40911 ;
  assign n41471 = ~n41469 & n41470 ;
  assign n41472 = ~n40880 & n40888 ;
  assign n41473 = n40861 & ~n40914 ;
  assign n41474 = ~n41472 & n41473 ;
  assign n41475 = ~n41471 & ~n41474 ;
  assign n41468 = n40867 & n40911 ;
  assign n41476 = ~n40855 & ~n41468 ;
  assign n41477 = n40931 & n41476 ;
  assign n41478 = ~n41475 & n41477 ;
  assign n41479 = ~n40881 & n40928 ;
  assign n41480 = ~n40919 & ~n41479 ;
  assign n41481 = ~n40861 & ~n41480 ;
  assign n41482 = n40855 & ~n40932 ;
  assign n41483 = ~n41464 & n41482 ;
  assign n41484 = ~n41481 & n41483 ;
  assign n41485 = ~n41478 & ~n41484 ;
  assign n41486 = ~n41467 & ~n41485 ;
  assign n41487 = ~\u1_L5_reg[1]/NET0131  & ~n41486 ;
  assign n41488 = \u1_L5_reg[1]/NET0131  & n41486 ;
  assign n41489 = ~n41487 & ~n41488 ;
  assign n41496 = ~n41101 & ~n41115 ;
  assign n41497 = n41105 & n41496 ;
  assign n41503 = ~n41130 & ~n41497 ;
  assign n41504 = ~n41137 & n41503 ;
  assign n41501 = n41094 & n41104 ;
  assign n41502 = ~n41409 & n41501 ;
  assign n41505 = ~n41147 & ~n41502 ;
  assign n41506 = n41504 & n41505 ;
  assign n41492 = n41088 & ~n41101 ;
  assign n41493 = ~n41115 & n41139 ;
  assign n41494 = ~n41492 & ~n41493 ;
  assign n41495 = n41082 & ~n41494 ;
  assign n41498 = n41101 & n41105 ;
  assign n41499 = ~n41120 & ~n41498 ;
  assign n41500 = n41115 & ~n41499 ;
  assign n41507 = ~n41495 & ~n41500 ;
  assign n41508 = n41506 & n41507 ;
  assign n41509 = ~n41107 & ~n41115 ;
  assign n41510 = ~n41413 & n41509 ;
  assign n41512 = ~n41102 & n41115 ;
  assign n41511 = n41094 & n41117 ;
  assign n41513 = ~n41154 & ~n41511 ;
  assign n41514 = n41512 & n41513 ;
  assign n41515 = ~n41510 & ~n41514 ;
  assign n41516 = ~n41094 & ~n41492 ;
  assign n41517 = n41082 & ~n41119 ;
  assign n41518 = n41516 & n41517 ;
  assign n41519 = n41130 & ~n41423 ;
  assign n41520 = ~n41518 & n41519 ;
  assign n41521 = ~n41515 & n41520 ;
  assign n41522 = ~n41508 & ~n41521 ;
  assign n41490 = n41115 & n41118 ;
  assign n41491 = n41095 & n41132 ;
  assign n41523 = ~n41490 & ~n41491 ;
  assign n41524 = ~n41522 & n41523 ;
  assign n41525 = ~\u1_L5_reg[21]/NET0131  & ~n41524 ;
  assign n41526 = \u1_L5_reg[21]/NET0131  & n41524 ;
  assign n41527 = ~n41525 & ~n41526 ;
  assign n41546 = ~n40567 & ~n40599 ;
  assign n41547 = ~n40565 & ~n41546 ;
  assign n41548 = ~n40593 & ~n41547 ;
  assign n41549 = n40584 & ~n41548 ;
  assign n41550 = n40825 & n40833 ;
  assign n41551 = ~n40610 & ~n41550 ;
  assign n41552 = ~n40832 & n41551 ;
  assign n41553 = ~n41549 & n41552 ;
  assign n41554 = ~n40537 & ~n41553 ;
  assign n41528 = ~n40599 & ~n40607 ;
  assign n41529 = n40572 & ~n41528 ;
  assign n41535 = ~n40558 & ~n40584 ;
  assign n41534 = n40586 & n40825 ;
  assign n41536 = ~n40831 & ~n41534 ;
  assign n41537 = n41535 & n41536 ;
  assign n41530 = n40537 & n40599 ;
  assign n41531 = ~n40537 & n40565 ;
  assign n41532 = ~n40551 & n41531 ;
  assign n41533 = ~n40833 & n41532 ;
  assign n41538 = ~n41530 & ~n41533 ;
  assign n41539 = n41537 & n41538 ;
  assign n41540 = n40537 & ~n40574 ;
  assign n41541 = n40590 & n41540 ;
  assign n41542 = n40584 & ~n40835 ;
  assign n41543 = ~n40606 & n41542 ;
  assign n41544 = ~n41541 & n41543 ;
  assign n41545 = ~n41539 & ~n41544 ;
  assign n41555 = ~n41529 & ~n41545 ;
  assign n41556 = ~n41554 & n41555 ;
  assign n41557 = \u1_L5_reg[23]/NET0131  & ~n41556 ;
  assign n41558 = ~\u1_L5_reg[23]/NET0131  & n41556 ;
  assign n41559 = ~n41557 & ~n41558 ;
  assign n41566 = ~n41315 & ~n41333 ;
  assign n41565 = n41315 & ~n41389 ;
  assign n41567 = n41303 & ~n41322 ;
  assign n41568 = ~n41565 & ~n41567 ;
  assign n41569 = ~n41566 & n41568 ;
  assign n41562 = n41303 & ~n41331 ;
  assign n41560 = ~n41315 & ~n41329 ;
  assign n41561 = ~n41303 & ~n41560 ;
  assign n41563 = ~n41309 & ~n41561 ;
  assign n41564 = ~n41562 & n41563 ;
  assign n41570 = ~n41362 & ~n41564 ;
  assign n41571 = ~n41569 & n41570 ;
  assign n41573 = ~n41315 & n41342 ;
  assign n41574 = ~n41303 & ~n41573 ;
  assign n41575 = ~n41345 & n41574 ;
  assign n41576 = ~n41334 & ~n41389 ;
  assign n41577 = ~n41322 & ~n41576 ;
  assign n41578 = n41315 & n41342 ;
  assign n41579 = n41303 & ~n41560 ;
  assign n41580 = ~n41578 & n41579 ;
  assign n41581 = ~n41577 & n41580 ;
  assign n41582 = ~n41575 & ~n41581 ;
  assign n41572 = n41329 & n41332 ;
  assign n41583 = ~n41323 & n41362 ;
  assign n41584 = ~n41572 & n41583 ;
  assign n41585 = ~n41582 & n41584 ;
  assign n41586 = ~n41571 & ~n41585 ;
  assign n41589 = ~n41385 & ~n41572 ;
  assign n41590 = n41334 & n41336 ;
  assign n41591 = n41589 & ~n41590 ;
  assign n41592 = n41303 & ~n41591 ;
  assign n41587 = n41329 & n41343 ;
  assign n41588 = ~n41303 & n41587 ;
  assign n41593 = ~n41330 & ~n41588 ;
  assign n41594 = ~n41592 & n41593 ;
  assign n41595 = ~n41586 & n41594 ;
  assign n41596 = ~\u1_L5_reg[25]/NET0131  & ~n41595 ;
  assign n41597 = \u1_L5_reg[25]/NET0131  & n41595 ;
  assign n41598 = ~n41596 & ~n41597 ;
  assign n41602 = n40867 & n40881 ;
  assign n41601 = ~n40867 & ~n40881 ;
  assign n41603 = ~n40887 & ~n40918 ;
  assign n41604 = ~n41601 & n41603 ;
  assign n41605 = ~n41602 & n41604 ;
  assign n41599 = ~n40895 & ~n40932 ;
  assign n41600 = ~n40855 & ~n41599 ;
  assign n41606 = ~n40861 & ~n41600 ;
  assign n41607 = ~n41605 & n41606 ;
  assign n41608 = n40861 & ~n40899 ;
  assign n41609 = ~n40930 & n41608 ;
  assign n41610 = ~n41607 & ~n41609 ;
  assign n41615 = ~n40919 & ~n40923 ;
  assign n41616 = ~n41602 & n41615 ;
  assign n41617 = n40887 & ~n41616 ;
  assign n41612 = n40888 & n40891 ;
  assign n41613 = ~n40926 & ~n41612 ;
  assign n41614 = ~n40861 & ~n41613 ;
  assign n41611 = ~n40887 & n40903 ;
  assign n41618 = n40855 & ~n40901 ;
  assign n41619 = ~n41611 & n41618 ;
  assign n41620 = ~n41614 & n41619 ;
  assign n41621 = ~n41617 & n41620 ;
  assign n41624 = ~n40855 & ~n40898 ;
  assign n41625 = ~n40935 & n41624 ;
  assign n41622 = n40867 & ~n40918 ;
  assign n41623 = n41197 & n41622 ;
  assign n41626 = ~n40930 & ~n41623 ;
  assign n41627 = n41625 & n41626 ;
  assign n41628 = ~n41621 & ~n41627 ;
  assign n41629 = ~n41610 & ~n41628 ;
  assign n41630 = ~\u1_L5_reg[26]/NET0131  & ~n41629 ;
  assign n41631 = \u1_L5_reg[26]/NET0131  & n41629 ;
  assign n41632 = ~n41630 & ~n41631 ;
  assign n41636 = ~n40985 & ~n40986 ;
  assign n41637 = n40978 & n41636 ;
  assign n41635 = n40985 & n41023 ;
  assign n41638 = n40953 & ~n41021 ;
  assign n41639 = ~n41635 & n41638 ;
  assign n41640 = ~n41637 & n41639 ;
  assign n41642 = ~n40953 & ~n40979 ;
  assign n41641 = ~n40993 & ~n41287 ;
  assign n41643 = ~n41266 & n41641 ;
  assign n41644 = n41642 & n41643 ;
  assign n41645 = ~n41640 & ~n41644 ;
  assign n41633 = ~n41021 & ~n41023 ;
  assign n41634 = n40986 & ~n41633 ;
  assign n41646 = n41009 & ~n41634 ;
  assign n41647 = ~n41645 & n41646 ;
  assign n41648 = n40953 & n41641 ;
  assign n41649 = ~n40981 & ~n40987 ;
  assign n41650 = ~n41260 & n41649 ;
  assign n41651 = n41642 & n41650 ;
  assign n41652 = ~n41648 & ~n41651 ;
  assign n41653 = n40971 & n41272 ;
  assign n41654 = ~n41009 & ~n41266 ;
  assign n41655 = ~n41653 & n41654 ;
  assign n41656 = ~n41652 & n41655 ;
  assign n41657 = ~n41647 & ~n41656 ;
  assign n41658 = ~\u1_L5_reg[28]/NET0131  & n41657 ;
  assign n41659 = \u1_L5_reg[28]/NET0131  & ~n41657 ;
  assign n41660 = ~n41658 & ~n41659 ;
  assign n41673 = n41334 & n41347 ;
  assign n41674 = ~n41573 & ~n41673 ;
  assign n41675 = n41303 & ~n41674 ;
  assign n41676 = n41329 & n41373 ;
  assign n41677 = n41391 & ~n41676 ;
  assign n41678 = ~n41675 & n41677 ;
  assign n41679 = n41362 & ~n41678 ;
  assign n41662 = n41336 & ~n41343 ;
  assign n41663 = n41574 & ~n41662 ;
  assign n41664 = n41303 & ~n41335 ;
  assign n41665 = ~n41578 & n41664 ;
  assign n41666 = ~n41663 & ~n41665 ;
  assign n41667 = ~n41345 & n41589 ;
  assign n41668 = ~n41666 & n41667 ;
  assign n41669 = ~n41362 & ~n41668 ;
  assign n41661 = ~n41322 & n41588 ;
  assign n41670 = n41336 & ~n41364 ;
  assign n41671 = ~n41332 & ~n41670 ;
  assign n41672 = n41303 & ~n41671 ;
  assign n41680 = ~n41661 & ~n41672 ;
  assign n41681 = ~n41669 & n41680 ;
  assign n41682 = ~n41679 & n41681 ;
  assign n41683 = ~\u1_L5_reg[8]/NET0131  & ~n41682 ;
  assign n41684 = \u1_L5_reg[8]/NET0131  & n41682 ;
  assign n41685 = ~n41683 & ~n41684 ;
  assign n41702 = ~n41102 & ~n41118 ;
  assign n41703 = ~n41498 & n41702 ;
  assign n41704 = ~n41115 & ~n41703 ;
  assign n41705 = ~n41103 & ~n41511 ;
  assign n41693 = n41094 & n41101 ;
  assign n41698 = ~n41408 & ~n41693 ;
  assign n41699 = n41088 & n41115 ;
  assign n41700 = ~n41134 & n41699 ;
  assign n41701 = ~n41698 & n41700 ;
  assign n41706 = ~n41147 & ~n41701 ;
  assign n41707 = n41705 & n41706 ;
  assign n41708 = ~n41704 & n41707 ;
  assign n41709 = n41130 & ~n41708 ;
  assign n41686 = ~n41406 & ~n41516 ;
  assign n41687 = n41115 & ~n41399 ;
  assign n41688 = ~n41686 & n41687 ;
  assign n41689 = ~n41141 & ~n41688 ;
  assign n41690 = ~n41130 & ~n41689 ;
  assign n41691 = ~n41136 & ~n41143 ;
  assign n41692 = ~n41115 & ~n41691 ;
  assign n41694 = n41411 & n41693 ;
  assign n41695 = ~n41497 & ~n41694 ;
  assign n41696 = ~n41130 & ~n41695 ;
  assign n41697 = n41134 & n41409 ;
  assign n41710 = ~n41133 & ~n41697 ;
  assign n41711 = ~n41696 & n41710 ;
  assign n41712 = ~n41692 & n41711 ;
  assign n41713 = ~n41690 & n41712 ;
  assign n41714 = ~n41709 & n41713 ;
  assign n41715 = ~\u1_L5_reg[27]/NET0131  & ~n41714 ;
  assign n41716 = \u1_L5_reg[27]/NET0131  & n41714 ;
  assign n41717 = ~n41715 & ~n41716 ;
  assign n41723 = ~n40779 & ~n40800 ;
  assign n41725 = ~n40766 & n41238 ;
  assign n41726 = n41723 & ~n41725 ;
  assign n41724 = ~n40766 & ~n41723 ;
  assign n41727 = ~n40758 & ~n41724 ;
  assign n41728 = ~n41726 & n41727 ;
  assign n41718 = n40768 & n40800 ;
  assign n41719 = n40731 & ~n40800 ;
  assign n41720 = n40789 & ~n41719 ;
  assign n41721 = ~n40751 & ~n41720 ;
  assign n41722 = n40758 & ~n41721 ;
  assign n41729 = ~n41718 & ~n41722 ;
  assign n41730 = ~n41728 & n41729 ;
  assign n41731 = n40725 & ~n41730 ;
  assign n41733 = ~n41230 & ~n41238 ;
  assign n41734 = ~n40758 & ~n41733 ;
  assign n41735 = ~n40737 & n40782 ;
  assign n41736 = n40758 & ~n41230 ;
  assign n41737 = ~n41735 & n41736 ;
  assign n41738 = ~n41734 & ~n41737 ;
  assign n41732 = n40737 & ~n41232 ;
  assign n41739 = n40799 & ~n41732 ;
  assign n41740 = ~n41738 & n41739 ;
  assign n41741 = ~n40725 & ~n41740 ;
  assign n41742 = n40758 & n40781 ;
  assign n41743 = ~n40769 & n40796 ;
  assign n41744 = n40762 & n41743 ;
  assign n41745 = ~n41742 & ~n41744 ;
  assign n41746 = ~n41741 & n41745 ;
  assign n41747 = ~n41731 & n41746 ;
  assign n41748 = \u1_L5_reg[32]/NET0131  & n41747 ;
  assign n41749 = ~\u1_L5_reg[32]/NET0131  & ~n41747 ;
  assign n41750 = ~n41748 & ~n41749 ;
  assign n41751 = ~n41322 & n41587 ;
  assign n41752 = n41362 & ~n41751 ;
  assign n41753 = ~n41330 & ~n41374 ;
  assign n41754 = n41752 & n41753 ;
  assign n41755 = ~n41333 & n41343 ;
  assign n41756 = ~n41362 & ~n41755 ;
  assign n41757 = ~n41347 & ~n41349 ;
  assign n41758 = ~n41573 & n41757 ;
  assign n41759 = n41756 & n41758 ;
  assign n41760 = ~n41754 & ~n41759 ;
  assign n41761 = ~n41303 & ~n41344 ;
  assign n41762 = ~n41673 & n41761 ;
  assign n41763 = ~n41384 & n41762 ;
  assign n41764 = ~n41760 & n41763 ;
  assign n41765 = ~n41309 & n41336 ;
  assign n41766 = ~n41367 & ~n41765 ;
  assign n41767 = n41756 & n41766 ;
  assign n41768 = ~n41329 & n41331 ;
  assign n41769 = ~n41366 & ~n41768 ;
  assign n41770 = n41752 & n41769 ;
  assign n41771 = ~n41767 & ~n41770 ;
  assign n41772 = ~n41388 & n41664 ;
  assign n41773 = ~n41771 & n41772 ;
  assign n41774 = ~n41764 & ~n41773 ;
  assign n41775 = ~\u1_L5_reg[3]/NET0131  & n41774 ;
  assign n41776 = \u1_L5_reg[3]/NET0131  & ~n41774 ;
  assign n41777 = ~n41775 & ~n41776 ;
  assign n41778 = decrypt_pad & ~\u1_uk_K_r5_reg[25]/NET0131  ;
  assign n41779 = ~decrypt_pad & ~\u1_uk_K_r5_reg[3]/NET0131  ;
  assign n41780 = ~n41778 & ~n41779 ;
  assign n41781 = \u1_R5_reg[13]/NET0131  & ~n41780 ;
  assign n41782 = ~\u1_R5_reg[13]/NET0131  & n41780 ;
  assign n41783 = ~n41781 & ~n41782 ;
  assign n41791 = decrypt_pad & ~\u1_uk_K_r5_reg[20]/NET0131  ;
  assign n41792 = ~decrypt_pad & ~\u1_uk_K_r5_reg[55]/NET0131  ;
  assign n41793 = ~n41791 & ~n41792 ;
  assign n41794 = \u1_R5_reg[9]/NET0131  & ~n41793 ;
  assign n41795 = ~\u1_R5_reg[9]/NET0131  & n41793 ;
  assign n41796 = ~n41794 & ~n41795 ;
  assign n41805 = ~n41783 & n41796 ;
  assign n41806 = decrypt_pad & ~\u1_uk_K_r5_reg[54]/NET0131  ;
  assign n41807 = ~decrypt_pad & ~\u1_uk_K_r5_reg[32]/NET0131  ;
  assign n41808 = ~n41806 & ~n41807 ;
  assign n41809 = \u1_R5_reg[11]/NET0131  & ~n41808 ;
  assign n41810 = ~\u1_R5_reg[11]/NET0131  & n41808 ;
  assign n41811 = ~n41809 & ~n41810 ;
  assign n41812 = ~n41805 & ~n41811 ;
  assign n41797 = decrypt_pad & ~\u1_uk_K_r5_reg[53]/NET0131  ;
  assign n41798 = ~decrypt_pad & ~\u1_uk_K_r5_reg[6]/NET0131  ;
  assign n41799 = ~n41797 & ~n41798 ;
  assign n41800 = \u1_R5_reg[10]/NET0131  & ~n41799 ;
  assign n41801 = ~\u1_R5_reg[10]/NET0131  & n41799 ;
  assign n41802 = ~n41800 & ~n41801 ;
  assign n41813 = n41796 & ~n41802 ;
  assign n41784 = decrypt_pad & ~\u1_uk_K_r5_reg[48]/NET0131  ;
  assign n41785 = ~decrypt_pad & ~\u1_uk_K_r5_reg[26]/NET0131  ;
  assign n41786 = ~n41784 & ~n41785 ;
  assign n41787 = \u1_R5_reg[8]/NET0131  & ~n41786 ;
  assign n41788 = ~\u1_R5_reg[8]/NET0131  & n41786 ;
  assign n41789 = ~n41787 & ~n41788 ;
  assign n41814 = n41783 & ~n41796 ;
  assign n41815 = n41789 & ~n41814 ;
  assign n41816 = ~n41813 & ~n41815 ;
  assign n41817 = n41812 & ~n41816 ;
  assign n41790 = ~n41783 & ~n41789 ;
  assign n41803 = n41796 & n41802 ;
  assign n41804 = n41790 & n41803 ;
  assign n41818 = decrypt_pad & ~\u1_uk_K_r5_reg[12]/P0001  ;
  assign n41819 = ~decrypt_pad & ~\u1_uk_K_r5_reg[47]/NET0131  ;
  assign n41820 = ~n41818 & ~n41819 ;
  assign n41821 = \u1_R5_reg[12]/NET0131  & ~n41820 ;
  assign n41822 = ~\u1_R5_reg[12]/NET0131  & n41820 ;
  assign n41823 = ~n41821 & ~n41822 ;
  assign n41824 = ~n41804 & n41823 ;
  assign n41825 = ~n41817 & n41824 ;
  assign n41829 = n41783 & n41789 ;
  assign n41830 = ~n41790 & ~n41829 ;
  assign n41826 = ~n41789 & n41811 ;
  assign n41828 = ~n41796 & ~n41802 ;
  assign n41837 = ~n41826 & n41828 ;
  assign n41838 = n41830 & n41837 ;
  assign n41839 = ~n41783 & n41789 ;
  assign n41840 = n41803 & n41839 ;
  assign n41827 = n41813 & n41826 ;
  assign n41841 = ~n41823 & ~n41827 ;
  assign n41842 = ~n41840 & n41841 ;
  assign n41843 = ~n41838 & n41842 ;
  assign n41831 = ~n41828 & ~n41830 ;
  assign n41832 = ~n41803 & n41831 ;
  assign n41833 = n41783 & ~n41789 ;
  assign n41834 = n41802 & n41833 ;
  assign n41835 = n41796 & n41834 ;
  assign n41836 = ~n41811 & n41835 ;
  assign n41844 = ~n41832 & ~n41836 ;
  assign n41845 = n41843 & n41844 ;
  assign n41846 = ~n41825 & ~n41845 ;
  assign n41848 = n41796 & n41839 ;
  assign n41849 = ~n41834 & ~n41848 ;
  assign n41850 = ~n41814 & n41849 ;
  assign n41851 = n41823 & ~n41850 ;
  assign n41847 = n41802 & n41814 ;
  assign n41852 = n41790 & ~n41802 ;
  assign n41853 = ~n41796 & n41852 ;
  assign n41854 = ~n41847 & ~n41853 ;
  assign n41855 = ~n41851 & n41854 ;
  assign n41856 = n41811 & ~n41855 ;
  assign n41857 = ~n41846 & ~n41856 ;
  assign n41858 = ~\u1_L5_reg[6]/NET0131  & ~n41857 ;
  assign n41859 = \u1_L5_reg[6]/NET0131  & n41857 ;
  assign n41860 = ~n41858 & ~n41859 ;
  assign n41878 = ~n40750 & ~n41236 ;
  assign n41861 = n40737 & ~n41723 ;
  assign n41879 = n40731 & n40800 ;
  assign n41880 = ~n41861 & ~n41879 ;
  assign n41881 = ~n41878 & n41880 ;
  assign n41882 = ~n40758 & ~n41881 ;
  assign n41862 = ~n41735 & ~n41861 ;
  assign n41863 = n40731 & ~n41862 ;
  assign n41872 = ~n40731 & ~n40744 ;
  assign n41873 = n41723 & n41872 ;
  assign n41883 = n40758 & n41873 ;
  assign n41884 = ~n41863 & ~n41883 ;
  assign n41885 = ~n41882 & n41884 ;
  assign n41886 = n40725 & ~n41885 ;
  assign n41864 = ~n40758 & n41863 ;
  assign n41865 = n40725 & ~n40758 ;
  assign n41866 = n40788 & ~n41723 ;
  assign n41867 = n40743 & ~n41248 ;
  assign n41868 = n40758 & n41719 ;
  assign n41869 = ~n41867 & n41868 ;
  assign n41870 = ~n41866 & ~n41869 ;
  assign n41871 = ~n40725 & ~n41870 ;
  assign n41874 = ~n40758 & n41873 ;
  assign n41875 = ~n40752 & ~n41874 ;
  assign n41876 = ~n41871 & n41875 ;
  assign n41877 = ~n41865 & ~n41876 ;
  assign n41887 = ~n41864 & ~n41877 ;
  assign n41888 = ~n41886 & n41887 ;
  assign n41889 = ~\u1_L5_reg[7]/NET0131  & ~n41888 ;
  assign n41890 = \u1_L5_reg[7]/NET0131  & n41888 ;
  assign n41891 = ~n41889 & ~n41890 ;
  assign n41894 = ~n40813 & n41546 ;
  assign n41895 = n40537 & ~n41894 ;
  assign n41896 = n40557 & n40815 ;
  assign n41892 = ~n40551 & ~n40826 ;
  assign n41893 = ~n40537 & ~n41892 ;
  assign n41897 = ~n40557 & n40609 ;
  assign n41898 = ~n41893 & ~n41897 ;
  assign n41899 = ~n41896 & n41898 ;
  assign n41900 = ~n41895 & n41899 ;
  assign n41901 = ~n40584 & ~n41900 ;
  assign n41902 = n40812 & n40825 ;
  assign n41903 = ~n41897 & ~n41902 ;
  assign n41904 = ~n40537 & ~n41903 ;
  assign n41906 = n40557 & ~n40590 ;
  assign n41907 = ~n40815 & n41906 ;
  assign n41905 = n40572 & ~n41892 ;
  assign n41908 = ~n40832 & ~n41905 ;
  assign n41909 = ~n41907 & n41908 ;
  assign n41910 = n40584 & ~n41909 ;
  assign n41911 = ~n41904 & ~n41910 ;
  assign n41912 = ~n41901 & n41911 ;
  assign n41913 = ~\u1_L5_reg[9]/NET0131  & ~n41912 ;
  assign n41914 = \u1_L5_reg[9]/NET0131  & n41912 ;
  assign n41915 = ~n41913 & ~n41914 ;
  assign n41916 = n41796 & n41829 ;
  assign n41917 = ~n41796 & n41833 ;
  assign n41918 = ~n41916 & ~n41917 ;
  assign n41919 = ~n41796 & n41839 ;
  assign n41920 = n41805 & n41826 ;
  assign n41921 = ~n41919 & ~n41920 ;
  assign n41922 = n41918 & n41921 ;
  assign n41923 = ~n41802 & ~n41922 ;
  assign n41924 = n41790 & n41802 ;
  assign n41925 = ~n41802 & n41839 ;
  assign n41926 = ~n41924 & ~n41925 ;
  assign n41927 = ~n41811 & ~n41926 ;
  assign n41928 = n41823 & ~n41835 ;
  assign n41929 = ~n41927 & n41928 ;
  assign n41930 = ~n41923 & n41929 ;
  assign n41935 = ~n41852 & n41918 ;
  assign n41936 = ~n41811 & ~n41935 ;
  assign n41931 = ~n41796 & ~n41829 ;
  assign n41932 = ~n41790 & n41811 ;
  assign n41933 = ~n41916 & n41932 ;
  assign n41934 = ~n41931 & n41933 ;
  assign n41937 = ~n41823 & ~n41853 ;
  assign n41938 = ~n41934 & n41937 ;
  assign n41939 = ~n41936 & n41938 ;
  assign n41940 = ~n41930 & ~n41939 ;
  assign n41941 = ~n41796 & n41924 ;
  assign n41942 = ~n41840 & ~n41941 ;
  assign n41943 = n41811 & ~n41942 ;
  assign n41944 = n41789 & n41802 ;
  assign n41945 = ~n41796 & n41944 ;
  assign n41946 = ~n41811 & n41945 ;
  assign n41947 = ~n41943 & ~n41946 ;
  assign n41948 = ~n41940 & n41947 ;
  assign n41949 = ~\u1_L5_reg[16]/NET0131  & ~n41948 ;
  assign n41950 = \u1_L5_reg[16]/NET0131  & n41948 ;
  assign n41951 = ~n41949 & ~n41950 ;
  assign n41956 = n40953 & ~n40988 ;
  assign n41953 = ~n40965 & n41014 ;
  assign n41954 = ~n41022 & ~n41953 ;
  assign n41955 = ~n40953 & ~n41954 ;
  assign n41957 = ~n40980 & ~n41955 ;
  assign n41958 = ~n41956 & n41957 ;
  assign n41959 = n41009 & ~n41958 ;
  assign n41966 = n40965 & ~n41015 ;
  assign n41967 = n41033 & ~n41966 ;
  assign n41965 = n40998 & ~n41636 ;
  assign n41963 = n40953 & n40959 ;
  assign n41964 = n40981 & n41963 ;
  assign n41968 = ~n41027 & ~n41964 ;
  assign n41969 = ~n41965 & n41968 ;
  assign n41970 = ~n41967 & n41969 ;
  assign n41971 = ~n41009 & ~n41970 ;
  assign n41952 = ~n40953 & n40993 ;
  assign n41960 = n40959 & n40998 ;
  assign n41961 = ~n41288 & ~n41960 ;
  assign n41962 = n40953 & ~n41961 ;
  assign n41972 = ~n41952 & ~n41962 ;
  assign n41973 = ~n41971 & n41972 ;
  assign n41974 = ~n41959 & n41973 ;
  assign n41975 = \u1_L5_reg[18]/NET0131  & n41974 ;
  assign n41976 = ~\u1_L5_reg[18]/NET0131  & ~n41974 ;
  assign n41977 = ~n41975 & ~n41976 ;
  assign n41988 = n41789 & n41803 ;
  assign n41987 = n41828 & ~n41833 ;
  assign n41989 = ~n41834 & ~n41987 ;
  assign n41990 = ~n41988 & n41989 ;
  assign n41991 = n41811 & ~n41990 ;
  assign n41992 = ~n41838 & ~n41991 ;
  assign n41993 = n41823 & ~n41992 ;
  assign n41978 = ~n41802 & n41833 ;
  assign n41979 = ~n41924 & ~n41978 ;
  assign n41980 = ~n41789 & n41805 ;
  assign n41981 = ~n41945 & ~n41980 ;
  assign n41982 = n41979 & n41981 ;
  assign n41983 = n41811 & ~n41982 ;
  assign n41984 = n41802 & n41919 ;
  assign n41985 = ~n41983 & ~n41984 ;
  assign n41986 = ~n41823 & ~n41985 ;
  assign n41994 = n41828 & ~n41830 ;
  assign n41995 = ~n41823 & n41849 ;
  assign n41996 = ~n41994 & n41995 ;
  assign n41997 = n41823 & ~n41831 ;
  assign n41998 = ~n41811 & ~n41997 ;
  assign n41999 = ~n41996 & n41998 ;
  assign n42000 = n41802 & ~n41811 ;
  assign n42001 = n41916 & n42000 ;
  assign n42002 = n41811 & ~n41814 ;
  assign n42003 = ~n41802 & ~n41805 ;
  assign n42004 = n41830 & n42003 ;
  assign n42005 = n42002 & n42004 ;
  assign n42006 = ~n42001 & ~n42005 ;
  assign n42007 = ~n41999 & n42006 ;
  assign n42008 = ~n41986 & n42007 ;
  assign n42009 = ~n41993 & n42008 ;
  assign n42010 = ~\u1_L5_reg[24]/NET0131  & ~n42009 ;
  assign n42011 = \u1_L5_reg[24]/NET0131  & n42009 ;
  assign n42012 = ~n42010 & ~n42011 ;
  assign n42028 = ~n41783 & n41813 ;
  assign n42027 = ~n41805 & n41944 ;
  assign n42029 = ~n41823 & ~n42027 ;
  assign n42030 = ~n42028 & n42029 ;
  assign n42024 = n41828 & n41839 ;
  assign n42025 = n41823 & ~n42024 ;
  assign n42026 = n41979 & n42025 ;
  assign n42031 = n41811 & ~n42026 ;
  assign n42032 = ~n42030 & n42031 ;
  assign n42018 = ~n41802 & ~n41917 ;
  assign n42019 = ~n41834 & ~n42018 ;
  assign n42020 = ~n41796 & ~n41839 ;
  assign n42021 = ~n41812 & ~n42020 ;
  assign n42022 = ~n41823 & ~n42021 ;
  assign n42023 = ~n42019 & n42022 ;
  assign n42033 = ~n41789 & n41823 ;
  assign n42034 = ~n41802 & ~n42033 ;
  assign n42035 = n41805 & ~n41811 ;
  assign n42036 = ~n42034 & n42035 ;
  assign n42013 = ~n41811 & ~n41823 ;
  assign n42014 = n41944 & ~n42013 ;
  assign n42015 = ~n42002 & n42014 ;
  assign n42016 = n41803 & n41823 ;
  assign n42017 = ~n41829 & n42016 ;
  assign n42037 = ~n42015 & ~n42017 ;
  assign n42038 = ~n42036 & n42037 ;
  assign n42039 = ~n42023 & n42038 ;
  assign n42040 = ~n42032 & n42039 ;
  assign n42041 = \u1_L5_reg[30]/NET0131  & ~n42040 ;
  assign n42042 = ~\u1_L5_reg[30]/NET0131  & n42040 ;
  assign n42043 = ~n42041 & ~n42042 ;
  assign n42044 = decrypt_pad & ~\u1_uk_K_r4_reg[50]/NET0131  ;
  assign n42045 = ~decrypt_pad & ~\u1_uk_K_r4_reg[31]/P0001  ;
  assign n42046 = ~n42044 & ~n42045 ;
  assign n42047 = \u1_R4_reg[28]/NET0131  & ~n42046 ;
  assign n42048 = ~\u1_R4_reg[28]/NET0131  & n42046 ;
  assign n42049 = ~n42047 & ~n42048 ;
  assign n42063 = decrypt_pad & ~\u1_uk_K_r4_reg[38]/NET0131  ;
  assign n42064 = ~decrypt_pad & ~\u1_uk_K_r4_reg[42]/NET0131  ;
  assign n42065 = ~n42063 & ~n42064 ;
  assign n42066 = \u1_R4_reg[24]/NET0131  & ~n42065 ;
  assign n42067 = ~\u1_R4_reg[24]/NET0131  & n42065 ;
  assign n42068 = ~n42066 & ~n42067 ;
  assign n42069 = decrypt_pad & ~\u1_uk_K_r4_reg[30]/NET0131  ;
  assign n42070 = ~decrypt_pad & ~\u1_uk_K_r4_reg[7]/NET0131  ;
  assign n42071 = ~n42069 & ~n42070 ;
  assign n42072 = \u1_R4_reg[26]/NET0131  & ~n42071 ;
  assign n42073 = ~\u1_R4_reg[26]/NET0131  & n42071 ;
  assign n42074 = ~n42072 & ~n42073 ;
  assign n42056 = decrypt_pad & ~\u1_uk_K_r4_reg[14]/NET0131  ;
  assign n42057 = ~decrypt_pad & ~\u1_uk_K_r4_reg[22]/NET0131  ;
  assign n42058 = ~n42056 & ~n42057 ;
  assign n42059 = \u1_R4_reg[25]/NET0131  & ~n42058 ;
  assign n42060 = ~\u1_R4_reg[25]/NET0131  & n42058 ;
  assign n42061 = ~n42059 & ~n42060 ;
  assign n42077 = decrypt_pad & ~\u1_uk_K_r4_reg[8]/NET0131  ;
  assign n42078 = ~decrypt_pad & ~\u1_uk_K_r4_reg[16]/NET0131  ;
  assign n42079 = ~n42077 & ~n42078 ;
  assign n42080 = \u1_R4_reg[27]/NET0131  & ~n42079 ;
  assign n42081 = ~\u1_R4_reg[27]/NET0131  & n42079 ;
  assign n42082 = ~n42080 & ~n42081 ;
  assign n42084 = ~n42061 & n42082 ;
  assign n42085 = ~n42074 & n42084 ;
  assign n42050 = decrypt_pad & ~\u1_uk_K_r4_reg[42]/NET0131  ;
  assign n42051 = ~decrypt_pad & ~\u1_uk_K_r4_reg[50]/NET0131  ;
  assign n42052 = ~n42050 & ~n42051 ;
  assign n42053 = \u1_R4_reg[29]/NET0131  & ~n42052 ;
  assign n42054 = ~\u1_R4_reg[29]/NET0131  & n42052 ;
  assign n42055 = ~n42053 & ~n42054 ;
  assign n42087 = n42055 & ~n42074 ;
  assign n42086 = ~n42061 & n42074 ;
  assign n42088 = ~n42082 & ~n42086 ;
  assign n42089 = ~n42087 & n42088 ;
  assign n42090 = ~n42085 & ~n42089 ;
  assign n42091 = n42068 & ~n42090 ;
  assign n42062 = ~n42055 & ~n42061 ;
  assign n42075 = ~n42068 & n42074 ;
  assign n42076 = n42062 & n42075 ;
  assign n42083 = n42076 & ~n42082 ;
  assign n42092 = ~n42068 & ~n42074 ;
  assign n42093 = n42068 & n42074 ;
  assign n42094 = ~n42092 & ~n42093 ;
  assign n42095 = n42055 & ~n42084 ;
  assign n42096 = ~n42094 & n42095 ;
  assign n42097 = ~n42083 & ~n42096 ;
  assign n42098 = ~n42091 & n42097 ;
  assign n42099 = ~n42049 & ~n42098 ;
  assign n42100 = ~n42055 & n42085 ;
  assign n42101 = n42061 & ~n42082 ;
  assign n42102 = ~n42094 & n42101 ;
  assign n42128 = ~n42100 & ~n42102 ;
  assign n42129 = ~n42099 & n42128 ;
  assign n42103 = ~n42061 & ~n42074 ;
  assign n42104 = n42061 & n42074 ;
  assign n42105 = ~n42103 & ~n42104 ;
  assign n42106 = ~n42055 & n42061 ;
  assign n42107 = n42049 & ~n42106 ;
  assign n42108 = n42105 & n42107 ;
  assign n42109 = ~n42062 & ~n42108 ;
  assign n42110 = n42068 & ~n42109 ;
  assign n42111 = n42055 & ~n42061 ;
  assign n42112 = ~n42106 & ~n42111 ;
  assign n42113 = n42075 & ~n42112 ;
  assign n42114 = ~n42110 & ~n42113 ;
  assign n42115 = n42082 & ~n42114 ;
  assign n42118 = n42055 & ~n42068 ;
  assign n42119 = n42061 & n42118 ;
  assign n42122 = n42074 & ~n42119 ;
  assign n42120 = n42068 & n42111 ;
  assign n42121 = ~n42119 & ~n42120 ;
  assign n42123 = ~n42082 & ~n42121 ;
  assign n42124 = ~n42122 & n42123 ;
  assign n42116 = n42075 & n42111 ;
  assign n42117 = n42062 & n42092 ;
  assign n42125 = ~n42116 & ~n42117 ;
  assign n42126 = ~n42124 & n42125 ;
  assign n42127 = n42049 & ~n42126 ;
  assign n42130 = ~n42115 & ~n42127 ;
  assign n42131 = n42129 & n42130 ;
  assign n42132 = ~\u1_L4_reg[22]/NET0131  & ~n42131 ;
  assign n42133 = \u1_L4_reg[22]/NET0131  & n42131 ;
  assign n42134 = ~n42132 & ~n42133 ;
  assign n42135 = decrypt_pad & ~\u1_uk_K_r4_reg[19]/NET0131  ;
  assign n42136 = ~decrypt_pad & ~\u1_uk_K_r4_reg[25]/NET0131  ;
  assign n42137 = ~n42135 & ~n42136 ;
  assign n42138 = \u1_R4_reg[4]/NET0131  & ~n42137 ;
  assign n42139 = ~\u1_R4_reg[4]/NET0131  & n42137 ;
  assign n42140 = ~n42138 & ~n42139 ;
  assign n42141 = decrypt_pad & ~\u1_uk_K_r4_reg[41]/NET0131  ;
  assign n42142 = ~decrypt_pad & ~\u1_uk_K_r4_reg[47]/NET0131  ;
  assign n42143 = ~n42141 & ~n42142 ;
  assign n42144 = \u1_R4_reg[3]/NET0131  & ~n42143 ;
  assign n42145 = ~\u1_R4_reg[3]/NET0131  & n42143 ;
  assign n42146 = ~n42144 & ~n42145 ;
  assign n42160 = decrypt_pad & ~\u1_uk_K_r4_reg[47]/NET0131  ;
  assign n42161 = ~decrypt_pad & ~\u1_uk_K_r4_reg[53]/NET0131  ;
  assign n42162 = ~n42160 & ~n42161 ;
  assign n42163 = \u1_R4_reg[5]/NET0131  & ~n42162 ;
  assign n42164 = ~\u1_R4_reg[5]/NET0131  & n42162 ;
  assign n42165 = ~n42163 & ~n42164 ;
  assign n42169 = decrypt_pad & ~\u1_uk_K_r4_reg[17]/NET0131  ;
  assign n42170 = ~decrypt_pad & ~\u1_uk_K_r4_reg[55]/NET0131  ;
  assign n42171 = ~n42169 & ~n42170 ;
  assign n42172 = \u1_R4_reg[1]/NET0131  & ~n42171 ;
  assign n42173 = ~\u1_R4_reg[1]/NET0131  & n42171 ;
  assign n42174 = ~n42172 & ~n42173 ;
  assign n42180 = n42165 & ~n42174 ;
  assign n42147 = decrypt_pad & ~\u1_uk_K_r4_reg[32]/NET0131  ;
  assign n42148 = ~decrypt_pad & ~\u1_uk_K_r4_reg[13]/NET0131  ;
  assign n42149 = ~n42147 & ~n42148 ;
  assign n42150 = \u1_R4_reg[2]/NET0131  & ~n42149 ;
  assign n42151 = ~\u1_R4_reg[2]/NET0131  & n42149 ;
  assign n42152 = ~n42150 & ~n42151 ;
  assign n42154 = decrypt_pad & ~\u1_uk_K_r4_reg[53]/NET0131  ;
  assign n42155 = ~decrypt_pad & ~\u1_uk_K_r4_reg[34]/NET0131  ;
  assign n42156 = ~n42154 & ~n42155 ;
  assign n42157 = \u1_R4_reg[32]/NET0131  & ~n42156 ;
  assign n42158 = ~\u1_R4_reg[32]/NET0131  & n42156 ;
  assign n42159 = ~n42157 & ~n42158 ;
  assign n42166 = ~n42159 & ~n42165 ;
  assign n42195 = n42152 & n42166 ;
  assign n42196 = ~n42180 & ~n42195 ;
  assign n42197 = n42146 & ~n42196 ;
  assign n42201 = ~n42159 & n42165 ;
  assign n42202 = n42146 & ~n42152 ;
  assign n42203 = n42174 & ~n42202 ;
  assign n42204 = n42201 & ~n42203 ;
  assign n42199 = n42152 & ~n42174 ;
  assign n42200 = ~n42159 & n42199 ;
  assign n42177 = ~n42165 & ~n42174 ;
  assign n42193 = ~n42152 & n42159 ;
  assign n42194 = n42177 & n42193 ;
  assign n42186 = ~n42146 & n42174 ;
  assign n42198 = n42159 & n42186 ;
  assign n42205 = ~n42194 & ~n42198 ;
  assign n42206 = ~n42200 & n42205 ;
  assign n42207 = ~n42204 & n42206 ;
  assign n42208 = ~n42197 & n42207 ;
  assign n42209 = n42140 & ~n42208 ;
  assign n42178 = n42159 & n42177 ;
  assign n42179 = n42152 & n42178 ;
  assign n42181 = ~n42152 & ~n42159 ;
  assign n42182 = ~n42180 & n42181 ;
  assign n42183 = ~n42179 & ~n42182 ;
  assign n42184 = ~n42146 & ~n42183 ;
  assign n42153 = n42146 & n42152 ;
  assign n42167 = n42159 & n42165 ;
  assign n42168 = ~n42166 & ~n42167 ;
  assign n42175 = n42168 & n42174 ;
  assign n42176 = n42153 & n42175 ;
  assign n42185 = n42166 & n42174 ;
  assign n42187 = n42167 & ~n42186 ;
  assign n42188 = ~n42185 & ~n42187 ;
  assign n42189 = ~n42152 & ~n42188 ;
  assign n42190 = ~n42176 & ~n42189 ;
  assign n42191 = ~n42184 & n42190 ;
  assign n42192 = ~n42140 & ~n42191 ;
  assign n42215 = n42167 & n42174 ;
  assign n42216 = n42152 & n42215 ;
  assign n42212 = n42165 & n42200 ;
  assign n42213 = ~n42152 & ~n42165 ;
  assign n42214 = n42174 & n42213 ;
  assign n42217 = ~n42212 & ~n42214 ;
  assign n42218 = ~n42216 & n42217 ;
  assign n42219 = ~n42146 & ~n42218 ;
  assign n42210 = n42146 & ~n42174 ;
  assign n42211 = n42193 & n42210 ;
  assign n42220 = n42146 & ~n42165 ;
  assign n42221 = n42200 & n42220 ;
  assign n42222 = ~n42211 & ~n42221 ;
  assign n42223 = ~n42219 & n42222 ;
  assign n42224 = ~n42192 & n42223 ;
  assign n42225 = ~n42209 & n42224 ;
  assign n42226 = ~\u1_L4_reg[31]/NET0131  & ~n42225 ;
  assign n42227 = \u1_L4_reg[31]/NET0131  & n42225 ;
  assign n42228 = ~n42226 & ~n42227 ;
  assign n42229 = decrypt_pad & ~\u1_uk_K_r4_reg[43]/NET0131  ;
  assign n42230 = ~decrypt_pad & ~\u1_uk_K_r4_reg[51]/NET0131  ;
  assign n42231 = ~n42229 & ~n42230 ;
  assign n42232 = \u1_R4_reg[24]/NET0131  & ~n42231 ;
  assign n42233 = ~\u1_R4_reg[24]/NET0131  & n42231 ;
  assign n42234 = ~n42232 & ~n42233 ;
  assign n42248 = decrypt_pad & ~\u1_uk_K_r4_reg[28]/NET0131  ;
  assign n42249 = ~decrypt_pad & ~\u1_uk_K_r4_reg[36]/NET0131  ;
  assign n42250 = ~n42248 & ~n42249 ;
  assign n42251 = \u1_R4_reg[22]/NET0131  & ~n42250 ;
  assign n42252 = ~\u1_R4_reg[22]/NET0131  & n42250 ;
  assign n42253 = ~n42251 & ~n42252 ;
  assign n42235 = decrypt_pad & ~\u1_uk_K_r4_reg[22]/NET0131  ;
  assign n42236 = ~decrypt_pad & ~\u1_uk_K_r4_reg[30]/NET0131  ;
  assign n42237 = ~n42235 & ~n42236 ;
  assign n42238 = \u1_R4_reg[20]/NET0131  & ~n42237 ;
  assign n42239 = ~\u1_R4_reg[20]/NET0131  & n42237 ;
  assign n42240 = ~n42238 & ~n42239 ;
  assign n42254 = decrypt_pad & ~\u1_uk_K_r4_reg[37]/NET0131  ;
  assign n42255 = ~decrypt_pad & ~\u1_uk_K_r4_reg[14]/NET0131  ;
  assign n42256 = ~n42254 & ~n42255 ;
  assign n42257 = \u1_R4_reg[21]/NET0131  & ~n42256 ;
  assign n42258 = ~\u1_R4_reg[21]/NET0131  & n42256 ;
  assign n42259 = ~n42257 & ~n42258 ;
  assign n42274 = ~n42240 & n42259 ;
  assign n42241 = decrypt_pad & ~\u1_uk_K_r4_reg[7]/NET0131  ;
  assign n42242 = ~decrypt_pad & ~\u1_uk_K_r4_reg[15]/NET0131  ;
  assign n42243 = ~n42241 & ~n42242 ;
  assign n42244 = \u1_R4_reg[25]/NET0131  & ~n42243 ;
  assign n42245 = ~\u1_R4_reg[25]/NET0131  & n42243 ;
  assign n42246 = ~n42244 & ~n42245 ;
  assign n42281 = n42240 & n42246 ;
  assign n42312 = ~n42274 & ~n42281 ;
  assign n42313 = n42253 & ~n42312 ;
  assign n42266 = decrypt_pad & ~\u1_uk_K_r4_reg[45]/NET0131  ;
  assign n42267 = ~decrypt_pad & ~\u1_uk_K_r4_reg[49]/NET0131  ;
  assign n42268 = ~n42266 & ~n42267 ;
  assign n42269 = \u1_R4_reg[23]/NET0131  & ~n42268 ;
  assign n42270 = ~\u1_R4_reg[23]/NET0131  & n42268 ;
  assign n42271 = ~n42269 & ~n42270 ;
  assign n42309 = n42246 & n42259 ;
  assign n42310 = ~n42240 & n42309 ;
  assign n42311 = ~n42253 & ~n42310 ;
  assign n42314 = ~n42271 & ~n42311 ;
  assign n42315 = ~n42313 & n42314 ;
  assign n42247 = n42240 & ~n42246 ;
  assign n42301 = n42247 & ~n42259 ;
  assign n42302 = ~n42253 & n42301 ;
  assign n42275 = n42253 & n42274 ;
  assign n42303 = n42259 & n42281 ;
  assign n42304 = ~n42275 & ~n42303 ;
  assign n42305 = ~n42302 & n42304 ;
  assign n42306 = n42271 & ~n42305 ;
  assign n42279 = ~n42253 & ~n42271 ;
  assign n42307 = n42279 & n42281 ;
  assign n42308 = ~n42259 & n42307 ;
  assign n42316 = ~n42306 & ~n42308 ;
  assign n42317 = ~n42315 & n42316 ;
  assign n42318 = n42234 & ~n42317 ;
  assign n42260 = ~n42253 & n42259 ;
  assign n42276 = n42240 & n42260 ;
  assign n42277 = ~n42275 & ~n42276 ;
  assign n42278 = ~n42271 & ~n42277 ;
  assign n42263 = ~n42240 & ~n42246 ;
  assign n42264 = ~n42259 & ~n42263 ;
  assign n42265 = n42253 & ~n42264 ;
  assign n42262 = n42240 & ~n42253 ;
  assign n42272 = ~n42262 & n42271 ;
  assign n42273 = ~n42265 & n42272 ;
  assign n42261 = n42247 & n42260 ;
  assign n42280 = n42247 & n42279 ;
  assign n42282 = n42253 & ~n42259 ;
  assign n42283 = n42281 & n42282 ;
  assign n42284 = ~n42280 & ~n42283 ;
  assign n42285 = ~n42261 & n42284 ;
  assign n42286 = ~n42273 & n42285 ;
  assign n42287 = ~n42278 & n42286 ;
  assign n42288 = ~n42234 & ~n42287 ;
  assign n42291 = ~n42240 & n42246 ;
  assign n42292 = ~n42253 & n42291 ;
  assign n42293 = ~n42259 & n42292 ;
  assign n42294 = n42271 & n42293 ;
  assign n42295 = n42259 & n42280 ;
  assign n42296 = ~n42294 & ~n42295 ;
  assign n42289 = n42263 & n42279 ;
  assign n42290 = ~n42259 & n42289 ;
  assign n42298 = n42271 & ~n42291 ;
  assign n42297 = ~n42246 & ~n42260 ;
  assign n42299 = ~n42262 & ~n42297 ;
  assign n42300 = n42298 & n42299 ;
  assign n42319 = ~n42290 & ~n42300 ;
  assign n42320 = n42296 & n42319 ;
  assign n42321 = ~n42288 & n42320 ;
  assign n42322 = ~n42318 & n42321 ;
  assign n42323 = \u1_L4_reg[11]/P0001  & ~n42322 ;
  assign n42324 = ~\u1_L4_reg[11]/P0001  & n42322 ;
  assign n42325 = ~n42323 & ~n42324 ;
  assign n42339 = decrypt_pad & ~\u1_uk_K_r4_reg[4]/NET0131  ;
  assign n42340 = ~decrypt_pad & ~\u1_uk_K_r4_reg[10]/NET0131  ;
  assign n42341 = ~n42339 & ~n42340 ;
  assign n42342 = \u1_R4_reg[13]/NET0131  & ~n42341 ;
  assign n42343 = ~\u1_R4_reg[13]/NET0131  & n42341 ;
  assign n42344 = ~n42342 & ~n42343 ;
  assign n42326 = decrypt_pad & ~\u1_uk_K_r4_reg[26]/NET0131  ;
  assign n42327 = ~decrypt_pad & ~\u1_uk_K_r4_reg[32]/NET0131  ;
  assign n42328 = ~n42326 & ~n42327 ;
  assign n42329 = \u1_R4_reg[17]/NET0131  & ~n42328 ;
  assign n42330 = ~\u1_R4_reg[17]/NET0131  & n42328 ;
  assign n42331 = ~n42329 & ~n42330 ;
  assign n42332 = decrypt_pad & ~\u1_uk_K_r4_reg[10]/NET0131  ;
  assign n42333 = ~decrypt_pad & ~\u1_uk_K_r4_reg[48]/NET0131  ;
  assign n42334 = ~n42332 & ~n42333 ;
  assign n42335 = \u1_R4_reg[12]/NET0131  & ~n42334 ;
  assign n42336 = ~\u1_R4_reg[12]/NET0131  & n42334 ;
  assign n42337 = ~n42335 & ~n42336 ;
  assign n42371 = n42331 & n42337 ;
  assign n42372 = n42344 & n42371 ;
  assign n42363 = ~n42331 & ~n42344 ;
  assign n42364 = ~n42337 & n42363 ;
  assign n42365 = decrypt_pad & ~\u1_uk_K_r4_reg[13]/NET0131  ;
  assign n42366 = ~decrypt_pad & ~\u1_uk_K_r4_reg[19]/NET0131  ;
  assign n42367 = ~n42365 & ~n42366 ;
  assign n42368 = \u1_R4_reg[15]/NET0131  & ~n42367 ;
  assign n42369 = ~\u1_R4_reg[15]/NET0131  & n42367 ;
  assign n42370 = ~n42368 & ~n42369 ;
  assign n42373 = ~n42364 & n42370 ;
  assign n42374 = ~n42372 & n42373 ;
  assign n42346 = decrypt_pad & ~\u1_uk_K_r4_reg[5]/NET0131  ;
  assign n42347 = ~decrypt_pad & ~\u1_uk_K_r4_reg[11]/NET0131  ;
  assign n42348 = ~n42346 & ~n42347 ;
  assign n42349 = \u1_R4_reg[14]/NET0131  & ~n42348 ;
  assign n42350 = ~\u1_R4_reg[14]/NET0131  & n42348 ;
  assign n42351 = ~n42349 & ~n42350 ;
  assign n42376 = ~n42331 & n42337 ;
  assign n42377 = n42351 & n42376 ;
  assign n42375 = n42331 & ~n42344 ;
  assign n42378 = ~n42370 & ~n42375 ;
  assign n42379 = ~n42377 & n42378 ;
  assign n42380 = ~n42374 & ~n42379 ;
  assign n42338 = ~n42331 & ~n42337 ;
  assign n42345 = n42338 & n42344 ;
  assign n42352 = n42345 & n42351 ;
  assign n42353 = ~n42331 & ~n42351 ;
  assign n42354 = ~n42337 & n42353 ;
  assign n42355 = ~n42344 & n42354 ;
  assign n42356 = ~n42352 & ~n42355 ;
  assign n42384 = n42337 & ~n42351 ;
  assign n42385 = ~n42344 & n42384 ;
  assign n42386 = n42331 & n42385 ;
  assign n42357 = decrypt_pad & ~\u1_uk_K_r4_reg[46]/NET0131  ;
  assign n42358 = ~decrypt_pad & ~\u1_uk_K_r4_reg[27]/P0001  ;
  assign n42359 = ~n42357 & ~n42358 ;
  assign n42360 = \u1_R4_reg[16]/NET0131  & ~n42359 ;
  assign n42361 = ~\u1_R4_reg[16]/NET0131  & n42359 ;
  assign n42362 = ~n42360 & ~n42361 ;
  assign n42381 = n42344 & n42370 ;
  assign n42382 = n42351 & n42381 ;
  assign n42383 = ~n42337 & n42382 ;
  assign n42387 = ~n42362 & ~n42383 ;
  assign n42388 = ~n42386 & n42387 ;
  assign n42389 = n42356 & n42388 ;
  assign n42390 = ~n42380 & n42389 ;
  assign n42391 = n42364 & ~n42370 ;
  assign n42392 = n42351 & n42391 ;
  assign n42393 = n42331 & ~n42337 ;
  assign n42405 = ~n42344 & n42370 ;
  assign n42406 = n42393 & n42405 ;
  assign n42404 = n42376 & n42381 ;
  assign n42407 = n42362 & ~n42404 ;
  assign n42408 = ~n42406 & n42407 ;
  assign n42394 = n42344 & ~n42351 ;
  assign n42395 = n42393 & n42394 ;
  assign n42396 = n42337 & n42344 ;
  assign n42397 = n42331 & n42351 ;
  assign n42398 = n42396 & n42397 ;
  assign n42399 = ~n42395 & ~n42398 ;
  assign n42400 = ~n42351 & ~n42370 ;
  assign n42401 = ~n42337 & ~n42344 ;
  assign n42402 = ~n42396 & ~n42401 ;
  assign n42403 = n42400 & n42402 ;
  assign n42409 = n42399 & ~n42403 ;
  assign n42410 = n42408 & n42409 ;
  assign n42411 = ~n42392 & n42410 ;
  assign n42412 = ~n42390 & ~n42411 ;
  assign n42413 = ~n42370 & ~n42395 ;
  assign n42414 = ~n42344 & n42377 ;
  assign n42415 = n42370 & ~n42414 ;
  assign n42416 = ~n42355 & n42415 ;
  assign n42417 = ~n42413 & ~n42416 ;
  assign n42418 = ~n42351 & n42404 ;
  assign n42419 = ~n42417 & ~n42418 ;
  assign n42420 = ~n42412 & n42419 ;
  assign n42421 = ~\u1_L4_reg[20]/NET0131  & ~n42420 ;
  assign n42422 = \u1_L4_reg[20]/NET0131  & n42420 ;
  assign n42423 = ~n42421 & ~n42422 ;
  assign n42424 = decrypt_pad & ~\u1_uk_K_r4_reg[52]/NET0131  ;
  assign n42425 = ~decrypt_pad & ~\u1_uk_K_r4_reg[1]/NET0131  ;
  assign n42426 = ~n42424 & ~n42425 ;
  assign n42427 = \u1_R4_reg[28]/NET0131  & ~n42426 ;
  assign n42428 = ~\u1_R4_reg[28]/NET0131  & n42426 ;
  assign n42429 = ~n42427 & ~n42428 ;
  assign n42437 = decrypt_pad & ~\u1_uk_K_r4_reg[21]/NET0131  ;
  assign n42438 = ~decrypt_pad & ~\u1_uk_K_r4_reg[29]/NET0131  ;
  assign n42439 = ~n42437 & ~n42438 ;
  assign n42440 = \u1_R4_reg[30]/NET0131  & ~n42439 ;
  assign n42441 = ~\u1_R4_reg[30]/NET0131  & n42439 ;
  assign n42442 = ~n42440 & ~n42441 ;
  assign n42430 = decrypt_pad & ~\u1_uk_K_r4_reg[51]/NET0131  ;
  assign n42431 = ~decrypt_pad & ~\u1_uk_K_r4_reg[28]/NET0131  ;
  assign n42432 = ~n42430 & ~n42431 ;
  assign n42433 = \u1_R4_reg[29]/NET0131  & ~n42432 ;
  assign n42434 = ~\u1_R4_reg[29]/NET0131  & n42432 ;
  assign n42435 = ~n42433 & ~n42434 ;
  assign n42444 = decrypt_pad & ~\u1_uk_K_r4_reg[36]/NET0131  ;
  assign n42445 = ~decrypt_pad & ~\u1_uk_K_r4_reg[44]/NET0131  ;
  assign n42446 = ~n42444 & ~n42445 ;
  assign n42447 = \u1_R4_reg[1]/NET0131  & ~n42446 ;
  assign n42448 = ~\u1_R4_reg[1]/NET0131  & n42446 ;
  assign n42449 = ~n42447 & ~n42448 ;
  assign n42469 = n42435 & ~n42449 ;
  assign n42470 = ~n42442 & n42469 ;
  assign n42454 = decrypt_pad & ~\u1_uk_K_r4_reg[9]/NET0131  ;
  assign n42455 = ~decrypt_pad & ~\u1_uk_K_r4_reg[45]/NET0131  ;
  assign n42456 = ~n42454 & ~n42455 ;
  assign n42457 = \u1_R4_reg[31]/P0001  & ~n42456 ;
  assign n42458 = ~\u1_R4_reg[31]/P0001  & n42456 ;
  assign n42459 = ~n42457 & ~n42458 ;
  assign n42466 = ~n42442 & ~n42459 ;
  assign n42467 = n42442 & n42449 ;
  assign n42468 = n42435 & n42467 ;
  assign n42471 = ~n42466 & ~n42468 ;
  assign n42472 = ~n42470 & n42471 ;
  assign n42473 = n42429 & ~n42472 ;
  assign n42436 = n42429 & ~n42435 ;
  assign n42443 = n42436 & n42442 ;
  assign n42450 = n42443 & ~n42449 ;
  assign n42451 = ~n42429 & n42449 ;
  assign n42452 = ~n42435 & n42451 ;
  assign n42453 = ~n42450 & ~n42452 ;
  assign n42460 = ~n42453 & n42459 ;
  assign n42461 = ~n42429 & n42442 ;
  assign n42462 = ~n42449 & ~n42461 ;
  assign n42463 = ~n42435 & n42449 ;
  assign n42464 = ~n42459 & ~n42463 ;
  assign n42465 = ~n42462 & n42464 ;
  assign n42474 = ~n42460 & ~n42465 ;
  assign n42475 = ~n42473 & n42474 ;
  assign n42476 = decrypt_pad & ~\u1_uk_K_r4_reg[15]/NET0131  ;
  assign n42477 = ~decrypt_pad & ~\u1_uk_K_r4_reg[23]/P0001  ;
  assign n42478 = ~n42476 & ~n42477 ;
  assign n42479 = \u1_R4_reg[32]/NET0131  & ~n42478 ;
  assign n42480 = ~\u1_R4_reg[32]/NET0131  & n42478 ;
  assign n42481 = ~n42479 & ~n42480 ;
  assign n42482 = ~n42475 & ~n42481 ;
  assign n42502 = n42429 & n42470 ;
  assign n42489 = n42429 & ~n42442 ;
  assign n42490 = ~n42469 & ~n42489 ;
  assign n42503 = n42459 & ~n42490 ;
  assign n42504 = ~n42502 & n42503 ;
  assign n42505 = ~n42429 & n42468 ;
  assign n42506 = ~n42435 & ~n42442 ;
  assign n42507 = ~n42429 & n42506 ;
  assign n42508 = ~n42459 & n42507 ;
  assign n42509 = ~n42505 & ~n42508 ;
  assign n42510 = ~n42504 & n42509 ;
  assign n42511 = n42481 & ~n42510 ;
  assign n42487 = n42429 & ~n42449 ;
  assign n42488 = n42435 & ~n42442 ;
  assign n42491 = ~n42487 & ~n42488 ;
  assign n42492 = ~n42490 & n42491 ;
  assign n42483 = ~n42435 & ~n42449 ;
  assign n42484 = ~n42429 & n42483 ;
  assign n42485 = ~n42442 & n42484 ;
  assign n42486 = n42461 & n42463 ;
  assign n42493 = ~n42485 & ~n42486 ;
  assign n42494 = ~n42492 & n42493 ;
  assign n42495 = n42459 & ~n42494 ;
  assign n42496 = n42429 & n42435 ;
  assign n42497 = ~n42449 & n42496 ;
  assign n42498 = n42466 & n42497 ;
  assign n42499 = n42442 & ~n42459 ;
  assign n42500 = n42436 & n42481 ;
  assign n42501 = n42499 & n42500 ;
  assign n42512 = ~n42498 & ~n42501 ;
  assign n42513 = ~n42495 & n42512 ;
  assign n42514 = ~n42511 & n42513 ;
  assign n42515 = ~n42482 & n42514 ;
  assign n42516 = \u1_L4_reg[5]/NET0131  & ~n42515 ;
  assign n42517 = ~\u1_L4_reg[5]/NET0131  & n42515 ;
  assign n42518 = ~n42516 & ~n42517 ;
  assign n42519 = n42376 & ~n42394 ;
  assign n42520 = n42413 & ~n42519 ;
  assign n42521 = n42370 & ~n42386 ;
  assign n42522 = ~n42345 & n42521 ;
  assign n42523 = ~n42520 & ~n42522 ;
  assign n42524 = n42397 & ~n42402 ;
  assign n42525 = ~n42523 & ~n42524 ;
  assign n42526 = n42362 & ~n42525 ;
  assign n42527 = n42371 & n42400 ;
  assign n42533 = n42344 & n42384 ;
  assign n42534 = ~n42527 & ~n42533 ;
  assign n42535 = ~n42391 & n42534 ;
  assign n42528 = n42370 & n42393 ;
  assign n42529 = ~n42351 & n42528 ;
  assign n42530 = n42331 & ~n42351 ;
  assign n42531 = n42337 & n42405 ;
  assign n42532 = ~n42530 & n42531 ;
  assign n42536 = ~n42529 & ~n42532 ;
  assign n42537 = n42535 & n42536 ;
  assign n42538 = n42356 & n42537 ;
  assign n42539 = ~n42362 & ~n42538 ;
  assign n42540 = ~n42355 & ~n42524 ;
  assign n42541 = ~n42370 & ~n42540 ;
  assign n42542 = ~n42383 & ~n42418 ;
  assign n42543 = ~n42541 & n42542 ;
  assign n42544 = ~n42539 & n42543 ;
  assign n42545 = ~n42526 & n42544 ;
  assign n42546 = ~\u1_L4_reg[10]/NET0131  & ~n42545 ;
  assign n42547 = \u1_L4_reg[10]/NET0131  & n42545 ;
  assign n42548 = ~n42546 & ~n42547 ;
  assign n42559 = ~n42082 & n42112 ;
  assign n42549 = ~n42068 & n42106 ;
  assign n42550 = ~n42074 & n42549 ;
  assign n42557 = ~n42084 & ~n42104 ;
  assign n42558 = n42118 & ~n42557 ;
  assign n42562 = ~n42550 & ~n42558 ;
  assign n42563 = ~n42559 & n42562 ;
  assign n42551 = ~n42055 & n42068 ;
  assign n42552 = ~n42074 & n42551 ;
  assign n42553 = n42055 & n42093 ;
  assign n42554 = ~n42552 & ~n42553 ;
  assign n42555 = ~n42061 & ~n42554 ;
  assign n42556 = ~n42082 & n42093 ;
  assign n42560 = ~n42049 & ~n42076 ;
  assign n42561 = ~n42556 & n42560 ;
  assign n42564 = ~n42555 & n42561 ;
  assign n42565 = n42563 & n42564 ;
  assign n42568 = ~n42118 & ~n42551 ;
  assign n42567 = ~n42068 & n42082 ;
  assign n42569 = n42086 & ~n42567 ;
  assign n42570 = ~n42568 & n42569 ;
  assign n42566 = n42074 & n42549 ;
  assign n42575 = n42049 & ~n42566 ;
  assign n42576 = ~n42570 & n42575 ;
  assign n42571 = ~n42074 & ~n42121 ;
  assign n42572 = n42061 & n42068 ;
  assign n42573 = ~n42117 & ~n42572 ;
  assign n42574 = n42082 & ~n42573 ;
  assign n42577 = ~n42571 & ~n42574 ;
  assign n42578 = n42576 & n42577 ;
  assign n42579 = ~n42565 & ~n42578 ;
  assign n42580 = \u1_L4_reg[12]/NET0131  & n42579 ;
  assign n42581 = ~\u1_L4_reg[12]/NET0131  & ~n42579 ;
  assign n42582 = ~n42580 & ~n42581 ;
  assign n42583 = decrypt_pad & ~\u1_uk_K_r4_reg[0]/P0001  ;
  assign n42584 = ~decrypt_pad & ~\u1_uk_K_r4_reg[8]/NET0131  ;
  assign n42585 = ~n42583 & ~n42584 ;
  assign n42586 = \u1_R4_reg[20]/NET0131  & ~n42585 ;
  assign n42587 = ~\u1_R4_reg[20]/NET0131  & n42585 ;
  assign n42588 = ~n42586 & ~n42587 ;
  assign n42625 = decrypt_pad & ~\u1_uk_K_r4_reg[16]/NET0131  ;
  assign n42626 = ~decrypt_pad & ~\u1_uk_K_r4_reg[52]/NET0131  ;
  assign n42627 = ~n42625 & ~n42626 ;
  assign n42628 = \u1_R4_reg[19]/NET0131  & ~n42627 ;
  assign n42629 = ~\u1_R4_reg[19]/NET0131  & n42627 ;
  assign n42630 = ~n42628 & ~n42629 ;
  assign n42602 = decrypt_pad & ~\u1_uk_K_r4_reg[29]/NET0131  ;
  assign n42603 = ~decrypt_pad & ~\u1_uk_K_r4_reg[37]/NET0131  ;
  assign n42604 = ~n42602 & ~n42603 ;
  assign n42605 = \u1_R4_reg[18]/NET0131  & ~n42604 ;
  assign n42606 = ~\u1_R4_reg[18]/NET0131  & n42604 ;
  assign n42607 = ~n42605 & ~n42606 ;
  assign n42589 = decrypt_pad & ~\u1_uk_K_r4_reg[44]/NET0131  ;
  assign n42590 = ~decrypt_pad & ~\u1_uk_K_r4_reg[21]/NET0131  ;
  assign n42591 = ~n42589 & ~n42590 ;
  assign n42592 = \u1_R4_reg[16]/NET0131  & ~n42591 ;
  assign n42593 = ~\u1_R4_reg[16]/NET0131  & n42591 ;
  assign n42594 = ~n42592 & ~n42593 ;
  assign n42595 = decrypt_pad & ~\u1_uk_K_r4_reg[1]/NET0131  ;
  assign n42596 = ~decrypt_pad & ~\u1_uk_K_r4_reg[9]/NET0131  ;
  assign n42597 = ~n42595 & ~n42596 ;
  assign n42598 = \u1_R4_reg[21]/NET0131  & ~n42597 ;
  assign n42599 = ~\u1_R4_reg[21]/NET0131  & n42597 ;
  assign n42600 = ~n42598 & ~n42599 ;
  assign n42601 = n42594 & ~n42600 ;
  assign n42608 = decrypt_pad & ~\u1_uk_K_r4_reg[35]/NET0131  ;
  assign n42609 = ~decrypt_pad & ~\u1_uk_K_r4_reg[43]/NET0131  ;
  assign n42610 = ~n42608 & ~n42609 ;
  assign n42611 = \u1_R4_reg[17]/NET0131  & ~n42610 ;
  assign n42612 = ~\u1_R4_reg[17]/NET0131  & n42610 ;
  assign n42613 = ~n42611 & ~n42612 ;
  assign n42662 = n42601 & ~n42613 ;
  assign n42663 = ~n42607 & n42662 ;
  assign n42614 = ~n42607 & n42613 ;
  assign n42632 = n42594 & n42600 ;
  assign n42664 = n42614 & n42632 ;
  assign n42646 = ~n42594 & n42600 ;
  assign n42647 = ~n42613 & n42646 ;
  assign n42622 = ~n42600 & n42613 ;
  assign n42661 = n42607 & n42622 ;
  assign n42665 = ~n42647 & ~n42661 ;
  assign n42666 = ~n42664 & n42665 ;
  assign n42667 = ~n42663 & n42666 ;
  assign n42668 = ~n42630 & ~n42667 ;
  assign n42618 = ~n42594 & n42614 ;
  assign n42619 = n42594 & n42607 ;
  assign n42620 = n42600 & ~n42619 ;
  assign n42657 = ~n42601 & ~n42622 ;
  assign n42658 = ~n42620 & n42657 ;
  assign n42659 = ~n42618 & ~n42658 ;
  assign n42660 = n42630 & ~n42659 ;
  assign n42669 = n42600 & ~n42607 ;
  assign n42670 = ~n42601 & ~n42669 ;
  assign n42640 = ~n42594 & ~n42613 ;
  assign n42671 = n42607 & n42613 ;
  assign n42672 = ~n42640 & ~n42671 ;
  assign n42673 = n42670 & n42672 ;
  assign n42674 = ~n42660 & ~n42673 ;
  assign n42675 = ~n42668 & n42674 ;
  assign n42676 = ~n42588 & ~n42675 ;
  assign n42621 = ~n42618 & n42620 ;
  assign n42623 = n42594 & n42622 ;
  assign n42624 = ~n42621 & ~n42623 ;
  assign n42631 = ~n42624 & n42630 ;
  assign n42615 = n42607 & ~n42613 ;
  assign n42616 = ~n42614 & ~n42615 ;
  assign n42617 = n42601 & ~n42616 ;
  assign n42633 = n42607 & n42630 ;
  assign n42634 = n42632 & ~n42633 ;
  assign n42635 = n42616 & n42634 ;
  assign n42636 = ~n42617 & ~n42635 ;
  assign n42637 = ~n42631 & n42636 ;
  assign n42638 = n42588 & ~n42637 ;
  assign n42641 = ~n42600 & n42640 ;
  assign n42642 = n42607 & n42641 ;
  assign n42639 = ~n42607 & n42623 ;
  assign n42643 = n42630 & ~n42639 ;
  assign n42644 = ~n42642 & n42643 ;
  assign n42650 = n42613 & n42646 ;
  assign n42651 = ~n42641 & ~n42650 ;
  assign n42652 = n42588 & ~n42607 ;
  assign n42653 = ~n42651 & n42652 ;
  assign n42645 = ~n42594 & n42622 ;
  assign n42648 = ~n42645 & ~n42647 ;
  assign n42649 = n42607 & ~n42648 ;
  assign n42654 = ~n42630 & ~n42649 ;
  assign n42655 = ~n42653 & n42654 ;
  assign n42656 = ~n42644 & ~n42655 ;
  assign n42677 = ~n42638 & ~n42656 ;
  assign n42678 = ~n42676 & n42677 ;
  assign n42679 = ~\u1_L4_reg[14]/NET0131  & ~n42678 ;
  assign n42680 = \u1_L4_reg[14]/NET0131  & n42678 ;
  assign n42681 = ~n42679 & ~n42680 ;
  assign n42682 = ~n42470 & ~n42496 ;
  assign n42683 = ~n42452 & n42682 ;
  assign n42684 = n42459 & ~n42683 ;
  assign n42685 = n42483 & n42489 ;
  assign n42686 = ~n42684 & ~n42685 ;
  assign n42687 = ~n42481 & ~n42686 ;
  assign n42691 = n42463 & n42499 ;
  assign n42688 = n42429 & n42488 ;
  assign n42690 = n42461 & n42469 ;
  assign n42693 = ~n42688 & ~n42690 ;
  assign n42694 = ~n42691 & n42693 ;
  assign n42689 = n42459 & n42484 ;
  assign n42692 = n42443 & n42449 ;
  assign n42695 = ~n42689 & ~n42692 ;
  assign n42696 = n42694 & n42695 ;
  assign n42697 = n42481 & ~n42696 ;
  assign n42699 = n42436 & ~n42481 ;
  assign n42698 = n42451 & n42488 ;
  assign n42701 = ~n42690 & ~n42698 ;
  assign n42702 = ~n42699 & n42701 ;
  assign n42700 = ~n42443 & ~n42459 ;
  assign n42703 = ~n42485 & n42700 ;
  assign n42704 = n42702 & n42703 ;
  assign n42705 = ~n42442 & n42452 ;
  assign n42706 = n42459 & ~n42505 ;
  assign n42707 = ~n42705 & n42706 ;
  assign n42708 = ~n42704 & ~n42707 ;
  assign n42709 = ~n42697 & ~n42708 ;
  assign n42710 = ~n42687 & n42709 ;
  assign n42711 = \u1_L4_reg[15]/P0001  & n42710 ;
  assign n42712 = ~\u1_L4_reg[15]/P0001  & ~n42710 ;
  assign n42713 = ~n42711 & ~n42712 ;
  assign n42729 = ~n42353 & ~n42375 ;
  assign n42730 = n42337 & ~n42729 ;
  assign n42731 = ~n42370 & ~n42730 ;
  assign n42732 = ~n42354 & n42415 ;
  assign n42733 = ~n42731 & ~n42732 ;
  assign n42734 = n42376 & n42394 ;
  assign n42735 = n42399 & ~n42734 ;
  assign n42736 = ~n42733 & n42735 ;
  assign n42737 = ~n42362 & ~n42736 ;
  assign n42721 = n42344 & n42393 ;
  assign n42722 = ~n42376 & n42394 ;
  assign n42723 = ~n42721 & ~n42722 ;
  assign n42724 = ~n42370 & ~n42723 ;
  assign n42719 = n42344 & n42377 ;
  assign n42725 = n42351 & n42401 ;
  assign n42726 = ~n42719 & ~n42725 ;
  assign n42727 = ~n42724 & n42726 ;
  assign n42728 = n42362 & ~n42727 ;
  assign n42714 = ~n42352 & ~n42524 ;
  assign n42715 = n42370 & ~n42714 ;
  assign n42720 = ~n42370 & n42719 ;
  assign n42716 = ~n42375 & ~n42385 ;
  assign n42717 = n42362 & n42370 ;
  assign n42718 = ~n42716 & n42717 ;
  assign n42738 = ~n42392 & ~n42718 ;
  assign n42739 = ~n42720 & n42738 ;
  assign n42740 = ~n42715 & n42739 ;
  assign n42741 = ~n42728 & n42740 ;
  assign n42742 = ~n42737 & n42741 ;
  assign n42743 = ~\u1_L4_reg[1]/NET0131  & ~n42742 ;
  assign n42744 = \u1_L4_reg[1]/NET0131  & n42742 ;
  assign n42745 = ~n42743 & ~n42744 ;
  assign n42748 = ~n42152 & ~n42174 ;
  assign n42749 = ~n42159 & ~n42748 ;
  assign n42753 = n42167 & n42748 ;
  assign n42754 = ~n42749 & ~n42753 ;
  assign n42755 = n42146 & ~n42754 ;
  assign n42752 = n42159 & n42214 ;
  assign n42750 = ~n42146 & ~n42193 ;
  assign n42751 = ~n42749 & n42750 ;
  assign n42746 = n42152 & n42174 ;
  assign n42747 = n42165 & n42746 ;
  assign n42756 = n42140 & ~n42747 ;
  assign n42757 = ~n42751 & n42756 ;
  assign n42758 = ~n42752 & n42757 ;
  assign n42759 = ~n42755 & n42758 ;
  assign n42762 = n42159 & ~n42180 ;
  assign n42763 = ~n42201 & ~n42746 ;
  assign n42764 = ~n42762 & n42763 ;
  assign n42765 = ~n42146 & ~n42764 ;
  assign n42766 = n42152 & n42185 ;
  assign n42770 = n42146 & ~n42766 ;
  assign n42767 = n42174 & n42201 ;
  assign n42768 = ~n42152 & n42767 ;
  assign n42769 = ~n42178 & ~n42215 ;
  assign n42771 = ~n42768 & n42769 ;
  assign n42772 = n42770 & n42771 ;
  assign n42773 = ~n42765 & ~n42772 ;
  assign n42760 = ~n42165 & n42746 ;
  assign n42761 = n42159 & n42760 ;
  assign n42774 = ~n42140 & ~n42212 ;
  assign n42775 = ~n42761 & n42774 ;
  assign n42776 = ~n42773 & n42775 ;
  assign n42777 = ~n42759 & ~n42776 ;
  assign n42778 = ~\u1_L4_reg[17]/NET0131  & n42777 ;
  assign n42779 = \u1_L4_reg[17]/NET0131  & ~n42777 ;
  assign n42780 = ~n42778 & ~n42779 ;
  assign n42783 = ~n42463 & n42489 ;
  assign n42784 = ~n42459 & ~n42783 ;
  assign n42785 = ~n42692 & n42784 ;
  assign n42787 = ~n42496 & ~n42506 ;
  assign n42788 = ~n42783 & ~n42787 ;
  assign n42786 = n42435 & n42451 ;
  assign n42789 = n42459 & ~n42786 ;
  assign n42790 = ~n42788 & n42789 ;
  assign n42791 = ~n42785 & ~n42790 ;
  assign n42781 = ~n42484 & ~n42497 ;
  assign n42782 = n42442 & ~n42781 ;
  assign n42792 = n42481 & ~n42705 ;
  assign n42793 = ~n42782 & n42792 ;
  assign n42794 = ~n42791 & n42793 ;
  assign n42795 = ~n42497 & ~n42507 ;
  assign n42796 = ~n42443 & n42795 ;
  assign n42797 = n42459 & ~n42796 ;
  assign n42801 = n42435 & n42461 ;
  assign n42805 = ~n42481 & ~n42801 ;
  assign n42806 = ~n42450 & n42805 ;
  assign n42802 = n42429 & n42449 ;
  assign n42803 = ~n42466 & ~n42488 ;
  assign n42804 = n42802 & ~n42803 ;
  assign n42798 = ~n42429 & ~n42459 ;
  assign n42799 = ~n42467 & ~n42469 ;
  assign n42800 = n42798 & ~n42799 ;
  assign n42807 = ~n42485 & ~n42800 ;
  assign n42808 = ~n42804 & n42807 ;
  assign n42809 = n42806 & n42808 ;
  assign n42810 = ~n42797 & n42809 ;
  assign n42811 = ~n42794 & ~n42810 ;
  assign n42812 = ~\u1_L4_reg[21]/NET0131  & n42811 ;
  assign n42813 = \u1_L4_reg[21]/NET0131  & ~n42811 ;
  assign n42814 = ~n42812 & ~n42813 ;
  assign n42827 = ~n42600 & ~n42614 ;
  assign n42828 = ~n42619 & n42827 ;
  assign n42826 = n42613 & n42632 ;
  assign n42829 = ~n42640 & ~n42826 ;
  assign n42830 = ~n42828 & n42829 ;
  assign n42831 = n42630 & ~n42830 ;
  assign n42833 = ~n42613 & n42632 ;
  assign n42834 = ~n42618 & ~n42833 ;
  assign n42835 = ~n42630 & ~n42834 ;
  assign n42832 = n42613 & n42669 ;
  assign n42836 = n42619 & n42622 ;
  assign n42837 = ~n42832 & ~n42836 ;
  assign n42838 = ~n42835 & n42837 ;
  assign n42839 = ~n42831 & n42838 ;
  assign n42840 = n42588 & ~n42839 ;
  assign n42820 = ~n42622 & n42630 ;
  assign n42819 = ~n42630 & ~n42640 ;
  assign n42821 = ~n42607 & ~n42819 ;
  assign n42822 = ~n42820 & n42821 ;
  assign n42815 = n42607 & n42650 ;
  assign n42816 = ~n42594 & n42671 ;
  assign n42817 = ~n42662 & ~n42816 ;
  assign n42818 = ~n42630 & ~n42817 ;
  assign n42823 = ~n42815 & ~n42818 ;
  assign n42824 = ~n42822 & n42823 ;
  assign n42825 = ~n42588 & ~n42824 ;
  assign n42843 = ~n42642 & ~n42836 ;
  assign n42844 = ~n42607 & n42646 ;
  assign n42845 = ~n42613 & n42844 ;
  assign n42846 = n42843 & ~n42845 ;
  assign n42847 = n42630 & ~n42846 ;
  assign n42841 = n42594 & ~n42630 ;
  assign n42842 = n42615 & n42841 ;
  assign n42848 = ~n42664 & ~n42842 ;
  assign n42849 = ~n42847 & n42848 ;
  assign n42850 = ~n42825 & n42849 ;
  assign n42851 = ~n42840 & n42850 ;
  assign n42852 = ~\u1_L4_reg[25]/NET0131  & ~n42851 ;
  assign n42853 = \u1_L4_reg[25]/NET0131  & n42851 ;
  assign n42854 = ~n42852 & ~n42853 ;
  assign n42855 = decrypt_pad & ~\u1_uk_K_r4_reg[20]/NET0131  ;
  assign n42856 = ~decrypt_pad & ~\u1_uk_K_r4_reg[26]/NET0131  ;
  assign n42857 = ~n42855 & ~n42856 ;
  assign n42858 = \u1_R4_reg[8]/NET0131  & ~n42857 ;
  assign n42859 = ~\u1_R4_reg[8]/NET0131  & n42857 ;
  assign n42860 = ~n42858 & ~n42859 ;
  assign n42861 = decrypt_pad & ~\u1_uk_K_r4_reg[54]/NET0131  ;
  assign n42862 = ~decrypt_pad & ~\u1_uk_K_r4_reg[3]/NET0131  ;
  assign n42863 = ~n42861 & ~n42862 ;
  assign n42864 = \u1_R4_reg[7]/NET0131  & ~n42863 ;
  assign n42865 = ~\u1_R4_reg[7]/NET0131  & n42863 ;
  assign n42866 = ~n42864 & ~n42865 ;
  assign n42880 = decrypt_pad & ~\u1_uk_K_r4_reg[12]/NET0131  ;
  assign n42881 = ~decrypt_pad & ~\u1_uk_K_r4_reg[18]/NET0131  ;
  assign n42882 = ~n42880 & ~n42881 ;
  assign n42883 = \u1_R4_reg[5]/NET0131  & ~n42882 ;
  assign n42884 = ~\u1_R4_reg[5]/NET0131  & n42882 ;
  assign n42885 = ~n42883 & ~n42884 ;
  assign n42867 = decrypt_pad & ~\u1_uk_K_r4_reg[33]/NET0131  ;
  assign n42868 = ~decrypt_pad & ~\u1_uk_K_r4_reg[39]/NET0131  ;
  assign n42869 = ~n42867 & ~n42868 ;
  assign n42870 = \u1_R4_reg[4]/NET0131  & ~n42869 ;
  assign n42871 = ~\u1_R4_reg[4]/NET0131  & n42869 ;
  assign n42872 = ~n42870 & ~n42871 ;
  assign n42873 = decrypt_pad & ~\u1_uk_K_r4_reg[25]/NET0131  ;
  assign n42874 = ~decrypt_pad & ~\u1_uk_K_r4_reg[6]/NET0131  ;
  assign n42875 = ~n42873 & ~n42874 ;
  assign n42876 = \u1_R4_reg[9]/NET0131  & ~n42875 ;
  assign n42877 = ~\u1_R4_reg[9]/NET0131  & n42875 ;
  assign n42878 = ~n42876 & ~n42877 ;
  assign n42895 = ~n42872 & n42878 ;
  assign n42896 = ~n42885 & n42895 ;
  assign n42887 = decrypt_pad & ~\u1_uk_K_r4_reg[3]/NET0131  ;
  assign n42888 = ~decrypt_pad & ~\u1_uk_K_r4_reg[41]/NET0131  ;
  assign n42889 = ~n42887 & ~n42888 ;
  assign n42890 = \u1_R4_reg[6]/NET0131  & ~n42889 ;
  assign n42891 = ~\u1_R4_reg[6]/NET0131  & n42889 ;
  assign n42892 = ~n42890 & ~n42891 ;
  assign n42897 = n42872 & n42885 ;
  assign n42898 = n42872 & ~n42878 ;
  assign n42899 = ~n42897 & ~n42898 ;
  assign n42900 = n42892 & ~n42899 ;
  assign n42901 = ~n42896 & ~n42900 ;
  assign n42902 = ~n42866 & ~n42901 ;
  assign n42903 = ~n42878 & n42885 ;
  assign n42904 = ~n42896 & ~n42903 ;
  assign n42905 = ~n42892 & ~n42904 ;
  assign n42879 = n42872 & n42878 ;
  assign n42886 = n42879 & ~n42885 ;
  assign n42893 = n42886 & n42892 ;
  assign n42894 = n42866 & n42893 ;
  assign n42906 = ~n42866 & ~n42885 ;
  assign n42907 = n42878 & ~n42892 ;
  assign n42908 = n42906 & n42907 ;
  assign n42909 = n42885 & n42892 ;
  assign n42910 = n42895 & n42909 ;
  assign n42911 = ~n42908 & ~n42910 ;
  assign n42912 = ~n42894 & n42911 ;
  assign n42913 = ~n42905 & n42912 ;
  assign n42914 = ~n42902 & n42913 ;
  assign n42915 = ~n42860 & ~n42914 ;
  assign n42932 = ~n42872 & ~n42878 ;
  assign n42933 = ~n42893 & ~n42932 ;
  assign n42934 = n42860 & ~n42933 ;
  assign n42925 = ~n42885 & n42892 ;
  assign n42935 = n42895 & ~n42925 ;
  assign n42936 = ~n42934 & ~n42935 ;
  assign n42927 = n42885 & ~n42892 ;
  assign n42937 = ~n42866 & ~n42927 ;
  assign n42938 = ~n42936 & n42937 ;
  assign n42916 = ~n42885 & n42898 ;
  assign n42917 = ~n42892 & n42916 ;
  assign n42918 = n42866 & n42885 ;
  assign n42919 = ~n42872 & n42892 ;
  assign n42920 = n42918 & ~n42919 ;
  assign n42921 = n42897 & n42907 ;
  assign n42922 = ~n42920 & ~n42921 ;
  assign n42923 = ~n42917 & n42922 ;
  assign n42924 = n42860 & ~n42923 ;
  assign n42928 = n42872 & ~n42927 ;
  assign n42926 = ~n42872 & ~n42925 ;
  assign n42929 = n42866 & ~n42895 ;
  assign n42930 = ~n42926 & n42929 ;
  assign n42931 = ~n42928 & n42930 ;
  assign n42939 = ~n42924 & ~n42931 ;
  assign n42940 = ~n42938 & n42939 ;
  assign n42941 = ~n42915 & n42940 ;
  assign n42942 = \u1_L4_reg[2]/NET0131  & n42941 ;
  assign n42943 = ~\u1_L4_reg[2]/NET0131  & ~n42941 ;
  assign n42944 = ~n42942 & ~n42943 ;
  assign n42945 = ~n42395 & n42521 ;
  assign n42946 = ~n42331 & n42402 ;
  assign n42947 = ~n42372 & ~n42946 ;
  assign n42948 = ~n42351 & ~n42947 ;
  assign n42949 = ~n42363 & ~n42725 ;
  assign n42950 = ~n42362 & ~n42949 ;
  assign n42951 = ~n42370 & ~n42950 ;
  assign n42952 = ~n42948 & n42951 ;
  assign n42953 = ~n42945 & ~n42952 ;
  assign n42954 = ~n42394 & ~n42405 ;
  assign n42955 = n42338 & ~n42954 ;
  assign n42962 = n42362 & ~n42719 ;
  assign n42963 = ~n42955 & n42962 ;
  assign n42956 = ~n42344 & n42530 ;
  assign n42957 = ~n42371 & ~n42956 ;
  assign n42958 = ~n42370 & ~n42384 ;
  assign n42959 = ~n42957 & n42958 ;
  assign n42960 = ~n42528 & ~n42721 ;
  assign n42961 = n42351 & ~n42960 ;
  assign n42964 = ~n42959 & ~n42961 ;
  assign n42965 = n42963 & n42964 ;
  assign n42966 = n42382 & ~n42393 ;
  assign n42967 = ~n42362 & ~n42385 ;
  assign n42968 = ~n42395 & ~n42404 ;
  assign n42969 = n42967 & n42968 ;
  assign n42970 = ~n42966 & n42969 ;
  assign n42971 = ~n42965 & ~n42970 ;
  assign n42972 = ~n42953 & ~n42971 ;
  assign n42973 = ~\u1_L4_reg[26]/NET0131  & ~n42972 ;
  assign n42974 = \u1_L4_reg[26]/NET0131  & n42972 ;
  assign n42975 = ~n42973 & ~n42974 ;
  assign n42989 = ~n42895 & ~n42898 ;
  assign n42998 = ~n42872 & ~n42892 ;
  assign n42999 = n42885 & ~n42998 ;
  assign n43000 = n42989 & n42999 ;
  assign n43001 = ~n42916 & ~n43000 ;
  assign n43002 = n42866 & ~n43001 ;
  assign n42980 = n42885 & n42895 ;
  assign n42981 = ~n42892 & n42932 ;
  assign n42982 = ~n42980 & ~n42981 ;
  assign n42997 = ~n42866 & ~n42982 ;
  assign n42994 = n42866 & n42872 ;
  assign n42995 = ~n42886 & ~n42994 ;
  assign n42996 = ~n42892 & ~n42995 ;
  assign n43003 = n42895 & n42925 ;
  assign n43004 = ~n42996 & ~n43003 ;
  assign n43005 = ~n42997 & n43004 ;
  assign n43006 = ~n43002 & n43005 ;
  assign n43007 = n42860 & ~n43006 ;
  assign n42976 = n42898 & n42909 ;
  assign n42977 = ~n42885 & n42919 ;
  assign n42978 = ~n42976 & ~n42977 ;
  assign n42979 = ~n42866 & ~n42978 ;
  assign n42983 = n42866 & n42982 ;
  assign n42984 = ~n42892 & n42898 ;
  assign n42985 = ~n42866 & ~n42897 ;
  assign n42986 = ~n42896 & n42985 ;
  assign n42987 = ~n42984 & n42986 ;
  assign n42988 = ~n42983 & ~n42987 ;
  assign n42990 = n42925 & n42989 ;
  assign n42991 = ~n42976 & ~n42990 ;
  assign n42992 = ~n42988 & n42991 ;
  assign n42993 = ~n42860 & ~n42992 ;
  assign n43008 = ~n42979 & ~n42993 ;
  assign n43009 = ~n43007 & n43008 ;
  assign n43010 = ~\u1_L4_reg[28]/NET0131  & ~n43009 ;
  assign n43011 = \u1_L4_reg[28]/NET0131  & n43009 ;
  assign n43012 = ~n43010 & ~n43011 ;
  assign n43035 = ~n42301 & ~n42303 ;
  assign n43036 = n42253 & ~n42274 ;
  assign n43037 = n42297 & ~n43036 ;
  assign n43038 = n43035 & ~n43037 ;
  assign n43039 = n42271 & ~n43038 ;
  assign n43018 = n42247 & n42259 ;
  assign n43019 = n42253 & n43018 ;
  assign n43032 = ~n42253 & ~n42312 ;
  assign n43033 = ~n43019 & ~n43032 ;
  assign n43034 = ~n42271 & ~n43033 ;
  assign n43040 = n42282 & n42291 ;
  assign n43041 = ~n43034 & ~n43040 ;
  assign n43042 = ~n43039 & n43041 ;
  assign n43043 = ~n42234 & ~n43042 ;
  assign n43020 = ~n42246 & n42253 ;
  assign n43021 = n42274 & ~n43020 ;
  assign n43022 = ~n43019 & ~n43021 ;
  assign n43023 = n42271 & ~n43022 ;
  assign n43013 = ~n42259 & n42263 ;
  assign n43014 = ~n42247 & n42253 ;
  assign n43015 = ~n42291 & n43014 ;
  assign n43016 = ~n43013 & ~n43015 ;
  assign n43017 = ~n42271 & ~n43016 ;
  assign n43024 = n42263 & n42282 ;
  assign n43025 = n42284 & ~n43024 ;
  assign n43026 = ~n42293 & n43025 ;
  assign n43027 = ~n43017 & n43026 ;
  assign n43028 = ~n43023 & n43027 ;
  assign n43029 = n42234 & ~n43028 ;
  assign n43030 = ~n42253 & n42271 ;
  assign n43031 = n42309 & n43030 ;
  assign n43044 = ~n42302 & ~n43031 ;
  assign n43045 = ~n43029 & n43044 ;
  assign n43046 = ~n43043 & n43045 ;
  assign n43047 = \u1_L4_reg[29]/NET0131  & ~n43046 ;
  assign n43048 = ~\u1_L4_reg[29]/NET0131  & n43046 ;
  assign n43049 = ~n43047 & ~n43048 ;
  assign n43056 = ~n42246 & n42260 ;
  assign n43058 = ~n42279 & ~n43056 ;
  assign n43059 = ~n42240 & ~n43058 ;
  assign n43057 = ~n42271 & n43056 ;
  assign n43061 = n42253 & n42309 ;
  assign n43060 = n42281 & n43030 ;
  assign n43062 = n42234 & ~n43060 ;
  assign n43063 = ~n43061 & n43062 ;
  assign n43064 = ~n43057 & n43063 ;
  assign n43065 = ~n43059 & n43064 ;
  assign n43051 = n42271 & ~n43018 ;
  assign n43066 = ~n42283 & ~n42292 ;
  assign n43067 = n43051 & n43066 ;
  assign n43068 = n42259 & n42263 ;
  assign n43069 = ~n42271 & ~n43040 ;
  assign n43070 = ~n43068 & n43069 ;
  assign n43071 = ~n43067 & ~n43070 ;
  assign n43072 = ~n42234 & ~n42307 ;
  assign n43073 = ~n42302 & n43072 ;
  assign n43074 = ~n43071 & n43073 ;
  assign n43075 = ~n43065 & ~n43074 ;
  assign n43052 = ~n42310 & ~n43013 ;
  assign n43053 = n43051 & n43052 ;
  assign n43050 = ~n42271 & n43035 ;
  assign n43054 = n42253 & ~n43050 ;
  assign n43055 = ~n43053 & n43054 ;
  assign n43076 = ~n42289 & ~n43055 ;
  assign n43077 = ~n43075 & n43076 ;
  assign n43078 = ~\u1_L4_reg[4]/NET0131  & ~n43077 ;
  assign n43079 = \u1_L4_reg[4]/NET0131  & n43077 ;
  assign n43080 = ~n43078 & ~n43079 ;
  assign n43082 = ~n42878 & ~n42885 ;
  assign n43083 = n42892 & n43082 ;
  assign n43084 = ~n42866 & ~n42886 ;
  assign n43085 = ~n43083 & n43084 ;
  assign n43087 = n42878 & n42919 ;
  assign n43086 = ~n42892 & n43082 ;
  assign n43088 = n42866 & ~n43086 ;
  assign n43089 = ~n43087 & n43088 ;
  assign n43090 = ~n43085 & ~n43089 ;
  assign n43081 = n42903 & n42998 ;
  assign n43091 = n42860 & ~n43081 ;
  assign n43092 = n42911 & n43091 ;
  assign n43093 = ~n43090 & n43092 ;
  assign n43096 = n42878 & ~n42906 ;
  assign n43097 = n42998 & n43096 ;
  assign n43094 = n42892 & ~n42903 ;
  assign n43095 = n42994 & n43094 ;
  assign n43098 = ~n42860 & ~n43095 ;
  assign n43099 = ~n43097 & n43098 ;
  assign n43100 = n42885 & n42932 ;
  assign n43101 = ~n42866 & ~n43003 ;
  assign n43102 = ~n43100 & n43101 ;
  assign n43103 = ~n42917 & n43102 ;
  assign n43104 = n43099 & n43103 ;
  assign n43105 = ~n43093 & ~n43104 ;
  assign n43106 = ~n42921 & ~n42976 ;
  assign n43107 = ~n43105 & n43106 ;
  assign n43108 = n42885 & ~n42984 ;
  assign n43109 = ~n42896 & ~n42916 ;
  assign n43110 = ~n43108 & n43109 ;
  assign n43111 = n42866 & ~n43110 ;
  assign n43112 = n43099 & n43111 ;
  assign n43113 = ~n43107 & ~n43112 ;
  assign n43114 = ~\u1_L4_reg[13]/NET0131  & ~n43113 ;
  assign n43115 = \u1_L4_reg[13]/NET0131  & n43113 ;
  assign n43116 = ~n43114 & ~n43115 ;
  assign n43118 = n42253 & ~n43052 ;
  assign n43122 = n42234 & ~n43056 ;
  assign n43123 = ~n42293 & n43122 ;
  assign n43117 = n42271 & n42276 ;
  assign n43119 = ~n42240 & ~n42271 ;
  assign n43120 = ~n42259 & ~n43119 ;
  assign n43121 = ~n42298 & n43120 ;
  assign n43124 = ~n43117 & ~n43121 ;
  assign n43125 = n43123 & n43124 ;
  assign n43126 = ~n43118 & n43125 ;
  assign n43129 = n42240 & ~n42260 ;
  assign n43130 = ~n43068 & ~n43129 ;
  assign n43131 = n42271 & ~n43130 ;
  assign n43128 = ~n42271 & ~n43052 ;
  assign n43127 = n42253 & n42303 ;
  assign n43132 = ~n42234 & ~n43127 ;
  assign n43133 = ~n43128 & n43132 ;
  assign n43134 = ~n43131 & n43133 ;
  assign n43135 = ~n43126 & ~n43134 ;
  assign n43136 = n42296 & ~n42308 ;
  assign n43137 = ~n43135 & n43136 ;
  assign n43138 = ~\u1_L4_reg[19]/P0001  & ~n43137 ;
  assign n43139 = \u1_L4_reg[19]/P0001  & n43137 ;
  assign n43140 = ~n43138 & ~n43139 ;
  assign n43143 = ~n42180 & ~n42185 ;
  assign n43144 = ~n42159 & ~n43143 ;
  assign n43145 = ~n42179 & ~n43144 ;
  assign n43146 = ~n42146 & ~n43145 ;
  assign n43147 = n42140 & ~n43146 ;
  assign n43149 = ~n42152 & n42177 ;
  assign n43153 = ~n42747 & ~n43149 ;
  assign n43150 = n42153 & n42201 ;
  assign n43141 = ~n42146 & n42152 ;
  assign n43151 = n42167 & n43141 ;
  assign n43154 = ~n43150 & ~n43151 ;
  assign n43155 = n43153 & n43154 ;
  assign n43148 = n42146 & n42185 ;
  assign n43152 = ~n42140 & ~n42198 ;
  assign n43156 = ~n43148 & n43152 ;
  assign n43157 = n43155 & n43156 ;
  assign n43158 = ~n43147 & ~n43157 ;
  assign n43159 = n42146 & ~n42213 ;
  assign n43160 = n42175 & n43159 ;
  assign n43161 = ~n42221 & ~n42753 ;
  assign n43162 = ~n43160 & n43161 ;
  assign n43163 = n42140 & ~n43162 ;
  assign n43164 = n42201 & n42748 ;
  assign n43165 = ~n42752 & ~n43164 ;
  assign n43166 = ~n42146 & ~n43165 ;
  assign n43167 = ~n42152 & n43148 ;
  assign n43142 = n42215 & n43141 ;
  assign n43168 = ~n42211 & ~n43142 ;
  assign n43169 = ~n43167 & n43168 ;
  assign n43170 = ~n43166 & n43169 ;
  assign n43171 = ~n43163 & n43170 ;
  assign n43172 = ~n43158 & n43171 ;
  assign n43173 = \u1_L4_reg[23]/NET0131  & ~n43172 ;
  assign n43174 = ~\u1_L4_reg[23]/NET0131  & n43172 ;
  assign n43175 = ~n43173 & ~n43174 ;
  assign n43179 = ~n42786 & n42795 ;
  assign n43180 = ~n42459 & ~n43179 ;
  assign n43177 = n42459 & ~n42487 ;
  assign n43178 = ~n42682 & n43177 ;
  assign n43176 = ~n42442 & n42463 ;
  assign n43181 = ~n42450 & ~n43176 ;
  assign n43182 = ~n42505 & n43181 ;
  assign n43183 = ~n43178 & n43182 ;
  assign n43184 = ~n43180 & n43183 ;
  assign n43185 = n42481 & ~n43184 ;
  assign n43189 = n42459 & ~n42470 ;
  assign n43188 = n42449 & ~n42488 ;
  assign n43190 = ~n42801 & ~n43188 ;
  assign n43191 = n43189 & n43190 ;
  assign n43187 = n42499 & n42802 ;
  assign n43186 = n42469 & n42798 ;
  assign n43192 = ~n42486 & ~n43186 ;
  assign n43193 = ~n43187 & n43192 ;
  assign n43194 = ~n43191 & n43193 ;
  assign n43195 = ~n42481 & ~n43194 ;
  assign n43198 = ~n42459 & n42492 ;
  assign n43196 = n42442 & n42459 ;
  assign n43197 = n42483 & n43196 ;
  assign n43199 = ~n42498 & ~n43197 ;
  assign n43200 = ~n43198 & n43199 ;
  assign n43201 = ~n43195 & n43200 ;
  assign n43202 = ~n43185 & n43201 ;
  assign n43203 = ~\u1_L4_reg[27]/NET0131  & ~n43202 ;
  assign n43204 = \u1_L4_reg[27]/NET0131  & n43202 ;
  assign n43205 = ~n43203 & ~n43204 ;
  assign n43217 = n42093 & n42106 ;
  assign n43218 = ~n42074 & n42568 ;
  assign n43219 = ~n42103 & ~n42120 ;
  assign n43220 = ~n43218 & ~n43219 ;
  assign n43221 = ~n42082 & ~n42549 ;
  assign n43222 = ~n43220 & n43221 ;
  assign n43224 = ~n42104 & ~n42551 ;
  assign n43225 = n42112 & n43224 ;
  assign n43223 = n42074 & n42551 ;
  assign n43226 = n42082 & ~n43223 ;
  assign n43227 = ~n43225 & n43226 ;
  assign n43228 = ~n43222 & ~n43227 ;
  assign n43229 = ~n43217 & ~n43228 ;
  assign n43230 = n42049 & ~n43229 ;
  assign n43206 = n42061 & ~n42554 ;
  assign n43210 = ~n42113 & ~n43206 ;
  assign n43207 = ~n42552 & n42559 ;
  assign n43208 = ~n42120 & ~n42552 ;
  assign n43209 = n42082 & ~n43208 ;
  assign n43211 = ~n43207 & ~n43209 ;
  assign n43212 = n43210 & n43211 ;
  assign n43213 = ~n42049 & ~n43212 ;
  assign n43214 = n42082 & n42116 ;
  assign n43215 = n42101 & ~n42551 ;
  assign n43216 = n42094 & n43215 ;
  assign n43231 = ~n43214 & ~n43216 ;
  assign n43232 = ~n43213 & n43231 ;
  assign n43233 = ~n43230 & n43232 ;
  assign n43234 = \u1_L4_reg[32]/NET0131  & n43233 ;
  assign n43235 = ~\u1_L4_reg[32]/NET0131  & ~n43233 ;
  assign n43236 = ~n43234 & ~n43235 ;
  assign n43243 = decrypt_pad & ~\u1_uk_K_r4_reg[40]/NET0131  ;
  assign n43244 = ~decrypt_pad & ~\u1_uk_K_r4_reg[46]/NET0131  ;
  assign n43245 = ~n43243 & ~n43244 ;
  assign n43246 = \u1_R4_reg[11]/P0001  & ~n43245 ;
  assign n43247 = ~\u1_R4_reg[11]/P0001  & n43245 ;
  assign n43248 = ~n43246 & ~n43247 ;
  assign n43237 = decrypt_pad & ~\u1_uk_K_r4_reg[55]/NET0131  ;
  assign n43238 = ~decrypt_pad & ~\u1_uk_K_r4_reg[4]/NET0131  ;
  assign n43239 = ~n43237 & ~n43238 ;
  assign n43240 = \u1_R4_reg[12]/NET0131  & ~n43239 ;
  assign n43241 = ~\u1_R4_reg[12]/NET0131  & n43239 ;
  assign n43242 = ~n43240 & ~n43241 ;
  assign n43249 = decrypt_pad & ~\u1_uk_K_r4_reg[11]/NET0131  ;
  assign n43250 = ~decrypt_pad & ~\u1_uk_K_r4_reg[17]/NET0131  ;
  assign n43251 = ~n43249 & ~n43250 ;
  assign n43252 = \u1_R4_reg[13]/NET0131  & ~n43251 ;
  assign n43253 = ~\u1_R4_reg[13]/NET0131  & n43251 ;
  assign n43254 = ~n43252 & ~n43253 ;
  assign n43262 = decrypt_pad & ~\u1_uk_K_r4_reg[6]/NET0131  ;
  assign n43263 = ~decrypt_pad & ~\u1_uk_K_r4_reg[12]/NET0131  ;
  assign n43264 = ~n43262 & ~n43263 ;
  assign n43265 = \u1_R4_reg[9]/NET0131  & ~n43264 ;
  assign n43266 = ~\u1_R4_reg[9]/NET0131  & n43264 ;
  assign n43267 = ~n43265 & ~n43266 ;
  assign n43307 = n43254 & ~n43267 ;
  assign n43255 = decrypt_pad & ~\u1_uk_K_r4_reg[34]/NET0131  ;
  assign n43256 = ~decrypt_pad & ~\u1_uk_K_r4_reg[40]/NET0131  ;
  assign n43257 = ~n43255 & ~n43256 ;
  assign n43258 = \u1_R4_reg[8]/NET0131  & ~n43257 ;
  assign n43259 = ~\u1_R4_reg[8]/NET0131  & n43257 ;
  assign n43260 = ~n43258 & ~n43259 ;
  assign n43287 = ~n43254 & n43267 ;
  assign n43288 = n43260 & n43287 ;
  assign n43261 = n43254 & ~n43260 ;
  assign n43269 = decrypt_pad & ~\u1_uk_K_r4_reg[39]/NET0131  ;
  assign n43270 = ~decrypt_pad & ~\u1_uk_K_r4_reg[20]/NET0131  ;
  assign n43271 = ~n43269 & ~n43270 ;
  assign n43272 = \u1_R4_reg[10]/NET0131  & ~n43271 ;
  assign n43273 = ~\u1_R4_reg[10]/NET0131  & n43271 ;
  assign n43274 = ~n43272 & ~n43273 ;
  assign n43309 = n43261 & n43274 ;
  assign n43310 = ~n43288 & ~n43309 ;
  assign n43311 = ~n43307 & n43310 ;
  assign n43312 = n43242 & ~n43311 ;
  assign n43308 = n43274 & n43307 ;
  assign n43279 = ~n43254 & ~n43260 ;
  assign n43313 = ~n43274 & n43279 ;
  assign n43314 = ~n43267 & n43313 ;
  assign n43315 = ~n43308 & ~n43314 ;
  assign n43316 = ~n43312 & n43315 ;
  assign n43317 = n43248 & ~n43316 ;
  assign n43280 = n43254 & n43260 ;
  assign n43281 = ~n43279 & ~n43280 ;
  assign n43278 = ~n43267 & ~n43274 ;
  assign n43284 = n43248 & ~n43260 ;
  assign n43290 = n43278 & ~n43284 ;
  assign n43291 = n43281 & n43290 ;
  assign n43285 = n43267 & ~n43274 ;
  assign n43286 = n43284 & n43285 ;
  assign n43289 = n43274 & n43288 ;
  assign n43292 = ~n43286 & ~n43289 ;
  assign n43293 = ~n43291 & n43292 ;
  assign n43268 = n43261 & n43267 ;
  assign n43275 = n43268 & n43274 ;
  assign n43276 = ~n43248 & n43275 ;
  assign n43277 = n43267 & n43274 ;
  assign n43282 = ~n43278 & ~n43281 ;
  assign n43283 = ~n43277 & n43282 ;
  assign n43294 = ~n43276 & ~n43283 ;
  assign n43295 = n43293 & n43294 ;
  assign n43296 = ~n43242 & ~n43295 ;
  assign n43297 = n43242 & n43277 ;
  assign n43298 = n43279 & n43297 ;
  assign n43299 = n43254 & n43285 ;
  assign n43300 = n43260 & ~n43267 ;
  assign n43301 = ~n43254 & n43300 ;
  assign n43302 = n43267 & n43280 ;
  assign n43303 = ~n43301 & ~n43302 ;
  assign n43304 = ~n43299 & n43303 ;
  assign n43305 = n43242 & ~n43248 ;
  assign n43306 = ~n43304 & n43305 ;
  assign n43318 = ~n43298 & ~n43306 ;
  assign n43319 = ~n43296 & n43318 ;
  assign n43320 = ~n43317 & n43319 ;
  assign n43321 = ~\u1_L4_reg[6]/NET0131  & ~n43320 ;
  assign n43322 = \u1_L4_reg[6]/NET0131  & n43320 ;
  assign n43323 = ~n43321 & ~n43322 ;
  assign n43327 = ~n42062 & n43218 ;
  assign n43328 = n42082 & ~n43327 ;
  assign n43329 = ~n42068 & ~n42105 ;
  assign n43324 = n42061 & ~n42568 ;
  assign n43330 = ~n42082 & ~n43223 ;
  assign n43331 = ~n43324 & n43330 ;
  assign n43332 = ~n43329 & n43331 ;
  assign n43333 = ~n43328 & ~n43332 ;
  assign n43325 = ~n42120 & ~n43324 ;
  assign n43326 = n42074 & ~n43325 ;
  assign n43334 = n42049 & ~n43326 ;
  assign n43335 = ~n43333 & n43334 ;
  assign n43336 = n42104 & ~n42568 ;
  assign n43337 = n42082 & ~n42120 ;
  assign n43338 = ~n43218 & n43337 ;
  assign n43339 = ~n43336 & n43338 ;
  assign n43340 = ~n42049 & ~n43339 ;
  assign n43341 = ~n43335 & ~n43340 ;
  assign n43342 = ~n42082 & n43326 ;
  assign n43343 = ~n42082 & n43327 ;
  assign n43344 = ~n42076 & ~n43343 ;
  assign n43345 = n42049 & ~n42082 ;
  assign n43346 = ~n43344 & ~n43345 ;
  assign n43347 = ~n43342 & ~n43346 ;
  assign n43348 = ~n43341 & n43347 ;
  assign n43349 = ~\u1_L4_reg[7]/NET0131  & ~n43348 ;
  assign n43350 = \u1_L4_reg[7]/NET0131  & n43348 ;
  assign n43351 = ~n43349 & ~n43350 ;
  assign n43366 = ~n42607 & n42641 ;
  assign n43367 = ~n42833 & ~n43366 ;
  assign n43368 = n42630 & ~n43367 ;
  assign n43369 = ~n42607 & n42841 ;
  assign n43370 = ~n42649 & ~n43369 ;
  assign n43371 = ~n43368 & n43370 ;
  assign n43372 = n42588 & ~n43371 ;
  assign n43352 = n42630 & n42826 ;
  assign n43357 = ~n42618 & ~n43352 ;
  assign n43358 = n42843 & n43357 ;
  assign n43353 = ~n42615 & n42646 ;
  assign n43354 = ~n42833 & ~n43353 ;
  assign n43355 = ~n42630 & ~n43354 ;
  assign n43356 = n42630 & n42663 ;
  assign n43359 = ~n43355 & ~n43356 ;
  assign n43360 = n43358 & n43359 ;
  assign n43361 = ~n42588 & ~n43360 ;
  assign n43362 = ~n42600 & n42842 ;
  assign n43363 = ~n42616 & n42646 ;
  assign n43364 = ~n42661 & ~n43363 ;
  assign n43365 = n42630 & ~n43364 ;
  assign n43373 = ~n43362 & ~n43365 ;
  assign n43374 = ~n43361 & n43373 ;
  assign n43375 = ~n43372 & n43374 ;
  assign n43376 = ~\u1_L4_reg[8]/NET0131  & ~n43375 ;
  assign n43377 = \u1_L4_reg[8]/NET0131  & n43375 ;
  assign n43378 = ~n43376 & ~n43377 ;
  assign n43379 = n43261 & ~n43267 ;
  assign n43396 = n43284 & n43287 ;
  assign n43397 = ~n43379 & ~n43396 ;
  assign n43398 = n43303 & n43397 ;
  assign n43399 = ~n43274 & ~n43398 ;
  assign n43390 = n43274 & n43279 ;
  assign n43400 = n43260 & ~n43274 ;
  assign n43401 = ~n43254 & n43400 ;
  assign n43402 = ~n43390 & ~n43401 ;
  assign n43403 = ~n43248 & ~n43402 ;
  assign n43404 = ~n43275 & ~n43403 ;
  assign n43405 = ~n43399 & n43404 ;
  assign n43406 = n43242 & ~n43405 ;
  assign n43380 = ~n43302 & ~n43313 ;
  assign n43381 = ~n43379 & n43380 ;
  assign n43382 = ~n43248 & ~n43381 ;
  assign n43383 = ~n43267 & ~n43280 ;
  assign n43384 = n43248 & ~n43279 ;
  assign n43385 = ~n43302 & n43384 ;
  assign n43386 = ~n43383 & n43385 ;
  assign n43387 = ~n43314 & ~n43386 ;
  assign n43388 = ~n43382 & n43387 ;
  assign n43389 = ~n43242 & ~n43388 ;
  assign n43391 = ~n43267 & n43390 ;
  assign n43392 = ~n43289 & ~n43391 ;
  assign n43393 = n43248 & ~n43392 ;
  assign n43394 = ~n43248 & n43274 ;
  assign n43395 = n43300 & n43394 ;
  assign n43407 = ~n43393 & ~n43395 ;
  assign n43408 = ~n43389 & n43407 ;
  assign n43409 = ~n43406 & n43408 ;
  assign n43410 = ~\u1_L4_reg[16]/NET0131  & ~n43409 ;
  assign n43411 = \u1_L4_reg[16]/NET0131  & n43409 ;
  assign n43412 = ~n43410 & ~n43411 ;
  assign n43429 = ~n43248 & n43282 ;
  assign n43423 = n43260 & n43277 ;
  assign n43424 = ~n43309 & ~n43423 ;
  assign n43425 = n43248 & ~n43424 ;
  assign n43426 = n43248 & ~n43274 ;
  assign n43427 = ~n43261 & ~n43267 ;
  assign n43428 = n43426 & n43427 ;
  assign n43430 = ~n43291 & ~n43428 ;
  assign n43431 = ~n43425 & n43430 ;
  assign n43432 = ~n43429 & n43431 ;
  assign n43433 = n43242 & ~n43432 ;
  assign n43413 = n43261 & ~n43274 ;
  assign n43414 = ~n43390 & ~n43413 ;
  assign n43415 = n43267 & n43279 ;
  assign n43416 = n43274 & n43300 ;
  assign n43417 = ~n43415 & ~n43416 ;
  assign n43418 = n43414 & n43417 ;
  assign n43419 = n43248 & ~n43418 ;
  assign n43420 = n43274 & n43301 ;
  assign n43421 = ~n43419 & ~n43420 ;
  assign n43422 = ~n43242 & ~n43421 ;
  assign n43437 = n43278 & ~n43281 ;
  assign n43438 = n43310 & ~n43437 ;
  assign n43439 = ~n43242 & ~n43248 ;
  assign n43440 = ~n43438 & n43439 ;
  assign n43434 = n43302 & n43394 ;
  assign n43435 = ~n43268 & ~n43301 ;
  assign n43436 = n43426 & ~n43435 ;
  assign n43441 = ~n43434 & ~n43436 ;
  assign n43442 = ~n43440 & n43441 ;
  assign n43443 = ~n43422 & n43442 ;
  assign n43444 = ~n43433 & n43443 ;
  assign n43445 = ~\u1_L4_reg[24]/NET0131  & ~n43444 ;
  assign n43446 = \u1_L4_reg[24]/NET0131  & n43444 ;
  assign n43447 = ~n43445 & ~n43446 ;
  assign n43453 = n43274 & n43379 ;
  assign n43457 = ~n43242 & ~n43437 ;
  assign n43458 = ~n43453 & n43457 ;
  assign n43448 = n43260 & n43274 ;
  assign n43449 = ~n43287 & n43448 ;
  assign n43450 = ~n43254 & n43285 ;
  assign n43451 = ~n43449 & ~n43450 ;
  assign n43452 = n43248 & ~n43451 ;
  assign n43454 = ~n43287 & n43400 ;
  assign n43455 = ~n43268 & ~n43454 ;
  assign n43456 = ~n43248 & ~n43455 ;
  assign n43459 = ~n43452 & ~n43456 ;
  assign n43460 = n43458 & n43459 ;
  assign n43463 = ~n43274 & n43301 ;
  assign n43464 = n43414 & ~n43463 ;
  assign n43465 = n43248 & ~n43464 ;
  assign n43461 = ~n43415 & ~n43448 ;
  assign n43462 = ~n43248 & ~n43461 ;
  assign n43466 = n43242 & ~n43462 ;
  assign n43467 = ~n43465 & n43466 ;
  assign n43468 = ~n43460 & ~n43467 ;
  assign n43471 = n43248 & n43307 ;
  assign n43472 = n43448 & n43471 ;
  assign n43469 = ~n43280 & n43297 ;
  assign n43470 = n43287 & n43394 ;
  assign n43473 = ~n43469 & ~n43470 ;
  assign n43474 = ~n43472 & n43473 ;
  assign n43475 = ~n43468 & n43474 ;
  assign n43476 = \u1_L4_reg[30]/NET0131  & ~n43475 ;
  assign n43477 = ~\u1_L4_reg[30]/NET0131  & n43475 ;
  assign n43478 = ~n43476 & ~n43477 ;
  assign n43489 = n42594 & n42669 ;
  assign n43490 = ~n42645 & ~n43489 ;
  assign n43491 = n42630 & ~n43490 ;
  assign n43492 = ~n42630 & n42650 ;
  assign n43488 = n42607 & n42662 ;
  assign n43493 = ~n42664 & ~n43488 ;
  assign n43494 = ~n43492 & n43493 ;
  assign n43495 = ~n43491 & n43494 ;
  assign n43496 = n42588 & ~n43495 ;
  assign n43483 = ~n42623 & ~n42844 ;
  assign n43484 = n42630 & ~n43483 ;
  assign n43480 = ~n42601 & n42615 ;
  assign n43481 = ~n42670 & ~n42833 ;
  assign n43482 = ~n42630 & ~n43481 ;
  assign n43485 = ~n43480 & ~n43482 ;
  assign n43486 = ~n43484 & n43485 ;
  assign n43487 = ~n42588 & ~n43486 ;
  assign n43497 = n42615 & n42632 ;
  assign n43498 = ~n42639 & ~n43497 ;
  assign n43499 = ~n43366 & n43498 ;
  assign n43500 = ~n42630 & ~n43499 ;
  assign n43479 = n42633 & n42647 ;
  assign n43501 = ~n43356 & ~n43479 ;
  assign n43502 = ~n43500 & n43501 ;
  assign n43503 = ~n43487 & n43502 ;
  assign n43504 = ~n43496 & n43503 ;
  assign n43505 = ~\u1_L4_reg[3]/NET0131  & ~n43504 ;
  assign n43506 = \u1_L4_reg[3]/NET0131  & n43504 ;
  assign n43507 = ~n43505 & ~n43506 ;
  assign n43521 = n42769 & ~n43144 ;
  assign n43522 = n42152 & ~n43521 ;
  assign n43512 = ~n42177 & ~n42767 ;
  assign n43523 = n42202 & ~n43512 ;
  assign n43524 = ~n42752 & ~n43523 ;
  assign n43525 = ~n43522 & n43524 ;
  assign n43526 = n42140 & ~n43525 ;
  assign n43508 = ~n42152 & n42215 ;
  assign n43509 = n42152 & n42767 ;
  assign n43510 = ~n43508 & ~n43509 ;
  assign n43511 = ~n42146 & ~n43510 ;
  assign n43513 = ~n42146 & n43512 ;
  assign n43514 = n42146 & ~n42760 ;
  assign n43515 = n43143 & n43514 ;
  assign n43516 = ~n43513 & ~n43515 ;
  assign n43517 = ~n42168 & n42199 ;
  assign n43518 = ~n43508 & ~n43517 ;
  assign n43519 = ~n43516 & n43518 ;
  assign n43520 = ~n42140 & ~n43519 ;
  assign n43527 = ~n43511 & ~n43520 ;
  assign n43528 = ~n43526 & n43527 ;
  assign n43529 = ~\u1_L4_reg[9]/NET0131  & ~n43528 ;
  assign n43530 = \u1_L4_reg[9]/NET0131  & n43528 ;
  assign n43531 = ~n43529 & ~n43530 ;
  assign n43541 = n42866 & ~n42904 ;
  assign n43542 = ~n42907 & ~n43082 ;
  assign n43543 = ~n42994 & ~n42998 ;
  assign n43544 = ~n43542 & n43543 ;
  assign n43545 = ~n43541 & ~n43544 ;
  assign n43546 = n42860 & ~n43545 ;
  assign n43533 = n42879 & n42918 ;
  assign n43536 = ~n42976 & ~n43086 ;
  assign n43537 = ~n43533 & n43536 ;
  assign n43534 = ~n42918 & ~n42927 ;
  assign n43535 = n42926 & n43534 ;
  assign n43538 = ~n42893 & ~n43535 ;
  assign n43539 = n43537 & n43538 ;
  assign n43540 = ~n42860 & ~n43539 ;
  assign n43532 = ~n42866 & n42980 ;
  assign n43547 = n42879 & n42892 ;
  assign n43548 = ~n43081 & ~n43547 ;
  assign n43549 = n42866 & ~n43548 ;
  assign n43550 = ~n43532 & ~n43549 ;
  assign n43551 = ~n43540 & n43550 ;
  assign n43552 = ~n43546 & n43551 ;
  assign n43553 = \u1_L4_reg[18]/NET0131  & n43552 ;
  assign n43554 = ~\u1_L4_reg[18]/NET0131  & ~n43552 ;
  assign n43555 = ~n43553 & ~n43554 ;
  assign n43569 = n5844 & n5856 ;
  assign n43570 = ~n5868 & ~n43569 ;
  assign n43571 = ~n5865 & ~n43570 ;
  assign n43577 = n5853 & n5865 ;
  assign n43576 = n5844 & ~n5865 ;
  assign n43578 = n5838 & ~n43576 ;
  assign n43579 = ~n43577 & n43578 ;
  assign n43572 = ~n5844 & n5865 ;
  assign n43573 = ~n5899 & ~n43572 ;
  assign n43574 = n5898 & ~n43573 ;
  assign n43575 = n5865 & n5877 ;
  assign n43580 = ~n43574 & ~n43575 ;
  assign n43581 = ~n43579 & n43580 ;
  assign n43582 = ~n43571 & n43581 ;
  assign n43583 = ~n5883 & ~n43582 ;
  assign n43561 = n5865 & n5869 ;
  assign n43562 = ~n5856 & ~n43561 ;
  assign n43563 = ~n5844 & ~n43562 ;
  assign n43556 = ~n5837 & n5850 ;
  assign n43557 = ~n5831 & n5875 ;
  assign n43558 = ~n43556 & ~n43557 ;
  assign n43559 = n5865 & ~n43558 ;
  assign n43560 = ~n5852 & n5884 ;
  assign n43564 = n5857 & ~n5865 ;
  assign n43565 = ~n43560 & ~n43564 ;
  assign n43566 = ~n43559 & n43565 ;
  assign n43567 = ~n43563 & n43566 ;
  assign n43568 = n5883 & ~n43567 ;
  assign n43586 = ~n5857 & ~n5884 ;
  assign n43587 = n5851 & ~n43586 ;
  assign n43588 = ~n5889 & ~n43587 ;
  assign n43589 = ~n5865 & ~n43588 ;
  assign n43584 = n5865 & n5875 ;
  assign n43585 = n5884 & n43584 ;
  assign n43590 = n5831 & n5865 ;
  assign n43591 = n5899 & n43590 ;
  assign n43592 = ~n43585 & ~n43591 ;
  assign n43593 = ~n43589 & n43592 ;
  assign n43594 = ~n43568 & n43593 ;
  assign n43595 = ~n43583 & n43594 ;
  assign n43596 = ~\u1_L3_reg[31]/NET0131  & ~n43595 ;
  assign n43597 = \u1_L3_reg[31]/NET0131  & n43595 ;
  assign n43598 = ~n43596 & ~n43597 ;
  assign n43599 = decrypt_pad & ~\u1_uk_K_r3_reg[29]/NET0131  ;
  assign n43600 = ~decrypt_pad & ~\u1_uk_K_r3_reg[38]/NET0131  ;
  assign n43601 = ~n43599 & ~n43600 ;
  assign n43602 = \u1_R3_reg[24]/NET0131  & ~n43601 ;
  assign n43603 = ~\u1_R3_reg[24]/NET0131  & n43601 ;
  assign n43604 = ~n43602 & ~n43603 ;
  assign n43618 = decrypt_pad & ~\u1_uk_K_r3_reg[14]/NET0131  ;
  assign n43619 = ~decrypt_pad & ~\u1_uk_K_r3_reg[50]/NET0131  ;
  assign n43620 = ~n43618 & ~n43619 ;
  assign n43621 = \u1_R3_reg[22]/NET0131  & ~n43620 ;
  assign n43622 = ~\u1_R3_reg[22]/NET0131  & n43620 ;
  assign n43623 = ~n43621 & ~n43622 ;
  assign n43624 = decrypt_pad & ~\u1_uk_K_r3_reg[23]/NET0131  ;
  assign n43625 = ~decrypt_pad & ~\u1_uk_K_r3_reg[28]/NET0131  ;
  assign n43626 = ~n43624 & ~n43625 ;
  assign n43627 = \u1_R3_reg[21]/NET0131  & ~n43626 ;
  assign n43628 = ~\u1_R3_reg[21]/NET0131  & n43626 ;
  assign n43629 = ~n43627 & ~n43628 ;
  assign n43605 = decrypt_pad & ~\u1_uk_K_r3_reg[8]/NET0131  ;
  assign n43606 = ~decrypt_pad & ~\u1_uk_K_r3_reg[44]/NET0131  ;
  assign n43607 = ~n43605 & ~n43606 ;
  assign n43608 = \u1_R3_reg[20]/NET0131  & ~n43607 ;
  assign n43609 = ~\u1_R3_reg[20]/NET0131  & n43607 ;
  assign n43610 = ~n43608 & ~n43609 ;
  assign n43611 = decrypt_pad & ~\u1_uk_K_r3_reg[52]/NET0131  ;
  assign n43612 = ~decrypt_pad & ~\u1_uk_K_r3_reg[29]/NET0131  ;
  assign n43613 = ~n43611 & ~n43612 ;
  assign n43614 = \u1_R3_reg[25]/NET0131  & ~n43613 ;
  assign n43615 = ~\u1_R3_reg[25]/NET0131  & n43613 ;
  assign n43616 = ~n43614 & ~n43615 ;
  assign n43636 = ~n43610 & n43616 ;
  assign n43681 = n43629 & n43636 ;
  assign n43682 = ~n43623 & ~n43681 ;
  assign n43659 = n43610 & n43616 ;
  assign n43660 = n43623 & n43659 ;
  assign n43639 = decrypt_pad & ~\u1_uk_K_r3_reg[31]/NET0131  ;
  assign n43640 = ~decrypt_pad & ~\u1_uk_K_r3_reg[8]/NET0131  ;
  assign n43641 = ~n43639 & ~n43640 ;
  assign n43642 = \u1_R3_reg[23]/NET0131  & ~n43641 ;
  assign n43643 = ~\u1_R3_reg[23]/NET0131  & n43641 ;
  assign n43644 = ~n43642 & ~n43643 ;
  assign n43650 = n43623 & n43629 ;
  assign n43651 = ~n43610 & n43650 ;
  assign n43683 = ~n43644 & ~n43651 ;
  assign n43684 = ~n43660 & n43683 ;
  assign n43685 = ~n43682 & n43684 ;
  assign n43617 = n43610 & ~n43616 ;
  assign n43674 = n43617 & ~n43629 ;
  assign n43675 = ~n43623 & n43674 ;
  assign n43673 = n43629 & n43659 ;
  assign n43676 = ~n43651 & ~n43673 ;
  assign n43677 = ~n43675 & n43676 ;
  assign n43678 = n43644 & ~n43677 ;
  assign n43646 = ~n43623 & ~n43644 ;
  assign n43679 = n43646 & n43659 ;
  assign n43680 = ~n43629 & n43679 ;
  assign n43686 = ~n43678 & ~n43680 ;
  assign n43687 = ~n43685 & n43686 ;
  assign n43688 = n43604 & ~n43687 ;
  assign n43632 = n43610 & ~n43629 ;
  assign n43633 = n43623 & n43632 ;
  assign n43634 = ~n43610 & ~n43623 ;
  assign n43635 = ~n43633 & ~n43634 ;
  assign n43637 = ~n43629 & n43636 ;
  assign n43638 = n43635 & ~n43637 ;
  assign n43645 = ~n43638 & n43644 ;
  assign n43630 = ~n43623 & n43629 ;
  assign n43652 = n43610 & n43630 ;
  assign n43653 = ~n43651 & ~n43652 ;
  assign n43654 = ~n43644 & ~n43653 ;
  assign n43631 = n43617 & n43630 ;
  assign n43647 = n43617 & n43646 ;
  assign n43648 = n43616 & n43633 ;
  assign n43649 = ~n43647 & ~n43648 ;
  assign n43655 = ~n43631 & n43649 ;
  assign n43656 = ~n43654 & n43655 ;
  assign n43657 = ~n43645 & n43656 ;
  assign n43658 = ~n43604 & ~n43657 ;
  assign n43661 = n43629 & n43634 ;
  assign n43662 = ~n43616 & n43661 ;
  assign n43663 = ~n43660 & ~n43662 ;
  assign n43664 = n43644 & ~n43663 ;
  assign n43665 = ~n43610 & ~n43616 ;
  assign n43666 = ~n43629 & n43665 ;
  assign n43667 = n43646 & n43666 ;
  assign n43668 = ~n43623 & n43644 ;
  assign n43669 = n43637 & n43668 ;
  assign n43670 = n43617 & n43629 ;
  assign n43671 = n43646 & n43670 ;
  assign n43672 = ~n43669 & ~n43671 ;
  assign n43689 = ~n43667 & n43672 ;
  assign n43690 = ~n43664 & n43689 ;
  assign n43691 = ~n43658 & n43690 ;
  assign n43692 = ~n43688 & n43691 ;
  assign n43693 = ~\u1_L3_reg[11]/NET0131  & n43692 ;
  assign n43694 = \u1_L3_reg[11]/NET0131  & ~n43692 ;
  assign n43695 = ~n43693 & ~n43694 ;
  assign n43696 = decrypt_pad & ~\u1_uk_K_r3_reg[36]/NET0131  ;
  assign n43697 = ~decrypt_pad & ~\u1_uk_K_r3_reg[45]/NET0131  ;
  assign n43698 = ~n43696 & ~n43697 ;
  assign n43699 = \u1_R3_reg[28]/NET0131  & ~n43698 ;
  assign n43700 = ~\u1_R3_reg[28]/NET0131  & n43698 ;
  assign n43701 = ~n43699 & ~n43700 ;
  assign n43702 = decrypt_pad & ~\u1_uk_K_r3_reg[16]/NET0131  ;
  assign n43703 = ~decrypt_pad & ~\u1_uk_K_r3_reg[21]/NET0131  ;
  assign n43704 = ~n43702 & ~n43703 ;
  assign n43705 = \u1_R3_reg[26]/NET0131  & ~n43704 ;
  assign n43706 = ~\u1_R3_reg[26]/NET0131  & n43704 ;
  assign n43707 = ~n43705 & ~n43706 ;
  assign n43708 = decrypt_pad & ~\u1_uk_K_r3_reg[0]/NET0131  ;
  assign n43709 = ~decrypt_pad & ~\u1_uk_K_r3_reg[36]/NET0131  ;
  assign n43710 = ~n43708 & ~n43709 ;
  assign n43711 = \u1_R3_reg[25]/NET0131  & ~n43710 ;
  assign n43712 = ~\u1_R3_reg[25]/NET0131  & n43710 ;
  assign n43713 = ~n43711 & ~n43712 ;
  assign n43742 = ~n43707 & ~n43713 ;
  assign n43714 = decrypt_pad & ~\u1_uk_K_r3_reg[28]/NET0131  ;
  assign n43715 = ~decrypt_pad & ~\u1_uk_K_r3_reg[9]/NET0131  ;
  assign n43716 = ~n43714 & ~n43715 ;
  assign n43717 = \u1_R3_reg[29]/NET0131  & ~n43716 ;
  assign n43718 = ~\u1_R3_reg[29]/NET0131  & n43716 ;
  assign n43719 = ~n43717 & ~n43718 ;
  assign n43745 = ~n43707 & ~n43719 ;
  assign n43765 = ~n43742 & ~n43745 ;
  assign n43721 = decrypt_pad & ~\u1_uk_K_r3_reg[51]/NET0131  ;
  assign n43722 = ~decrypt_pad & ~\u1_uk_K_r3_reg[1]/NET0131  ;
  assign n43723 = ~n43721 & ~n43722 ;
  assign n43724 = \u1_R3_reg[24]/NET0131  & ~n43723 ;
  assign n43725 = ~\u1_R3_reg[24]/NET0131  & n43723 ;
  assign n43726 = ~n43724 & ~n43725 ;
  assign n43729 = decrypt_pad & ~\u1_uk_K_r3_reg[49]/NET0131  ;
  assign n43730 = ~decrypt_pad & ~\u1_uk_K_r3_reg[30]/NET0131  ;
  assign n43731 = ~n43729 & ~n43730 ;
  assign n43732 = \u1_R3_reg[27]/NET0131  & ~n43731 ;
  assign n43733 = ~\u1_R3_reg[27]/NET0131  & n43731 ;
  assign n43734 = ~n43732 & ~n43733 ;
  assign n43744 = n43707 & n43713 ;
  assign n43764 = n43734 & ~n43744 ;
  assign n43766 = n43726 & n43764 ;
  assign n43767 = n43765 & n43766 ;
  assign n43758 = n43719 & n43726 ;
  assign n43759 = n43742 & n43758 ;
  assign n43760 = n43713 & n43719 ;
  assign n43761 = ~n43726 & n43760 ;
  assign n43762 = ~n43759 & ~n43761 ;
  assign n43763 = ~n43734 & ~n43762 ;
  assign n43753 = ~n43719 & ~n43726 ;
  assign n43754 = n43742 & n43753 ;
  assign n43755 = n43719 & ~n43726 ;
  assign n43756 = n43707 & ~n43713 ;
  assign n43757 = n43755 & n43756 ;
  assign n43768 = ~n43754 & ~n43757 ;
  assign n43769 = ~n43763 & n43768 ;
  assign n43770 = ~n43767 & n43769 ;
  assign n43771 = n43701 & ~n43770 ;
  assign n43746 = ~n43734 & ~n43744 ;
  assign n43747 = ~n43745 & n43746 ;
  assign n43743 = n43734 & ~n43742 ;
  assign n43748 = n43726 & ~n43743 ;
  assign n43749 = ~n43747 & n43748 ;
  assign n43720 = ~n43713 & ~n43719 ;
  assign n43727 = n43720 & ~n43726 ;
  assign n43728 = n43707 & n43727 ;
  assign n43735 = n43728 & ~n43734 ;
  assign n43736 = ~n43707 & ~n43726 ;
  assign n43737 = n43707 & n43726 ;
  assign n43738 = ~n43736 & ~n43737 ;
  assign n43739 = ~n43713 & n43734 ;
  assign n43740 = n43719 & ~n43739 ;
  assign n43741 = ~n43738 & n43740 ;
  assign n43750 = ~n43735 & ~n43741 ;
  assign n43751 = ~n43749 & n43750 ;
  assign n43752 = ~n43701 & ~n43751 ;
  assign n43774 = n43744 & n43753 ;
  assign n43775 = ~n43757 & ~n43774 ;
  assign n43776 = ~n43719 & n43726 ;
  assign n43777 = ~n43713 & n43776 ;
  assign n43778 = n43775 & ~n43777 ;
  assign n43779 = n43734 & ~n43778 ;
  assign n43772 = n43713 & ~n43734 ;
  assign n43773 = ~n43738 & n43772 ;
  assign n43780 = n43739 & n43745 ;
  assign n43781 = ~n43773 & ~n43780 ;
  assign n43782 = ~n43779 & n43781 ;
  assign n43783 = ~n43752 & n43782 ;
  assign n43784 = ~n43771 & n43783 ;
  assign n43785 = ~\u1_L3_reg[22]/NET0131  & ~n43784 ;
  assign n43786 = \u1_L3_reg[22]/NET0131  & n43784 ;
  assign n43787 = ~n43785 & ~n43786 ;
  assign n43844 = decrypt_pad & ~\u1_uk_K_r3_reg[32]/NET0131  ;
  assign n43845 = ~decrypt_pad & ~\u1_uk_K_r3_reg[41]/NET0131  ;
  assign n43846 = ~n43844 & ~n43845 ;
  assign n43847 = \u1_R3_reg[16]/NET0131  & ~n43846 ;
  assign n43848 = ~\u1_R3_reg[16]/NET0131  & n43846 ;
  assign n43849 = ~n43847 & ~n43848 ;
  assign n43788 = decrypt_pad & ~\u1_uk_K_r3_reg[53]/NET0131  ;
  assign n43789 = ~decrypt_pad & ~\u1_uk_K_r3_reg[5]/NET0131  ;
  assign n43790 = ~n43788 & ~n43789 ;
  assign n43791 = \u1_R3_reg[12]/NET0131  & ~n43790 ;
  assign n43792 = ~\u1_R3_reg[12]/NET0131  & n43790 ;
  assign n43793 = ~n43791 & ~n43792 ;
  assign n43814 = decrypt_pad & ~\u1_uk_K_r3_reg[12]/NET0131  ;
  assign n43815 = ~decrypt_pad & ~\u1_uk_K_r3_reg[46]/NET0131  ;
  assign n43816 = ~n43814 & ~n43815 ;
  assign n43817 = \u1_R3_reg[17]/NET0131  & ~n43816 ;
  assign n43818 = ~\u1_R3_reg[17]/NET0131  & n43816 ;
  assign n43819 = ~n43817 & ~n43818 ;
  assign n43822 = n43793 & ~n43819 ;
  assign n43794 = decrypt_pad & ~\u1_uk_K_r3_reg[47]/NET0131  ;
  assign n43795 = ~decrypt_pad & ~\u1_uk_K_r3_reg[24]/NET0131  ;
  assign n43796 = ~n43794 & ~n43795 ;
  assign n43797 = \u1_R3_reg[13]/NET0131  & ~n43796 ;
  assign n43798 = ~\u1_R3_reg[13]/NET0131  & n43796 ;
  assign n43799 = ~n43797 & ~n43798 ;
  assign n43801 = decrypt_pad & ~\u1_uk_K_r3_reg[24]/NET0131  ;
  assign n43802 = ~decrypt_pad & ~\u1_uk_K_r3_reg[33]/NET0131  ;
  assign n43803 = ~n43801 & ~n43802 ;
  assign n43804 = \u1_R3_reg[15]/NET0131  & ~n43803 ;
  assign n43805 = ~\u1_R3_reg[15]/NET0131  & n43803 ;
  assign n43806 = ~n43804 & ~n43805 ;
  assign n43830 = n43799 & n43806 ;
  assign n43851 = n43822 & n43830 ;
  assign n43807 = decrypt_pad & ~\u1_uk_K_r3_reg[48]/NET0131  ;
  assign n43808 = ~decrypt_pad & ~\u1_uk_K_r3_reg[25]/NET0131  ;
  assign n43809 = ~n43807 & ~n43808 ;
  assign n43810 = \u1_R3_reg[14]/NET0131  & ~n43809 ;
  assign n43811 = ~\u1_R3_reg[14]/NET0131  & n43809 ;
  assign n43812 = ~n43810 & ~n43811 ;
  assign n43852 = ~n43793 & n43819 ;
  assign n43853 = n43799 & n43852 ;
  assign n43854 = ~n43812 & n43853 ;
  assign n43855 = ~n43851 & ~n43854 ;
  assign n43856 = n43806 & n43852 ;
  assign n43857 = ~n43799 & n43856 ;
  assign n43829 = n43793 & n43819 ;
  assign n43858 = n43812 & n43829 ;
  assign n43859 = n43799 & n43858 ;
  assign n43864 = ~n43857 & ~n43859 ;
  assign n43834 = ~n43799 & ~n43819 ;
  assign n43835 = ~n43793 & n43834 ;
  assign n43836 = ~n43806 & n43812 ;
  assign n43860 = n43835 & n43836 ;
  assign n43813 = ~n43806 & ~n43812 ;
  assign n43800 = ~n43793 & n43799 ;
  assign n43861 = n43793 & ~n43799 ;
  assign n43862 = ~n43800 & ~n43861 ;
  assign n43863 = n43813 & ~n43862 ;
  assign n43865 = ~n43860 & ~n43863 ;
  assign n43866 = n43864 & n43865 ;
  assign n43867 = n43855 & n43866 ;
  assign n43868 = n43849 & ~n43867 ;
  assign n43823 = n43812 & n43822 ;
  assign n43824 = ~n43799 & n43819 ;
  assign n43825 = ~n43823 & ~n43824 ;
  assign n43826 = ~n43806 & ~n43825 ;
  assign n43827 = n43800 & ~n43819 ;
  assign n43828 = n43812 & n43827 ;
  assign n43838 = n43806 & n43812 ;
  assign n43839 = n43800 & n43838 ;
  assign n43840 = ~n43828 & ~n43839 ;
  assign n43831 = ~n43799 & ~n43812 ;
  assign n43832 = ~n43830 & ~n43831 ;
  assign n43833 = n43829 & ~n43832 ;
  assign n43837 = n43835 & ~n43836 ;
  assign n43841 = ~n43833 & ~n43837 ;
  assign n43842 = n43840 & n43841 ;
  assign n43843 = ~n43826 & n43842 ;
  assign n43850 = ~n43843 & ~n43849 ;
  assign n43869 = ~n43812 & ~n43819 ;
  assign n43870 = ~n43793 & n43869 ;
  assign n43871 = ~n43799 & n43870 ;
  assign n43872 = ~n43819 & n43861 ;
  assign n43873 = n43812 & n43872 ;
  assign n43874 = ~n43871 & ~n43873 ;
  assign n43875 = n43806 & ~n43874 ;
  assign n43820 = n43813 & n43819 ;
  assign n43821 = n43800 & n43820 ;
  assign n43876 = ~n43812 & n43851 ;
  assign n43877 = ~n43821 & ~n43876 ;
  assign n43878 = ~n43875 & n43877 ;
  assign n43879 = ~n43850 & n43878 ;
  assign n43880 = ~n43868 & n43879 ;
  assign n43881 = ~\u1_L3_reg[20]/NET0131  & ~n43880 ;
  assign n43882 = \u1_L3_reg[20]/NET0131  & n43880 ;
  assign n43883 = ~n43881 & ~n43882 ;
  assign n43890 = n43617 & n43650 ;
  assign n43891 = ~n43661 & ~n43890 ;
  assign n43901 = ~n43681 & n43891 ;
  assign n43902 = n43644 & ~n43901 ;
  assign n43903 = ~n43630 & n43665 ;
  assign n43904 = ~n43660 & ~n43903 ;
  assign n43905 = ~n43644 & ~n43904 ;
  assign n43885 = ~n43623 & ~n43629 ;
  assign n43900 = n43636 & n43885 ;
  assign n43906 = n43623 & n43666 ;
  assign n43907 = ~n43900 & ~n43906 ;
  assign n43908 = n43649 & n43907 ;
  assign n43909 = ~n43905 & n43908 ;
  assign n43910 = ~n43902 & n43909 ;
  assign n43911 = n43604 & ~n43910 ;
  assign n43884 = ~n43673 & ~n43674 ;
  assign n43886 = ~n43651 & ~n43885 ;
  assign n43887 = ~n43616 & ~n43886 ;
  assign n43888 = n43884 & ~n43887 ;
  assign n43889 = n43644 & ~n43888 ;
  assign n43892 = ~n43644 & ~n43891 ;
  assign n43893 = n43623 & n43637 ;
  assign n43894 = ~n43679 & ~n43893 ;
  assign n43895 = ~n43892 & n43894 ;
  assign n43896 = ~n43889 & n43895 ;
  assign n43897 = ~n43604 & ~n43896 ;
  assign n43898 = n43616 & n43629 ;
  assign n43899 = n43668 & n43898 ;
  assign n43912 = ~n43675 & ~n43899 ;
  assign n43913 = ~n43897 & n43912 ;
  assign n43914 = ~n43911 & n43913 ;
  assign n43915 = \u1_L3_reg[29]/NET0131  & ~n43914 ;
  assign n43916 = ~\u1_L3_reg[29]/NET0131  & n43914 ;
  assign n43917 = ~n43915 & ~n43916 ;
  assign n43918 = decrypt_pad & ~\u1_uk_K_r3_reg[6]/NET0131  ;
  assign n43919 = ~decrypt_pad & ~\u1_uk_K_r3_reg[40]/NET0131  ;
  assign n43920 = ~n43918 & ~n43919 ;
  assign n43921 = \u1_R3_reg[8]/NET0131  & ~n43920 ;
  assign n43922 = ~\u1_R3_reg[8]/NET0131  & n43920 ;
  assign n43923 = ~n43921 & ~n43922 ;
  assign n43924 = decrypt_pad & ~\u1_uk_K_r3_reg[40]/NET0131  ;
  assign n43925 = ~decrypt_pad & ~\u1_uk_K_r3_reg[17]/NET0131  ;
  assign n43926 = ~n43924 & ~n43925 ;
  assign n43927 = \u1_R3_reg[7]/NET0131  & ~n43926 ;
  assign n43928 = ~\u1_R3_reg[7]/NET0131  & n43926 ;
  assign n43929 = ~n43927 & ~n43928 ;
  assign n43943 = decrypt_pad & ~\u1_uk_K_r3_reg[55]/NET0131  ;
  assign n43944 = ~decrypt_pad & ~\u1_uk_K_r3_reg[32]/NET0131  ;
  assign n43945 = ~n43943 & ~n43944 ;
  assign n43946 = \u1_R3_reg[5]/NET0131  & ~n43945 ;
  assign n43947 = ~\u1_R3_reg[5]/NET0131  & n43945 ;
  assign n43948 = ~n43946 & ~n43947 ;
  assign n43930 = decrypt_pad & ~\u1_uk_K_r3_reg[19]/NET0131  ;
  assign n43931 = ~decrypt_pad & ~\u1_uk_K_r3_reg[53]/NET0131  ;
  assign n43932 = ~n43930 & ~n43931 ;
  assign n43933 = \u1_R3_reg[4]/NET0131  & ~n43932 ;
  assign n43934 = ~\u1_R3_reg[4]/NET0131  & n43932 ;
  assign n43935 = ~n43933 & ~n43934 ;
  assign n43936 = decrypt_pad & ~\u1_uk_K_r3_reg[11]/NET0131  ;
  assign n43937 = ~decrypt_pad & ~\u1_uk_K_r3_reg[20]/NET0131  ;
  assign n43938 = ~n43936 & ~n43937 ;
  assign n43939 = \u1_R3_reg[9]/NET0131  & ~n43938 ;
  assign n43940 = ~\u1_R3_reg[9]/NET0131  & n43938 ;
  assign n43941 = ~n43939 & ~n43940 ;
  assign n43958 = ~n43935 & n43941 ;
  assign n43959 = ~n43948 & n43958 ;
  assign n43950 = decrypt_pad & ~\u1_uk_K_r3_reg[46]/NET0131  ;
  assign n43951 = ~decrypt_pad & ~\u1_uk_K_r3_reg[55]/NET0131  ;
  assign n43952 = ~n43950 & ~n43951 ;
  assign n43953 = \u1_R3_reg[6]/NET0131  & ~n43952 ;
  assign n43954 = ~\u1_R3_reg[6]/NET0131  & n43952 ;
  assign n43955 = ~n43953 & ~n43954 ;
  assign n43960 = n43935 & n43948 ;
  assign n43961 = n43935 & ~n43941 ;
  assign n43962 = ~n43960 & ~n43961 ;
  assign n43963 = n43955 & ~n43962 ;
  assign n43964 = ~n43959 & ~n43963 ;
  assign n43965 = ~n43929 & ~n43964 ;
  assign n43966 = ~n43941 & n43948 ;
  assign n43967 = ~n43959 & ~n43966 ;
  assign n43968 = ~n43955 & ~n43967 ;
  assign n43942 = n43935 & n43941 ;
  assign n43949 = n43942 & ~n43948 ;
  assign n43956 = n43949 & n43955 ;
  assign n43957 = n43929 & n43956 ;
  assign n43969 = ~n43929 & ~n43948 ;
  assign n43970 = n43941 & ~n43955 ;
  assign n43971 = n43969 & n43970 ;
  assign n43972 = n43948 & n43955 ;
  assign n43973 = n43958 & n43972 ;
  assign n43974 = ~n43971 & ~n43973 ;
  assign n43975 = ~n43957 & n43974 ;
  assign n43976 = ~n43968 & n43975 ;
  assign n43977 = ~n43965 & n43976 ;
  assign n43978 = ~n43923 & ~n43977 ;
  assign n43995 = ~n43935 & ~n43941 ;
  assign n43996 = ~n43956 & ~n43995 ;
  assign n43997 = n43923 & ~n43996 ;
  assign n43979 = ~n43948 & n43955 ;
  assign n43998 = n43958 & ~n43979 ;
  assign n43999 = ~n43997 & ~n43998 ;
  assign n43994 = n43948 & ~n43955 ;
  assign n44000 = ~n43929 & ~n43994 ;
  assign n44001 = ~n43999 & n44000 ;
  assign n43980 = ~n43941 & n43979 ;
  assign n43981 = ~n43935 & n43980 ;
  assign n43982 = ~n43955 & n43960 ;
  assign n43983 = ~n43981 & ~n43982 ;
  assign n43984 = n43929 & ~n43983 ;
  assign n43985 = ~n43948 & n43961 ;
  assign n43986 = n43942 & n43948 ;
  assign n43987 = ~n43985 & ~n43986 ;
  assign n43988 = ~n43955 & ~n43987 ;
  assign n43989 = ~n43935 & n43955 ;
  assign n43990 = n43929 & n43948 ;
  assign n43991 = ~n43989 & n43990 ;
  assign n43992 = ~n43988 & ~n43991 ;
  assign n43993 = n43923 & ~n43992 ;
  assign n44002 = ~n43984 & ~n43993 ;
  assign n44003 = ~n44001 & n44002 ;
  assign n44004 = ~n43978 & n44003 ;
  assign n44005 = \u1_L3_reg[2]/NET0131  & n44004 ;
  assign n44006 = ~\u1_L3_reg[2]/NET0131  & ~n44004 ;
  assign n44007 = ~n44005 & ~n44006 ;
  assign n44019 = n43659 & n43668 ;
  assign n44018 = n43623 & n43898 ;
  assign n44020 = n43604 & ~n44018 ;
  assign n44021 = ~n44019 & n44020 ;
  assign n44022 = ~n43662 & n44021 ;
  assign n44023 = n43616 & ~n43635 ;
  assign n44024 = ~n43670 & ~n44023 ;
  assign n44025 = n43644 & ~n44024 ;
  assign n44026 = ~n43604 & ~n43679 ;
  assign n44027 = ~n43675 & n44026 ;
  assign n44028 = ~n44025 & n44027 ;
  assign n44029 = ~n44022 & ~n44028 ;
  assign n44009 = n43629 & n43665 ;
  assign n44010 = ~n43893 & ~n44009 ;
  assign n44011 = ~n43604 & ~n44010 ;
  assign n44008 = ~n43623 & n43665 ;
  assign n44012 = ~n43616 & n43630 ;
  assign n44013 = ~n43634 & ~n44012 ;
  assign n44014 = n43604 & ~n44013 ;
  assign n44015 = ~n44008 & ~n44014 ;
  assign n44016 = ~n44011 & n44015 ;
  assign n44017 = ~n43644 & ~n44016 ;
  assign n44033 = ~n43644 & n43884 ;
  assign n44030 = ~n43666 & ~n43681 ;
  assign n44031 = n43644 & ~n43670 ;
  assign n44032 = n44030 & n44031 ;
  assign n44034 = n43623 & ~n44032 ;
  assign n44035 = ~n44033 & n44034 ;
  assign n44036 = ~n44017 & ~n44035 ;
  assign n44037 = ~n44029 & n44036 ;
  assign n44038 = ~\u1_L3_reg[4]/NET0131  & ~n44037 ;
  assign n44039 = \u1_L3_reg[4]/NET0131  & n44037 ;
  assign n44040 = ~n44038 & ~n44039 ;
  assign n44060 = decrypt_pad & ~\u1_uk_K_r3_reg[37]/NET0131  ;
  assign n44061 = ~decrypt_pad & ~\u1_uk_K_r3_reg[42]/NET0131  ;
  assign n44062 = ~n44060 & ~n44061 ;
  assign n44063 = \u1_R3_reg[29]/NET0131  & ~n44062 ;
  assign n44064 = ~\u1_R3_reg[29]/NET0131  & n44062 ;
  assign n44065 = ~n44063 & ~n44064 ;
  assign n44053 = decrypt_pad & ~\u1_uk_K_r3_reg[22]/NET0131  ;
  assign n44054 = ~decrypt_pad & ~\u1_uk_K_r3_reg[31]/NET0131  ;
  assign n44055 = ~n44053 & ~n44054 ;
  assign n44056 = \u1_R3_reg[1]/NET0131  & ~n44055 ;
  assign n44057 = ~\u1_R3_reg[1]/NET0131  & n44055 ;
  assign n44058 = ~n44056 & ~n44057 ;
  assign n44041 = decrypt_pad & ~\u1_uk_K_r3_reg[7]/NET0131  ;
  assign n44042 = ~decrypt_pad & ~\u1_uk_K_r3_reg[43]/NET0131  ;
  assign n44043 = ~n44041 & ~n44042 ;
  assign n44044 = \u1_R3_reg[30]/NET0131  & ~n44043 ;
  assign n44045 = ~\u1_R3_reg[30]/NET0131  & n44043 ;
  assign n44046 = ~n44044 & ~n44045 ;
  assign n44047 = decrypt_pad & ~\u1_uk_K_r3_reg[38]/NET0131  ;
  assign n44048 = ~decrypt_pad & ~\u1_uk_K_r3_reg[15]/NET0131  ;
  assign n44049 = ~n44047 & ~n44048 ;
  assign n44050 = \u1_R3_reg[28]/NET0131  & ~n44049 ;
  assign n44051 = ~\u1_R3_reg[28]/NET0131  & n44049 ;
  assign n44052 = ~n44050 & ~n44051 ;
  assign n44068 = ~n44046 & n44052 ;
  assign n44071 = ~n44058 & n44068 ;
  assign n44072 = n44065 & n44071 ;
  assign n44069 = ~n44058 & n44065 ;
  assign n44070 = ~n44068 & ~n44069 ;
  assign n44073 = decrypt_pad & ~\u1_uk_K_r3_reg[50]/NET0131  ;
  assign n44074 = ~decrypt_pad & ~\u1_uk_K_r3_reg[0]/NET0131  ;
  assign n44075 = ~n44073 & ~n44074 ;
  assign n44076 = \u1_R3_reg[31]/P0001  & ~n44075 ;
  assign n44077 = ~\u1_R3_reg[31]/P0001  & n44075 ;
  assign n44078 = ~n44076 & ~n44077 ;
  assign n44079 = ~n44070 & n44078 ;
  assign n44080 = ~n44072 & n44079 ;
  assign n44087 = ~n44046 & ~n44065 ;
  assign n44088 = ~n44052 & n44087 ;
  assign n44089 = ~n44078 & n44088 ;
  assign n44059 = ~n44052 & n44058 ;
  assign n44066 = n44059 & n44065 ;
  assign n44067 = n44046 & n44066 ;
  assign n44081 = decrypt_pad & ~\u1_uk_K_r3_reg[1]/NET0131  ;
  assign n44082 = ~decrypt_pad & ~\u1_uk_K_r3_reg[37]/NET0131  ;
  assign n44083 = ~n44081 & ~n44082 ;
  assign n44084 = \u1_R3_reg[32]/NET0131  & ~n44083 ;
  assign n44085 = ~\u1_R3_reg[32]/NET0131  & n44083 ;
  assign n44086 = ~n44084 & ~n44085 ;
  assign n44090 = ~n44067 & n44086 ;
  assign n44091 = ~n44089 & n44090 ;
  assign n44092 = ~n44080 & n44091 ;
  assign n44099 = n44052 & ~n44065 ;
  assign n44100 = n44046 & n44099 ;
  assign n44101 = ~n44058 & n44100 ;
  assign n44098 = n44059 & ~n44065 ;
  assign n44102 = n44078 & ~n44098 ;
  assign n44103 = ~n44101 & n44102 ;
  assign n44105 = n44046 & ~n44058 ;
  assign n44106 = ~n44052 & n44105 ;
  assign n44104 = n44058 & n44065 ;
  assign n44107 = ~n44078 & ~n44104 ;
  assign n44108 = ~n44106 & n44107 ;
  assign n44109 = ~n44103 & ~n44108 ;
  assign n44096 = ~n44069 & n44078 ;
  assign n44097 = n44068 & ~n44096 ;
  assign n44093 = n44052 & n44065 ;
  assign n44094 = n44046 & n44093 ;
  assign n44095 = n44058 & n44094 ;
  assign n44110 = ~n44086 & ~n44095 ;
  assign n44111 = ~n44097 & n44110 ;
  assign n44112 = ~n44109 & n44111 ;
  assign n44113 = ~n44092 & ~n44112 ;
  assign n44114 = ~n44078 & ~n44100 ;
  assign n44115 = ~n44078 & ~n44086 ;
  assign n44116 = ~n44114 & ~n44115 ;
  assign n44117 = ~n44072 & ~n44116 ;
  assign n44118 = n44065 & n44106 ;
  assign n44119 = ~n44058 & n44088 ;
  assign n44120 = ~n44118 & ~n44119 ;
  assign n44121 = n44046 & n44098 ;
  assign n44122 = n44058 & ~n44065 ;
  assign n44123 = n44068 & n44122 ;
  assign n44124 = n44078 & ~n44123 ;
  assign n44125 = ~n44121 & n44124 ;
  assign n44126 = n44120 & n44125 ;
  assign n44127 = ~n44117 & ~n44126 ;
  assign n44128 = ~n44113 & ~n44127 ;
  assign n44129 = \u1_L3_reg[5]/NET0131  & ~n44128 ;
  assign n44130 = ~\u1_L3_reg[5]/NET0131  & n44128 ;
  assign n44131 = ~n44129 & ~n44130 ;
  assign n44135 = n43799 & ~n43812 ;
  assign n44150 = n43822 & ~n44135 ;
  assign n44151 = ~n43854 & ~n44150 ;
  assign n44152 = ~n43806 & ~n44151 ;
  assign n44132 = ~n43799 & n43812 ;
  assign n44144 = n43852 & n44132 ;
  assign n44145 = ~n43859 & ~n44144 ;
  assign n44146 = n43793 & n43831 ;
  assign n44147 = n43819 & n44146 ;
  assign n44148 = ~n43827 & ~n44147 ;
  assign n44149 = n43806 & ~n44148 ;
  assign n44153 = n44145 & ~n44149 ;
  assign n44154 = ~n44152 & n44153 ;
  assign n44155 = n43849 & ~n44154 ;
  assign n44133 = ~n43834 & ~n44132 ;
  assign n44134 = n43806 & ~n44133 ;
  assign n44136 = ~n43820 & ~n44135 ;
  assign n44137 = ~n44134 & n44136 ;
  assign n44138 = n43793 & ~n44137 ;
  assign n44139 = ~n43835 & ~n43856 ;
  assign n44140 = ~n43838 & ~n44139 ;
  assign n44141 = ~n43828 & ~n44140 ;
  assign n44142 = ~n44138 & n44141 ;
  assign n44143 = ~n43849 & ~n44142 ;
  assign n44156 = ~n43871 & n44145 ;
  assign n44157 = ~n43806 & ~n44156 ;
  assign n44158 = ~n43839 & ~n43876 ;
  assign n44159 = ~n44157 & n44158 ;
  assign n44160 = ~n44143 & n44159 ;
  assign n44161 = ~n44155 & n44160 ;
  assign n44162 = ~\u1_L3_reg[10]/NET0131  & ~n44161 ;
  assign n44163 = \u1_L3_reg[10]/NET0131  & n44161 ;
  assign n44164 = ~n44162 & ~n44163 ;
  assign n44171 = ~n43742 & ~n43744 ;
  assign n44172 = n43753 & n44171 ;
  assign n44169 = ~n43739 & ~n43744 ;
  assign n44170 = n43755 & ~n44169 ;
  assign n44176 = ~n43701 & ~n44170 ;
  assign n44177 = ~n44172 & n44176 ;
  assign n44165 = n43726 & n43745 ;
  assign n44166 = n43719 & n43737 ;
  assign n44167 = ~n44165 & ~n44166 ;
  assign n44168 = ~n43713 & ~n44167 ;
  assign n44173 = ~n43720 & ~n43760 ;
  assign n44174 = ~n43737 & n44173 ;
  assign n44175 = ~n43734 & ~n44174 ;
  assign n44178 = ~n44168 & ~n44175 ;
  assign n44179 = n44177 & n44178 ;
  assign n44180 = ~n43734 & n43757 ;
  assign n44186 = n43701 & ~n43759 ;
  assign n44187 = ~n43774 & n44186 ;
  assign n44188 = ~n44180 & n44187 ;
  assign n44181 = ~n43736 & ~n43777 ;
  assign n44182 = n43765 & ~n44181 ;
  assign n44183 = n43713 & n43726 ;
  assign n44184 = ~n43754 & ~n44183 ;
  assign n44185 = n43734 & ~n44184 ;
  assign n44189 = ~n44182 & ~n44185 ;
  assign n44190 = n44188 & n44189 ;
  assign n44191 = ~n44179 & ~n44190 ;
  assign n44192 = \u1_L3_reg[12]/NET0131  & n44191 ;
  assign n44193 = ~\u1_L3_reg[12]/NET0131  & ~n44191 ;
  assign n44194 = ~n44192 & ~n44193 ;
  assign n44222 = decrypt_pad & ~\u1_uk_K_r3_reg[2]/NET0131  ;
  assign n44223 = ~decrypt_pad & ~\u1_uk_K_r3_reg[7]/NET0131  ;
  assign n44224 = ~n44222 & ~n44223 ;
  assign n44225 = \u1_R3_reg[19]/NET0131  & ~n44224 ;
  assign n44226 = ~\u1_R3_reg[19]/NET0131  & n44224 ;
  assign n44227 = ~n44225 & ~n44226 ;
  assign n44208 = decrypt_pad & ~\u1_uk_K_r3_reg[15]/NET0131  ;
  assign n44209 = ~decrypt_pad & ~\u1_uk_K_r3_reg[51]/NET0131  ;
  assign n44210 = ~n44208 & ~n44209 ;
  assign n44211 = \u1_R3_reg[18]/NET0131  & ~n44210 ;
  assign n44212 = ~\u1_R3_reg[18]/NET0131  & n44210 ;
  assign n44213 = ~n44211 & ~n44212 ;
  assign n44201 = decrypt_pad & ~\u1_uk_K_r3_reg[42]/NET0131  ;
  assign n44202 = ~decrypt_pad & ~\u1_uk_K_r3_reg[23]/NET0131  ;
  assign n44203 = ~n44201 & ~n44202 ;
  assign n44204 = \u1_R3_reg[21]/NET0131  & ~n44203 ;
  assign n44205 = ~\u1_R3_reg[21]/NET0131  & n44203 ;
  assign n44206 = ~n44204 & ~n44205 ;
  assign n44195 = decrypt_pad & ~\u1_uk_K_r3_reg[30]/NET0131  ;
  assign n44196 = ~decrypt_pad & ~\u1_uk_K_r3_reg[35]/NET0131  ;
  assign n44197 = ~n44195 & ~n44196 ;
  assign n44198 = \u1_R3_reg[16]/NET0131  & ~n44197 ;
  assign n44199 = ~\u1_R3_reg[16]/NET0131  & n44197 ;
  assign n44200 = ~n44198 & ~n44199 ;
  assign n44215 = decrypt_pad & ~\u1_uk_K_r3_reg[21]/NET0131  ;
  assign n44216 = ~decrypt_pad & ~\u1_uk_K_r3_reg[2]/NET0131  ;
  assign n44217 = ~n44215 & ~n44216 ;
  assign n44218 = \u1_R3_reg[17]/NET0131  & ~n44217 ;
  assign n44219 = ~\u1_R3_reg[17]/NET0131  & n44217 ;
  assign n44220 = ~n44218 & ~n44219 ;
  assign n44228 = ~n44200 & ~n44220 ;
  assign n44229 = n44206 & n44228 ;
  assign n44230 = n44213 & n44229 ;
  assign n44231 = ~n44200 & ~n44206 ;
  assign n44232 = n44213 & n44231 ;
  assign n44233 = n44220 & n44232 ;
  assign n44234 = ~n44230 & ~n44233 ;
  assign n44235 = ~n44227 & n44234 ;
  assign n44207 = ~n44200 & n44206 ;
  assign n44214 = n44207 & ~n44213 ;
  assign n44221 = n44214 & n44220 ;
  assign n44236 = ~n44213 & ~n44220 ;
  assign n44237 = n44231 & n44236 ;
  assign n44238 = ~n44221 & ~n44237 ;
  assign n44239 = n44235 & n44238 ;
  assign n44240 = n44200 & n44220 ;
  assign n44241 = ~n44206 & n44240 ;
  assign n44245 = ~n44213 & n44241 ;
  assign n44246 = ~n44220 & n44232 ;
  assign n44247 = ~n44245 & ~n44246 ;
  assign n44242 = n44227 & ~n44241 ;
  assign n44243 = n44200 & n44206 ;
  assign n44244 = ~n44213 & n44243 ;
  assign n44248 = ~n44213 & n44220 ;
  assign n44249 = n44207 & ~n44248 ;
  assign n44250 = ~n44244 & ~n44249 ;
  assign n44251 = n44242 & n44250 ;
  assign n44252 = n44247 & n44251 ;
  assign n44253 = ~n44239 & ~n44252 ;
  assign n44254 = n44213 & n44220 ;
  assign n44255 = ~n44227 & n44254 ;
  assign n44256 = ~n44236 & ~n44255 ;
  assign n44257 = n44243 & ~n44256 ;
  assign n44258 = n44213 & ~n44220 ;
  assign n44259 = n44200 & ~n44206 ;
  assign n44260 = n44258 & n44259 ;
  assign n44261 = decrypt_pad & ~\u1_uk_K_r3_reg[45]/NET0131  ;
  assign n44262 = ~decrypt_pad & ~\u1_uk_K_r3_reg[22]/NET0131  ;
  assign n44263 = ~n44261 & ~n44262 ;
  assign n44264 = \u1_R3_reg[20]/NET0131  & ~n44263 ;
  assign n44265 = ~\u1_R3_reg[20]/NET0131  & n44263 ;
  assign n44266 = ~n44264 & ~n44265 ;
  assign n44267 = ~n44260 & n44266 ;
  assign n44268 = ~n44245 & n44267 ;
  assign n44269 = ~n44257 & n44268 ;
  assign n44270 = ~n44253 & n44269 ;
  assign n44271 = n44243 & n44248 ;
  assign n44274 = ~n44229 & ~n44271 ;
  assign n44272 = n44236 & n44259 ;
  assign n44273 = ~n44206 & n44254 ;
  assign n44275 = ~n44272 & ~n44273 ;
  assign n44276 = n44274 & n44275 ;
  assign n44277 = n44235 & n44276 ;
  assign n44279 = n44206 & n44213 ;
  assign n44280 = ~n44228 & ~n44279 ;
  assign n44281 = ~n44207 & ~n44280 ;
  assign n44278 = ~n44200 & n44248 ;
  assign n44282 = n44227 & ~n44278 ;
  assign n44283 = ~n44281 & n44282 ;
  assign n44284 = n44247 & n44283 ;
  assign n44285 = ~n44277 & ~n44284 ;
  assign n44287 = ~n44206 & n44278 ;
  assign n44286 = n44243 & n44258 ;
  assign n44288 = ~n44266 & ~n44286 ;
  assign n44289 = ~n44287 & n44288 ;
  assign n44290 = ~n44285 & n44289 ;
  assign n44291 = ~n44270 & ~n44290 ;
  assign n44292 = ~\u1_L3_reg[14]/NET0131  & n44291 ;
  assign n44293 = \u1_L3_reg[14]/NET0131  & ~n44291 ;
  assign n44294 = ~n44292 & ~n44293 ;
  assign n44303 = ~n44046 & n44069 ;
  assign n44304 = ~n44093 & ~n44098 ;
  assign n44305 = ~n44303 & n44304 ;
  assign n44306 = n44078 & ~n44305 ;
  assign n44307 = ~n44065 & n44071 ;
  assign n44308 = ~n44086 & ~n44307 ;
  assign n44309 = ~n44306 & n44308 ;
  assign n44310 = ~n44046 & n44065 ;
  assign n44311 = n44052 & n44310 ;
  assign n44318 = n44086 & ~n44311 ;
  assign n44312 = ~n44052 & ~n44058 ;
  assign n44313 = ~n44065 & n44078 ;
  assign n44314 = n44312 & n44313 ;
  assign n44315 = n44046 & ~n44078 ;
  assign n44316 = n44122 & n44315 ;
  assign n44319 = ~n44314 & ~n44316 ;
  assign n44320 = n44318 & n44319 ;
  assign n44317 = n44058 & n44100 ;
  assign n44321 = ~n44118 & ~n44317 ;
  assign n44322 = n44320 & n44321 ;
  assign n44323 = ~n44309 & ~n44322 ;
  assign n44295 = ~n44046 & n44066 ;
  assign n44296 = n44114 & ~n44295 ;
  assign n44297 = n44120 & n44296 ;
  assign n44298 = n44058 & n44088 ;
  assign n44299 = ~n44067 & n44078 ;
  assign n44300 = ~n44298 & n44299 ;
  assign n44301 = ~n44297 & ~n44300 ;
  assign n44302 = n44099 & n44115 ;
  assign n44324 = ~n44301 & ~n44302 ;
  assign n44325 = ~n44323 & n44324 ;
  assign n44326 = \u1_L3_reg[15]/P0001  & n44325 ;
  assign n44327 = ~\u1_L3_reg[15]/P0001  & ~n44325 ;
  assign n44328 = ~n44326 & ~n44327 ;
  assign n44333 = ~n43929 & ~n43949 ;
  assign n44334 = ~n43980 & n44333 ;
  assign n44337 = n43941 & n43989 ;
  assign n44335 = ~n43948 & ~n43955 ;
  assign n44336 = ~n43941 & n44335 ;
  assign n44338 = n43929 & ~n44336 ;
  assign n44339 = ~n44337 & n44338 ;
  assign n44340 = ~n44334 & ~n44339 ;
  assign n44331 = n43948 & n43995 ;
  assign n44332 = ~n43955 & n44331 ;
  assign n44341 = n43923 & n43974 ;
  assign n44342 = ~n44332 & n44341 ;
  assign n44343 = ~n44340 & n44342 ;
  assign n44347 = ~n43935 & ~n43969 ;
  assign n44348 = n43970 & n44347 ;
  assign n44344 = n43929 & n43935 ;
  assign n44345 = n43955 & ~n43966 ;
  assign n44346 = n44344 & n44345 ;
  assign n44349 = ~n43923 & ~n44346 ;
  assign n44350 = ~n44348 & n44349 ;
  assign n44353 = ~n43929 & ~n44331 ;
  assign n44351 = n43958 & n43979 ;
  assign n44352 = n43961 & n44335 ;
  assign n44354 = ~n44351 & ~n44352 ;
  assign n44355 = n44353 & n44354 ;
  assign n44356 = n44350 & n44355 ;
  assign n44357 = ~n44343 & ~n44356 ;
  assign n44329 = n43961 & n43972 ;
  assign n44330 = n43941 & n43982 ;
  assign n44358 = ~n44329 & ~n44330 ;
  assign n44359 = ~n44357 & n44358 ;
  assign n44362 = ~n43942 & ~n43995 ;
  assign n44363 = ~n43948 & ~n44362 ;
  assign n44360 = ~n43955 & n43961 ;
  assign n44361 = n43948 & n44360 ;
  assign n44364 = n43929 & ~n44361 ;
  assign n44365 = ~n44363 & n44364 ;
  assign n44366 = n44350 & n44365 ;
  assign n44367 = ~n44359 & ~n44366 ;
  assign n44368 = ~\u1_L3_reg[13]/NET0131  & ~n44367 ;
  assign n44369 = \u1_L3_reg[13]/NET0131  & n44367 ;
  assign n44370 = ~n44368 & ~n44369 ;
  assign n44382 = n43610 & ~n43630 ;
  assign n44383 = ~n44009 & ~n44382 ;
  assign n44384 = n43644 & ~n44383 ;
  assign n44380 = n43629 & n43660 ;
  assign n44381 = ~n43644 & ~n44030 ;
  assign n44385 = ~n44380 & ~n44381 ;
  assign n44386 = ~n44384 & n44385 ;
  assign n44387 = ~n43604 & ~n44386 ;
  assign n44374 = n43623 & ~n44030 ;
  assign n44371 = ~n43637 & ~n43652 ;
  assign n44372 = n43644 & ~n44371 ;
  assign n44373 = n43632 & ~n43644 ;
  assign n44375 = ~n43900 & ~n44012 ;
  assign n44376 = ~n44373 & n44375 ;
  assign n44377 = ~n44372 & n44376 ;
  assign n44378 = ~n44374 & n44377 ;
  assign n44379 = n43604 & ~n44378 ;
  assign n44388 = n43672 & ~n43680 ;
  assign n44389 = ~n44379 & n44388 ;
  assign n44390 = ~n44387 & n44389 ;
  assign n44391 = ~\u1_L3_reg[19]/NET0131  & ~n44390 ;
  assign n44392 = \u1_L3_reg[19]/NET0131  & n44390 ;
  assign n44393 = ~n44391 & ~n44392 ;
  assign n44408 = ~n43824 & ~n43869 ;
  assign n44409 = n43793 & ~n44408 ;
  assign n44410 = ~n43806 & ~n44409 ;
  assign n44411 = n43806 & ~n43870 ;
  assign n44412 = ~n43873 & n44411 ;
  assign n44413 = ~n44410 & ~n44412 ;
  assign n44414 = ~n43822 & ~n43852 ;
  assign n44415 = n44135 & ~n44414 ;
  assign n44416 = ~n43859 & ~n44415 ;
  assign n44417 = ~n44413 & n44416 ;
  assign n44418 = ~n43849 & ~n44417 ;
  assign n44401 = ~n43822 & n44135 ;
  assign n44402 = ~n43853 & ~n44401 ;
  assign n44403 = ~n43806 & ~n44402 ;
  assign n44396 = n43799 & n43823 ;
  assign n44404 = ~n43793 & n44132 ;
  assign n44405 = ~n44396 & ~n44404 ;
  assign n44406 = ~n44403 & n44405 ;
  assign n44407 = n43849 & ~n44406 ;
  assign n44394 = ~n43828 & n44145 ;
  assign n44395 = n43806 & ~n44394 ;
  assign n44398 = ~n43824 & ~n44146 ;
  assign n44399 = n43806 & n43849 ;
  assign n44400 = ~n44398 & n44399 ;
  assign n44397 = ~n43806 & n44396 ;
  assign n44419 = ~n43860 & ~n44397 ;
  assign n44420 = ~n44400 & n44419 ;
  assign n44421 = ~n44395 & n44420 ;
  assign n44422 = ~n44407 & n44421 ;
  assign n44423 = ~n44418 & n44422 ;
  assign n44424 = ~\u1_L3_reg[1]/NET0131  & ~n44423 ;
  assign n44425 = \u1_L3_reg[1]/NET0131  & n44423 ;
  assign n44426 = ~n44424 & ~n44425 ;
  assign n44437 = n5837 & n43561 ;
  assign n44438 = ~n5900 & ~n43585 ;
  assign n44439 = ~n44437 & n44438 ;
  assign n44440 = ~n43575 & n44439 ;
  assign n44441 = n5883 & ~n44440 ;
  assign n44428 = n5850 & ~n5893 ;
  assign n44429 = ~n5897 & n44428 ;
  assign n44430 = n5838 & ~n5850 ;
  assign n44431 = n5865 & n44430 ;
  assign n44427 = ~n5837 & n5852 ;
  assign n44432 = ~n5891 & ~n43564 ;
  assign n44433 = ~n44427 & n44432 ;
  assign n44434 = ~n44431 & n44433 ;
  assign n44435 = ~n44429 & n44434 ;
  assign n44436 = ~n5883 & ~n44435 ;
  assign n44447 = ~n43556 & ~n44430 ;
  assign n44448 = ~n5831 & ~n44447 ;
  assign n44449 = ~n43569 & ~n44448 ;
  assign n44450 = ~n5865 & n5883 ;
  assign n44451 = ~n44449 & n44450 ;
  assign n44443 = n5850 & n5894 ;
  assign n44444 = ~n5890 & ~n44443 ;
  assign n44445 = ~n5865 & ~n44444 ;
  assign n44446 = n5858 & n43576 ;
  assign n44442 = n43572 & n44430 ;
  assign n44452 = ~n43591 & ~n44442 ;
  assign n44453 = ~n44446 & n44452 ;
  assign n44454 = ~n44445 & n44453 ;
  assign n44455 = ~n44451 & n44454 ;
  assign n44456 = ~n44436 & n44455 ;
  assign n44457 = ~n44441 & n44456 ;
  assign n44458 = \u1_L3_reg[23]/NET0131  & ~n44457 ;
  assign n44459 = ~\u1_L3_reg[23]/NET0131  & n44457 ;
  assign n44460 = ~n44458 & ~n44459 ;
  assign n44479 = n43955 & n44331 ;
  assign n44480 = n43987 & ~n44479 ;
  assign n44481 = n43929 & ~n44480 ;
  assign n44464 = ~n43955 & n43995 ;
  assign n44465 = n43948 & n43958 ;
  assign n44466 = ~n44464 & ~n44465 ;
  assign n44478 = ~n43929 & ~n44466 ;
  assign n44476 = ~n43949 & ~n44344 ;
  assign n44477 = ~n43955 & ~n44476 ;
  assign n44482 = ~n44351 & ~n44477 ;
  assign n44483 = ~n44478 & n44482 ;
  assign n44484 = ~n44481 & n44483 ;
  assign n44485 = n43923 & ~n44484 ;
  assign n44461 = ~n43948 & n43989 ;
  assign n44462 = ~n44329 & ~n44461 ;
  assign n44463 = ~n43929 & ~n44462 ;
  assign n44467 = n43929 & n44466 ;
  assign n44468 = ~n43929 & ~n43960 ;
  assign n44469 = ~n43959 & n44468 ;
  assign n44470 = ~n44360 & n44469 ;
  assign n44471 = ~n44467 & ~n44470 ;
  assign n44472 = n43979 & ~n44362 ;
  assign n44473 = ~n44329 & ~n44472 ;
  assign n44474 = ~n44471 & n44473 ;
  assign n44475 = ~n43923 & ~n44474 ;
  assign n44486 = ~n44463 & ~n44475 ;
  assign n44487 = ~n44485 & n44486 ;
  assign n44488 = ~\u1_L3_reg[28]/NET0131  & ~n44487 ;
  assign n44489 = \u1_L3_reg[28]/NET0131  & n44487 ;
  assign n44490 = ~n44488 & ~n44489 ;
  assign n44491 = ~n44220 & n44243 ;
  assign n44492 = ~n44227 & ~n44491 ;
  assign n44493 = ~n44278 & n44492 ;
  assign n44494 = n44206 & n44240 ;
  assign n44495 = n44227 & ~n44494 ;
  assign n44496 = ~n44206 & n44236 ;
  assign n44497 = ~n44228 & ~n44232 ;
  assign n44498 = ~n44496 & n44497 ;
  assign n44499 = n44495 & n44498 ;
  assign n44500 = ~n44493 & ~n44499 ;
  assign n44501 = n44206 & n44248 ;
  assign n44502 = n44213 & n44241 ;
  assign n44503 = ~n44501 & ~n44502 ;
  assign n44504 = ~n44500 & n44503 ;
  assign n44505 = n44266 & ~n44504 ;
  assign n44513 = ~n44207 & n44227 ;
  assign n44512 = ~n44254 & ~n44259 ;
  assign n44514 = ~n44240 & ~n44512 ;
  assign n44515 = ~n44513 & n44514 ;
  assign n44517 = ~n44206 & n44220 ;
  assign n44518 = n44227 & ~n44517 ;
  assign n44516 = ~n44227 & ~n44228 ;
  assign n44519 = ~n44213 & ~n44516 ;
  assign n44520 = ~n44518 & n44519 ;
  assign n44521 = ~n44515 & ~n44520 ;
  assign n44522 = ~n44266 & ~n44521 ;
  assign n44506 = ~n44246 & ~n44502 ;
  assign n44507 = n44207 & n44236 ;
  assign n44508 = n44506 & ~n44507 ;
  assign n44509 = n44227 & ~n44508 ;
  assign n44510 = n44200 & ~n44227 ;
  assign n44511 = n44258 & n44510 ;
  assign n44523 = ~n44271 & ~n44511 ;
  assign n44524 = ~n44509 & n44523 ;
  assign n44525 = ~n44522 & n44524 ;
  assign n44526 = ~n44505 & n44525 ;
  assign n44527 = ~\u1_L3_reg[25]/NET0131  & ~n44526 ;
  assign n44528 = \u1_L3_reg[25]/NET0131  & n44526 ;
  assign n44529 = ~n44527 & ~n44528 ;
  assign n44538 = ~n44237 & ~n44491 ;
  assign n44539 = n44227 & ~n44538 ;
  assign n44540 = ~n44213 & n44510 ;
  assign n44541 = n44234 & ~n44540 ;
  assign n44542 = ~n44539 & n44541 ;
  assign n44543 = n44266 & ~n44542 ;
  assign n44531 = n44207 & ~n44258 ;
  assign n44532 = n44492 & ~n44531 ;
  assign n44533 = ~n44272 & n44495 ;
  assign n44534 = ~n44532 & ~n44533 ;
  assign n44535 = ~n44278 & n44506 ;
  assign n44536 = ~n44534 & n44535 ;
  assign n44537 = ~n44266 & ~n44536 ;
  assign n44530 = ~n44227 & n44260 ;
  assign n44544 = ~n44221 & ~n44273 ;
  assign n44545 = ~n44230 & n44544 ;
  assign n44546 = n44227 & ~n44545 ;
  assign n44547 = ~n44530 & ~n44546 ;
  assign n44548 = ~n44537 & n44547 ;
  assign n44549 = ~n44543 & n44548 ;
  assign n44550 = ~\u1_L3_reg[8]/NET0131  & ~n44549 ;
  assign n44551 = \u1_L3_reg[8]/NET0131  & n44549 ;
  assign n44552 = ~n44550 & ~n44551 ;
  assign n44558 = ~n44058 & n44093 ;
  assign n44559 = ~n44066 & ~n44088 ;
  assign n44560 = ~n44558 & n44559 ;
  assign n44561 = ~n44078 & ~n44560 ;
  assign n44555 = ~n44052 & ~n44303 ;
  assign n44554 = n44052 & ~n44104 ;
  assign n44556 = n44078 & ~n44554 ;
  assign n44557 = ~n44555 & n44556 ;
  assign n44553 = n44058 & n44087 ;
  assign n44562 = ~n44067 & ~n44553 ;
  assign n44563 = ~n44101 & n44562 ;
  assign n44564 = ~n44557 & n44563 ;
  assign n44565 = ~n44561 & n44564 ;
  assign n44566 = n44086 & ~n44565 ;
  assign n44581 = ~n44072 & ~n44123 ;
  assign n44582 = ~n44118 & n44581 ;
  assign n44583 = ~n44078 & ~n44582 ;
  assign n44568 = ~n44052 & n44065 ;
  assign n44569 = ~n44058 & ~n44568 ;
  assign n44570 = ~n44310 & ~n44569 ;
  assign n44571 = n44078 & ~n44303 ;
  assign n44572 = ~n44570 & n44571 ;
  assign n44573 = ~n44121 & ~n44572 ;
  assign n44574 = ~n44086 & ~n44573 ;
  assign n44567 = n44105 & n44313 ;
  assign n44575 = n44065 & ~n44078 ;
  assign n44576 = n44312 & n44575 ;
  assign n44577 = n44052 & n44058 ;
  assign n44578 = n44315 & n44577 ;
  assign n44579 = ~n44576 & ~n44578 ;
  assign n44580 = ~n44086 & ~n44579 ;
  assign n44584 = ~n44567 & ~n44580 ;
  assign n44585 = ~n44574 & n44584 ;
  assign n44586 = ~n44583 & n44585 ;
  assign n44587 = ~n44566 & n44586 ;
  assign n44588 = ~\u1_L3_reg[27]/NET0131  & ~n44587 ;
  assign n44589 = \u1_L3_reg[27]/NET0131  & n44587 ;
  assign n44590 = ~n44588 & ~n44589 ;
  assign n44596 = ~n43755 & ~n43776 ;
  assign n44598 = ~n43742 & n44173 ;
  assign n44599 = n44596 & ~n44598 ;
  assign n44597 = ~n43742 & ~n44596 ;
  assign n44600 = ~n43734 & ~n44597 ;
  assign n44601 = ~n44599 & n44600 ;
  assign n44591 = n43744 & n43776 ;
  assign n44592 = n43707 & ~n43776 ;
  assign n44593 = n43765 & ~n44592 ;
  assign n44594 = ~n43727 & ~n44593 ;
  assign n44595 = n43734 & ~n44594 ;
  assign n44602 = ~n44591 & ~n44595 ;
  assign n44603 = ~n44601 & n44602 ;
  assign n44604 = n43701 & ~n44603 ;
  assign n44606 = ~n44165 & ~n44173 ;
  assign n44607 = ~n43734 & ~n44606 ;
  assign n44608 = ~n43713 & n43758 ;
  assign n44609 = n43734 & ~n44165 ;
  assign n44610 = ~n44608 & n44609 ;
  assign n44611 = ~n44607 & ~n44610 ;
  assign n44605 = n43713 & ~n44167 ;
  assign n44612 = n43775 & ~n44605 ;
  assign n44613 = ~n44611 & n44612 ;
  assign n44614 = ~n43701 & ~n44613 ;
  assign n44615 = n43734 & n43757 ;
  assign n44616 = ~n43745 & n43772 ;
  assign n44617 = n43738 & n44616 ;
  assign n44618 = ~n44615 & ~n44617 ;
  assign n44619 = ~n44614 & n44618 ;
  assign n44620 = ~n44604 & n44619 ;
  assign n44621 = \u1_L3_reg[32]/NET0131  & n44620 ;
  assign n44622 = ~\u1_L3_reg[32]/NET0131  & ~n44620 ;
  assign n44623 = ~n44621 & ~n44622 ;
  assign n44625 = ~n44214 & n44242 ;
  assign n44626 = ~n44231 & ~n44279 ;
  assign n44627 = n44492 & n44626 ;
  assign n44628 = ~n44625 & ~n44627 ;
  assign n44624 = n44258 & ~n44259 ;
  assign n44629 = ~n44266 & ~n44624 ;
  assign n44630 = ~n44628 & n44629 ;
  assign n44634 = ~n44200 & n44517 ;
  assign n44635 = ~n44244 & ~n44634 ;
  assign n44636 = n44227 & ~n44635 ;
  assign n44631 = n44207 & ~n44227 ;
  assign n44632 = ~n44244 & ~n44631 ;
  assign n44633 = n44220 & ~n44632 ;
  assign n44637 = n44267 & ~n44633 ;
  assign n44638 = ~n44636 & n44637 ;
  assign n44639 = ~n44630 & ~n44638 ;
  assign n44640 = ~n44227 & ~n44237 ;
  assign n44641 = ~n44286 & n44640 ;
  assign n44642 = ~n44245 & n44641 ;
  assign n44643 = n44227 & ~n44272 ;
  assign n44644 = ~n44230 & n44643 ;
  assign n44645 = ~n44642 & ~n44644 ;
  assign n44646 = ~n44639 & ~n44645 ;
  assign n44647 = ~\u1_L3_reg[3]/NET0131  & ~n44646 ;
  assign n44648 = \u1_L3_reg[3]/NET0131  & n44646 ;
  assign n44649 = ~n44647 & ~n44648 ;
  assign n44667 = ~n43726 & ~n44171 ;
  assign n44650 = n43713 & ~n44596 ;
  assign n44668 = n43707 & n43776 ;
  assign n44669 = ~n44650 & ~n44668 ;
  assign n44670 = ~n44667 & n44669 ;
  assign n44671 = ~n43734 & ~n44670 ;
  assign n44651 = ~n44608 & ~n44650 ;
  assign n44652 = n43707 & ~n44651 ;
  assign n44661 = ~n43707 & ~n43720 ;
  assign n44662 = n44596 & n44661 ;
  assign n44672 = n43734 & n44662 ;
  assign n44673 = ~n44652 & ~n44672 ;
  assign n44674 = ~n44671 & n44673 ;
  assign n44675 = n43701 & ~n44674 ;
  assign n44653 = ~n43734 & n44652 ;
  assign n44654 = n43701 & ~n43734 ;
  assign n44655 = n43764 & ~n44596 ;
  assign n44656 = n43719 & ~n44183 ;
  assign n44657 = n43734 & n44592 ;
  assign n44658 = ~n44656 & n44657 ;
  assign n44659 = ~n44655 & ~n44658 ;
  assign n44660 = ~n43701 & ~n44659 ;
  assign n44663 = ~n43734 & n44662 ;
  assign n44664 = ~n43728 & ~n44663 ;
  assign n44665 = ~n44660 & n44664 ;
  assign n44666 = ~n44654 & ~n44665 ;
  assign n44676 = ~n44653 & ~n44666 ;
  assign n44677 = ~n44675 & n44676 ;
  assign n44678 = ~\u1_L3_reg[7]/NET0131  & ~n44677 ;
  assign n44679 = \u1_L3_reg[7]/NET0131  & n44677 ;
  assign n44680 = ~n44678 & ~n44679 ;
  assign n44700 = decrypt_pad & ~\u1_uk_K_r3_reg[26]/NET0131  ;
  assign n44701 = ~decrypt_pad & ~\u1_uk_K_r3_reg[3]/NET0131  ;
  assign n44702 = ~n44700 & ~n44701 ;
  assign n44703 = \u1_R3_reg[11]/NET0131  & ~n44702 ;
  assign n44704 = ~\u1_R3_reg[11]/NET0131  & n44702 ;
  assign n44705 = ~n44703 & ~n44704 ;
  assign n44681 = decrypt_pad & ~\u1_uk_K_r3_reg[41]/NET0131  ;
  assign n44682 = ~decrypt_pad & ~\u1_uk_K_r3_reg[18]/NET0131  ;
  assign n44683 = ~n44681 & ~n44682 ;
  assign n44684 = \u1_R3_reg[12]/NET0131  & ~n44683 ;
  assign n44685 = ~\u1_R3_reg[12]/NET0131  & n44683 ;
  assign n44686 = ~n44684 & ~n44685 ;
  assign n44687 = decrypt_pad & ~\u1_uk_K_r3_reg[54]/NET0131  ;
  assign n44688 = ~decrypt_pad & ~\u1_uk_K_r3_reg[6]/NET0131  ;
  assign n44689 = ~n44687 & ~n44688 ;
  assign n44690 = \u1_R3_reg[13]/NET0131  & ~n44689 ;
  assign n44691 = ~\u1_R3_reg[13]/NET0131  & n44689 ;
  assign n44692 = ~n44690 & ~n44691 ;
  assign n44693 = decrypt_pad & ~\u1_uk_K_r3_reg[17]/NET0131  ;
  assign n44694 = ~decrypt_pad & ~\u1_uk_K_r3_reg[26]/NET0131  ;
  assign n44695 = ~n44693 & ~n44694 ;
  assign n44696 = \u1_R3_reg[9]/NET0131  & ~n44695 ;
  assign n44697 = ~\u1_R3_reg[9]/NET0131  & n44695 ;
  assign n44698 = ~n44696 & ~n44697 ;
  assign n44714 = n44692 & ~n44698 ;
  assign n44707 = decrypt_pad & ~\u1_uk_K_r3_reg[25]/NET0131  ;
  assign n44708 = ~decrypt_pad & ~\u1_uk_K_r3_reg[34]/NET0131  ;
  assign n44709 = ~n44707 & ~n44708 ;
  assign n44710 = \u1_R3_reg[10]/NET0131  & ~n44709 ;
  assign n44711 = ~\u1_R3_reg[10]/NET0131  & n44709 ;
  assign n44712 = ~n44710 & ~n44711 ;
  assign n44715 = decrypt_pad & ~\u1_uk_K_r3_reg[20]/NET0131  ;
  assign n44716 = ~decrypt_pad & ~\u1_uk_K_r3_reg[54]/NET0131  ;
  assign n44717 = ~n44715 & ~n44716 ;
  assign n44718 = \u1_R3_reg[8]/NET0131  & ~n44717 ;
  assign n44719 = ~\u1_R3_reg[8]/NET0131  & n44717 ;
  assign n44720 = ~n44718 & ~n44719 ;
  assign n44742 = n44692 & ~n44720 ;
  assign n44743 = n44712 & n44742 ;
  assign n44699 = ~n44692 & n44698 ;
  assign n44744 = n44699 & n44720 ;
  assign n44745 = ~n44743 & ~n44744 ;
  assign n44746 = ~n44714 & n44745 ;
  assign n44747 = n44686 & ~n44746 ;
  assign n44741 = n44712 & n44714 ;
  assign n44724 = ~n44692 & ~n44720 ;
  assign n44748 = ~n44698 & n44724 ;
  assign n44749 = ~n44712 & n44748 ;
  assign n44750 = ~n44741 & ~n44749 ;
  assign n44751 = ~n44747 & n44750 ;
  assign n44752 = n44705 & ~n44751 ;
  assign n44706 = ~n44699 & ~n44705 ;
  assign n44713 = n44698 & ~n44712 ;
  assign n44721 = ~n44714 & n44720 ;
  assign n44722 = ~n44713 & ~n44721 ;
  assign n44723 = n44706 & ~n44722 ;
  assign n44725 = n44698 & n44712 ;
  assign n44726 = n44724 & n44725 ;
  assign n44727 = ~n44723 & ~n44726 ;
  assign n44728 = n44686 & ~n44727 ;
  assign n44731 = ~n44698 & ~n44712 ;
  assign n44732 = ~n44725 & ~n44731 ;
  assign n44729 = n44692 & n44720 ;
  assign n44730 = ~n44724 & ~n44729 ;
  assign n44733 = n44705 & ~n44720 ;
  assign n44737 = n44730 & ~n44733 ;
  assign n44738 = ~n44732 & ~n44737 ;
  assign n44734 = ~n44712 & n44733 ;
  assign n44735 = n44730 & n44732 ;
  assign n44736 = ~n44734 & n44735 ;
  assign n44739 = ~n44686 & ~n44736 ;
  assign n44740 = ~n44738 & n44739 ;
  assign n44753 = ~n44728 & ~n44740 ;
  assign n44754 = ~n44752 & n44753 ;
  assign n44755 = ~\u1_L3_reg[6]/NET0131  & ~n44754 ;
  assign n44756 = \u1_L3_reg[6]/NET0131  & n44754 ;
  assign n44757 = ~n44755 & ~n44756 ;
  assign n44773 = n5859 & ~n44448 ;
  assign n44774 = n5844 & ~n44773 ;
  assign n44765 = n5837 & ~n5869 ;
  assign n44766 = ~n43556 & ~n44765 ;
  assign n44772 = n43572 & n44766 ;
  assign n44775 = ~n5890 & ~n44772 ;
  assign n44776 = ~n44774 & n44775 ;
  assign n44777 = n5883 & ~n44776 ;
  assign n44758 = ~n5844 & n5858 ;
  assign n44759 = ~n5831 & n5891 ;
  assign n44760 = ~n44758 & ~n44759 ;
  assign n44761 = ~n5865 & ~n44760 ;
  assign n44763 = ~n5876 & n44447 ;
  assign n44764 = n5865 & ~n44763 ;
  assign n44767 = ~n5865 & n44766 ;
  assign n44762 = n5844 & n5871 ;
  assign n44768 = ~n44758 & ~n44762 ;
  assign n44769 = ~n44767 & n44768 ;
  assign n44770 = ~n44764 & n44769 ;
  assign n44771 = ~n5883 & ~n44770 ;
  assign n44778 = ~n44761 & ~n44771 ;
  assign n44779 = ~n44777 & n44778 ;
  assign n44780 = ~\u1_L3_reg[9]/NET0131  & ~n44779 ;
  assign n44781 = \u1_L3_reg[9]/NET0131  & n44779 ;
  assign n44782 = ~n44780 & ~n44781 ;
  assign n44785 = n44698 & n44729 ;
  assign n44786 = ~n44698 & n44742 ;
  assign n44787 = ~n44785 & ~n44786 ;
  assign n44788 = ~n44692 & n44720 ;
  assign n44789 = ~n44698 & n44788 ;
  assign n44790 = n44699 & n44733 ;
  assign n44791 = ~n44789 & ~n44790 ;
  assign n44792 = n44787 & n44791 ;
  assign n44793 = ~n44712 & ~n44792 ;
  assign n44794 = n44712 & n44724 ;
  assign n44795 = ~n44712 & n44788 ;
  assign n44796 = ~n44794 & ~n44795 ;
  assign n44797 = ~n44705 & ~n44796 ;
  assign n44783 = n44698 & n44742 ;
  assign n44784 = n44712 & n44783 ;
  assign n44798 = n44686 & ~n44784 ;
  assign n44799 = ~n44797 & n44798 ;
  assign n44800 = ~n44793 & n44799 ;
  assign n44801 = ~n44712 & n44724 ;
  assign n44802 = n44787 & ~n44801 ;
  assign n44803 = ~n44705 & ~n44802 ;
  assign n44804 = ~n44698 & ~n44729 ;
  assign n44805 = n44705 & ~n44724 ;
  assign n44806 = ~n44785 & n44805 ;
  assign n44807 = ~n44804 & n44806 ;
  assign n44808 = ~n44686 & ~n44749 ;
  assign n44809 = ~n44807 & n44808 ;
  assign n44810 = ~n44803 & n44809 ;
  assign n44811 = ~n44800 & ~n44810 ;
  assign n44816 = n44705 & ~n44744 ;
  assign n44817 = ~n44748 & n44816 ;
  assign n44812 = n44712 & n44720 ;
  assign n44813 = ~n44698 & n44812 ;
  assign n44814 = ~n44705 & ~n44813 ;
  assign n44815 = n44705 & ~n44712 ;
  assign n44818 = ~n44814 & ~n44815 ;
  assign n44819 = ~n44817 & n44818 ;
  assign n44820 = ~n44811 & ~n44819 ;
  assign n44821 = ~\u1_L3_reg[16]/NET0131  & ~n44820 ;
  assign n44822 = \u1_L3_reg[16]/NET0131  & n44820 ;
  assign n44823 = ~n44821 & ~n44822 ;
  assign n44825 = n43935 & n43970 ;
  assign n44826 = ~n43985 & ~n44825 ;
  assign n44827 = ~n43929 & ~n44826 ;
  assign n44824 = n43929 & ~n43967 ;
  assign n44828 = n43923 & ~n43981 ;
  assign n44829 = ~n44824 & n44828 ;
  assign n44830 = ~n44827 & n44829 ;
  assign n44832 = ~n43929 & n43972 ;
  assign n44833 = ~n44335 & ~n44832 ;
  assign n44834 = ~n43935 & ~n44833 ;
  assign n44835 = ~n43923 & ~n44329 ;
  assign n44836 = ~n44336 & n44835 ;
  assign n44831 = n43929 & n43986 ;
  assign n44837 = ~n43956 & ~n44831 ;
  assign n44838 = n44836 & n44837 ;
  assign n44839 = ~n44834 & n44838 ;
  assign n44840 = ~n44830 & ~n44839 ;
  assign n44841 = ~n43929 & n44465 ;
  assign n44842 = n43942 & n43955 ;
  assign n44843 = ~n44332 & ~n44842 ;
  assign n44844 = n43929 & ~n44843 ;
  assign n44845 = ~n44841 & ~n44844 ;
  assign n44846 = ~n44840 & n44845 ;
  assign n44847 = \u1_L3_reg[18]/NET0131  & n44846 ;
  assign n44848 = ~\u1_L3_reg[18]/NET0131  & ~n44846 ;
  assign n44849 = ~n44847 & ~n44848 ;
  assign n44864 = ~n44712 & n44742 ;
  assign n44865 = ~n44794 & ~n44864 ;
  assign n44866 = n44698 & n44724 ;
  assign n44867 = ~n44813 & ~n44866 ;
  assign n44868 = n44865 & n44867 ;
  assign n44869 = n44705 & ~n44868 ;
  assign n44870 = n44712 & n44789 ;
  assign n44871 = ~n44869 & ~n44870 ;
  assign n44872 = ~n44686 & ~n44871 ;
  assign n44853 = ~n44705 & ~n44731 ;
  assign n44854 = ~n44788 & n44853 ;
  assign n44855 = ~n44698 & n44815 ;
  assign n44856 = ~n44854 & ~n44855 ;
  assign n44857 = ~n44742 & ~n44856 ;
  assign n44852 = n44731 & n44737 ;
  assign n44858 = n44720 & n44725 ;
  assign n44859 = ~n44743 & ~n44858 ;
  assign n44860 = n44705 & ~n44859 ;
  assign n44861 = ~n44852 & ~n44860 ;
  assign n44862 = ~n44857 & n44861 ;
  assign n44863 = n44686 & ~n44862 ;
  assign n44875 = ~n44730 & n44731 ;
  assign n44876 = n44745 & ~n44875 ;
  assign n44877 = ~n44686 & ~n44705 ;
  assign n44878 = ~n44876 & n44877 ;
  assign n44850 = ~n44705 & n44712 ;
  assign n44851 = n44785 & n44850 ;
  assign n44873 = ~n44783 & ~n44789 ;
  assign n44874 = n44815 & ~n44873 ;
  assign n44879 = ~n44851 & ~n44874 ;
  assign n44880 = ~n44878 & n44879 ;
  assign n44881 = ~n44863 & n44880 ;
  assign n44882 = ~n44872 & n44881 ;
  assign n44883 = ~\u1_L3_reg[24]/NET0131  & ~n44882 ;
  assign n44884 = \u1_L3_reg[24]/NET0131  & n44882 ;
  assign n44885 = ~n44883 & ~n44884 ;
  assign n44887 = ~n44705 & ~n44812 ;
  assign n44888 = ~n44866 & n44887 ;
  assign n44889 = n44731 & n44788 ;
  assign n44890 = n44705 & ~n44889 ;
  assign n44891 = n44865 & n44890 ;
  assign n44892 = ~n44888 & ~n44891 ;
  assign n44893 = n44686 & ~n44892 ;
  assign n44894 = ~n44712 & ~n44786 ;
  assign n44895 = ~n44743 & ~n44894 ;
  assign n44896 = ~n44698 & ~n44788 ;
  assign n44897 = ~n44706 & ~n44896 ;
  assign n44898 = ~n44895 & ~n44897 ;
  assign n44899 = ~n44699 & n44812 ;
  assign n44900 = ~n44692 & n44713 ;
  assign n44901 = ~n44899 & ~n44900 ;
  assign n44902 = n44705 & ~n44901 ;
  assign n44903 = ~n44686 & ~n44902 ;
  assign n44904 = ~n44898 & n44903 ;
  assign n44905 = ~n44893 & ~n44904 ;
  assign n44908 = n44705 & n44714 ;
  assign n44909 = n44812 & n44908 ;
  assign n44886 = n44699 & n44850 ;
  assign n44906 = n44686 & n44725 ;
  assign n44907 = ~n44729 & n44906 ;
  assign n44910 = ~n44886 & ~n44907 ;
  assign n44911 = ~n44909 & n44910 ;
  assign n44912 = ~n44905 & n44911 ;
  assign n44913 = \u1_L3_reg[30]/NET0131  & ~n44912 ;
  assign n44914 = ~\u1_L3_reg[30]/NET0131  & n44912 ;
  assign n44915 = ~n44913 & ~n44914 ;
  assign n44916 = decrypt_pad & ~\u1_uk_K_r2_reg[22]/NET0131  ;
  assign n44917 = ~decrypt_pad & ~\u1_uk_K_r2_reg[0]/NET0131  ;
  assign n44918 = ~n44916 & ~n44917 ;
  assign n44919 = \u1_R2_reg[28]/NET0131  & ~n44918 ;
  assign n44920 = ~\u1_R2_reg[28]/NET0131  & n44918 ;
  assign n44921 = ~n44919 & ~n44920 ;
  assign n44922 = decrypt_pad & ~\u1_uk_K_r2_reg[2]/NET0131  ;
  assign n44923 = ~decrypt_pad & ~\u1_uk_K_r2_reg[35]/NET0131  ;
  assign n44924 = ~n44922 & ~n44923 ;
  assign n44925 = \u1_R2_reg[26]/NET0131  & ~n44924 ;
  assign n44926 = ~\u1_R2_reg[26]/NET0131  & n44924 ;
  assign n44927 = ~n44925 & ~n44926 ;
  assign n44928 = decrypt_pad & ~\u1_uk_K_r2_reg[45]/NET0131  ;
  assign n44929 = ~decrypt_pad & ~\u1_uk_K_r2_reg[50]/NET0131  ;
  assign n44930 = ~n44928 & ~n44929 ;
  assign n44931 = \u1_R2_reg[25]/NET0131  & ~n44930 ;
  assign n44932 = ~\u1_R2_reg[25]/NET0131  & n44930 ;
  assign n44933 = ~n44931 & ~n44932 ;
  assign n44962 = ~n44927 & ~n44933 ;
  assign n44934 = decrypt_pad & ~\u1_uk_K_r2_reg[14]/NET0131  ;
  assign n44935 = ~decrypt_pad & ~\u1_uk_K_r2_reg[23]/NET0131  ;
  assign n44936 = ~n44934 & ~n44935 ;
  assign n44937 = \u1_R2_reg[29]/NET0131  & ~n44936 ;
  assign n44938 = ~\u1_R2_reg[29]/NET0131  & n44936 ;
  assign n44939 = ~n44937 & ~n44938 ;
  assign n44965 = ~n44927 & ~n44939 ;
  assign n44985 = ~n44962 & ~n44965 ;
  assign n44941 = decrypt_pad & ~\u1_uk_K_r2_reg[37]/NET0131  ;
  assign n44942 = ~decrypt_pad & ~\u1_uk_K_r2_reg[15]/NET0131  ;
  assign n44943 = ~n44941 & ~n44942 ;
  assign n44944 = \u1_R2_reg[24]/NET0131  & ~n44943 ;
  assign n44945 = ~\u1_R2_reg[24]/NET0131  & n44943 ;
  assign n44946 = ~n44944 & ~n44945 ;
  assign n44949 = decrypt_pad & ~\u1_uk_K_r2_reg[35]/NET0131  ;
  assign n44950 = ~decrypt_pad & ~\u1_uk_K_r2_reg[44]/NET0131  ;
  assign n44951 = ~n44949 & ~n44950 ;
  assign n44952 = \u1_R2_reg[27]/NET0131  & ~n44951 ;
  assign n44953 = ~\u1_R2_reg[27]/NET0131  & n44951 ;
  assign n44954 = ~n44952 & ~n44953 ;
  assign n44964 = n44927 & n44933 ;
  assign n44984 = n44954 & ~n44964 ;
  assign n44986 = n44946 & n44984 ;
  assign n44987 = n44985 & n44986 ;
  assign n44978 = n44939 & n44946 ;
  assign n44979 = n44962 & n44978 ;
  assign n44980 = n44933 & n44939 ;
  assign n44981 = ~n44946 & n44980 ;
  assign n44982 = ~n44979 & ~n44981 ;
  assign n44983 = ~n44954 & ~n44982 ;
  assign n44973 = ~n44939 & ~n44946 ;
  assign n44974 = n44962 & n44973 ;
  assign n44975 = n44939 & ~n44946 ;
  assign n44976 = n44927 & ~n44933 ;
  assign n44977 = n44975 & n44976 ;
  assign n44988 = ~n44974 & ~n44977 ;
  assign n44989 = ~n44983 & n44988 ;
  assign n44990 = ~n44987 & n44989 ;
  assign n44991 = n44921 & ~n44990 ;
  assign n44966 = ~n44954 & ~n44964 ;
  assign n44967 = ~n44965 & n44966 ;
  assign n44963 = n44954 & ~n44962 ;
  assign n44968 = n44946 & ~n44963 ;
  assign n44969 = ~n44967 & n44968 ;
  assign n44940 = ~n44933 & ~n44939 ;
  assign n44947 = n44940 & ~n44946 ;
  assign n44948 = n44927 & n44947 ;
  assign n44955 = n44948 & ~n44954 ;
  assign n44956 = ~n44927 & ~n44946 ;
  assign n44957 = n44927 & n44946 ;
  assign n44958 = ~n44956 & ~n44957 ;
  assign n44959 = ~n44933 & n44954 ;
  assign n44960 = n44939 & ~n44959 ;
  assign n44961 = ~n44958 & n44960 ;
  assign n44970 = ~n44955 & ~n44961 ;
  assign n44971 = ~n44969 & n44970 ;
  assign n44972 = ~n44921 & ~n44971 ;
  assign n44994 = n44964 & n44973 ;
  assign n44995 = ~n44977 & ~n44994 ;
  assign n44996 = ~n44939 & n44946 ;
  assign n44997 = ~n44933 & n44996 ;
  assign n44998 = n44995 & ~n44997 ;
  assign n44999 = n44954 & ~n44998 ;
  assign n44992 = n44933 & ~n44954 ;
  assign n44993 = ~n44958 & n44992 ;
  assign n45000 = n44959 & n44965 ;
  assign n45001 = ~n44993 & ~n45000 ;
  assign n45002 = ~n44999 & n45001 ;
  assign n45003 = ~n44972 & n45002 ;
  assign n45004 = ~n44991 & n45003 ;
  assign n45005 = ~\u1_L2_reg[22]/NET0131  & ~n45004 ;
  assign n45006 = \u1_L2_reg[22]/NET0131  & n45004 ;
  assign n45007 = ~n45005 & ~n45006 ;
  assign n45008 = decrypt_pad & ~\u1_uk_K_r2_reg[48]/NET0131  ;
  assign n45009 = ~decrypt_pad & ~\u1_uk_K_r2_reg[53]/P0001  ;
  assign n45010 = ~n45008 & ~n45009 ;
  assign n45011 = \u1_R2_reg[4]/NET0131  & ~n45010 ;
  assign n45012 = ~\u1_R2_reg[4]/NET0131  & n45010 ;
  assign n45013 = ~n45011 & ~n45012 ;
  assign n45033 = decrypt_pad & ~\u1_uk_K_r2_reg[25]/NET0131  ;
  assign n45034 = ~decrypt_pad & ~\u1_uk_K_r2_reg[5]/NET0131  ;
  assign n45035 = ~n45033 & ~n45034 ;
  assign n45036 = \u1_R2_reg[32]/NET0131  & ~n45035 ;
  assign n45037 = ~\u1_R2_reg[32]/NET0131  & n45035 ;
  assign n45038 = ~n45036 & ~n45037 ;
  assign n45042 = decrypt_pad & ~\u1_uk_K_r2_reg[46]/NET0131  ;
  assign n45043 = ~decrypt_pad & ~\u1_uk_K_r2_reg[26]/NET0131  ;
  assign n45044 = ~n45042 & ~n45043 ;
  assign n45045 = \u1_R2_reg[1]/NET0131  & ~n45044 ;
  assign n45046 = ~\u1_R2_reg[1]/NET0131  & n45044 ;
  assign n45047 = ~n45045 & ~n45046 ;
  assign n45014 = decrypt_pad & ~\u1_uk_K_r2_reg[4]/NET0131  ;
  assign n45015 = ~decrypt_pad & ~\u1_uk_K_r2_reg[41]/NET0131  ;
  assign n45016 = ~n45014 & ~n45015 ;
  assign n45017 = \u1_R2_reg[2]/NET0131  & ~n45016 ;
  assign n45018 = ~\u1_R2_reg[2]/NET0131  & n45016 ;
  assign n45019 = ~n45017 & ~n45018 ;
  assign n45027 = decrypt_pad & ~\u1_uk_K_r2_reg[19]/NET0131  ;
  assign n45028 = ~decrypt_pad & ~\u1_uk_K_r2_reg[24]/NET0131  ;
  assign n45029 = ~n45027 & ~n45028 ;
  assign n45030 = \u1_R2_reg[5]/NET0131  & ~n45029 ;
  assign n45031 = ~\u1_R2_reg[5]/NET0131  & n45029 ;
  assign n45032 = ~n45030 & ~n45031 ;
  assign n45075 = ~n45019 & ~n45032 ;
  assign n45076 = ~n45047 & n45075 ;
  assign n45077 = n45038 & ~n45076 ;
  assign n45040 = ~n45032 & ~n45038 ;
  assign n45020 = decrypt_pad & ~\u1_uk_K_r2_reg[13]/NET0131  ;
  assign n45021 = ~decrypt_pad & ~\u1_uk_K_r2_reg[18]/NET0131  ;
  assign n45022 = ~n45020 & ~n45021 ;
  assign n45023 = \u1_R2_reg[3]/NET0131  & ~n45022 ;
  assign n45024 = ~\u1_R2_reg[3]/NET0131  & n45022 ;
  assign n45025 = ~n45023 & ~n45024 ;
  assign n45073 = ~n45019 & n45025 ;
  assign n45074 = n45047 & ~n45073 ;
  assign n45078 = ~n45040 & ~n45074 ;
  assign n45079 = ~n45077 & n45078 ;
  assign n45056 = n45032 & ~n45047 ;
  assign n45066 = n45019 & ~n45038 ;
  assign n45067 = ~n45032 & n45066 ;
  assign n45068 = ~n45056 & ~n45067 ;
  assign n45069 = n45025 & ~n45068 ;
  assign n45070 = ~n45038 & n45047 ;
  assign n45050 = ~n45025 & n45047 ;
  assign n45071 = ~n45050 & ~n45066 ;
  assign n45072 = ~n45070 & ~n45071 ;
  assign n45080 = ~n45069 & ~n45072 ;
  assign n45081 = ~n45079 & n45080 ;
  assign n45082 = n45013 & ~n45081 ;
  assign n45057 = ~n45019 & ~n45038 ;
  assign n45058 = n45038 & ~n45047 ;
  assign n45059 = n45019 & n45058 ;
  assign n45060 = ~n45057 & ~n45059 ;
  assign n45061 = ~n45025 & ~n45056 ;
  assign n45062 = ~n45060 & n45061 ;
  assign n45026 = n45019 & n45025 ;
  assign n45039 = n45032 & n45038 ;
  assign n45041 = ~n45039 & ~n45040 ;
  assign n45048 = n45041 & n45047 ;
  assign n45049 = n45026 & n45048 ;
  assign n45051 = n45039 & ~n45050 ;
  assign n45052 = ~n45032 & n45047 ;
  assign n45053 = ~n45038 & n45052 ;
  assign n45054 = ~n45051 & ~n45053 ;
  assign n45055 = ~n45019 & ~n45054 ;
  assign n45063 = ~n45049 & ~n45055 ;
  assign n45064 = ~n45062 & n45063 ;
  assign n45065 = ~n45013 & ~n45064 ;
  assign n45083 = n45025 & ~n45047 ;
  assign n45084 = ~n45019 & n45038 ;
  assign n45085 = ~n45067 & ~n45084 ;
  assign n45086 = n45083 & ~n45085 ;
  assign n45088 = n45019 & n45032 ;
  assign n45089 = n45047 & n45088 ;
  assign n45090 = n45038 & n45089 ;
  assign n45087 = n45056 & n45066 ;
  assign n45091 = n45047 & n45075 ;
  assign n45092 = ~n45087 & ~n45091 ;
  assign n45093 = ~n45090 & n45092 ;
  assign n45094 = ~n45025 & ~n45093 ;
  assign n45095 = ~n45086 & ~n45094 ;
  assign n45096 = ~n45065 & n45095 ;
  assign n45097 = ~n45082 & n45096 ;
  assign n45098 = ~\u1_L2_reg[31]/NET0131  & ~n45097 ;
  assign n45099 = \u1_L2_reg[31]/NET0131  & n45097 ;
  assign n45100 = ~n45098 & ~n45099 ;
  assign n45155 = decrypt_pad & ~\u1_uk_K_r2_reg[15]/NET0131  ;
  assign n45156 = ~decrypt_pad & ~\u1_uk_K_r2_reg[52]/NET0131  ;
  assign n45157 = ~n45155 & ~n45156 ;
  assign n45158 = \u1_R2_reg[24]/NET0131  & ~n45157 ;
  assign n45159 = ~\u1_R2_reg[24]/NET0131  & n45157 ;
  assign n45160 = ~n45158 & ~n45159 ;
  assign n45124 = decrypt_pad & ~\u1_uk_K_r2_reg[44]/NET0131  ;
  assign n45125 = ~decrypt_pad & ~\u1_uk_K_r2_reg[22]/NET0131  ;
  assign n45126 = ~n45124 & ~n45125 ;
  assign n45127 = \u1_R2_reg[23]/NET0131  & ~n45126 ;
  assign n45128 = ~\u1_R2_reg[23]/NET0131  & n45126 ;
  assign n45129 = ~n45127 & ~n45128 ;
  assign n45101 = decrypt_pad & ~\u1_uk_K_r2_reg[9]/NET0131  ;
  assign n45102 = ~decrypt_pad & ~\u1_uk_K_r2_reg[42]/NET0131  ;
  assign n45103 = ~n45101 & ~n45102 ;
  assign n45104 = \u1_R2_reg[21]/NET0131  & ~n45103 ;
  assign n45105 = ~\u1_R2_reg[21]/NET0131  & n45103 ;
  assign n45106 = ~n45104 & ~n45105 ;
  assign n45107 = decrypt_pad & ~\u1_uk_K_r2_reg[49]/NET0131  ;
  assign n45108 = ~decrypt_pad & ~\u1_uk_K_r2_reg[31]/NET0131  ;
  assign n45109 = ~n45107 & ~n45108 ;
  assign n45110 = \u1_R2_reg[20]/NET0131  & ~n45109 ;
  assign n45111 = ~\u1_R2_reg[20]/NET0131  & n45109 ;
  assign n45112 = ~n45110 & ~n45111 ;
  assign n45113 = n45106 & ~n45112 ;
  assign n45114 = decrypt_pad & ~\u1_uk_K_r2_reg[0]/NET0131  ;
  assign n45115 = ~decrypt_pad & ~\u1_uk_K_r2_reg[9]/NET0131  ;
  assign n45116 = ~n45114 & ~n45115 ;
  assign n45117 = \u1_R2_reg[22]/NET0131  & ~n45116 ;
  assign n45118 = ~\u1_R2_reg[22]/NET0131  & n45116 ;
  assign n45119 = ~n45117 & ~n45118 ;
  assign n45120 = n45113 & n45119 ;
  assign n45132 = decrypt_pad & ~\u1_uk_K_r2_reg[38]/NET0131  ;
  assign n45133 = ~decrypt_pad & ~\u1_uk_K_r2_reg[43]/NET0131  ;
  assign n45134 = ~n45132 & ~n45133 ;
  assign n45135 = \u1_R2_reg[25]/NET0131  & ~n45134 ;
  assign n45136 = ~\u1_R2_reg[25]/NET0131  & n45134 ;
  assign n45137 = ~n45135 & ~n45136 ;
  assign n45180 = n45106 & ~n45137 ;
  assign n45181 = n45112 & ~n45180 ;
  assign n45138 = ~n45119 & ~n45137 ;
  assign n45182 = ~n45106 & ~n45138 ;
  assign n45183 = n45181 & ~n45182 ;
  assign n45184 = ~n45120 & ~n45183 ;
  assign n45185 = n45129 & ~n45184 ;
  assign n45143 = n45112 & n45137 ;
  assign n45176 = ~n45113 & ~n45143 ;
  assign n45177 = n45119 & ~n45176 ;
  assign n45148 = ~n45112 & n45137 ;
  assign n45174 = n45106 & n45148 ;
  assign n45175 = ~n45119 & ~n45174 ;
  assign n45178 = ~n45129 & ~n45175 ;
  assign n45179 = ~n45177 & n45178 ;
  assign n45170 = ~n45119 & ~n45129 ;
  assign n45186 = n45143 & n45170 ;
  assign n45187 = ~n45106 & n45186 ;
  assign n45188 = ~n45179 & ~n45187 ;
  assign n45189 = ~n45185 & n45188 ;
  assign n45190 = n45160 & ~n45189 ;
  assign n45121 = n45106 & n45112 ;
  assign n45122 = ~n45119 & n45121 ;
  assign n45123 = ~n45120 & ~n45122 ;
  assign n45130 = ~n45123 & ~n45129 ;
  assign n45139 = ~n45106 & n45129 ;
  assign n45149 = n45139 & n45148 ;
  assign n45146 = n45121 & n45138 ;
  assign n45131 = ~n45119 & n45129 ;
  assign n45147 = ~n45112 & n45131 ;
  assign n45150 = ~n45146 & ~n45147 ;
  assign n45151 = ~n45149 & n45150 ;
  assign n45140 = ~n45138 & ~n45139 ;
  assign n45141 = n45112 & ~n45131 ;
  assign n45142 = ~n45140 & n45141 ;
  assign n45144 = n45119 & n45143 ;
  assign n45145 = ~n45106 & n45144 ;
  assign n45152 = ~n45142 & ~n45145 ;
  assign n45153 = n45151 & n45152 ;
  assign n45154 = ~n45130 & n45153 ;
  assign n45161 = ~n45154 & ~n45160 ;
  assign n45166 = n45121 & ~n45137 ;
  assign n45167 = ~n45129 & n45166 ;
  assign n45168 = ~n45149 & ~n45167 ;
  assign n45169 = ~n45119 & ~n45168 ;
  assign n45162 = n45113 & ~n45137 ;
  assign n45163 = ~n45119 & n45162 ;
  assign n45164 = ~n45144 & ~n45163 ;
  assign n45165 = n45129 & ~n45164 ;
  assign n45171 = ~n45112 & ~n45137 ;
  assign n45172 = n45170 & n45171 ;
  assign n45173 = ~n45106 & n45172 ;
  assign n45191 = ~n45165 & ~n45173 ;
  assign n45192 = ~n45169 & n45191 ;
  assign n45193 = ~n45161 & n45192 ;
  assign n45194 = ~n45190 & n45193 ;
  assign n45195 = \u1_L2_reg[11]/NET0131  & ~n45194 ;
  assign n45196 = ~\u1_L2_reg[11]/NET0131  & n45194 ;
  assign n45197 = ~n45195 & ~n45196 ;
  assign n45210 = decrypt_pad & ~\u1_uk_K_r2_reg[33]/NET0131  ;
  assign n45211 = ~decrypt_pad & ~\u1_uk_K_r2_reg[13]/NET0131  ;
  assign n45212 = ~n45210 & ~n45211 ;
  assign n45213 = \u1_R2_reg[13]/NET0131  & ~n45212 ;
  assign n45214 = ~\u1_R2_reg[13]/NET0131  & n45212 ;
  assign n45215 = ~n45213 & ~n45214 ;
  assign n45204 = decrypt_pad & ~\u1_uk_K_r2_reg[39]/NET0131  ;
  assign n45205 = ~decrypt_pad & ~\u1_uk_K_r2_reg[19]/NET0131  ;
  assign n45206 = ~n45204 & ~n45205 ;
  assign n45207 = \u1_R2_reg[12]/NET0131  & ~n45206 ;
  assign n45208 = ~\u1_R2_reg[12]/NET0131  & n45206 ;
  assign n45209 = ~n45207 & ~n45208 ;
  assign n45223 = decrypt_pad & ~\u1_uk_K_r2_reg[55]/NET0131  ;
  assign n45224 = ~decrypt_pad & ~\u1_uk_K_r2_reg[3]/NET0131  ;
  assign n45225 = ~n45223 & ~n45224 ;
  assign n45226 = \u1_R2_reg[17]/NET0131  & ~n45225 ;
  assign n45227 = ~\u1_R2_reg[17]/NET0131  & n45225 ;
  assign n45228 = ~n45226 & ~n45227 ;
  assign n45255 = n45209 & n45228 ;
  assign n45256 = n45215 & n45255 ;
  assign n45198 = decrypt_pad & ~\u1_uk_K_r2_reg[10]/NET0131  ;
  assign n45199 = ~decrypt_pad & ~\u1_uk_K_r2_reg[47]/NET0131  ;
  assign n45200 = ~n45198 & ~n45199 ;
  assign n45201 = \u1_R2_reg[15]/NET0131  & ~n45200 ;
  assign n45202 = ~\u1_R2_reg[15]/NET0131  & n45200 ;
  assign n45203 = ~n45201 & ~n45202 ;
  assign n45253 = ~n45215 & ~n45228 ;
  assign n45254 = ~n45209 & n45253 ;
  assign n45257 = n45203 & ~n45254 ;
  assign n45258 = ~n45256 & n45257 ;
  assign n45217 = decrypt_pad & ~\u1_uk_K_r2_reg[34]/NET0131  ;
  assign n45218 = ~decrypt_pad & ~\u1_uk_K_r2_reg[39]/NET0131  ;
  assign n45219 = ~n45217 & ~n45218 ;
  assign n45220 = \u1_R2_reg[14]/NET0131  & ~n45219 ;
  assign n45221 = ~\u1_R2_reg[14]/NET0131  & n45219 ;
  assign n45222 = ~n45220 & ~n45221 ;
  assign n45235 = n45209 & ~n45228 ;
  assign n45259 = n45222 & n45235 ;
  assign n45260 = ~n45215 & n45228 ;
  assign n45261 = ~n45203 & ~n45260 ;
  assign n45262 = ~n45259 & n45261 ;
  assign n45263 = ~n45258 & ~n45262 ;
  assign n45232 = ~n45222 & ~n45228 ;
  assign n45233 = ~n45209 & n45232 ;
  assign n45234 = ~n45215 & n45233 ;
  assign n45216 = ~n45209 & n45215 ;
  assign n45244 = n45216 & ~n45228 ;
  assign n45245 = n45222 & n45244 ;
  assign n45246 = ~n45234 & ~n45245 ;
  assign n45266 = n45209 & ~n45222 ;
  assign n45267 = ~n45215 & n45266 ;
  assign n45268 = n45228 & n45267 ;
  assign n45247 = decrypt_pad & ~\u1_uk_K_r2_reg[18]/NET0131  ;
  assign n45248 = ~decrypt_pad & ~\u1_uk_K_r2_reg[55]/NET0131  ;
  assign n45249 = ~n45247 & ~n45248 ;
  assign n45250 = \u1_R2_reg[16]/NET0131  & ~n45249 ;
  assign n45251 = ~\u1_R2_reg[16]/NET0131  & n45249 ;
  assign n45252 = ~n45250 & ~n45251 ;
  assign n45241 = n45203 & n45215 ;
  assign n45264 = n45222 & n45241 ;
  assign n45265 = ~n45209 & n45264 ;
  assign n45269 = ~n45252 & ~n45265 ;
  assign n45270 = ~n45268 & n45269 ;
  assign n45271 = n45246 & n45270 ;
  assign n45272 = ~n45263 & n45271 ;
  assign n45273 = ~n45203 & n45254 ;
  assign n45274 = ~n45256 & ~n45273 ;
  assign n45275 = n45222 & ~n45274 ;
  assign n45276 = ~n45203 & ~n45222 ;
  assign n45277 = n45209 & ~n45215 ;
  assign n45278 = ~n45216 & ~n45277 ;
  assign n45279 = n45276 & ~n45278 ;
  assign n45284 = n45252 & ~n45279 ;
  assign n45229 = ~n45222 & n45228 ;
  assign n45230 = n45216 & n45229 ;
  assign n45242 = n45235 & n45241 ;
  assign n45280 = ~n45230 & ~n45242 ;
  assign n45281 = ~n45209 & n45228 ;
  assign n45282 = n45203 & n45281 ;
  assign n45283 = ~n45215 & n45282 ;
  assign n45285 = n45280 & ~n45283 ;
  assign n45286 = n45284 & n45285 ;
  assign n45287 = ~n45275 & n45286 ;
  assign n45288 = ~n45272 & ~n45287 ;
  assign n45231 = ~n45203 & ~n45230 ;
  assign n45236 = ~n45215 & n45222 ;
  assign n45237 = n45235 & n45236 ;
  assign n45238 = n45203 & ~n45237 ;
  assign n45239 = ~n45234 & n45238 ;
  assign n45240 = ~n45231 & ~n45239 ;
  assign n45243 = ~n45222 & n45242 ;
  assign n45289 = ~n45240 & ~n45243 ;
  assign n45290 = ~n45288 & n45289 ;
  assign n45291 = ~\u1_L2_reg[20]/NET0131  & ~n45290 ;
  assign n45292 = \u1_L2_reg[20]/NET0131  & n45290 ;
  assign n45293 = ~n45291 & ~n45292 ;
  assign n45294 = decrypt_pad & ~\u1_uk_K_r2_reg[42]/NET0131  ;
  assign n45295 = ~decrypt_pad & ~\u1_uk_K_r2_reg[51]/NET0131  ;
  assign n45296 = ~n45294 & ~n45295 ;
  assign n45297 = \u1_R2_reg[32]/NET0131  & ~n45296 ;
  assign n45298 = ~\u1_R2_reg[32]/NET0131  & n45296 ;
  assign n45299 = ~n45297 & ~n45298 ;
  assign n45325 = decrypt_pad & ~\u1_uk_K_r2_reg[52]/NET0131  ;
  assign n45326 = ~decrypt_pad & ~\u1_uk_K_r2_reg[2]/NET0131  ;
  assign n45327 = ~n45325 & ~n45326 ;
  assign n45328 = \u1_R2_reg[30]/NET0131  & ~n45327 ;
  assign n45329 = ~\u1_R2_reg[30]/NET0131  & n45327 ;
  assign n45330 = ~n45328 & ~n45329 ;
  assign n45318 = decrypt_pad & ~\u1_uk_K_r2_reg[51]/NET0131  ;
  assign n45319 = ~decrypt_pad & ~\u1_uk_K_r2_reg[29]/NET0131  ;
  assign n45320 = ~n45318 & ~n45319 ;
  assign n45321 = \u1_R2_reg[28]/NET0131  & ~n45320 ;
  assign n45322 = ~\u1_R2_reg[28]/NET0131  & n45320 ;
  assign n45323 = ~n45321 & ~n45322 ;
  assign n45306 = decrypt_pad & ~\u1_uk_K_r2_reg[8]/NET0131  ;
  assign n45307 = ~decrypt_pad & ~\u1_uk_K_r2_reg[45]/NET0131  ;
  assign n45308 = ~n45306 & ~n45307 ;
  assign n45309 = \u1_R2_reg[1]/NET0131  & ~n45308 ;
  assign n45310 = ~\u1_R2_reg[1]/NET0131  & n45308 ;
  assign n45311 = ~n45309 & ~n45310 ;
  assign n45312 = decrypt_pad & ~\u1_uk_K_r2_reg[23]/NET0131  ;
  assign n45313 = ~decrypt_pad & ~\u1_uk_K_r2_reg[1]/NET0131  ;
  assign n45314 = ~n45312 & ~n45313 ;
  assign n45315 = \u1_R2_reg[29]/NET0131  & ~n45314 ;
  assign n45316 = ~\u1_R2_reg[29]/NET0131  & n45314 ;
  assign n45317 = ~n45315 & ~n45316 ;
  assign n45337 = n45311 & n45317 ;
  assign n45366 = ~n45323 & n45337 ;
  assign n45367 = n45330 & n45366 ;
  assign n45360 = ~n45317 & ~n45330 ;
  assign n45361 = ~n45323 & n45360 ;
  assign n45300 = decrypt_pad & ~\u1_uk_K_r2_reg[36]/NET0131  ;
  assign n45301 = ~decrypt_pad & ~\u1_uk_K_r2_reg[14]/NET0131  ;
  assign n45302 = ~n45300 & ~n45301 ;
  assign n45303 = \u1_R2_reg[31]/P0001  & ~n45302 ;
  assign n45304 = ~\u1_R2_reg[31]/P0001  & n45302 ;
  assign n45305 = ~n45303 & ~n45304 ;
  assign n45324 = ~n45317 & n45323 ;
  assign n45331 = n45324 & n45330 ;
  assign n45368 = ~n45305 & ~n45331 ;
  assign n45369 = ~n45361 & n45368 ;
  assign n45343 = n45323 & ~n45330 ;
  assign n45370 = ~n45311 & n45317 ;
  assign n45372 = ~n45343 & n45370 ;
  assign n45371 = n45343 & ~n45370 ;
  assign n45373 = n45305 & ~n45371 ;
  assign n45374 = ~n45372 & n45373 ;
  assign n45375 = ~n45369 & ~n45374 ;
  assign n45376 = ~n45367 & ~n45375 ;
  assign n45377 = n45299 & ~n45376 ;
  assign n45332 = ~n45311 & n45331 ;
  assign n45333 = n45311 & ~n45323 ;
  assign n45334 = ~n45317 & n45333 ;
  assign n45335 = n45305 & ~n45334 ;
  assign n45336 = ~n45332 & n45335 ;
  assign n45338 = ~n45311 & ~n45323 ;
  assign n45339 = n45330 & n45338 ;
  assign n45340 = ~n45305 & ~n45337 ;
  assign n45341 = ~n45339 & n45340 ;
  assign n45342 = ~n45336 & ~n45341 ;
  assign n45344 = ~n45305 & n45343 ;
  assign n45347 = ~n45311 & ~n45343 ;
  assign n45345 = n45323 & n45330 ;
  assign n45346 = n45311 & ~n45345 ;
  assign n45348 = n45317 & ~n45346 ;
  assign n45349 = ~n45347 & n45348 ;
  assign n45350 = ~n45344 & ~n45349 ;
  assign n45351 = ~n45342 & n45350 ;
  assign n45352 = ~n45299 & ~n45351 ;
  assign n45354 = n45317 & ~n45330 ;
  assign n45355 = n45317 & ~n45323 ;
  assign n45356 = ~n45311 & ~n45355 ;
  assign n45357 = ~n45354 & ~n45356 ;
  assign n45358 = n45311 & ~n45343 ;
  assign n45359 = n45357 & ~n45358 ;
  assign n45353 = n45330 & n45334 ;
  assign n45362 = ~n45311 & n45361 ;
  assign n45363 = ~n45353 & ~n45362 ;
  assign n45364 = ~n45359 & n45363 ;
  assign n45365 = n45305 & ~n45364 ;
  assign n45378 = n45344 & n45370 ;
  assign n45379 = ~n45365 & ~n45378 ;
  assign n45380 = ~n45352 & n45379 ;
  assign n45381 = ~n45377 & n45380 ;
  assign n45382 = \u1_L2_reg[5]/NET0131  & ~n45381 ;
  assign n45383 = ~\u1_L2_reg[5]/NET0131  & n45381 ;
  assign n45384 = ~n45382 & ~n45383 ;
  assign n45396 = n45203 & ~n45268 ;
  assign n45397 = ~n45244 & n45396 ;
  assign n45398 = n45215 & ~n45222 ;
  assign n45399 = n45235 & ~n45398 ;
  assign n45400 = n45231 & ~n45399 ;
  assign n45401 = ~n45397 & ~n45400 ;
  assign n45402 = n45222 & n45256 ;
  assign n45403 = ~n45209 & n45236 ;
  assign n45404 = n45228 & n45403 ;
  assign n45405 = ~n45402 & ~n45404 ;
  assign n45406 = ~n45401 & n45405 ;
  assign n45407 = n45252 & ~n45406 ;
  assign n45385 = n45215 & n45266 ;
  assign n45386 = n45255 & n45276 ;
  assign n45390 = ~n45385 & ~n45386 ;
  assign n45391 = ~n45273 & n45390 ;
  assign n45387 = n45203 & ~n45229 ;
  assign n45388 = n45277 & n45387 ;
  assign n45389 = ~n45222 & n45282 ;
  assign n45392 = ~n45388 & ~n45389 ;
  assign n45393 = n45391 & n45392 ;
  assign n45394 = n45246 & n45393 ;
  assign n45395 = ~n45252 & ~n45394 ;
  assign n45408 = ~n45234 & n45405 ;
  assign n45409 = ~n45203 & ~n45408 ;
  assign n45410 = ~n45243 & ~n45265 ;
  assign n45411 = ~n45409 & n45410 ;
  assign n45412 = ~n45395 & n45411 ;
  assign n45413 = ~n45407 & n45412 ;
  assign n45414 = ~\u1_L2_reg[10]/NET0131  & ~n45413 ;
  assign n45415 = \u1_L2_reg[10]/NET0131  & n45413 ;
  assign n45416 = ~n45414 & ~n45415 ;
  assign n45423 = ~n44962 & ~n44964 ;
  assign n45424 = n44973 & n45423 ;
  assign n45421 = ~n44959 & ~n44964 ;
  assign n45422 = n44975 & ~n45421 ;
  assign n45428 = ~n44921 & ~n45422 ;
  assign n45429 = ~n45424 & n45428 ;
  assign n45417 = n44946 & n44965 ;
  assign n45418 = n44939 & n44957 ;
  assign n45419 = ~n45417 & ~n45418 ;
  assign n45420 = ~n44933 & ~n45419 ;
  assign n45425 = ~n44940 & ~n44980 ;
  assign n45426 = ~n44957 & n45425 ;
  assign n45427 = ~n44954 & ~n45426 ;
  assign n45430 = ~n45420 & ~n45427 ;
  assign n45431 = n45429 & n45430 ;
  assign n45432 = ~n44954 & n44977 ;
  assign n45438 = n44921 & ~n44979 ;
  assign n45439 = ~n44994 & n45438 ;
  assign n45440 = ~n45432 & n45439 ;
  assign n45433 = ~n44956 & ~n44997 ;
  assign n45434 = n44985 & ~n45433 ;
  assign n45435 = n44933 & n44946 ;
  assign n45436 = ~n44974 & ~n45435 ;
  assign n45437 = n44954 & ~n45436 ;
  assign n45441 = ~n45434 & ~n45437 ;
  assign n45442 = n45440 & n45441 ;
  assign n45443 = ~n45431 & ~n45442 ;
  assign n45444 = \u1_L2_reg[12]/NET0131  & n45443 ;
  assign n45445 = ~\u1_L2_reg[12]/NET0131  & ~n45443 ;
  assign n45446 = ~n45444 & ~n45445 ;
  assign n45447 = decrypt_pad & ~\u1_uk_K_r2_reg[31]/NET0131  ;
  assign n45448 = ~decrypt_pad & ~\u1_uk_K_r2_reg[36]/NET0131  ;
  assign n45449 = ~n45447 & ~n45448 ;
  assign n45450 = \u1_R2_reg[20]/NET0131  & ~n45449 ;
  assign n45451 = ~\u1_R2_reg[20]/NET0131  & n45449 ;
  assign n45452 = ~n45450 & ~n45451 ;
  assign n45489 = decrypt_pad & ~\u1_uk_K_r2_reg[43]/NET0131  ;
  assign n45490 = ~decrypt_pad & ~\u1_uk_K_r2_reg[21]/NET0131  ;
  assign n45491 = ~n45489 & ~n45490 ;
  assign n45492 = \u1_R2_reg[19]/NET0131  & ~n45491 ;
  assign n45493 = ~\u1_R2_reg[19]/NET0131  & n45491 ;
  assign n45494 = ~n45492 & ~n45493 ;
  assign n45466 = decrypt_pad & ~\u1_uk_K_r2_reg[1]/NET0131  ;
  assign n45467 = ~decrypt_pad & ~\u1_uk_K_r2_reg[38]/NET0131  ;
  assign n45468 = ~n45466 & ~n45467 ;
  assign n45469 = \u1_R2_reg[18]/NET0131  & ~n45468 ;
  assign n45470 = ~\u1_R2_reg[18]/NET0131  & n45468 ;
  assign n45471 = ~n45469 & ~n45470 ;
  assign n45453 = decrypt_pad & ~\u1_uk_K_r2_reg[16]/NET0131  ;
  assign n45454 = ~decrypt_pad & ~\u1_uk_K_r2_reg[49]/NET0131  ;
  assign n45455 = ~n45453 & ~n45454 ;
  assign n45456 = \u1_R2_reg[16]/NET0131  & ~n45455 ;
  assign n45457 = ~\u1_R2_reg[16]/NET0131  & n45455 ;
  assign n45458 = ~n45456 & ~n45457 ;
  assign n45459 = decrypt_pad & ~\u1_uk_K_r2_reg[28]/NET0131  ;
  assign n45460 = ~decrypt_pad & ~\u1_uk_K_r2_reg[37]/NET0131  ;
  assign n45461 = ~n45459 & ~n45460 ;
  assign n45462 = \u1_R2_reg[21]/NET0131  & ~n45461 ;
  assign n45463 = ~\u1_R2_reg[21]/NET0131  & n45461 ;
  assign n45464 = ~n45462 & ~n45463 ;
  assign n45465 = n45458 & ~n45464 ;
  assign n45472 = decrypt_pad & ~\u1_uk_K_r2_reg[7]/NET0131  ;
  assign n45473 = ~decrypt_pad & ~\u1_uk_K_r2_reg[16]/NET0131  ;
  assign n45474 = ~n45472 & ~n45473 ;
  assign n45475 = \u1_R2_reg[17]/NET0131  & ~n45474 ;
  assign n45476 = ~\u1_R2_reg[17]/NET0131  & n45474 ;
  assign n45477 = ~n45475 & ~n45476 ;
  assign n45526 = n45465 & ~n45477 ;
  assign n45527 = ~n45471 & n45526 ;
  assign n45478 = ~n45471 & n45477 ;
  assign n45496 = n45458 & n45464 ;
  assign n45528 = n45478 & n45496 ;
  assign n45510 = ~n45458 & n45464 ;
  assign n45511 = ~n45477 & n45510 ;
  assign n45486 = ~n45464 & n45477 ;
  assign n45525 = n45471 & n45486 ;
  assign n45529 = ~n45511 & ~n45525 ;
  assign n45530 = ~n45528 & n45529 ;
  assign n45531 = ~n45527 & n45530 ;
  assign n45532 = ~n45494 & ~n45531 ;
  assign n45482 = ~n45458 & n45478 ;
  assign n45483 = n45458 & n45471 ;
  assign n45484 = n45464 & ~n45483 ;
  assign n45521 = ~n45465 & ~n45486 ;
  assign n45522 = ~n45484 & n45521 ;
  assign n45523 = ~n45482 & ~n45522 ;
  assign n45524 = n45494 & ~n45523 ;
  assign n45533 = n45464 & ~n45471 ;
  assign n45534 = ~n45465 & ~n45533 ;
  assign n45504 = ~n45458 & ~n45477 ;
  assign n45535 = n45471 & n45477 ;
  assign n45536 = ~n45504 & ~n45535 ;
  assign n45537 = n45534 & n45536 ;
  assign n45538 = ~n45524 & ~n45537 ;
  assign n45539 = ~n45532 & n45538 ;
  assign n45540 = ~n45452 & ~n45539 ;
  assign n45485 = ~n45482 & n45484 ;
  assign n45487 = n45458 & n45486 ;
  assign n45488 = ~n45485 & ~n45487 ;
  assign n45495 = ~n45488 & n45494 ;
  assign n45479 = n45471 & ~n45477 ;
  assign n45480 = ~n45478 & ~n45479 ;
  assign n45481 = n45465 & ~n45480 ;
  assign n45497 = n45471 & n45494 ;
  assign n45498 = n45496 & ~n45497 ;
  assign n45499 = n45480 & n45498 ;
  assign n45500 = ~n45481 & ~n45499 ;
  assign n45501 = ~n45495 & n45500 ;
  assign n45502 = n45452 & ~n45501 ;
  assign n45505 = ~n45464 & n45504 ;
  assign n45506 = n45471 & n45505 ;
  assign n45503 = ~n45471 & n45487 ;
  assign n45507 = n45494 & ~n45503 ;
  assign n45508 = ~n45506 & n45507 ;
  assign n45514 = n45477 & n45510 ;
  assign n45515 = ~n45505 & ~n45514 ;
  assign n45516 = n45452 & ~n45471 ;
  assign n45517 = ~n45515 & n45516 ;
  assign n45509 = ~n45458 & n45486 ;
  assign n45512 = ~n45509 & ~n45511 ;
  assign n45513 = n45471 & ~n45512 ;
  assign n45518 = ~n45494 & ~n45513 ;
  assign n45519 = ~n45517 & n45518 ;
  assign n45520 = ~n45508 & ~n45519 ;
  assign n45541 = ~n45502 & ~n45520 ;
  assign n45542 = ~n45540 & n45541 ;
  assign n45543 = ~\u1_L2_reg[14]/NET0131  & ~n45542 ;
  assign n45544 = \u1_L2_reg[14]/NET0131  & n45542 ;
  assign n45545 = ~n45543 & ~n45544 ;
  assign n45551 = ~n45041 & ~n45047 ;
  assign n45552 = ~n45032 & n45057 ;
  assign n45553 = ~n45551 & ~n45552 ;
  assign n45554 = ~n45025 & ~n45553 ;
  assign n45546 = ~n45052 & ~n45056 ;
  assign n45547 = n45025 & n45546 ;
  assign n45548 = n45019 & n45052 ;
  assign n45549 = ~n45547 & ~n45548 ;
  assign n45550 = n45038 & ~n45549 ;
  assign n45555 = ~n45013 & ~n45087 ;
  assign n45556 = ~n45550 & n45555 ;
  assign n45557 = ~n45554 & n45556 ;
  assign n45558 = ~n45066 & ~n45070 ;
  assign n45561 = n45056 & n45084 ;
  assign n45562 = n45558 & ~n45561 ;
  assign n45563 = n45025 & ~n45562 ;
  assign n45564 = n45038 & n45091 ;
  assign n45559 = ~n45025 & ~n45084 ;
  assign n45560 = n45558 & n45559 ;
  assign n45565 = n45013 & ~n45089 ;
  assign n45566 = ~n45560 & n45565 ;
  assign n45567 = ~n45564 & n45566 ;
  assign n45568 = ~n45563 & n45567 ;
  assign n45569 = ~n45557 & ~n45568 ;
  assign n45571 = n45047 & ~n45075 ;
  assign n45570 = n45025 & ~n45038 ;
  assign n45572 = ~n45088 & n45570 ;
  assign n45573 = n45571 & n45572 ;
  assign n45574 = ~n45569 & ~n45573 ;
  assign n45575 = ~\u1_L2_reg[17]/NET0131  & ~n45574 ;
  assign n45576 = \u1_L2_reg[17]/NET0131  & n45574 ;
  assign n45577 = ~n45575 & ~n45576 ;
  assign n45598 = ~n45260 & ~n45267 ;
  assign n45599 = n45252 & ~n45598 ;
  assign n45600 = ~n45245 & n45405 ;
  assign n45601 = ~n45599 & n45600 ;
  assign n45602 = n45203 & ~n45601 ;
  assign n45578 = ~n45232 & ~n45260 ;
  assign n45579 = n45209 & ~n45578 ;
  assign n45580 = ~n45203 & ~n45579 ;
  assign n45581 = ~n45233 & n45238 ;
  assign n45582 = ~n45580 & ~n45581 ;
  assign n45583 = ~n45235 & ~n45281 ;
  assign n45584 = n45398 & ~n45583 ;
  assign n45585 = ~n45402 & ~n45584 ;
  assign n45586 = ~n45582 & n45585 ;
  assign n45587 = ~n45252 & ~n45586 ;
  assign n45588 = ~n45235 & n45398 ;
  assign n45589 = n45215 & n45281 ;
  assign n45590 = ~n45588 & ~n45589 ;
  assign n45591 = ~n45203 & ~n45590 ;
  assign n45592 = n45215 & n45259 ;
  assign n45593 = ~n45403 & ~n45592 ;
  assign n45594 = ~n45591 & n45593 ;
  assign n45595 = n45252 & ~n45594 ;
  assign n45596 = ~n45203 & ~n45228 ;
  assign n45597 = ~n45593 & n45596 ;
  assign n45603 = ~n45595 & ~n45597 ;
  assign n45604 = ~n45587 & n45603 ;
  assign n45605 = ~n45602 & n45604 ;
  assign n45606 = ~\u1_L2_reg[1]/NET0131  & ~n45605 ;
  assign n45607 = \u1_L2_reg[1]/NET0131  & n45605 ;
  assign n45608 = ~n45606 & ~n45607 ;
  assign n45620 = ~n45317 & n45330 ;
  assign n45621 = ~n45305 & n45311 ;
  assign n45622 = n45620 & n45621 ;
  assign n45628 = n45299 & ~n45622 ;
  assign n45624 = n45317 & n45323 ;
  assign n45625 = ~n45330 & n45624 ;
  assign n45626 = n45305 & ~n45317 ;
  assign n45627 = n45338 & n45626 ;
  assign n45629 = ~n45625 & ~n45627 ;
  assign n45630 = n45628 & n45629 ;
  assign n45610 = n45317 & n45339 ;
  assign n45623 = n45311 & n45331 ;
  assign n45631 = ~n45610 & ~n45623 ;
  assign n45632 = n45630 & n45631 ;
  assign n45633 = ~n45330 & n45370 ;
  assign n45634 = ~n45334 & ~n45624 ;
  assign n45635 = ~n45633 & n45634 ;
  assign n45636 = n45305 & ~n45635 ;
  assign n45637 = ~n45311 & n45343 ;
  assign n45638 = ~n45317 & n45637 ;
  assign n45639 = ~n45299 & ~n45638 ;
  assign n45640 = ~n45636 & n45639 ;
  assign n45641 = ~n45632 & ~n45640 ;
  assign n45609 = n45333 & n45354 ;
  assign n45611 = ~n45362 & ~n45609 ;
  assign n45612 = n45368 & ~n45610 ;
  assign n45613 = n45611 & n45612 ;
  assign n45614 = ~n45330 & n45334 ;
  assign n45615 = n45305 & ~n45367 ;
  assign n45616 = ~n45614 & n45615 ;
  assign n45617 = ~n45613 & ~n45616 ;
  assign n45618 = ~n45299 & ~n45305 ;
  assign n45619 = n45324 & n45618 ;
  assign n45642 = ~n45617 & ~n45619 ;
  assign n45643 = ~n45641 & n45642 ;
  assign n45644 = \u1_L2_reg[15]/P0001  & n45643 ;
  assign n45645 = ~\u1_L2_reg[15]/P0001  & ~n45643 ;
  assign n45646 = ~n45644 & ~n45645 ;
  assign n45651 = n45305 & ~n45366 ;
  assign n45649 = n45330 & n45624 ;
  assign n45650 = n45311 & n45360 ;
  assign n45652 = ~n45649 & ~n45650 ;
  assign n45653 = n45651 & n45652 ;
  assign n45654 = ~n45305 & ~n45637 ;
  assign n45655 = ~n45623 & n45654 ;
  assign n45656 = ~n45653 & ~n45655 ;
  assign n45657 = ~n45324 & n45330 ;
  assign n45658 = n45356 & n45657 ;
  assign n45659 = n45299 & ~n45614 ;
  assign n45660 = ~n45658 & n45659 ;
  assign n45661 = ~n45656 & n45660 ;
  assign n45662 = n45305 & ~n45311 ;
  assign n45663 = ~n45333 & ~n45662 ;
  assign n45664 = ~n45330 & ~n45663 ;
  assign n45665 = ~n45345 & ~n45626 ;
  assign n45666 = ~n45356 & n45665 ;
  assign n45667 = ~n45664 & n45666 ;
  assign n45671 = ~n45299 & ~n45332 ;
  assign n45668 = n45323 & ~n45337 ;
  assign n45669 = n45305 & ~n45360 ;
  assign n45670 = n45668 & n45669 ;
  assign n45672 = ~n45362 & ~n45670 ;
  assign n45673 = n45671 & n45672 ;
  assign n45674 = ~n45667 & n45673 ;
  assign n45675 = ~n45661 & ~n45674 ;
  assign n45647 = n45305 & n45361 ;
  assign n45648 = n45621 & n45625 ;
  assign n45676 = ~n45647 & ~n45648 ;
  assign n45677 = ~n45675 & n45676 ;
  assign n45678 = ~\u1_L2_reg[21]/NET0131  & ~n45677 ;
  assign n45679 = \u1_L2_reg[21]/NET0131  & n45677 ;
  assign n45680 = ~n45678 & ~n45679 ;
  assign n45693 = ~n45464 & ~n45478 ;
  assign n45694 = ~n45483 & n45693 ;
  assign n45692 = n45477 & n45496 ;
  assign n45695 = ~n45504 & ~n45692 ;
  assign n45696 = ~n45694 & n45695 ;
  assign n45697 = n45494 & ~n45696 ;
  assign n45699 = ~n45477 & n45496 ;
  assign n45700 = ~n45482 & ~n45699 ;
  assign n45701 = ~n45494 & ~n45700 ;
  assign n45698 = n45477 & n45533 ;
  assign n45702 = n45483 & n45486 ;
  assign n45703 = ~n45698 & ~n45702 ;
  assign n45704 = ~n45701 & n45703 ;
  assign n45705 = ~n45697 & n45704 ;
  assign n45706 = n45452 & ~n45705 ;
  assign n45686 = ~n45486 & n45494 ;
  assign n45685 = ~n45494 & ~n45504 ;
  assign n45687 = ~n45471 & ~n45685 ;
  assign n45688 = ~n45686 & n45687 ;
  assign n45681 = n45471 & n45514 ;
  assign n45682 = ~n45458 & n45535 ;
  assign n45683 = ~n45526 & ~n45682 ;
  assign n45684 = ~n45494 & ~n45683 ;
  assign n45689 = ~n45681 & ~n45684 ;
  assign n45690 = ~n45688 & n45689 ;
  assign n45691 = ~n45452 & ~n45690 ;
  assign n45709 = ~n45506 & ~n45702 ;
  assign n45710 = ~n45471 & n45510 ;
  assign n45711 = ~n45477 & n45710 ;
  assign n45712 = n45709 & ~n45711 ;
  assign n45713 = n45494 & ~n45712 ;
  assign n45707 = n45458 & ~n45494 ;
  assign n45708 = n45479 & n45707 ;
  assign n45714 = ~n45528 & ~n45708 ;
  assign n45715 = ~n45713 & n45714 ;
  assign n45716 = ~n45691 & n45715 ;
  assign n45717 = ~n45706 & n45716 ;
  assign n45718 = ~\u1_L2_reg[25]/NET0131  & ~n45717 ;
  assign n45719 = \u1_L2_reg[25]/NET0131  & n45717 ;
  assign n45720 = ~n45718 & ~n45719 ;
  assign n45721 = ~n45230 & n45396 ;
  assign n45722 = ~n45228 & ~n45278 ;
  assign n45723 = ~n45256 & ~n45722 ;
  assign n45724 = ~n45222 & ~n45723 ;
  assign n45725 = ~n45253 & ~n45403 ;
  assign n45726 = ~n45252 & ~n45725 ;
  assign n45727 = ~n45203 & ~n45726 ;
  assign n45728 = ~n45724 & n45727 ;
  assign n45729 = ~n45721 & ~n45728 ;
  assign n45738 = n45252 & ~n45592 ;
  assign n45734 = n45203 & n45254 ;
  assign n45737 = ~n45222 & n45244 ;
  assign n45739 = ~n45734 & ~n45737 ;
  assign n45740 = n45738 & n45739 ;
  assign n45730 = ~n45215 & n45229 ;
  assign n45731 = ~n45255 & ~n45730 ;
  assign n45732 = ~n45203 & ~n45266 ;
  assign n45733 = ~n45731 & n45732 ;
  assign n45735 = ~n45282 & ~n45589 ;
  assign n45736 = n45222 & ~n45735 ;
  assign n45741 = ~n45733 & ~n45736 ;
  assign n45742 = n45740 & n45741 ;
  assign n45743 = n45264 & ~n45281 ;
  assign n45744 = ~n45252 & ~n45267 ;
  assign n45745 = n45280 & n45744 ;
  assign n45746 = ~n45743 & n45745 ;
  assign n45747 = ~n45742 & ~n45746 ;
  assign n45748 = ~n45729 & ~n45747 ;
  assign n45749 = ~\u1_L2_reg[26]/NET0131  & ~n45748 ;
  assign n45750 = \u1_L2_reg[26]/NET0131  & n45748 ;
  assign n45751 = ~n45749 & ~n45750 ;
  assign n45757 = ~n45106 & n45137 ;
  assign n45758 = n45181 & ~n45757 ;
  assign n45759 = ~n45106 & ~n45119 ;
  assign n45760 = ~n45120 & ~n45759 ;
  assign n45761 = ~n45137 & ~n45760 ;
  assign n45762 = ~n45758 & ~n45761 ;
  assign n45763 = n45129 & ~n45762 ;
  assign n45752 = ~n45119 & ~n45176 ;
  assign n45753 = n45119 & ~n45137 ;
  assign n45754 = n45121 & n45753 ;
  assign n45755 = ~n45752 & ~n45754 ;
  assign n45756 = ~n45129 & ~n45755 ;
  assign n45764 = ~n45112 & n45757 ;
  assign n45765 = n45119 & n45764 ;
  assign n45766 = ~n45756 & ~n45765 ;
  assign n45767 = ~n45763 & n45766 ;
  assign n45768 = ~n45160 & ~n45767 ;
  assign n45773 = n45113 & ~n45753 ;
  assign n45774 = ~n45754 & ~n45773 ;
  assign n45775 = n45129 & ~n45774 ;
  assign n45777 = n45119 & ~n45143 ;
  assign n45778 = ~n45171 & n45777 ;
  assign n45776 = n45129 & ~n45182 ;
  assign n45779 = ~n45752 & ~n45776 ;
  assign n45780 = ~n45778 & n45779 ;
  assign n45781 = ~n45775 & ~n45780 ;
  assign n45782 = n45160 & ~n45781 ;
  assign n45769 = ~n45106 & n45112 ;
  assign n45770 = n45138 & n45769 ;
  assign n45771 = n45106 & n45137 ;
  assign n45772 = n45131 & n45771 ;
  assign n45783 = ~n45770 & ~n45772 ;
  assign n45784 = ~n45782 & n45783 ;
  assign n45785 = ~n45768 & n45784 ;
  assign n45786 = \u1_L2_reg[29]/NET0131  & ~n45785 ;
  assign n45787 = ~\u1_L2_reg[29]/NET0131  & n45785 ;
  assign n45788 = ~n45786 & ~n45787 ;
  assign n45789 = decrypt_pad & ~\u1_uk_K_r2_reg[17]/NET0131  ;
  assign n45790 = ~decrypt_pad & ~\u1_uk_K_r2_reg[54]/NET0131  ;
  assign n45791 = ~n45789 & ~n45790 ;
  assign n45792 = \u1_R2_reg[8]/NET0131  & ~n45791 ;
  assign n45793 = ~\u1_R2_reg[8]/NET0131  & n45791 ;
  assign n45794 = ~n45792 & ~n45793 ;
  assign n45795 = decrypt_pad & ~\u1_uk_K_r2_reg[26]/NET0131  ;
  assign n45796 = ~decrypt_pad & ~\u1_uk_K_r2_reg[6]/NET0131  ;
  assign n45797 = ~n45795 & ~n45796 ;
  assign n45798 = \u1_R2_reg[7]/NET0131  & ~n45797 ;
  assign n45799 = ~\u1_R2_reg[7]/NET0131  & n45797 ;
  assign n45800 = ~n45798 & ~n45799 ;
  assign n45814 = decrypt_pad & ~\u1_uk_K_r2_reg[41]/NET0131  ;
  assign n45815 = ~decrypt_pad & ~\u1_uk_K_r2_reg[46]/NET0131  ;
  assign n45816 = ~n45814 & ~n45815 ;
  assign n45817 = \u1_R2_reg[5]/NET0131  & ~n45816 ;
  assign n45818 = ~\u1_R2_reg[5]/NET0131  & n45816 ;
  assign n45819 = ~n45817 & ~n45818 ;
  assign n45801 = decrypt_pad & ~\u1_uk_K_r2_reg[5]/NET0131  ;
  assign n45802 = ~decrypt_pad & ~\u1_uk_K_r2_reg[10]/NET0131  ;
  assign n45803 = ~n45801 & ~n45802 ;
  assign n45804 = \u1_R2_reg[4]/NET0131  & ~n45803 ;
  assign n45805 = ~\u1_R2_reg[4]/NET0131  & n45803 ;
  assign n45806 = ~n45804 & ~n45805 ;
  assign n45807 = decrypt_pad & ~\u1_uk_K_r2_reg[54]/NET0131  ;
  assign n45808 = ~decrypt_pad & ~\u1_uk_K_r2_reg[34]/NET0131  ;
  assign n45809 = ~n45807 & ~n45808 ;
  assign n45810 = \u1_R2_reg[9]/NET0131  & ~n45809 ;
  assign n45811 = ~\u1_R2_reg[9]/NET0131  & n45809 ;
  assign n45812 = ~n45810 & ~n45811 ;
  assign n45829 = ~n45806 & n45812 ;
  assign n45830 = ~n45819 & n45829 ;
  assign n45821 = decrypt_pad & ~\u1_uk_K_r2_reg[32]/NET0131  ;
  assign n45822 = ~decrypt_pad & ~\u1_uk_K_r2_reg[12]/NET0131  ;
  assign n45823 = ~n45821 & ~n45822 ;
  assign n45824 = \u1_R2_reg[6]/NET0131  & ~n45823 ;
  assign n45825 = ~\u1_R2_reg[6]/NET0131  & n45823 ;
  assign n45826 = ~n45824 & ~n45825 ;
  assign n45831 = n45806 & n45819 ;
  assign n45832 = n45806 & ~n45812 ;
  assign n45833 = ~n45831 & ~n45832 ;
  assign n45834 = n45826 & ~n45833 ;
  assign n45835 = ~n45830 & ~n45834 ;
  assign n45836 = ~n45800 & ~n45835 ;
  assign n45837 = ~n45812 & n45819 ;
  assign n45838 = ~n45830 & ~n45837 ;
  assign n45839 = ~n45826 & ~n45838 ;
  assign n45813 = n45806 & n45812 ;
  assign n45820 = n45813 & ~n45819 ;
  assign n45827 = n45820 & n45826 ;
  assign n45828 = n45800 & n45827 ;
  assign n45840 = ~n45800 & ~n45819 ;
  assign n45841 = n45812 & ~n45826 ;
  assign n45842 = n45840 & n45841 ;
  assign n45843 = n45819 & n45826 ;
  assign n45844 = n45829 & n45843 ;
  assign n45845 = ~n45842 & ~n45844 ;
  assign n45846 = ~n45828 & n45845 ;
  assign n45847 = ~n45839 & n45846 ;
  assign n45848 = ~n45836 & n45847 ;
  assign n45849 = ~n45794 & ~n45848 ;
  assign n45866 = ~n45806 & ~n45812 ;
  assign n45867 = ~n45827 & ~n45866 ;
  assign n45868 = n45794 & ~n45867 ;
  assign n45859 = ~n45819 & n45826 ;
  assign n45869 = n45829 & ~n45859 ;
  assign n45870 = ~n45868 & ~n45869 ;
  assign n45861 = n45819 & ~n45826 ;
  assign n45871 = ~n45800 & ~n45861 ;
  assign n45872 = ~n45870 & n45871 ;
  assign n45850 = ~n45819 & n45832 ;
  assign n45851 = ~n45826 & n45850 ;
  assign n45852 = n45800 & n45819 ;
  assign n45853 = ~n45806 & n45826 ;
  assign n45854 = n45852 & ~n45853 ;
  assign n45855 = n45831 & n45841 ;
  assign n45856 = ~n45854 & ~n45855 ;
  assign n45857 = ~n45851 & n45856 ;
  assign n45858 = n45794 & ~n45857 ;
  assign n45862 = n45806 & ~n45861 ;
  assign n45860 = ~n45806 & ~n45859 ;
  assign n45863 = n45800 & ~n45829 ;
  assign n45864 = ~n45860 & n45863 ;
  assign n45865 = ~n45862 & n45864 ;
  assign n45873 = ~n45858 & ~n45865 ;
  assign n45874 = ~n45872 & n45873 ;
  assign n45875 = ~n45849 & n45874 ;
  assign n45876 = \u1_L2_reg[2]/NET0131  & n45875 ;
  assign n45877 = ~\u1_L2_reg[2]/NET0131  & ~n45875 ;
  assign n45878 = ~n45876 & ~n45877 ;
  assign n45892 = ~n45829 & ~n45832 ;
  assign n45901 = ~n45806 & ~n45826 ;
  assign n45902 = n45819 & ~n45901 ;
  assign n45903 = n45892 & n45902 ;
  assign n45904 = ~n45850 & ~n45903 ;
  assign n45905 = n45800 & ~n45904 ;
  assign n45883 = n45819 & n45829 ;
  assign n45884 = ~n45826 & n45866 ;
  assign n45885 = ~n45883 & ~n45884 ;
  assign n45900 = ~n45800 & ~n45885 ;
  assign n45897 = n45800 & n45806 ;
  assign n45898 = ~n45820 & ~n45897 ;
  assign n45899 = ~n45826 & ~n45898 ;
  assign n45906 = n45829 & n45859 ;
  assign n45907 = ~n45899 & ~n45906 ;
  assign n45908 = ~n45900 & n45907 ;
  assign n45909 = ~n45905 & n45908 ;
  assign n45910 = n45794 & ~n45909 ;
  assign n45879 = n45832 & n45843 ;
  assign n45880 = ~n45819 & n45853 ;
  assign n45881 = ~n45879 & ~n45880 ;
  assign n45882 = ~n45800 & ~n45881 ;
  assign n45886 = n45800 & n45885 ;
  assign n45887 = ~n45826 & n45832 ;
  assign n45888 = ~n45800 & ~n45831 ;
  assign n45889 = ~n45830 & n45888 ;
  assign n45890 = ~n45887 & n45889 ;
  assign n45891 = ~n45886 & ~n45890 ;
  assign n45893 = n45859 & n45892 ;
  assign n45894 = ~n45879 & ~n45893 ;
  assign n45895 = ~n45891 & n45894 ;
  assign n45896 = ~n45794 & ~n45895 ;
  assign n45911 = ~n45882 & ~n45896 ;
  assign n45912 = ~n45910 & n45911 ;
  assign n45913 = ~\u1_L2_reg[28]/NET0131  & ~n45912 ;
  assign n45914 = \u1_L2_reg[28]/NET0131  & n45912 ;
  assign n45915 = ~n45913 & ~n45914 ;
  assign n45918 = n45131 & n45143 ;
  assign n45916 = n45119 & n45771 ;
  assign n45919 = n45160 & ~n45916 ;
  assign n45920 = ~n45918 & n45919 ;
  assign n45917 = n45170 & ~n45181 ;
  assign n45921 = ~n45163 & ~n45917 ;
  assign n45922 = n45920 & n45921 ;
  assign n45924 = n45129 & ~n45166 ;
  assign n45923 = ~n45119 & n45148 ;
  assign n45925 = ~n45145 & ~n45923 ;
  assign n45926 = n45924 & n45925 ;
  assign n45927 = ~n45129 & ~n45162 ;
  assign n45928 = ~n45765 & n45927 ;
  assign n45929 = ~n45926 & ~n45928 ;
  assign n45930 = ~n45160 & ~n45186 ;
  assign n45931 = ~n45770 & n45930 ;
  assign n45932 = ~n45929 & n45931 ;
  assign n45933 = ~n45922 & ~n45932 ;
  assign n45935 = ~n45112 & ~n45180 ;
  assign n45936 = ~n45757 & n45935 ;
  assign n45937 = n45924 & ~n45936 ;
  assign n45934 = ~n45129 & ~n45758 ;
  assign n45938 = n45119 & ~n45934 ;
  assign n45939 = ~n45937 & n45938 ;
  assign n45940 = ~n45172 & ~n45939 ;
  assign n45941 = ~n45933 & n45940 ;
  assign n45942 = ~\u1_L2_reg[4]/NET0131  & ~n45941 ;
  assign n45943 = \u1_L2_reg[4]/NET0131  & n45941 ;
  assign n45944 = ~n45942 & ~n45943 ;
  assign n45946 = ~n45812 & ~n45819 ;
  assign n45947 = n45826 & n45946 ;
  assign n45948 = ~n45800 & ~n45820 ;
  assign n45949 = ~n45947 & n45948 ;
  assign n45951 = n45812 & n45853 ;
  assign n45950 = ~n45826 & n45946 ;
  assign n45952 = n45800 & ~n45950 ;
  assign n45953 = ~n45951 & n45952 ;
  assign n45954 = ~n45949 & ~n45953 ;
  assign n45945 = n45837 & n45901 ;
  assign n45955 = n45794 & ~n45945 ;
  assign n45956 = n45845 & n45955 ;
  assign n45957 = ~n45954 & n45956 ;
  assign n45960 = n45812 & ~n45840 ;
  assign n45961 = n45901 & n45960 ;
  assign n45958 = n45826 & ~n45837 ;
  assign n45959 = n45897 & n45958 ;
  assign n45962 = ~n45794 & ~n45959 ;
  assign n45963 = ~n45961 & n45962 ;
  assign n45964 = n45819 & n45866 ;
  assign n45965 = ~n45800 & ~n45906 ;
  assign n45966 = ~n45964 & n45965 ;
  assign n45967 = ~n45851 & n45966 ;
  assign n45968 = n45963 & n45967 ;
  assign n45969 = ~n45957 & ~n45968 ;
  assign n45970 = ~n45855 & ~n45879 ;
  assign n45971 = ~n45969 & n45970 ;
  assign n45972 = n45819 & ~n45887 ;
  assign n45973 = ~n45830 & ~n45850 ;
  assign n45974 = ~n45972 & n45973 ;
  assign n45975 = n45800 & ~n45974 ;
  assign n45976 = n45963 & n45975 ;
  assign n45977 = ~n45971 & ~n45976 ;
  assign n45978 = ~\u1_L2_reg[13]/NET0131  & ~n45977 ;
  assign n45979 = \u1_L2_reg[13]/NET0131  & n45977 ;
  assign n45980 = ~n45978 & ~n45979 ;
  assign n45983 = ~n45129 & n45936 ;
  assign n45981 = ~n45122 & n45129 ;
  assign n45982 = ~n45935 & n45981 ;
  assign n45984 = n45112 & n45916 ;
  assign n45985 = ~n45160 & ~n45984 ;
  assign n45986 = ~n45982 & n45985 ;
  assign n45987 = ~n45983 & n45986 ;
  assign n45988 = n45119 & n45936 ;
  assign n45993 = ~n45149 & n45160 ;
  assign n45994 = ~n45988 & n45993 ;
  assign n45989 = ~n45180 & ~n45764 ;
  assign n45990 = ~n45119 & ~n45989 ;
  assign n45991 = ~n45129 & ~n45769 ;
  assign n45992 = ~n45981 & ~n45991 ;
  assign n45995 = ~n45990 & ~n45992 ;
  assign n45996 = n45994 & n45995 ;
  assign n45997 = ~n45987 & ~n45996 ;
  assign n45998 = ~n45169 & ~n45187 ;
  assign n45999 = ~n45997 & n45998 ;
  assign n46000 = ~\u1_L2_reg[19]/NET0131  & ~n45999 ;
  assign n46001 = \u1_L2_reg[19]/NET0131  & n45999 ;
  assign n46002 = ~n46000 & ~n46001 ;
  assign n46024 = ~n45038 & ~n45546 ;
  assign n46025 = ~n45032 & n45059 ;
  assign n46026 = ~n46024 & ~n46025 ;
  assign n46027 = n45013 & ~n46026 ;
  assign n46023 = n45056 & n45057 ;
  assign n46028 = ~n45564 & ~n46023 ;
  assign n46029 = ~n46027 & n46028 ;
  assign n46030 = ~n45025 & ~n46029 ;
  assign n46003 = ~n45053 & ~n45058 ;
  assign n46004 = n45025 & ~n46003 ;
  assign n46005 = ~n45090 & ~n46004 ;
  assign n46006 = ~n45026 & ~n46005 ;
  assign n46007 = n45025 & ~n45084 ;
  assign n46008 = n45048 & n46007 ;
  assign n46009 = n45067 & n45083 ;
  assign n46010 = n45013 & ~n45561 ;
  assign n46011 = ~n46009 & n46010 ;
  assign n46012 = ~n46008 & n46011 ;
  assign n46018 = ~n45013 & ~n45076 ;
  assign n46019 = ~n45089 & n46018 ;
  assign n46013 = ~n45052 & ~n45088 ;
  assign n46014 = n45570 & ~n46013 ;
  assign n46015 = ~n45047 & ~n45088 ;
  assign n46016 = ~n45025 & n45038 ;
  assign n46017 = ~n46015 & n46016 ;
  assign n46020 = ~n46014 & ~n46017 ;
  assign n46021 = n46019 & n46020 ;
  assign n46022 = ~n46012 & ~n46021 ;
  assign n46031 = ~n46006 & ~n46022 ;
  assign n46032 = ~n46030 & n46031 ;
  assign n46033 = \u1_L2_reg[23]/NET0131  & ~n46032 ;
  assign n46034 = ~\u1_L2_reg[23]/NET0131  & n46032 ;
  assign n46035 = ~n46033 & ~n46034 ;
  assign n46036 = n45323 & n45370 ;
  assign n46037 = ~n45361 & ~n45366 ;
  assign n46038 = ~n46036 & n46037 ;
  assign n46039 = ~n45305 & ~n46038 ;
  assign n46040 = ~n45323 & ~n45633 ;
  assign n46041 = n45305 & ~n45668 ;
  assign n46042 = ~n46040 & n46041 ;
  assign n46043 = ~n45332 & ~n45650 ;
  assign n46044 = ~n45367 & n46043 ;
  assign n46045 = ~n46042 & n46044 ;
  assign n46046 = ~n46039 & n46045 ;
  assign n46047 = n45299 & ~n46046 ;
  assign n46048 = n45305 & ~n45633 ;
  assign n46049 = ~n45357 & n46048 ;
  assign n46050 = ~n45353 & ~n46049 ;
  assign n46051 = ~n45299 & ~n46050 ;
  assign n46054 = ~n45305 & n45359 ;
  assign n46052 = ~n45346 & n45618 ;
  assign n46053 = ~n45356 & n46052 ;
  assign n46055 = n45620 & n45662 ;
  assign n46056 = ~n45378 & ~n46055 ;
  assign n46057 = ~n46053 & n46056 ;
  assign n46058 = ~n46054 & n46057 ;
  assign n46059 = ~n46051 & n46058 ;
  assign n46060 = ~n46047 & n46059 ;
  assign n46061 = ~\u1_L2_reg[27]/NET0131  & ~n46060 ;
  assign n46062 = \u1_L2_reg[27]/NET0131  & n46060 ;
  assign n46063 = ~n46061 & ~n46062 ;
  assign n46069 = ~n44975 & ~n44996 ;
  assign n46071 = ~n44962 & n45425 ;
  assign n46072 = n46069 & ~n46071 ;
  assign n46070 = ~n44962 & ~n46069 ;
  assign n46073 = ~n44954 & ~n46070 ;
  assign n46074 = ~n46072 & n46073 ;
  assign n46064 = n44964 & n44996 ;
  assign n46065 = n44927 & ~n44996 ;
  assign n46066 = n44985 & ~n46065 ;
  assign n46067 = ~n44947 & ~n46066 ;
  assign n46068 = n44954 & ~n46067 ;
  assign n46075 = ~n46064 & ~n46068 ;
  assign n46076 = ~n46074 & n46075 ;
  assign n46077 = n44921 & ~n46076 ;
  assign n46079 = ~n45417 & ~n45425 ;
  assign n46080 = ~n44954 & ~n46079 ;
  assign n46081 = ~n44933 & n44978 ;
  assign n46082 = n44954 & ~n45417 ;
  assign n46083 = ~n46081 & n46082 ;
  assign n46084 = ~n46080 & ~n46083 ;
  assign n46078 = n44933 & ~n45419 ;
  assign n46085 = n44995 & ~n46078 ;
  assign n46086 = ~n46084 & n46085 ;
  assign n46087 = ~n44921 & ~n46086 ;
  assign n46088 = n44954 & n44977 ;
  assign n46089 = ~n44965 & n44992 ;
  assign n46090 = n44958 & n46089 ;
  assign n46091 = ~n46088 & ~n46090 ;
  assign n46092 = ~n46087 & n46091 ;
  assign n46093 = ~n46077 & n46092 ;
  assign n46094 = \u1_L2_reg[32]/NET0131  & n46093 ;
  assign n46095 = ~\u1_L2_reg[32]/NET0131  & ~n46093 ;
  assign n46096 = ~n46094 & ~n46095 ;
  assign n46116 = decrypt_pad & ~\u1_uk_K_r2_reg[12]/NET0131  ;
  assign n46117 = ~decrypt_pad & ~\u1_uk_K_r2_reg[17]/NET0131  ;
  assign n46118 = ~n46116 & ~n46117 ;
  assign n46119 = \u1_R2_reg[11]/NET0131  & ~n46118 ;
  assign n46120 = ~\u1_R2_reg[11]/NET0131  & n46118 ;
  assign n46121 = ~n46119 & ~n46120 ;
  assign n46097 = decrypt_pad & ~\u1_uk_K_r2_reg[27]/NET0131  ;
  assign n46098 = ~decrypt_pad & ~\u1_uk_K_r2_reg[32]/NET0131  ;
  assign n46099 = ~n46097 & ~n46098 ;
  assign n46100 = \u1_R2_reg[12]/NET0131  & ~n46099 ;
  assign n46101 = ~\u1_R2_reg[12]/NET0131  & n46099 ;
  assign n46102 = ~n46100 & ~n46101 ;
  assign n46103 = decrypt_pad & ~\u1_uk_K_r2_reg[3]/NET0131  ;
  assign n46104 = ~decrypt_pad & ~\u1_uk_K_r2_reg[40]/NET0131  ;
  assign n46105 = ~n46103 & ~n46104 ;
  assign n46106 = \u1_R2_reg[9]/NET0131  & ~n46105 ;
  assign n46107 = ~\u1_R2_reg[9]/NET0131  & n46105 ;
  assign n46108 = ~n46106 & ~n46107 ;
  assign n46130 = decrypt_pad & ~\u1_uk_K_r2_reg[40]/NET0131  ;
  assign n46131 = ~decrypt_pad & ~\u1_uk_K_r2_reg[20]/NET0131  ;
  assign n46132 = ~n46130 & ~n46131 ;
  assign n46133 = \u1_R2_reg[13]/NET0131  & ~n46132 ;
  assign n46134 = ~\u1_R2_reg[13]/NET0131  & n46132 ;
  assign n46135 = ~n46133 & ~n46134 ;
  assign n46159 = ~n46108 & n46135 ;
  assign n46109 = decrypt_pad & ~\u1_uk_K_r2_reg[11]/NET0131  ;
  assign n46110 = ~decrypt_pad & ~\u1_uk_K_r2_reg[48]/NET0131  ;
  assign n46111 = ~n46109 & ~n46110 ;
  assign n46112 = \u1_R2_reg[10]/NET0131  & ~n46111 ;
  assign n46113 = ~\u1_R2_reg[10]/NET0131  & n46111 ;
  assign n46114 = ~n46112 & ~n46113 ;
  assign n46122 = decrypt_pad & ~\u1_uk_K_r2_reg[6]/NET0131  ;
  assign n46123 = ~decrypt_pad & ~\u1_uk_K_r2_reg[11]/NET0131  ;
  assign n46124 = ~n46122 & ~n46123 ;
  assign n46125 = \u1_R2_reg[8]/NET0131  & ~n46124 ;
  assign n46126 = ~\u1_R2_reg[8]/NET0131  & n46124 ;
  assign n46127 = ~n46125 & ~n46126 ;
  assign n46136 = ~n46127 & n46135 ;
  assign n46137 = n46114 & n46136 ;
  assign n46141 = n46127 & ~n46135 ;
  assign n46166 = n46108 & n46141 ;
  assign n46167 = ~n46137 & ~n46166 ;
  assign n46168 = ~n46159 & n46167 ;
  assign n46169 = n46102 & ~n46168 ;
  assign n46165 = n46114 & n46159 ;
  assign n46144 = ~n46127 & ~n46135 ;
  assign n46170 = ~n46114 & n46144 ;
  assign n46171 = ~n46108 & n46170 ;
  assign n46172 = ~n46165 & ~n46171 ;
  assign n46173 = ~n46169 & n46172 ;
  assign n46174 = n46121 & ~n46173 ;
  assign n46140 = n46108 & n46114 ;
  assign n46143 = ~n46108 & ~n46114 ;
  assign n46145 = n46127 & n46135 ;
  assign n46146 = ~n46144 & ~n46145 ;
  assign n46147 = ~n46143 & ~n46146 ;
  assign n46148 = ~n46140 & n46147 ;
  assign n46138 = n46108 & n46137 ;
  assign n46139 = ~n46121 & n46138 ;
  assign n46128 = n46121 & ~n46127 ;
  assign n46149 = ~n46128 & n46143 ;
  assign n46150 = n46146 & n46149 ;
  assign n46115 = n46108 & ~n46114 ;
  assign n46129 = n46115 & n46128 ;
  assign n46142 = n46140 & n46141 ;
  assign n46151 = ~n46129 & ~n46142 ;
  assign n46152 = ~n46150 & n46151 ;
  assign n46153 = ~n46139 & n46152 ;
  assign n46154 = ~n46148 & n46153 ;
  assign n46155 = ~n46102 & ~n46154 ;
  assign n46156 = n46102 & n46140 ;
  assign n46157 = n46144 & n46156 ;
  assign n46160 = ~n46115 & ~n46127 ;
  assign n46158 = n46108 & ~n46135 ;
  assign n46161 = n46102 & ~n46121 ;
  assign n46162 = ~n46158 & n46161 ;
  assign n46163 = ~n46159 & n46162 ;
  assign n46164 = ~n46160 & n46163 ;
  assign n46175 = ~n46157 & ~n46164 ;
  assign n46176 = ~n46155 & n46175 ;
  assign n46177 = ~n46174 & n46176 ;
  assign n46178 = ~\u1_L2_reg[6]/NET0131  & ~n46177 ;
  assign n46179 = \u1_L2_reg[6]/NET0131  & n46177 ;
  assign n46180 = ~n46178 & ~n46179 ;
  assign n46198 = ~n44946 & ~n45423 ;
  assign n46181 = n44933 & ~n46069 ;
  assign n46199 = n44927 & n44996 ;
  assign n46200 = ~n46181 & ~n46199 ;
  assign n46201 = ~n46198 & n46200 ;
  assign n46202 = ~n44954 & ~n46201 ;
  assign n46182 = ~n46081 & ~n46181 ;
  assign n46183 = n44927 & ~n46182 ;
  assign n46192 = ~n44927 & ~n44940 ;
  assign n46193 = n46069 & n46192 ;
  assign n46203 = n44954 & n46193 ;
  assign n46204 = ~n46183 & ~n46203 ;
  assign n46205 = ~n46202 & n46204 ;
  assign n46206 = n44921 & ~n46205 ;
  assign n46184 = ~n44954 & n46183 ;
  assign n46185 = n44921 & ~n44954 ;
  assign n46186 = n44984 & ~n46069 ;
  assign n46187 = n44939 & ~n45435 ;
  assign n46188 = n44954 & n46065 ;
  assign n46189 = ~n46187 & n46188 ;
  assign n46190 = ~n46186 & ~n46189 ;
  assign n46191 = ~n44921 & ~n46190 ;
  assign n46194 = ~n44954 & n46193 ;
  assign n46195 = ~n44948 & ~n46194 ;
  assign n46196 = ~n46191 & n46195 ;
  assign n46197 = ~n46185 & ~n46196 ;
  assign n46207 = ~n46184 & ~n46197 ;
  assign n46208 = ~n46206 & n46207 ;
  assign n46209 = ~\u1_L2_reg[7]/NET0131  & ~n46208 ;
  assign n46210 = \u1_L2_reg[7]/NET0131  & n46208 ;
  assign n46211 = ~n46209 & ~n46210 ;
  assign n46226 = ~n45471 & n45505 ;
  assign n46227 = ~n45699 & ~n46226 ;
  assign n46228 = n45494 & ~n46227 ;
  assign n46229 = ~n45471 & n45707 ;
  assign n46230 = ~n45513 & ~n46229 ;
  assign n46231 = ~n46228 & n46230 ;
  assign n46232 = n45452 & ~n46231 ;
  assign n46212 = n45494 & n45692 ;
  assign n46217 = ~n45482 & ~n46212 ;
  assign n46218 = n45709 & n46217 ;
  assign n46213 = ~n45479 & n45510 ;
  assign n46214 = ~n45699 & ~n46213 ;
  assign n46215 = ~n45494 & ~n46214 ;
  assign n46216 = n45494 & n45527 ;
  assign n46219 = ~n46215 & ~n46216 ;
  assign n46220 = n46218 & n46219 ;
  assign n46221 = ~n45452 & ~n46220 ;
  assign n46222 = ~n45464 & n45708 ;
  assign n46223 = ~n45480 & n45510 ;
  assign n46224 = ~n45525 & ~n46223 ;
  assign n46225 = n45494 & ~n46224 ;
  assign n46233 = ~n46222 & ~n46225 ;
  assign n46234 = ~n46221 & n46233 ;
  assign n46235 = ~n46232 & n46234 ;
  assign n46236 = ~\u1_L2_reg[8]/NET0131  & ~n46235 ;
  assign n46237 = \u1_L2_reg[8]/NET0131  & n46235 ;
  assign n46238 = ~n46236 & ~n46237 ;
  assign n46239 = n46108 & n46145 ;
  assign n46240 = ~n46108 & ~n46145 ;
  assign n46241 = ~n46239 & ~n46240 ;
  assign n46242 = ~n46144 & ~n46241 ;
  assign n46243 = n46128 & n46158 ;
  assign n46244 = ~n46242 & ~n46243 ;
  assign n46245 = ~n46114 & ~n46244 ;
  assign n46246 = n46114 & n46144 ;
  assign n46247 = ~n46114 & n46141 ;
  assign n46248 = ~n46246 & ~n46247 ;
  assign n46249 = ~n46121 & ~n46248 ;
  assign n46250 = n46102 & ~n46138 ;
  assign n46251 = ~n46249 & n46250 ;
  assign n46252 = ~n46245 & n46251 ;
  assign n46255 = ~n46108 & ~n46127 ;
  assign n46256 = n46135 & n46255 ;
  assign n46257 = ~n46170 & ~n46239 ;
  assign n46258 = ~n46256 & n46257 ;
  assign n46259 = ~n46121 & ~n46258 ;
  assign n46253 = n46121 & ~n46144 ;
  assign n46254 = n46241 & n46253 ;
  assign n46260 = ~n46102 & ~n46171 ;
  assign n46261 = ~n46254 & n46260 ;
  assign n46262 = ~n46259 & n46261 ;
  assign n46263 = ~n46252 & ~n46262 ;
  assign n46264 = n46114 & n46127 ;
  assign n46265 = ~n46108 & n46264 ;
  assign n46266 = ~n46121 & n46265 ;
  assign n46267 = ~n46108 & n46246 ;
  assign n46268 = ~n46142 & ~n46267 ;
  assign n46269 = n46121 & ~n46268 ;
  assign n46270 = ~n46266 & ~n46269 ;
  assign n46271 = ~n46263 & n46270 ;
  assign n46272 = ~\u1_L2_reg[16]/NET0131  & ~n46271 ;
  assign n46273 = \u1_L2_reg[16]/NET0131  & n46271 ;
  assign n46274 = ~n46272 & ~n46273 ;
  assign n46277 = ~n46121 & n46167 ;
  assign n46275 = ~n46135 & n46265 ;
  assign n46276 = n46143 & ~n46146 ;
  assign n46278 = ~n46275 & ~n46276 ;
  assign n46279 = n46277 & n46278 ;
  assign n46280 = ~n46114 & n46136 ;
  assign n46281 = ~n46246 & ~n46280 ;
  assign n46282 = n46108 & n46144 ;
  assign n46283 = n46121 & ~n46265 ;
  assign n46284 = ~n46282 & n46283 ;
  assign n46285 = n46281 & n46284 ;
  assign n46286 = ~n46279 & ~n46285 ;
  assign n46287 = ~n46102 & ~n46286 ;
  assign n46289 = ~n46114 & n46121 ;
  assign n46290 = ~n46108 & ~n46136 ;
  assign n46291 = n46289 & n46290 ;
  assign n46295 = n46102 & ~n46150 ;
  assign n46296 = ~n46291 & n46295 ;
  assign n46288 = ~n46121 & n46147 ;
  assign n46292 = n46108 & n46264 ;
  assign n46293 = ~n46137 & ~n46292 ;
  assign n46294 = n46121 & ~n46293 ;
  assign n46297 = ~n46288 & ~n46294 ;
  assign n46298 = n46296 & n46297 ;
  assign n46299 = ~n46287 & ~n46298 ;
  assign n46300 = n46114 & ~n46121 ;
  assign n46301 = n46239 & n46300 ;
  assign n46302 = ~n46158 & ~n46255 ;
  assign n46303 = ~n46145 & n46289 ;
  assign n46304 = n46302 & n46303 ;
  assign n46305 = ~n46301 & ~n46304 ;
  assign n46306 = ~n46299 & n46305 ;
  assign n46307 = ~\u1_L2_reg[24]/NET0131  & ~n46306 ;
  assign n46308 = \u1_L2_reg[24]/NET0131  & n46306 ;
  assign n46309 = ~n46307 & ~n46308 ;
  assign n46314 = n46141 & n46143 ;
  assign n46315 = n46281 & ~n46314 ;
  assign n46316 = n46121 & ~n46315 ;
  assign n46311 = n46140 & ~n46145 ;
  assign n46312 = ~n46264 & ~n46282 ;
  assign n46313 = ~n46121 & ~n46312 ;
  assign n46317 = ~n46311 & ~n46313 ;
  assign n46318 = ~n46316 & n46317 ;
  assign n46319 = n46102 & ~n46318 ;
  assign n46328 = ~n46121 & ~n46264 ;
  assign n46329 = n46302 & n46328 ;
  assign n46327 = ~n46127 & n46165 ;
  assign n46330 = ~n46276 & ~n46327 ;
  assign n46331 = ~n46329 & n46330 ;
  assign n46332 = ~n46102 & ~n46331 ;
  assign n46310 = n46158 & n46300 ;
  assign n46320 = ~n46158 & n46264 ;
  assign n46321 = n46115 & ~n46135 ;
  assign n46322 = ~n46320 & ~n46321 ;
  assign n46323 = ~n46102 & ~n46322 ;
  assign n46324 = n46127 & n46165 ;
  assign n46325 = ~n46323 & ~n46324 ;
  assign n46326 = n46121 & ~n46325 ;
  assign n46333 = ~n46310 & ~n46326 ;
  assign n46334 = ~n46332 & n46333 ;
  assign n46335 = ~n46319 & n46334 ;
  assign n46336 = \u1_L2_reg[30]/NET0131  & ~n46335 ;
  assign n46337 = ~\u1_L2_reg[30]/NET0131  & n46335 ;
  assign n46338 = ~n46336 & ~n46337 ;
  assign n46349 = n45458 & n45533 ;
  assign n46350 = ~n45509 & ~n46349 ;
  assign n46351 = n45494 & ~n46350 ;
  assign n46352 = ~n45494 & n45514 ;
  assign n46348 = n45471 & n45526 ;
  assign n46353 = ~n45528 & ~n46348 ;
  assign n46354 = ~n46352 & n46353 ;
  assign n46355 = ~n46351 & n46354 ;
  assign n46356 = n45452 & ~n46355 ;
  assign n46343 = ~n45487 & ~n45710 ;
  assign n46344 = n45494 & ~n46343 ;
  assign n46340 = ~n45465 & n45479 ;
  assign n46341 = ~n45534 & ~n45699 ;
  assign n46342 = ~n45494 & ~n46341 ;
  assign n46345 = ~n46340 & ~n46342 ;
  assign n46346 = ~n46344 & n46345 ;
  assign n46347 = ~n45452 & ~n46346 ;
  assign n46357 = n45479 & n45496 ;
  assign n46358 = ~n45503 & ~n46357 ;
  assign n46359 = ~n46226 & n46358 ;
  assign n46360 = ~n45494 & ~n46359 ;
  assign n46339 = n45497 & n45511 ;
  assign n46361 = ~n46216 & ~n46339 ;
  assign n46362 = ~n46360 & n46361 ;
  assign n46363 = ~n46347 & n46362 ;
  assign n46364 = ~n46356 & n46363 ;
  assign n46365 = ~\u1_L2_reg[3]/NET0131  & ~n46364 ;
  assign n46366 = \u1_L2_reg[3]/NET0131  & n46364 ;
  assign n46367 = ~n46365 & ~n46366 ;
  assign n46373 = ~n45053 & ~n45056 ;
  assign n46374 = ~n45548 & n46373 ;
  assign n46375 = n45025 & ~n46374 ;
  assign n46370 = n45019 & n45551 ;
  assign n46368 = ~n45039 & n45546 ;
  assign n46369 = ~n45025 & n46368 ;
  assign n46371 = ~n45019 & n45047 ;
  assign n46372 = n45039 & n46371 ;
  assign n46376 = ~n46369 & ~n46372 ;
  assign n46377 = ~n46370 & n46376 ;
  assign n46378 = ~n46375 & n46377 ;
  assign n46379 = ~n45013 & ~n46378 ;
  assign n46380 = n45070 & n45088 ;
  assign n46381 = ~n46372 & ~n46380 ;
  assign n46382 = ~n45025 & ~n46381 ;
  assign n46384 = n45019 & ~n45048 ;
  assign n46385 = ~n45551 & n46384 ;
  assign n46383 = n45073 & n46368 ;
  assign n46386 = ~n45564 & ~n46383 ;
  assign n46387 = ~n46385 & n46386 ;
  assign n46388 = n45013 & ~n46387 ;
  assign n46389 = ~n46382 & ~n46388 ;
  assign n46390 = ~n46379 & n46389 ;
  assign n46391 = ~\u1_L2_reg[9]/NET0131  & ~n46390 ;
  assign n46392 = \u1_L2_reg[9]/NET0131  & n46390 ;
  assign n46393 = ~n46391 & ~n46392 ;
  assign n46403 = n45800 & ~n45838 ;
  assign n46404 = ~n45841 & ~n45946 ;
  assign n46405 = ~n45897 & ~n45901 ;
  assign n46406 = ~n46404 & n46405 ;
  assign n46407 = ~n46403 & ~n46406 ;
  assign n46408 = n45794 & ~n46407 ;
  assign n46395 = n45813 & n45852 ;
  assign n46398 = ~n45879 & ~n45950 ;
  assign n46399 = ~n46395 & n46398 ;
  assign n46396 = ~n45852 & ~n45861 ;
  assign n46397 = n45860 & n46396 ;
  assign n46400 = ~n45827 & ~n46397 ;
  assign n46401 = n46399 & n46400 ;
  assign n46402 = ~n45794 & ~n46401 ;
  assign n46394 = ~n45800 & n45883 ;
  assign n46409 = n45813 & n45826 ;
  assign n46410 = ~n45945 & ~n46409 ;
  assign n46411 = n45800 & ~n46410 ;
  assign n46412 = ~n46394 & ~n46411 ;
  assign n46413 = ~n46402 & n46412 ;
  assign n46414 = ~n46408 & n46413 ;
  assign n46415 = \u1_L2_reg[18]/NET0131  & n46414 ;
  assign n46416 = ~\u1_L2_reg[18]/NET0131  & ~n46414 ;
  assign n46417 = ~n46415 & ~n46416 ;
  assign n46418 = decrypt_pad & ~\u1_uk_K_r1_reg[34]/NET0131  ;
  assign n46419 = ~decrypt_pad & ~\u1_uk_K_r1_reg[10]/P0001  ;
  assign n46420 = ~n46418 & ~n46419 ;
  assign n46421 = \u1_R1_reg[4]/NET0131  & ~n46420 ;
  assign n46422 = ~\u1_R1_reg[4]/NET0131  & n46420 ;
  assign n46423 = ~n46421 & ~n46422 ;
  assign n46443 = decrypt_pad & ~\u1_uk_K_r1_reg[11]/NET0131  ;
  assign n46444 = ~decrypt_pad & ~\u1_uk_K_r1_reg[19]/NET0131  ;
  assign n46445 = ~n46443 & ~n46444 ;
  assign n46446 = \u1_R1_reg[32]/NET0131  & ~n46445 ;
  assign n46447 = ~\u1_R1_reg[32]/NET0131  & n46445 ;
  assign n46448 = ~n46446 & ~n46447 ;
  assign n46452 = decrypt_pad & ~\u1_uk_K_r1_reg[32]/NET0131  ;
  assign n46453 = ~decrypt_pad & ~\u1_uk_K_r1_reg[40]/NET0131  ;
  assign n46454 = ~n46452 & ~n46453 ;
  assign n46455 = \u1_R1_reg[1]/NET0131  & ~n46454 ;
  assign n46456 = ~\u1_R1_reg[1]/NET0131  & n46454 ;
  assign n46457 = ~n46455 & ~n46456 ;
  assign n46424 = decrypt_pad & ~\u1_uk_K_r1_reg[47]/NET0131  ;
  assign n46425 = ~decrypt_pad & ~\u1_uk_K_r1_reg[55]/NET0131  ;
  assign n46426 = ~n46424 & ~n46425 ;
  assign n46427 = \u1_R1_reg[2]/NET0131  & ~n46426 ;
  assign n46428 = ~\u1_R1_reg[2]/NET0131  & n46426 ;
  assign n46429 = ~n46427 & ~n46428 ;
  assign n46437 = decrypt_pad & ~\u1_uk_K_r1_reg[5]/NET0131  ;
  assign n46438 = ~decrypt_pad & ~\u1_uk_K_r1_reg[13]/NET0131  ;
  assign n46439 = ~n46437 & ~n46438 ;
  assign n46440 = \u1_R1_reg[5]/NET0131  & ~n46439 ;
  assign n46441 = ~\u1_R1_reg[5]/NET0131  & n46439 ;
  assign n46442 = ~n46440 & ~n46441 ;
  assign n46485 = ~n46429 & ~n46442 ;
  assign n46486 = ~n46457 & n46485 ;
  assign n46487 = n46448 & ~n46486 ;
  assign n46450 = ~n46442 & ~n46448 ;
  assign n46430 = decrypt_pad & ~\u1_uk_K_r1_reg[24]/NET0131  ;
  assign n46431 = ~decrypt_pad & ~\u1_uk_K_r1_reg[32]/NET0131  ;
  assign n46432 = ~n46430 & ~n46431 ;
  assign n46433 = \u1_R1_reg[3]/NET0131  & ~n46432 ;
  assign n46434 = ~\u1_R1_reg[3]/NET0131  & n46432 ;
  assign n46435 = ~n46433 & ~n46434 ;
  assign n46483 = ~n46429 & n46435 ;
  assign n46484 = n46457 & ~n46483 ;
  assign n46488 = ~n46450 & ~n46484 ;
  assign n46489 = ~n46487 & n46488 ;
  assign n46466 = n46442 & ~n46457 ;
  assign n46476 = n46429 & ~n46448 ;
  assign n46477 = ~n46442 & n46476 ;
  assign n46478 = ~n46466 & ~n46477 ;
  assign n46479 = n46435 & ~n46478 ;
  assign n46480 = ~n46448 & n46457 ;
  assign n46460 = ~n46435 & n46457 ;
  assign n46481 = ~n46460 & ~n46476 ;
  assign n46482 = ~n46480 & ~n46481 ;
  assign n46490 = ~n46479 & ~n46482 ;
  assign n46491 = ~n46489 & n46490 ;
  assign n46492 = n46423 & ~n46491 ;
  assign n46467 = ~n46429 & ~n46448 ;
  assign n46468 = n46448 & ~n46457 ;
  assign n46469 = n46429 & n46468 ;
  assign n46470 = ~n46467 & ~n46469 ;
  assign n46471 = ~n46435 & ~n46466 ;
  assign n46472 = ~n46470 & n46471 ;
  assign n46436 = n46429 & n46435 ;
  assign n46449 = n46442 & n46448 ;
  assign n46451 = ~n46449 & ~n46450 ;
  assign n46458 = n46451 & n46457 ;
  assign n46459 = n46436 & n46458 ;
  assign n46461 = n46449 & ~n46460 ;
  assign n46462 = ~n46442 & n46457 ;
  assign n46463 = ~n46448 & n46462 ;
  assign n46464 = ~n46461 & ~n46463 ;
  assign n46465 = ~n46429 & ~n46464 ;
  assign n46473 = ~n46459 & ~n46465 ;
  assign n46474 = ~n46472 & n46473 ;
  assign n46475 = ~n46423 & ~n46474 ;
  assign n46493 = n46435 & ~n46457 ;
  assign n46494 = ~n46429 & n46448 ;
  assign n46495 = ~n46477 & ~n46494 ;
  assign n46496 = n46493 & ~n46495 ;
  assign n46498 = n46429 & n46442 ;
  assign n46499 = n46457 & n46498 ;
  assign n46500 = n46448 & n46499 ;
  assign n46497 = n46466 & n46476 ;
  assign n46501 = n46457 & n46485 ;
  assign n46502 = ~n46497 & ~n46501 ;
  assign n46503 = ~n46500 & n46502 ;
  assign n46504 = ~n46435 & ~n46503 ;
  assign n46505 = ~n46496 & ~n46504 ;
  assign n46506 = ~n46475 & n46505 ;
  assign n46507 = ~n46492 & n46506 ;
  assign n46508 = ~\u1_L1_reg[31]/NET0131  & ~n46507 ;
  assign n46509 = \u1_L1_reg[31]/NET0131  & n46507 ;
  assign n46510 = ~n46508 & ~n46509 ;
  assign n46511 = decrypt_pad & ~\u1_uk_K_r1_reg[1]/NET0131  ;
  assign n46512 = ~decrypt_pad & ~\u1_uk_K_r1_reg[7]/P0001  ;
  assign n46513 = ~n46511 & ~n46512 ;
  assign n46514 = \u1_R1_reg[24]/NET0131  & ~n46513 ;
  assign n46515 = ~\u1_R1_reg[24]/NET0131  & n46513 ;
  assign n46516 = ~n46514 & ~n46515 ;
  assign n46523 = decrypt_pad & ~\u1_uk_K_r1_reg[35]/NET0131  ;
  assign n46524 = ~decrypt_pad & ~\u1_uk_K_r1_reg[45]/NET0131  ;
  assign n46525 = ~n46523 & ~n46524 ;
  assign n46526 = \u1_R1_reg[20]/NET0131  & ~n46525 ;
  assign n46527 = ~\u1_R1_reg[20]/NET0131  & n46525 ;
  assign n46528 = ~n46526 & ~n46527 ;
  assign n46530 = decrypt_pad & ~\u1_uk_K_r1_reg[50]/NET0131  ;
  assign n46531 = ~decrypt_pad & ~\u1_uk_K_r1_reg[1]/NET0131  ;
  assign n46532 = ~n46530 & ~n46531 ;
  assign n46533 = \u1_R1_reg[21]/NET0131  & ~n46532 ;
  assign n46534 = ~\u1_R1_reg[21]/NET0131  & n46532 ;
  assign n46535 = ~n46533 & ~n46534 ;
  assign n46536 = decrypt_pad & ~\u1_uk_K_r1_reg[51]/NET0131  ;
  assign n46537 = ~decrypt_pad & ~\u1_uk_K_r1_reg[2]/NET0131  ;
  assign n46538 = ~n46536 & ~n46537 ;
  assign n46539 = \u1_R1_reg[25]/NET0131  & ~n46538 ;
  assign n46540 = ~\u1_R1_reg[25]/NET0131  & n46538 ;
  assign n46541 = ~n46539 & ~n46540 ;
  assign n46575 = n46535 & n46541 ;
  assign n46576 = ~n46528 & n46575 ;
  assign n46517 = decrypt_pad & ~\u1_uk_K_r1_reg[45]/NET0131  ;
  assign n46518 = ~decrypt_pad & ~\u1_uk_K_r1_reg[23]/NET0131  ;
  assign n46519 = ~n46517 & ~n46518 ;
  assign n46520 = \u1_R1_reg[22]/NET0131  & ~n46519 ;
  assign n46521 = ~\u1_R1_reg[22]/NET0131  & n46519 ;
  assign n46522 = ~n46520 & ~n46521 ;
  assign n46553 = n46528 & ~n46535 ;
  assign n46554 = n46541 & n46553 ;
  assign n46577 = ~n46522 & ~n46554 ;
  assign n46578 = ~n46576 & n46577 ;
  assign n46573 = n46528 & n46541 ;
  assign n46574 = n46522 & n46573 ;
  assign n46545 = decrypt_pad & ~\u1_uk_K_r1_reg[30]/NET0131  ;
  assign n46546 = ~decrypt_pad & ~\u1_uk_K_r1_reg[36]/NET0131  ;
  assign n46547 = ~n46545 & ~n46546 ;
  assign n46548 = \u1_R1_reg[23]/NET0131  & ~n46547 ;
  assign n46549 = ~\u1_R1_reg[23]/NET0131  & n46547 ;
  assign n46550 = ~n46548 & ~n46549 ;
  assign n46557 = ~n46528 & n46535 ;
  assign n46558 = n46522 & n46557 ;
  assign n46579 = ~n46550 & ~n46558 ;
  assign n46580 = ~n46574 & n46579 ;
  assign n46581 = ~n46578 & n46580 ;
  assign n46544 = n46528 & ~n46541 ;
  assign n46583 = ~n46522 & ~n46535 ;
  assign n46584 = n46544 & n46583 ;
  assign n46582 = n46535 & n46573 ;
  assign n46585 = ~n46558 & ~n46582 ;
  assign n46586 = ~n46584 & n46585 ;
  assign n46587 = n46550 & ~n46586 ;
  assign n46588 = ~n46581 & ~n46587 ;
  assign n46589 = n46516 & ~n46588 ;
  assign n46565 = n46522 & ~n46553 ;
  assign n46529 = ~n46522 & n46528 ;
  assign n46566 = ~n46529 & n46550 ;
  assign n46567 = ~n46565 & n46566 ;
  assign n46542 = n46535 & ~n46541 ;
  assign n46543 = n46529 & n46542 ;
  assign n46562 = ~n46528 & n46541 ;
  assign n46563 = ~n46535 & n46562 ;
  assign n46564 = n46550 & n46563 ;
  assign n46568 = ~n46543 & ~n46564 ;
  assign n46569 = ~n46567 & n46568 ;
  assign n46551 = ~n46522 & ~n46550 ;
  assign n46552 = n46544 & n46551 ;
  assign n46555 = n46522 & n46554 ;
  assign n46556 = ~n46552 & ~n46555 ;
  assign n46559 = n46529 & n46535 ;
  assign n46560 = ~n46558 & ~n46559 ;
  assign n46561 = ~n46550 & ~n46560 ;
  assign n46570 = n46556 & ~n46561 ;
  assign n46571 = n46569 & n46570 ;
  assign n46572 = ~n46516 & ~n46571 ;
  assign n46591 = ~n46541 & n46557 ;
  assign n46592 = ~n46522 & n46591 ;
  assign n46593 = ~n46574 & ~n46592 ;
  assign n46594 = n46550 & ~n46593 ;
  assign n46590 = ~n46522 & n46564 ;
  assign n46595 = ~n46528 & ~n46541 ;
  assign n46596 = ~n46535 & n46595 ;
  assign n46597 = n46528 & n46542 ;
  assign n46598 = ~n46596 & ~n46597 ;
  assign n46599 = n46551 & ~n46598 ;
  assign n46600 = ~n46590 & ~n46599 ;
  assign n46601 = ~n46594 & n46600 ;
  assign n46602 = ~n46572 & n46601 ;
  assign n46603 = ~n46589 & n46602 ;
  assign n46604 = \u1_L1_reg[11]/NET0131  & ~n46603 ;
  assign n46605 = ~\u1_L1_reg[11]/NET0131  & n46603 ;
  assign n46606 = ~n46604 & ~n46605 ;
  assign n46607 = decrypt_pad & ~\u1_uk_K_r1_reg[8]/NET0131  ;
  assign n46608 = ~decrypt_pad & ~\u1_uk_K_r1_reg[14]/NET0131  ;
  assign n46609 = ~n46607 & ~n46608 ;
  assign n46610 = \u1_R1_reg[28]/NET0131  & ~n46609 ;
  assign n46611 = ~\u1_R1_reg[28]/NET0131  & n46609 ;
  assign n46612 = ~n46610 & ~n46611 ;
  assign n46626 = decrypt_pad & ~\u1_uk_K_r1_reg[23]/NET0131  ;
  assign n46627 = ~decrypt_pad & ~\u1_uk_K_r1_reg[29]/NET0131  ;
  assign n46628 = ~n46626 & ~n46627 ;
  assign n46629 = \u1_R1_reg[24]/NET0131  & ~n46628 ;
  assign n46630 = ~\u1_R1_reg[24]/NET0131  & n46628 ;
  assign n46631 = ~n46629 & ~n46630 ;
  assign n46632 = decrypt_pad & ~\u1_uk_K_r1_reg[43]/NET0131  ;
  assign n46633 = ~decrypt_pad & ~\u1_uk_K_r1_reg[49]/NET0131  ;
  assign n46634 = ~n46632 & ~n46633 ;
  assign n46635 = \u1_R1_reg[26]/NET0131  & ~n46634 ;
  assign n46636 = ~\u1_R1_reg[26]/NET0131  & n46634 ;
  assign n46637 = ~n46635 & ~n46636 ;
  assign n46619 = decrypt_pad & ~\u1_uk_K_r1_reg[31]/NET0131  ;
  assign n46620 = ~decrypt_pad & ~\u1_uk_K_r1_reg[9]/NET0131  ;
  assign n46621 = ~n46619 & ~n46620 ;
  assign n46622 = \u1_R1_reg[25]/NET0131  & ~n46621 ;
  assign n46623 = ~\u1_R1_reg[25]/NET0131  & n46621 ;
  assign n46624 = ~n46622 & ~n46623 ;
  assign n46640 = decrypt_pad & ~\u1_uk_K_r1_reg[21]/NET0131  ;
  assign n46641 = ~decrypt_pad & ~\u1_uk_K_r1_reg[31]/NET0131  ;
  assign n46642 = ~n46640 & ~n46641 ;
  assign n46643 = \u1_R1_reg[27]/NET0131  & ~n46642 ;
  assign n46644 = ~\u1_R1_reg[27]/NET0131  & n46642 ;
  assign n46645 = ~n46643 & ~n46644 ;
  assign n46647 = ~n46624 & n46645 ;
  assign n46648 = ~n46637 & n46647 ;
  assign n46613 = decrypt_pad & ~\u1_uk_K_r1_reg[0]/NET0131  ;
  assign n46614 = ~decrypt_pad & ~\u1_uk_K_r1_reg[37]/NET0131  ;
  assign n46615 = ~n46613 & ~n46614 ;
  assign n46616 = \u1_R1_reg[29]/NET0131  & ~n46615 ;
  assign n46617 = ~\u1_R1_reg[29]/NET0131  & n46615 ;
  assign n46618 = ~n46616 & ~n46617 ;
  assign n46650 = n46618 & ~n46637 ;
  assign n46649 = ~n46624 & n46637 ;
  assign n46651 = ~n46645 & ~n46649 ;
  assign n46652 = ~n46650 & n46651 ;
  assign n46653 = ~n46648 & ~n46652 ;
  assign n46654 = n46631 & ~n46653 ;
  assign n46625 = ~n46618 & ~n46624 ;
  assign n46638 = ~n46631 & n46637 ;
  assign n46639 = n46625 & n46638 ;
  assign n46646 = n46639 & ~n46645 ;
  assign n46655 = ~n46631 & ~n46637 ;
  assign n46656 = n46631 & n46637 ;
  assign n46657 = ~n46655 & ~n46656 ;
  assign n46658 = n46618 & ~n46647 ;
  assign n46659 = ~n46657 & n46658 ;
  assign n46660 = ~n46646 & ~n46659 ;
  assign n46661 = ~n46654 & n46660 ;
  assign n46662 = ~n46612 & ~n46661 ;
  assign n46663 = ~n46618 & n46648 ;
  assign n46664 = n46624 & ~n46645 ;
  assign n46665 = ~n46657 & n46664 ;
  assign n46691 = ~n46663 & ~n46665 ;
  assign n46692 = ~n46662 & n46691 ;
  assign n46666 = ~n46624 & ~n46637 ;
  assign n46667 = n46624 & n46637 ;
  assign n46668 = ~n46666 & ~n46667 ;
  assign n46669 = ~n46618 & n46624 ;
  assign n46670 = n46612 & ~n46669 ;
  assign n46671 = n46668 & n46670 ;
  assign n46672 = ~n46625 & ~n46671 ;
  assign n46673 = n46631 & ~n46672 ;
  assign n46674 = n46618 & ~n46624 ;
  assign n46675 = ~n46669 & ~n46674 ;
  assign n46676 = n46638 & ~n46675 ;
  assign n46677 = ~n46673 & ~n46676 ;
  assign n46678 = n46645 & ~n46677 ;
  assign n46681 = n46618 & ~n46631 ;
  assign n46682 = n46624 & n46681 ;
  assign n46685 = n46637 & ~n46682 ;
  assign n46683 = n46631 & n46674 ;
  assign n46684 = ~n46682 & ~n46683 ;
  assign n46686 = ~n46645 & ~n46684 ;
  assign n46687 = ~n46685 & n46686 ;
  assign n46679 = n46638 & n46674 ;
  assign n46680 = n46625 & n46655 ;
  assign n46688 = ~n46679 & ~n46680 ;
  assign n46689 = ~n46687 & n46688 ;
  assign n46690 = n46612 & ~n46689 ;
  assign n46693 = ~n46678 & ~n46690 ;
  assign n46694 = n46692 & n46693 ;
  assign n46695 = ~\u1_L1_reg[22]/NET0131  & ~n46694 ;
  assign n46696 = \u1_L1_reg[22]/NET0131  & n46694 ;
  assign n46697 = ~n46695 & ~n46696 ;
  assign n46703 = ~n46451 & ~n46457 ;
  assign n46704 = ~n46442 & n46467 ;
  assign n46705 = ~n46703 & ~n46704 ;
  assign n46706 = ~n46435 & ~n46705 ;
  assign n46698 = ~n46462 & ~n46466 ;
  assign n46699 = n46435 & n46698 ;
  assign n46700 = n46429 & n46462 ;
  assign n46701 = ~n46699 & ~n46700 ;
  assign n46702 = n46448 & ~n46701 ;
  assign n46707 = ~n46423 & ~n46497 ;
  assign n46708 = ~n46702 & n46707 ;
  assign n46709 = ~n46706 & n46708 ;
  assign n46710 = ~n46476 & ~n46480 ;
  assign n46713 = n46466 & n46494 ;
  assign n46714 = n46710 & ~n46713 ;
  assign n46715 = n46435 & ~n46714 ;
  assign n46716 = n46448 & n46501 ;
  assign n46711 = ~n46435 & ~n46494 ;
  assign n46712 = n46710 & n46711 ;
  assign n46717 = n46423 & ~n46499 ;
  assign n46718 = ~n46712 & n46717 ;
  assign n46719 = ~n46716 & n46718 ;
  assign n46720 = ~n46715 & n46719 ;
  assign n46721 = ~n46709 & ~n46720 ;
  assign n46723 = n46457 & ~n46485 ;
  assign n46722 = n46435 & ~n46448 ;
  assign n46724 = ~n46498 & n46722 ;
  assign n46725 = n46723 & n46724 ;
  assign n46726 = ~n46721 & ~n46725 ;
  assign n46727 = ~\u1_L1_reg[17]/NET0131  & ~n46726 ;
  assign n46728 = \u1_L1_reg[17]/NET0131  & n46726 ;
  assign n46729 = ~n46727 & ~n46728 ;
  assign n46750 = ~n46535 & n46544 ;
  assign n46751 = ~n46582 & ~n46750 ;
  assign n46752 = ~n46558 & ~n46583 ;
  assign n46753 = ~n46541 & ~n46752 ;
  assign n46754 = n46751 & ~n46753 ;
  assign n46755 = n46550 & ~n46754 ;
  assign n46749 = n46522 & n46563 ;
  assign n46738 = n46522 & n46597 ;
  assign n46739 = ~n46522 & n46557 ;
  assign n46756 = n46529 & n46541 ;
  assign n46757 = ~n46739 & ~n46756 ;
  assign n46758 = ~n46738 & n46757 ;
  assign n46759 = ~n46550 & ~n46758 ;
  assign n46760 = ~n46749 & ~n46759 ;
  assign n46761 = ~n46755 & n46760 ;
  assign n46762 = ~n46516 & ~n46761 ;
  assign n46740 = ~n46576 & ~n46739 ;
  assign n46741 = ~n46738 & n46740 ;
  assign n46742 = n46550 & ~n46741 ;
  assign n46730 = n46522 & ~n46544 ;
  assign n46731 = ~n46562 & n46730 ;
  assign n46732 = ~n46596 & ~n46731 ;
  assign n46733 = ~n46550 & ~n46732 ;
  assign n46734 = ~n46522 & n46562 ;
  assign n46735 = n46522 & n46595 ;
  assign n46736 = ~n46734 & ~n46735 ;
  assign n46737 = ~n46535 & ~n46736 ;
  assign n46743 = n46556 & ~n46737 ;
  assign n46744 = ~n46733 & n46743 ;
  assign n46745 = ~n46742 & n46744 ;
  assign n46746 = n46516 & ~n46745 ;
  assign n46747 = ~n46522 & n46550 ;
  assign n46748 = n46575 & n46747 ;
  assign n46763 = ~n46584 & ~n46748 ;
  assign n46764 = ~n46746 & n46763 ;
  assign n46765 = ~n46762 & n46764 ;
  assign n46766 = \u1_L1_reg[29]/NET0131  & ~n46765 ;
  assign n46767 = ~\u1_L1_reg[29]/NET0131  & n46765 ;
  assign n46768 = ~n46766 & ~n46767 ;
  assign n46802 = decrypt_pad & ~\u1_uk_K_r1_reg[12]/NET0131  ;
  assign n46803 = ~decrypt_pad & ~\u1_uk_K_r1_reg[20]/NET0131  ;
  assign n46804 = ~n46802 & ~n46803 ;
  assign n46805 = \u1_R1_reg[7]/NET0131  & ~n46804 ;
  assign n46806 = ~\u1_R1_reg[7]/NET0131  & n46804 ;
  assign n46807 = ~n46805 & ~n46806 ;
  assign n46788 = decrypt_pad & ~\u1_uk_K_r1_reg[27]/NET0131  ;
  assign n46789 = ~decrypt_pad & ~\u1_uk_K_r1_reg[3]/NET0131  ;
  assign n46790 = ~n46788 & ~n46789 ;
  assign n46791 = \u1_R1_reg[5]/NET0131  & ~n46790 ;
  assign n46792 = ~\u1_R1_reg[5]/NET0131  & n46790 ;
  assign n46793 = ~n46791 & ~n46792 ;
  assign n46794 = decrypt_pad & ~\u1_uk_K_r1_reg[18]/NET0131  ;
  assign n46795 = ~decrypt_pad & ~\u1_uk_K_r1_reg[26]/NET0131  ;
  assign n46796 = ~n46794 & ~n46795 ;
  assign n46797 = \u1_R1_reg[6]/NET0131  & ~n46796 ;
  assign n46798 = ~\u1_R1_reg[6]/NET0131  & n46796 ;
  assign n46799 = ~n46797 & ~n46798 ;
  assign n46839 = n46793 & ~n46799 ;
  assign n46769 = decrypt_pad & ~\u1_uk_K_r1_reg[3]/NET0131  ;
  assign n46770 = ~decrypt_pad & ~\u1_uk_K_r1_reg[11]/NET0131  ;
  assign n46771 = ~n46769 & ~n46770 ;
  assign n46772 = \u1_R1_reg[8]/NET0131  & ~n46771 ;
  assign n46773 = ~\u1_R1_reg[8]/NET0131  & n46771 ;
  assign n46774 = ~n46772 & ~n46773 ;
  assign n46775 = decrypt_pad & ~\u1_uk_K_r1_reg[48]/NET0131  ;
  assign n46776 = ~decrypt_pad & ~\u1_uk_K_r1_reg[24]/NET0131  ;
  assign n46777 = ~n46775 & ~n46776 ;
  assign n46778 = \u1_R1_reg[4]/NET0131  & ~n46777 ;
  assign n46779 = ~\u1_R1_reg[4]/NET0131  & n46777 ;
  assign n46780 = ~n46778 & ~n46779 ;
  assign n46781 = decrypt_pad & ~\u1_uk_K_r1_reg[40]/NET0131  ;
  assign n46782 = ~decrypt_pad & ~\u1_uk_K_r1_reg[48]/NET0131  ;
  assign n46783 = ~n46781 & ~n46782 ;
  assign n46784 = \u1_R1_reg[9]/NET0131  & ~n46783 ;
  assign n46785 = ~\u1_R1_reg[9]/NET0131  & n46783 ;
  assign n46786 = ~n46784 & ~n46785 ;
  assign n46787 = n46780 & n46786 ;
  assign n46800 = ~n46793 & n46799 ;
  assign n46801 = n46787 & n46800 ;
  assign n46840 = ~n46780 & ~n46786 ;
  assign n46841 = ~n46801 & ~n46840 ;
  assign n46842 = n46774 & ~n46841 ;
  assign n46809 = ~n46780 & n46786 ;
  assign n46843 = ~n46800 & n46809 ;
  assign n46844 = ~n46842 & ~n46843 ;
  assign n46845 = ~n46839 & ~n46844 ;
  assign n46846 = ~n46807 & ~n46845 ;
  assign n46847 = ~n46786 & n46800 ;
  assign n46848 = ~n46780 & n46847 ;
  assign n46811 = n46780 & n46793 ;
  assign n46849 = ~n46799 & n46811 ;
  assign n46850 = n46807 & ~n46849 ;
  assign n46851 = ~n46848 & n46850 ;
  assign n46852 = ~n46846 & ~n46851 ;
  assign n46810 = ~n46793 & n46809 ;
  assign n46812 = n46780 & ~n46786 ;
  assign n46813 = ~n46811 & ~n46812 ;
  assign n46814 = n46799 & ~n46813 ;
  assign n46815 = ~n46810 & ~n46814 ;
  assign n46816 = ~n46807 & ~n46815 ;
  assign n46817 = ~n46786 & n46793 ;
  assign n46818 = ~n46810 & ~n46817 ;
  assign n46819 = ~n46799 & ~n46818 ;
  assign n46808 = n46801 & n46807 ;
  assign n46820 = ~n46793 & ~n46807 ;
  assign n46821 = n46786 & ~n46799 ;
  assign n46822 = n46820 & n46821 ;
  assign n46823 = n46793 & n46799 ;
  assign n46824 = n46809 & n46823 ;
  assign n46825 = ~n46822 & ~n46824 ;
  assign n46826 = ~n46808 & n46825 ;
  assign n46827 = ~n46819 & n46826 ;
  assign n46828 = ~n46816 & n46827 ;
  assign n46829 = ~n46774 & ~n46828 ;
  assign n46830 = ~n46793 & n46812 ;
  assign n46831 = n46787 & n46793 ;
  assign n46832 = ~n46830 & ~n46831 ;
  assign n46833 = ~n46799 & ~n46832 ;
  assign n46834 = ~n46780 & n46799 ;
  assign n46835 = n46793 & n46807 ;
  assign n46836 = ~n46834 & n46835 ;
  assign n46837 = ~n46833 & ~n46836 ;
  assign n46838 = n46774 & ~n46837 ;
  assign n46853 = ~n46829 & ~n46838 ;
  assign n46854 = ~n46852 & n46853 ;
  assign n46855 = \u1_L1_reg[2]/NET0131  & n46854 ;
  assign n46856 = ~\u1_L1_reg[2]/NET0131  & ~n46854 ;
  assign n46857 = ~n46855 & ~n46856 ;
  assign n46861 = ~n46591 & ~n46756 ;
  assign n46862 = ~n46749 & n46861 ;
  assign n46863 = ~n46550 & ~n46862 ;
  assign n46858 = ~n46597 & ~n46734 ;
  assign n46859 = ~n46555 & n46858 ;
  assign n46860 = n46550 & ~n46859 ;
  assign n46864 = ~n46584 & ~n46860 ;
  assign n46865 = ~n46863 & n46864 ;
  assign n46866 = ~n46516 & ~n46865 ;
  assign n46874 = n46522 & n46575 ;
  assign n46878 = ~n46592 & ~n46874 ;
  assign n46875 = n46528 & ~n46542 ;
  assign n46876 = n46551 & ~n46875 ;
  assign n46877 = n46550 & n46756 ;
  assign n46879 = ~n46876 & ~n46877 ;
  assign n46880 = n46878 & n46879 ;
  assign n46881 = n46516 & ~n46880 ;
  assign n46868 = ~n46576 & ~n46596 ;
  assign n46869 = n46550 & ~n46597 ;
  assign n46870 = n46868 & n46869 ;
  assign n46867 = ~n46550 & n46751 ;
  assign n46871 = n46522 & ~n46867 ;
  assign n46872 = ~n46870 & n46871 ;
  assign n46873 = n46551 & n46595 ;
  assign n46882 = ~n46872 & ~n46873 ;
  assign n46883 = ~n46881 & n46882 ;
  assign n46884 = ~n46866 & n46883 ;
  assign n46885 = ~\u1_L1_reg[4]/NET0131  & ~n46884 ;
  assign n46886 = \u1_L1_reg[4]/NET0131  & n46884 ;
  assign n46887 = ~n46885 & ~n46886 ;
  assign n46888 = decrypt_pad & ~\u1_uk_K_r1_reg[28]/NET0131  ;
  assign n46889 = ~decrypt_pad & ~\u1_uk_K_r1_reg[38]/NET0131  ;
  assign n46890 = ~n46888 & ~n46889 ;
  assign n46891 = \u1_R1_reg[32]/NET0131  & ~n46890 ;
  assign n46892 = ~\u1_R1_reg[32]/NET0131  & n46890 ;
  assign n46893 = ~n46891 & ~n46892 ;
  assign n46894 = decrypt_pad & ~\u1_uk_K_r1_reg[37]/NET0131  ;
  assign n46895 = ~decrypt_pad & ~\u1_uk_K_r1_reg[43]/NET0131  ;
  assign n46896 = ~n46894 & ~n46895 ;
  assign n46897 = \u1_R1_reg[28]/NET0131  & ~n46896 ;
  assign n46898 = ~\u1_R1_reg[28]/NET0131  & n46896 ;
  assign n46899 = ~n46897 & ~n46898 ;
  assign n46900 = decrypt_pad & ~\u1_uk_K_r1_reg[9]/NET0131  ;
  assign n46901 = ~decrypt_pad & ~\u1_uk_K_r1_reg[15]/NET0131  ;
  assign n46902 = ~n46900 & ~n46901 ;
  assign n46903 = \u1_R1_reg[29]/NET0131  & ~n46902 ;
  assign n46904 = ~\u1_R1_reg[29]/NET0131  & n46902 ;
  assign n46905 = ~n46903 & ~n46904 ;
  assign n46951 = n46899 & ~n46905 ;
  assign n46907 = decrypt_pad & ~\u1_uk_K_r1_reg[38]/NET0131  ;
  assign n46908 = ~decrypt_pad & ~\u1_uk_K_r1_reg[16]/NET0131  ;
  assign n46909 = ~n46907 & ~n46908 ;
  assign n46910 = \u1_R1_reg[30]/NET0131  & ~n46909 ;
  assign n46911 = ~\u1_R1_reg[30]/NET0131  & n46909 ;
  assign n46912 = ~n46910 & ~n46911 ;
  assign n46913 = decrypt_pad & ~\u1_uk_K_r1_reg[49]/NET0131  ;
  assign n46914 = ~decrypt_pad & ~\u1_uk_K_r1_reg[0]/NET0131  ;
  assign n46915 = ~n46913 & ~n46914 ;
  assign n46916 = \u1_R1_reg[1]/NET0131  & ~n46915 ;
  assign n46917 = ~\u1_R1_reg[1]/NET0131  & n46915 ;
  assign n46918 = ~n46916 & ~n46917 ;
  assign n46957 = n46912 & ~n46918 ;
  assign n46958 = n46951 & n46957 ;
  assign n46923 = decrypt_pad & ~\u1_uk_K_r1_reg[22]/NET0131  ;
  assign n46924 = ~decrypt_pad & ~\u1_uk_K_r1_reg[28]/NET0131  ;
  assign n46925 = ~n46923 & ~n46924 ;
  assign n46926 = \u1_R1_reg[31]/P0001  & ~n46925 ;
  assign n46927 = ~\u1_R1_reg[31]/P0001  & n46925 ;
  assign n46928 = ~n46926 & ~n46927 ;
  assign n46940 = ~n46899 & n46918 ;
  assign n46941 = ~n46905 & n46940 ;
  assign n46959 = n46928 & ~n46941 ;
  assign n46960 = ~n46958 & n46959 ;
  assign n46961 = n46905 & n46918 ;
  assign n46930 = n46899 & ~n46912 ;
  assign n46962 = ~n46928 & ~n46930 ;
  assign n46963 = ~n46961 & n46962 ;
  assign n46964 = ~n46960 & ~n46963 ;
  assign n46933 = ~n46918 & n46930 ;
  assign n46934 = n46905 & n46933 ;
  assign n46965 = ~n46899 & ~n46918 ;
  assign n46966 = ~n46928 & n46965 ;
  assign n46967 = n46899 & n46918 ;
  assign n46968 = n46905 & n46967 ;
  assign n46969 = ~n46966 & ~n46968 ;
  assign n46970 = n46912 & ~n46969 ;
  assign n46971 = ~n46934 & ~n46970 ;
  assign n46972 = ~n46964 & n46971 ;
  assign n46973 = ~n46893 & ~n46972 ;
  assign n46931 = n46905 & ~n46918 ;
  assign n46932 = ~n46930 & ~n46931 ;
  assign n46935 = n46928 & ~n46932 ;
  assign n46936 = ~n46934 & n46935 ;
  assign n46906 = ~n46899 & n46905 ;
  assign n46919 = n46912 & n46918 ;
  assign n46920 = n46906 & n46919 ;
  assign n46921 = ~n46905 & ~n46912 ;
  assign n46922 = ~n46899 & n46921 ;
  assign n46929 = n46922 & ~n46928 ;
  assign n46937 = ~n46920 & ~n46929 ;
  assign n46938 = ~n46936 & n46937 ;
  assign n46939 = n46893 & ~n46938 ;
  assign n46943 = n46906 & n46912 ;
  assign n46944 = ~n46922 & ~n46943 ;
  assign n46945 = ~n46918 & ~n46944 ;
  assign n46942 = n46912 & n46941 ;
  assign n46946 = ~n46905 & n46918 ;
  assign n46947 = n46930 & n46946 ;
  assign n46948 = n46928 & ~n46947 ;
  assign n46949 = ~n46942 & n46948 ;
  assign n46950 = ~n46945 & n46949 ;
  assign n46952 = n46893 & n46912 ;
  assign n46953 = n46951 & n46952 ;
  assign n46954 = ~n46928 & ~n46953 ;
  assign n46955 = ~n46934 & n46954 ;
  assign n46956 = ~n46950 & ~n46955 ;
  assign n46974 = ~n46939 & ~n46956 ;
  assign n46975 = ~n46973 & n46974 ;
  assign n46976 = \u1_L1_reg[5]/NET0131  & ~n46975 ;
  assign n46977 = ~\u1_L1_reg[5]/NET0131  & n46975 ;
  assign n46978 = ~n46976 & ~n46977 ;
  assign n46979 = decrypt_pad & ~\u1_uk_K_r1_reg[4]/NET0131  ;
  assign n46980 = ~decrypt_pad & ~\u1_uk_K_r1_reg[12]/NET0131  ;
  assign n46981 = ~n46979 & ~n46980 ;
  assign n46982 = \u1_R1_reg[16]/NET0131  & ~n46981 ;
  assign n46983 = ~\u1_R1_reg[16]/NET0131  & n46981 ;
  assign n46984 = ~n46982 & ~n46983 ;
  assign n47018 = decrypt_pad & ~\u1_uk_K_r1_reg[53]/NET0131  ;
  assign n47019 = ~decrypt_pad & ~\u1_uk_K_r1_reg[4]/NET0131  ;
  assign n47020 = ~n47018 & ~n47019 ;
  assign n47021 = \u1_R1_reg[15]/NET0131  & ~n47020 ;
  assign n47022 = ~\u1_R1_reg[15]/NET0131  & n47020 ;
  assign n47023 = ~n47021 & ~n47022 ;
  assign n46991 = decrypt_pad & ~\u1_uk_K_r1_reg[19]/NET0131  ;
  assign n46992 = ~decrypt_pad & ~\u1_uk_K_r1_reg[27]/NET0131  ;
  assign n46993 = ~n46991 & ~n46992 ;
  assign n46994 = \u1_R1_reg[13]/NET0131  & ~n46993 ;
  assign n46995 = ~\u1_R1_reg[13]/NET0131  & n46993 ;
  assign n46996 = ~n46994 & ~n46995 ;
  assign n46998 = decrypt_pad & ~\u1_uk_K_r1_reg[25]/NET0131  ;
  assign n46999 = ~decrypt_pad & ~\u1_uk_K_r1_reg[33]/NET0131  ;
  assign n47000 = ~n46998 & ~n46999 ;
  assign n47001 = \u1_R1_reg[12]/NET0131  & ~n47000 ;
  assign n47002 = ~\u1_R1_reg[12]/NET0131  & n47000 ;
  assign n47003 = ~n47001 & ~n47002 ;
  assign n47005 = decrypt_pad & ~\u1_uk_K_r1_reg[41]/NET0131  ;
  assign n47006 = ~decrypt_pad & ~\u1_uk_K_r1_reg[17]/NET0131  ;
  assign n47007 = ~n47005 & ~n47006 ;
  assign n47008 = \u1_R1_reg[17]/NET0131  & ~n47007 ;
  assign n47009 = ~\u1_R1_reg[17]/NET0131  & n47007 ;
  assign n47010 = ~n47008 & ~n47009 ;
  assign n47025 = ~n47003 & ~n47010 ;
  assign n47053 = n46996 & n47025 ;
  assign n46985 = decrypt_pad & ~\u1_uk_K_r1_reg[20]/NET0131  ;
  assign n46986 = ~decrypt_pad & ~\u1_uk_K_r1_reg[53]/NET0131  ;
  assign n46987 = ~n46985 & ~n46986 ;
  assign n46988 = \u1_R1_reg[14]/NET0131  & ~n46987 ;
  assign n46989 = ~\u1_R1_reg[14]/NET0131  & n46987 ;
  assign n46990 = ~n46988 & ~n46989 ;
  assign n47054 = ~n46996 & n47010 ;
  assign n47055 = n47003 & n47054 ;
  assign n47056 = ~n46990 & n47055 ;
  assign n47057 = ~n47053 & ~n47056 ;
  assign n47058 = n47023 & ~n47057 ;
  assign n47030 = n47003 & n47010 ;
  assign n47038 = n46996 & n47030 ;
  assign n47011 = ~n47003 & n47010 ;
  assign n47039 = ~n46996 & n47011 ;
  assign n47040 = ~n47038 & ~n47039 ;
  assign n47041 = n46990 & ~n47040 ;
  assign n46997 = ~n46990 & n46996 ;
  assign n47046 = n47003 & ~n47010 ;
  assign n47060 = ~n46997 & ~n47046 ;
  assign n47059 = n46997 & ~n47011 ;
  assign n47061 = ~n47023 & ~n47059 ;
  assign n47062 = ~n47060 & n47061 ;
  assign n47063 = ~n47041 & ~n47062 ;
  assign n47064 = ~n47058 & n47063 ;
  assign n47065 = n46984 & ~n47064 ;
  assign n47012 = ~n46990 & n47011 ;
  assign n47013 = n46990 & ~n46996 ;
  assign n47014 = ~n46996 & ~n47010 ;
  assign n47015 = ~n47013 & ~n47014 ;
  assign n47016 = n47003 & ~n47015 ;
  assign n47017 = ~n47012 & ~n47016 ;
  assign n47024 = ~n47017 & n47023 ;
  assign n47026 = ~n46997 & ~n47013 ;
  assign n47027 = n47025 & n47026 ;
  assign n47031 = ~n46990 & ~n47023 ;
  assign n47032 = n47030 & n47031 ;
  assign n47004 = n46997 & n47003 ;
  assign n47028 = ~n46996 & ~n47023 ;
  assign n47029 = n47025 & n47028 ;
  assign n47033 = ~n47004 & ~n47029 ;
  assign n47034 = ~n47032 & n47033 ;
  assign n47035 = ~n47027 & n47034 ;
  assign n47036 = ~n47024 & n47035 ;
  assign n47037 = ~n46984 & ~n47036 ;
  assign n47042 = ~n46990 & ~n46996 ;
  assign n47043 = n47025 & n47042 ;
  assign n47044 = ~n47041 & ~n47043 ;
  assign n47045 = ~n47023 & ~n47044 ;
  assign n47047 = n46996 & n47023 ;
  assign n47048 = n47046 & n47047 ;
  assign n47049 = ~n46990 & n47048 ;
  assign n47050 = n46990 & n47023 ;
  assign n47051 = n46996 & ~n47003 ;
  assign n47052 = n47050 & n47051 ;
  assign n47066 = ~n47049 & ~n47052 ;
  assign n47067 = ~n47045 & n47066 ;
  assign n47068 = ~n47037 & n47067 ;
  assign n47069 = ~n47065 & n47068 ;
  assign n47070 = ~\u1_L1_reg[10]/NET0131  & ~n47069 ;
  assign n47071 = \u1_L1_reg[10]/NET0131  & n47069 ;
  assign n47072 = ~n47070 & ~n47071 ;
  assign n47083 = ~n46645 & n46675 ;
  assign n47073 = ~n46631 & n46669 ;
  assign n47074 = ~n46637 & n47073 ;
  assign n47081 = ~n46647 & ~n46667 ;
  assign n47082 = n46681 & ~n47081 ;
  assign n47086 = ~n47074 & ~n47082 ;
  assign n47087 = ~n47083 & n47086 ;
  assign n47075 = ~n46618 & n46631 ;
  assign n47076 = ~n46637 & n47075 ;
  assign n47077 = n46618 & n46656 ;
  assign n47078 = ~n47076 & ~n47077 ;
  assign n47079 = ~n46624 & ~n47078 ;
  assign n47080 = ~n46645 & n46656 ;
  assign n47084 = ~n46612 & ~n46639 ;
  assign n47085 = ~n47080 & n47084 ;
  assign n47088 = ~n47079 & n47085 ;
  assign n47089 = n47087 & n47088 ;
  assign n47092 = ~n46681 & ~n47075 ;
  assign n47091 = ~n46631 & n46645 ;
  assign n47093 = n46649 & ~n47091 ;
  assign n47094 = ~n47092 & n47093 ;
  assign n47090 = n46637 & n47073 ;
  assign n47099 = n46612 & ~n47090 ;
  assign n47100 = ~n47094 & n47099 ;
  assign n47095 = ~n46637 & ~n46684 ;
  assign n47096 = n46624 & n46631 ;
  assign n47097 = ~n46680 & ~n47096 ;
  assign n47098 = n46645 & ~n47097 ;
  assign n47101 = ~n47095 & ~n47098 ;
  assign n47102 = n47100 & n47101 ;
  assign n47103 = ~n47089 & ~n47102 ;
  assign n47104 = \u1_L1_reg[12]/NET0131  & n47103 ;
  assign n47105 = ~\u1_L1_reg[12]/NET0131  & ~n47103 ;
  assign n47106 = ~n47104 & ~n47105 ;
  assign n47111 = n46787 & ~n46793 ;
  assign n47112 = ~n46807 & ~n46847 ;
  assign n47113 = ~n47111 & n47112 ;
  assign n47116 = n46786 & n46834 ;
  assign n47114 = ~n46793 & ~n46799 ;
  assign n47115 = ~n46786 & n47114 ;
  assign n47117 = n46807 & ~n47115 ;
  assign n47118 = ~n47116 & n47117 ;
  assign n47119 = ~n47113 & ~n47118 ;
  assign n47109 = ~n46780 & n46817 ;
  assign n47110 = ~n46799 & n47109 ;
  assign n47120 = n46774 & n46825 ;
  assign n47121 = ~n47110 & n47120 ;
  assign n47122 = ~n47119 & n47121 ;
  assign n47126 = ~n46780 & ~n46820 ;
  assign n47127 = n46821 & n47126 ;
  assign n47123 = n46780 & n46807 ;
  assign n47124 = n46799 & ~n46817 ;
  assign n47125 = n47123 & n47124 ;
  assign n47128 = ~n46774 & ~n47125 ;
  assign n47129 = ~n47127 & n47128 ;
  assign n47131 = n46799 & n46810 ;
  assign n47130 = ~n46799 & n46830 ;
  assign n47132 = ~n46807 & ~n47109 ;
  assign n47133 = ~n47130 & n47132 ;
  assign n47134 = ~n47131 & n47133 ;
  assign n47135 = n47129 & n47134 ;
  assign n47136 = ~n47122 & ~n47135 ;
  assign n47107 = n46812 & n46823 ;
  assign n47108 = n46811 & n46821 ;
  assign n47137 = ~n47107 & ~n47108 ;
  assign n47138 = ~n47136 & n47137 ;
  assign n47141 = ~n46787 & ~n46840 ;
  assign n47142 = ~n46793 & ~n47141 ;
  assign n47139 = ~n46799 & n46812 ;
  assign n47140 = n46793 & n47139 ;
  assign n47143 = n46807 & ~n47140 ;
  assign n47144 = ~n47142 & n47143 ;
  assign n47145 = n47129 & n47144 ;
  assign n47146 = ~n47138 & ~n47145 ;
  assign n47147 = ~\u1_L1_reg[13]/NET0131  & ~n47146 ;
  assign n47148 = \u1_L1_reg[13]/NET0131  & n47146 ;
  assign n47149 = ~n47147 & ~n47148 ;
  assign n47169 = n26881 & n26909 ;
  assign n47150 = n26861 & ~n26886 ;
  assign n47179 = ~n26892 & n47150 ;
  assign n47180 = ~n47169 & ~n47179 ;
  assign n47181 = n26875 & ~n47180 ;
  assign n47171 = ~n26855 & ~n26875 ;
  assign n47157 = n26861 & ~n26881 ;
  assign n47172 = n26868 & n47157 ;
  assign n47173 = ~n26918 & ~n47172 ;
  assign n47174 = n47171 & ~n47173 ;
  assign n47182 = n26855 & n26904 ;
  assign n47170 = ~n26855 & n47169 ;
  assign n47175 = n26855 & ~n26875 ;
  assign n47176 = n26868 & ~n47175 ;
  assign n47177 = n26883 & ~n26915 ;
  assign n47178 = ~n47176 & n47177 ;
  assign n47183 = ~n47170 & ~n47178 ;
  assign n47184 = ~n47182 & n47183 ;
  assign n47185 = ~n47174 & n47184 ;
  assign n47186 = ~n47181 & n47185 ;
  assign n47187 = n26849 & ~n47186 ;
  assign n47156 = ~n26855 & n26904 ;
  assign n47155 = n26855 & n26909 ;
  assign n47158 = ~n26868 & n47157 ;
  assign n47159 = ~n47155 & ~n47158 ;
  assign n47160 = ~n26924 & n47159 ;
  assign n47161 = ~n47156 & n47160 ;
  assign n47162 = ~n26875 & ~n47161 ;
  assign n47151 = ~n26897 & ~n26909 ;
  assign n47152 = ~n47150 & n47151 ;
  assign n47153 = ~n26892 & ~n47152 ;
  assign n47154 = n26875 & ~n47153 ;
  assign n47163 = ~n26862 & ~n26897 ;
  assign n47164 = ~n26882 & ~n26896 ;
  assign n47165 = n47163 & n47164 ;
  assign n47166 = ~n47154 & ~n47165 ;
  assign n47167 = ~n47162 & n47166 ;
  assign n47168 = ~n26849 & ~n47167 ;
  assign n47188 = ~n26919 & ~n47170 ;
  assign n47189 = n26875 & ~n47188 ;
  assign n47190 = n26855 & n47158 ;
  assign n47191 = ~n26861 & n26903 ;
  assign n47192 = ~n47190 & ~n47191 ;
  assign n47193 = ~n26875 & ~n47192 ;
  assign n47194 = ~n47189 & ~n47193 ;
  assign n47195 = ~n47168 & n47194 ;
  assign n47196 = ~n47187 & n47195 ;
  assign n47197 = ~\u1_L1_reg[14]/NET0131  & ~n47196 ;
  assign n47198 = \u1_L1_reg[14]/NET0131  & n47196 ;
  assign n47199 = ~n47197 & ~n47198 ;
  assign n47200 = n46990 & ~n47011 ;
  assign n47201 = ~n47046 & ~n47200 ;
  assign n47202 = ~n47023 & ~n47201 ;
  assign n47203 = n47003 & n47042 ;
  assign n47204 = n47023 & ~n47054 ;
  assign n47205 = ~n47203 & n47204 ;
  assign n47206 = ~n47028 & ~n47205 ;
  assign n47207 = ~n47202 & n47206 ;
  assign n47208 = n46990 & n47046 ;
  assign n47209 = n46996 & n47208 ;
  assign n47210 = ~n47003 & n47013 ;
  assign n47211 = n46984 & ~n47210 ;
  assign n47212 = ~n47209 & n47211 ;
  assign n47213 = ~n47207 & n47212 ;
  assign n47214 = ~n46990 & n47046 ;
  assign n47215 = ~n47023 & ~n47055 ;
  assign n47216 = ~n47214 & n47215 ;
  assign n47218 = ~n46996 & n47208 ;
  assign n47217 = ~n46990 & n47025 ;
  assign n47219 = n47023 & ~n47217 ;
  assign n47220 = ~n47218 & n47219 ;
  assign n47221 = ~n47216 & ~n47220 ;
  assign n47222 = n46990 & n47030 ;
  assign n47223 = ~n47012 & ~n47222 ;
  assign n47224 = n46996 & ~n47223 ;
  assign n47225 = n47004 & ~n47010 ;
  assign n47226 = ~n46984 & ~n47225 ;
  assign n47227 = ~n47224 & n47226 ;
  assign n47228 = ~n47221 & n47227 ;
  assign n47229 = ~n47213 & ~n47228 ;
  assign n47231 = n47040 & ~n47053 ;
  assign n47232 = n47050 & ~n47231 ;
  assign n47230 = ~n47023 & n47209 ;
  assign n47233 = n46990 & n47029 ;
  assign n47234 = ~n47230 & ~n47233 ;
  assign n47235 = ~n47232 & n47234 ;
  assign n47236 = ~n47229 & n47235 ;
  assign n47237 = ~\u1_L1_reg[1]/NET0131  & ~n47236 ;
  assign n47238 = \u1_L1_reg[1]/NET0131  & n47236 ;
  assign n47239 = ~n47237 & ~n47238 ;
  assign n47261 = ~n46448 & ~n46698 ;
  assign n47262 = ~n46442 & n46469 ;
  assign n47263 = ~n47261 & ~n47262 ;
  assign n47264 = n46423 & ~n47263 ;
  assign n47260 = n46466 & n46467 ;
  assign n47265 = ~n46716 & ~n47260 ;
  assign n47266 = ~n47264 & n47265 ;
  assign n47267 = ~n46435 & ~n47266 ;
  assign n47240 = ~n46463 & ~n46468 ;
  assign n47241 = n46435 & ~n47240 ;
  assign n47242 = ~n46500 & ~n47241 ;
  assign n47243 = ~n46436 & ~n47242 ;
  assign n47244 = n46435 & ~n46494 ;
  assign n47245 = n46458 & n47244 ;
  assign n47246 = n46477 & n46493 ;
  assign n47247 = n46423 & ~n46713 ;
  assign n47248 = ~n47246 & n47247 ;
  assign n47249 = ~n47245 & n47248 ;
  assign n47255 = ~n46423 & ~n46486 ;
  assign n47256 = ~n46499 & n47255 ;
  assign n47250 = ~n46462 & ~n46498 ;
  assign n47251 = n46722 & ~n47250 ;
  assign n47252 = ~n46457 & ~n46498 ;
  assign n47253 = ~n46435 & n46448 ;
  assign n47254 = ~n47252 & n47253 ;
  assign n47257 = ~n47251 & ~n47254 ;
  assign n47258 = n47256 & n47257 ;
  assign n47259 = ~n47249 & ~n47258 ;
  assign n47268 = ~n47243 & ~n47259 ;
  assign n47269 = ~n47267 & n47268 ;
  assign n47270 = \u1_L1_reg[23]/NET0131  & ~n47269 ;
  assign n47271 = ~\u1_L1_reg[23]/NET0131  & n47269 ;
  assign n47272 = ~n47270 & ~n47271 ;
  assign n47273 = n47011 & n47042 ;
  assign n47274 = ~n47222 & ~n47273 ;
  assign n47275 = ~n47023 & ~n47274 ;
  assign n47277 = ~n47208 & ~n47217 ;
  assign n47278 = n46996 & ~n47277 ;
  assign n47276 = n46990 & n47011 ;
  assign n47279 = ~n46996 & n47025 ;
  assign n47280 = ~n47276 & ~n47279 ;
  assign n47281 = ~n47278 & n47280 ;
  assign n47282 = ~n47028 & ~n47281 ;
  assign n47283 = ~n47275 & ~n47282 ;
  assign n47284 = n46984 & ~n47283 ;
  assign n47291 = n47047 & ~n47201 ;
  assign n47292 = n46997 & n47011 ;
  assign n47293 = ~n47203 & ~n47292 ;
  assign n47294 = ~n47291 & n47293 ;
  assign n47295 = ~n46984 & ~n47294 ;
  assign n47286 = ~n47014 & ~n47210 ;
  assign n47287 = ~n46984 & ~n47286 ;
  assign n47288 = ~n47046 & n47059 ;
  assign n47289 = ~n47287 & ~n47288 ;
  assign n47290 = ~n47023 & ~n47289 ;
  assign n47285 = n47028 & n47214 ;
  assign n47296 = n46997 & ~n47003 ;
  assign n47297 = ~n47203 & ~n47296 ;
  assign n47298 = n47010 & n47023 ;
  assign n47299 = ~n47297 & n47298 ;
  assign n47300 = ~n47285 & ~n47299 ;
  assign n47301 = ~n47290 & n47300 ;
  assign n47302 = ~n47295 & n47301 ;
  assign n47303 = ~n47284 & n47302 ;
  assign n47304 = ~\u1_L1_reg[26]/NET0131  & ~n47303 ;
  assign n47305 = \u1_L1_reg[26]/NET0131  & n47303 ;
  assign n47306 = ~n47304 & ~n47305 ;
  assign n47325 = n46799 & n47109 ;
  assign n47326 = n46832 & ~n47325 ;
  assign n47327 = n46807 & ~n47326 ;
  assign n47323 = ~n47111 & ~n47123 ;
  assign n47324 = ~n46799 & ~n47323 ;
  assign n47310 = n46793 & n46809 ;
  assign n47311 = ~n46799 & n46840 ;
  assign n47312 = ~n47310 & ~n47311 ;
  assign n47322 = ~n46807 & ~n47312 ;
  assign n47328 = ~n47131 & ~n47322 ;
  assign n47329 = ~n47324 & n47328 ;
  assign n47330 = ~n47327 & n47329 ;
  assign n47331 = n46774 & ~n47330 ;
  assign n47307 = ~n46793 & n46834 ;
  assign n47308 = ~n47107 & ~n47307 ;
  assign n47309 = ~n46807 & ~n47308 ;
  assign n47313 = n46807 & n47312 ;
  assign n47314 = ~n46807 & ~n46811 ;
  assign n47315 = ~n46810 & n47314 ;
  assign n47316 = ~n47139 & n47315 ;
  assign n47317 = ~n47313 & ~n47316 ;
  assign n47318 = n46800 & ~n47141 ;
  assign n47319 = ~n47107 & ~n47318 ;
  assign n47320 = ~n47317 & n47319 ;
  assign n47321 = ~n46774 & ~n47320 ;
  assign n47332 = ~n47309 & ~n47321 ;
  assign n47333 = ~n47331 & n47332 ;
  assign n47334 = ~\u1_L1_reg[28]/NET0131  & ~n47333 ;
  assign n47335 = \u1_L1_reg[28]/NET0131  & n47333 ;
  assign n47336 = ~n47334 & ~n47335 ;
  assign n47350 = ~n26884 & ~n47156 ;
  assign n47351 = n26875 & ~n47350 ;
  assign n47352 = ~n26915 & n47157 ;
  assign n47353 = ~n26893 & ~n47352 ;
  assign n47354 = ~n26875 & ~n47353 ;
  assign n47355 = ~n26892 & n26920 ;
  assign n47356 = ~n47354 & n47355 ;
  assign n47357 = ~n47351 & n47356 ;
  assign n47358 = ~n26849 & ~n47357 ;
  assign n47337 = ~n26855 & n26918 ;
  assign n47338 = ~n26893 & ~n47337 ;
  assign n47339 = n26875 & ~n47338 ;
  assign n47340 = n26881 & n47171 ;
  assign n47341 = n47192 & ~n47340 ;
  assign n47342 = ~n47339 & n47341 ;
  assign n47343 = n26849 & ~n47342 ;
  assign n47344 = ~n26875 & ~n47182 ;
  assign n47345 = n26875 & ~n47190 ;
  assign n47346 = n26861 & n26892 ;
  assign n47347 = ~n47155 & ~n47346 ;
  assign n47348 = n47345 & n47347 ;
  assign n47349 = ~n47344 & ~n47348 ;
  assign n47359 = ~n47343 & ~n47349 ;
  assign n47360 = ~n47358 & n47359 ;
  assign n47361 = ~\u1_L1_reg[8]/NET0131  & ~n47360 ;
  assign n47362 = \u1_L1_reg[8]/NET0131  & n47360 ;
  assign n47363 = ~n47361 & ~n47362 ;
  assign n47364 = ~n46905 & n46933 ;
  assign n47365 = ~n46906 & ~n46951 ;
  assign n47366 = ~n46965 & n47365 ;
  assign n47367 = n46905 & ~n46912 ;
  assign n47368 = ~n46918 & n47367 ;
  assign n47369 = ~n47366 & ~n47368 ;
  assign n47370 = n46928 & ~n47369 ;
  assign n47371 = ~n47364 & ~n47370 ;
  assign n47372 = ~n46893 & ~n47371 ;
  assign n47376 = ~n46918 & n46943 ;
  assign n47373 = n46912 & ~n46928 ;
  assign n47374 = n46946 & n47373 ;
  assign n47375 = n46919 & n46951 ;
  assign n47380 = ~n47374 & ~n47375 ;
  assign n47377 = ~n46905 & n46928 ;
  assign n47378 = n46965 & n47377 ;
  assign n47379 = n46905 & n46930 ;
  assign n47381 = ~n47378 & ~n47379 ;
  assign n47382 = n47380 & n47381 ;
  assign n47383 = ~n47376 & n47382 ;
  assign n47384 = n46893 & ~n47383 ;
  assign n47385 = n46918 & ~n46944 ;
  assign n47386 = n46928 & ~n47385 ;
  assign n47388 = n46893 & ~n46912 ;
  assign n47389 = n46951 & ~n47388 ;
  assign n47387 = n46940 & n47367 ;
  assign n47390 = ~n46928 & ~n47387 ;
  assign n47391 = ~n47389 & n47390 ;
  assign n47392 = ~n46945 & n47391 ;
  assign n47393 = ~n47386 & ~n47392 ;
  assign n47394 = ~n47384 & ~n47393 ;
  assign n47395 = ~n47372 & n47394 ;
  assign n47396 = \u1_L1_reg[15]/P0001  & n47395 ;
  assign n47397 = ~\u1_L1_reg[15]/P0001  & ~n47395 ;
  assign n47398 = ~n47396 & ~n47397 ;
  assign n47403 = n46940 & n47373 ;
  assign n47402 = n46921 & n46965 ;
  assign n47411 = ~n46958 & ~n47402 ;
  assign n47412 = ~n47403 & n47411 ;
  assign n47404 = n46905 & n46966 ;
  assign n47410 = ~n46893 & ~n46943 ;
  assign n47413 = ~n47404 & n47410 ;
  assign n47405 = n46918 & n46930 ;
  assign n47406 = ~n47377 & n47405 ;
  assign n47407 = ~n46921 & ~n46961 ;
  assign n47408 = n46899 & n46928 ;
  assign n47409 = n47407 & n47408 ;
  assign n47414 = ~n47406 & ~n47409 ;
  assign n47415 = n47413 & n47414 ;
  assign n47416 = n47412 & n47415 ;
  assign n47420 = n46905 & ~n46930 ;
  assign n47421 = ~n46965 & n47420 ;
  assign n47417 = n46918 & n46921 ;
  assign n47422 = n46928 & ~n47417 ;
  assign n47423 = ~n47421 & n47422 ;
  assign n47424 = ~n46928 & ~n46933 ;
  assign n47425 = ~n47375 & n47424 ;
  assign n47426 = ~n47423 & ~n47425 ;
  assign n47418 = ~n46957 & ~n47417 ;
  assign n47419 = n47365 & ~n47418 ;
  assign n47427 = n46893 & ~n47419 ;
  assign n47428 = ~n47426 & n47427 ;
  assign n47429 = ~n47416 & ~n47428 ;
  assign n47399 = ~n46928 & n46930 ;
  assign n47400 = n46961 & n47399 ;
  assign n47401 = n46922 & n46928 ;
  assign n47430 = ~n47400 & ~n47401 ;
  assign n47431 = ~n47429 & n47430 ;
  assign n47432 = ~\u1_L1_reg[21]/NET0131  & ~n47431 ;
  assign n47433 = \u1_L1_reg[21]/NET0131  & n47431 ;
  assign n47434 = ~n47432 & ~n47433 ;
  assign n47444 = ~n46899 & n47368 ;
  assign n47445 = ~n46968 & ~n47444 ;
  assign n47446 = n46928 & ~n47445 ;
  assign n47447 = ~n46899 & n47407 ;
  assign n47448 = n46899 & ~n46931 ;
  assign n47449 = ~n46928 & ~n47448 ;
  assign n47450 = ~n47447 & n47449 ;
  assign n47451 = ~n46920 & ~n46958 ;
  assign n47452 = ~n47417 & n47451 ;
  assign n47453 = ~n47450 & n47452 ;
  assign n47454 = ~n47446 & n47453 ;
  assign n47455 = n46893 & ~n47454 ;
  assign n47437 = n46928 & ~n46943 ;
  assign n47436 = n46918 & ~n47367 ;
  assign n47438 = ~n47368 & ~n47436 ;
  assign n47439 = n47437 & n47438 ;
  assign n47435 = n46967 & n47373 ;
  assign n47440 = ~n46942 & ~n47435 ;
  assign n47441 = ~n47404 & n47440 ;
  assign n47442 = ~n47439 & n47441 ;
  assign n47443 = ~n46893 & ~n47442 ;
  assign n47456 = n46957 & n47377 ;
  assign n47457 = ~n46934 & ~n46947 ;
  assign n47458 = ~n47376 & n47457 ;
  assign n47459 = ~n46928 & ~n47458 ;
  assign n47460 = ~n47456 & ~n47459 ;
  assign n47461 = ~n47443 & n47460 ;
  assign n47462 = ~n47455 & n47461 ;
  assign n47463 = ~\u1_L1_reg[27]/NET0131  & ~n47462 ;
  assign n47464 = \u1_L1_reg[27]/NET0131  & n47462 ;
  assign n47465 = ~n47463 & ~n47464 ;
  assign n47477 = n46656 & n46669 ;
  assign n47478 = ~n46637 & n47092 ;
  assign n47479 = ~n46666 & ~n46683 ;
  assign n47480 = ~n47478 & ~n47479 ;
  assign n47481 = ~n46645 & ~n47073 ;
  assign n47482 = ~n47480 & n47481 ;
  assign n47484 = ~n46667 & ~n47075 ;
  assign n47485 = n46675 & n47484 ;
  assign n47483 = n46637 & n47075 ;
  assign n47486 = n46645 & ~n47483 ;
  assign n47487 = ~n47485 & n47486 ;
  assign n47488 = ~n47482 & ~n47487 ;
  assign n47489 = ~n47477 & ~n47488 ;
  assign n47490 = n46612 & ~n47489 ;
  assign n47466 = n46624 & ~n47078 ;
  assign n47470 = ~n46676 & ~n47466 ;
  assign n47467 = ~n47076 & n47083 ;
  assign n47468 = ~n46683 & ~n47076 ;
  assign n47469 = n46645 & ~n47468 ;
  assign n47471 = ~n47467 & ~n47469 ;
  assign n47472 = n47470 & n47471 ;
  assign n47473 = ~n46612 & ~n47472 ;
  assign n47474 = n46645 & n46679 ;
  assign n47475 = n46664 & ~n47075 ;
  assign n47476 = n46657 & n47475 ;
  assign n47491 = ~n47474 & ~n47476 ;
  assign n47492 = ~n47473 & n47491 ;
  assign n47493 = ~n47490 & n47492 ;
  assign n47494 = \u1_L1_reg[32]/NET0131  & n47493 ;
  assign n47495 = ~\u1_L1_reg[32]/NET0131  & ~n47493 ;
  assign n47496 = ~n47494 & ~n47495 ;
  assign n47514 = ~n26862 & n26881 ;
  assign n47513 = ~n26881 & ~n26909 ;
  assign n47515 = n26875 & ~n47513 ;
  assign n47516 = ~n47514 & n47515 ;
  assign n47512 = ~n26875 & n47172 ;
  assign n47517 = ~n26924 & ~n47182 ;
  assign n47518 = ~n47512 & n47517 ;
  assign n47519 = ~n47516 & n47518 ;
  assign n47520 = n26849 & ~n47519 ;
  assign n47501 = ~n26893 & ~n47163 ;
  assign n47502 = ~n26875 & ~n47501 ;
  assign n47497 = ~n26897 & n26915 ;
  assign n47498 = n26862 & ~n26881 ;
  assign n47499 = ~n47169 & ~n47498 ;
  assign n47500 = n26875 & ~n47499 ;
  assign n47503 = ~n47497 & ~n47500 ;
  assign n47504 = ~n47502 & n47503 ;
  assign n47505 = ~n26849 & ~n47504 ;
  assign n47506 = ~n47156 & n47345 ;
  assign n47507 = n26883 & n26915 ;
  assign n47508 = ~n26875 & ~n47507 ;
  assign n47509 = ~n47170 & n47508 ;
  assign n47510 = ~n47337 & n47509 ;
  assign n47511 = ~n47506 & ~n47510 ;
  assign n47521 = ~n47505 & ~n47511 ;
  assign n47522 = ~n47520 & n47521 ;
  assign n47523 = ~\u1_L1_reg[3]/NET0131  & ~n47522 ;
  assign n47524 = \u1_L1_reg[3]/NET0131  & n47522 ;
  assign n47525 = ~n47523 & ~n47524 ;
  assign n47532 = decrypt_pad & ~\u1_uk_K_r1_reg[55]/NET0131  ;
  assign n47533 = ~decrypt_pad & ~\u1_uk_K_r1_reg[6]/NET0131  ;
  assign n47534 = ~n47532 & ~n47533 ;
  assign n47535 = \u1_R1_reg[11]/NET0131  & ~n47534 ;
  assign n47536 = ~\u1_R1_reg[11]/NET0131  & n47534 ;
  assign n47537 = ~n47535 & ~n47536 ;
  assign n47526 = decrypt_pad & ~\u1_uk_K_r1_reg[13]/NET0131  ;
  assign n47527 = ~decrypt_pad & ~\u1_uk_K_r1_reg[46]/NET0131  ;
  assign n47528 = ~n47526 & ~n47527 ;
  assign n47529 = \u1_R1_reg[12]/NET0131  & ~n47528 ;
  assign n47530 = ~\u1_R1_reg[12]/NET0131  & n47528 ;
  assign n47531 = ~n47529 & ~n47530 ;
  assign n47538 = decrypt_pad & ~\u1_uk_K_r1_reg[26]/NET0131  ;
  assign n47539 = ~decrypt_pad & ~\u1_uk_K_r1_reg[34]/NET0131  ;
  assign n47540 = ~n47538 & ~n47539 ;
  assign n47541 = \u1_R1_reg[13]/NET0131  & ~n47540 ;
  assign n47542 = ~\u1_R1_reg[13]/NET0131  & n47540 ;
  assign n47543 = ~n47541 & ~n47542 ;
  assign n47551 = decrypt_pad & ~\u1_uk_K_r1_reg[46]/NET0131  ;
  assign n47552 = ~decrypt_pad & ~\u1_uk_K_r1_reg[54]/NET0131  ;
  assign n47553 = ~n47551 & ~n47552 ;
  assign n47554 = \u1_R1_reg[9]/NET0131  & ~n47553 ;
  assign n47555 = ~\u1_R1_reg[9]/NET0131  & n47553 ;
  assign n47556 = ~n47554 & ~n47555 ;
  assign n47596 = n47543 & ~n47556 ;
  assign n47544 = decrypt_pad & ~\u1_uk_K_r1_reg[17]/NET0131  ;
  assign n47545 = ~decrypt_pad & ~\u1_uk_K_r1_reg[25]/NET0131  ;
  assign n47546 = ~n47544 & ~n47545 ;
  assign n47547 = \u1_R1_reg[8]/NET0131  & ~n47546 ;
  assign n47548 = ~\u1_R1_reg[8]/NET0131  & n47546 ;
  assign n47549 = ~n47547 & ~n47548 ;
  assign n47576 = ~n47543 & n47556 ;
  assign n47577 = n47549 & n47576 ;
  assign n47550 = n47543 & ~n47549 ;
  assign n47558 = decrypt_pad & ~\u1_uk_K_r1_reg[54]/NET0131  ;
  assign n47559 = ~decrypt_pad & ~\u1_uk_K_r1_reg[5]/NET0131  ;
  assign n47560 = ~n47558 & ~n47559 ;
  assign n47561 = \u1_R1_reg[10]/NET0131  & ~n47560 ;
  assign n47562 = ~\u1_R1_reg[10]/NET0131  & n47560 ;
  assign n47563 = ~n47561 & ~n47562 ;
  assign n47598 = n47550 & n47563 ;
  assign n47599 = ~n47577 & ~n47598 ;
  assign n47600 = ~n47596 & n47599 ;
  assign n47601 = n47531 & ~n47600 ;
  assign n47597 = n47563 & n47596 ;
  assign n47568 = ~n47543 & ~n47549 ;
  assign n47602 = ~n47563 & n47568 ;
  assign n47603 = ~n47556 & n47602 ;
  assign n47604 = ~n47597 & ~n47603 ;
  assign n47605 = ~n47601 & n47604 ;
  assign n47606 = n47537 & ~n47605 ;
  assign n47569 = n47543 & n47549 ;
  assign n47570 = ~n47568 & ~n47569 ;
  assign n47567 = ~n47556 & ~n47563 ;
  assign n47573 = n47537 & ~n47549 ;
  assign n47579 = n47567 & ~n47573 ;
  assign n47580 = n47570 & n47579 ;
  assign n47574 = n47556 & ~n47563 ;
  assign n47575 = n47573 & n47574 ;
  assign n47578 = n47563 & n47577 ;
  assign n47581 = ~n47575 & ~n47578 ;
  assign n47582 = ~n47580 & n47581 ;
  assign n47557 = n47550 & n47556 ;
  assign n47564 = n47557 & n47563 ;
  assign n47565 = ~n47537 & n47564 ;
  assign n47566 = n47556 & n47563 ;
  assign n47571 = ~n47567 & ~n47570 ;
  assign n47572 = ~n47566 & n47571 ;
  assign n47583 = ~n47565 & ~n47572 ;
  assign n47584 = n47582 & n47583 ;
  assign n47585 = ~n47531 & ~n47584 ;
  assign n47586 = n47531 & n47566 ;
  assign n47587 = n47568 & n47586 ;
  assign n47588 = n47543 & n47574 ;
  assign n47589 = n47549 & ~n47556 ;
  assign n47590 = ~n47543 & n47589 ;
  assign n47591 = n47556 & n47569 ;
  assign n47592 = ~n47590 & ~n47591 ;
  assign n47593 = ~n47588 & n47592 ;
  assign n47594 = n47531 & ~n47537 ;
  assign n47595 = ~n47593 & n47594 ;
  assign n47607 = ~n47587 & ~n47595 ;
  assign n47608 = ~n47585 & n47607 ;
  assign n47609 = ~n47606 & n47608 ;
  assign n47610 = ~\u1_L1_reg[6]/NET0131  & ~n47609 ;
  assign n47611 = \u1_L1_reg[6]/NET0131  & n47609 ;
  assign n47612 = ~n47610 & ~n47611 ;
  assign n47616 = ~n46625 & n47478 ;
  assign n47617 = n46645 & ~n47616 ;
  assign n47618 = ~n46631 & ~n46668 ;
  assign n47613 = n46624 & ~n47092 ;
  assign n47619 = ~n46645 & ~n47483 ;
  assign n47620 = ~n47613 & n47619 ;
  assign n47621 = ~n47618 & n47620 ;
  assign n47622 = ~n47617 & ~n47621 ;
  assign n47614 = ~n46683 & ~n47613 ;
  assign n47615 = n46637 & ~n47614 ;
  assign n47623 = n46612 & ~n47615 ;
  assign n47624 = ~n47622 & n47623 ;
  assign n47625 = n46667 & ~n47092 ;
  assign n47626 = n46645 & ~n46683 ;
  assign n47627 = ~n47478 & n47626 ;
  assign n47628 = ~n47625 & n47627 ;
  assign n47629 = ~n46612 & ~n47628 ;
  assign n47630 = ~n47624 & ~n47629 ;
  assign n47631 = ~n46645 & n47615 ;
  assign n47632 = ~n46645 & n47616 ;
  assign n47633 = ~n46639 & ~n47632 ;
  assign n47634 = n46612 & ~n46645 ;
  assign n47635 = ~n47633 & ~n47634 ;
  assign n47636 = ~n47631 & ~n47635 ;
  assign n47637 = ~n47630 & n47636 ;
  assign n47638 = ~\u1_L1_reg[7]/NET0131  & ~n47637 ;
  assign n47639 = \u1_L1_reg[7]/NET0131  & n47637 ;
  assign n47640 = ~n47638 & ~n47639 ;
  assign n47646 = ~n46463 & ~n46466 ;
  assign n47647 = ~n46700 & n47646 ;
  assign n47648 = n46435 & ~n47647 ;
  assign n47643 = n46429 & n46703 ;
  assign n47641 = ~n46449 & n46698 ;
  assign n47642 = ~n46435 & n47641 ;
  assign n47644 = ~n46429 & n46457 ;
  assign n47645 = n46449 & n47644 ;
  assign n47649 = ~n47642 & ~n47645 ;
  assign n47650 = ~n47643 & n47649 ;
  assign n47651 = ~n47648 & n47650 ;
  assign n47652 = ~n46423 & ~n47651 ;
  assign n47653 = n46480 & n46498 ;
  assign n47654 = ~n47645 & ~n47653 ;
  assign n47655 = ~n46435 & ~n47654 ;
  assign n47657 = n46429 & ~n46458 ;
  assign n47658 = ~n46703 & n47657 ;
  assign n47656 = n46483 & n47641 ;
  assign n47659 = ~n46716 & ~n47656 ;
  assign n47660 = ~n47658 & n47659 ;
  assign n47661 = n46423 & ~n47660 ;
  assign n47662 = ~n47655 & ~n47661 ;
  assign n47663 = ~n47652 & n47662 ;
  assign n47664 = ~\u1_L1_reg[9]/NET0131  & ~n47663 ;
  assign n47665 = \u1_L1_reg[9]/NET0131  & n47663 ;
  assign n47666 = ~n47664 & ~n47665 ;
  assign n47667 = n47550 & ~n47556 ;
  assign n47684 = n47573 & n47576 ;
  assign n47685 = ~n47667 & ~n47684 ;
  assign n47686 = n47592 & n47685 ;
  assign n47687 = ~n47563 & ~n47686 ;
  assign n47678 = n47563 & n47568 ;
  assign n47688 = n47549 & ~n47563 ;
  assign n47689 = ~n47543 & n47688 ;
  assign n47690 = ~n47678 & ~n47689 ;
  assign n47691 = ~n47537 & ~n47690 ;
  assign n47692 = ~n47564 & ~n47691 ;
  assign n47693 = ~n47687 & n47692 ;
  assign n47694 = n47531 & ~n47693 ;
  assign n47668 = ~n47591 & ~n47602 ;
  assign n47669 = ~n47667 & n47668 ;
  assign n47670 = ~n47537 & ~n47669 ;
  assign n47671 = ~n47556 & ~n47569 ;
  assign n47672 = n47537 & ~n47568 ;
  assign n47673 = ~n47591 & n47672 ;
  assign n47674 = ~n47671 & n47673 ;
  assign n47675 = ~n47603 & ~n47674 ;
  assign n47676 = ~n47670 & n47675 ;
  assign n47677 = ~n47531 & ~n47676 ;
  assign n47679 = ~n47556 & n47678 ;
  assign n47680 = ~n47578 & ~n47679 ;
  assign n47681 = n47537 & ~n47680 ;
  assign n47682 = ~n47537 & n47563 ;
  assign n47683 = n47589 & n47682 ;
  assign n47695 = ~n47681 & ~n47683 ;
  assign n47696 = ~n47677 & n47695 ;
  assign n47697 = ~n47694 & n47696 ;
  assign n47698 = ~\u1_L1_reg[16]/NET0131  & ~n47697 ;
  assign n47699 = \u1_L1_reg[16]/NET0131  & n47697 ;
  assign n47700 = ~n47698 & ~n47699 ;
  assign n47704 = n46807 & ~n46818 ;
  assign n47701 = n46780 & n46821 ;
  assign n47702 = ~n46830 & ~n47701 ;
  assign n47703 = ~n46807 & ~n47702 ;
  assign n47705 = n46774 & ~n46848 ;
  assign n47706 = ~n47703 & n47705 ;
  assign n47707 = ~n47704 & n47706 ;
  assign n47709 = ~n46807 & n46823 ;
  assign n47710 = ~n47114 & ~n47709 ;
  assign n47711 = ~n46780 & ~n47710 ;
  assign n47708 = n46807 & n46831 ;
  assign n47712 = ~n46774 & ~n46801 ;
  assign n47713 = ~n47107 & ~n47115 ;
  assign n47714 = n47712 & n47713 ;
  assign n47715 = ~n47708 & n47714 ;
  assign n47716 = ~n47711 & n47715 ;
  assign n47717 = ~n47707 & ~n47716 ;
  assign n47718 = ~n46807 & n47310 ;
  assign n47719 = n46787 & n46799 ;
  assign n47720 = ~n47110 & ~n47719 ;
  assign n47721 = n46807 & ~n47720 ;
  assign n47722 = ~n47718 & ~n47721 ;
  assign n47723 = ~n47717 & n47722 ;
  assign n47724 = \u1_L1_reg[18]/NET0131  & n47723 ;
  assign n47725 = ~\u1_L1_reg[18]/NET0131  & ~n47723 ;
  assign n47726 = ~n47724 & ~n47725 ;
  assign n47743 = ~n47537 & n47571 ;
  assign n47737 = n47549 & n47566 ;
  assign n47738 = ~n47598 & ~n47737 ;
  assign n47739 = n47537 & ~n47738 ;
  assign n47740 = n47537 & ~n47563 ;
  assign n47741 = ~n47550 & ~n47556 ;
  assign n47742 = n47740 & n47741 ;
  assign n47744 = ~n47580 & ~n47742 ;
  assign n47745 = ~n47739 & n47744 ;
  assign n47746 = ~n47743 & n47745 ;
  assign n47747 = n47531 & ~n47746 ;
  assign n47727 = n47550 & ~n47563 ;
  assign n47728 = ~n47678 & ~n47727 ;
  assign n47729 = n47556 & n47568 ;
  assign n47730 = n47563 & n47589 ;
  assign n47731 = ~n47729 & ~n47730 ;
  assign n47732 = n47728 & n47731 ;
  assign n47733 = n47537 & ~n47732 ;
  assign n47734 = n47563 & n47590 ;
  assign n47735 = ~n47733 & ~n47734 ;
  assign n47736 = ~n47531 & ~n47735 ;
  assign n47751 = n47567 & ~n47570 ;
  assign n47752 = n47599 & ~n47751 ;
  assign n47753 = ~n47531 & ~n47537 ;
  assign n47754 = ~n47752 & n47753 ;
  assign n47748 = n47591 & n47682 ;
  assign n47749 = ~n47557 & ~n47590 ;
  assign n47750 = n47740 & ~n47749 ;
  assign n47755 = ~n47748 & ~n47750 ;
  assign n47756 = ~n47754 & n47755 ;
  assign n47757 = ~n47736 & n47756 ;
  assign n47758 = ~n47747 & n47757 ;
  assign n47759 = ~\u1_L1_reg[24]/NET0131  & ~n47758 ;
  assign n47760 = \u1_L1_reg[24]/NET0131  & n47758 ;
  assign n47761 = ~n47759 & ~n47760 ;
  assign n47767 = n47563 & n47667 ;
  assign n47771 = ~n47531 & ~n47751 ;
  assign n47772 = ~n47767 & n47771 ;
  assign n47762 = n47549 & n47563 ;
  assign n47763 = ~n47576 & n47762 ;
  assign n47764 = ~n47543 & n47574 ;
  assign n47765 = ~n47763 & ~n47764 ;
  assign n47766 = n47537 & ~n47765 ;
  assign n47768 = ~n47576 & n47688 ;
  assign n47769 = ~n47557 & ~n47768 ;
  assign n47770 = ~n47537 & ~n47769 ;
  assign n47773 = ~n47766 & ~n47770 ;
  assign n47774 = n47772 & n47773 ;
  assign n47777 = ~n47563 & n47590 ;
  assign n47778 = n47728 & ~n47777 ;
  assign n47779 = n47537 & ~n47778 ;
  assign n47775 = ~n47729 & ~n47762 ;
  assign n47776 = ~n47537 & ~n47775 ;
  assign n47780 = n47531 & ~n47776 ;
  assign n47781 = ~n47779 & n47780 ;
  assign n47782 = ~n47774 & ~n47781 ;
  assign n47785 = n47537 & n47596 ;
  assign n47786 = n47762 & n47785 ;
  assign n47783 = ~n47569 & n47586 ;
  assign n47784 = n47576 & n47682 ;
  assign n47787 = ~n47783 & ~n47784 ;
  assign n47788 = ~n47786 & n47787 ;
  assign n47789 = ~n47782 & n47788 ;
  assign n47790 = \u1_L1_reg[30]/NET0131  & ~n47789 ;
  assign n47791 = ~\u1_L1_reg[30]/NET0131  & n47789 ;
  assign n47792 = ~n47790 & ~n47791 ;
  assign n47829 = decrypt_pad & ~\u1_uk_K_r0_reg[7]/NET0131  ;
  assign n47830 = ~decrypt_pad & ~\u1_uk_K_r0_reg[45]/NET0131  ;
  assign n47831 = ~n47829 & ~n47830 ;
  assign n47832 = \u1_R0_reg[27]/NET0131  & ~n47831 ;
  assign n47833 = ~\u1_R0_reg[27]/NET0131  & n47831 ;
  assign n47834 = ~n47832 & ~n47833 ;
  assign n47812 = decrypt_pad & ~\u1_uk_K_r0_reg[9]/NET0131  ;
  assign n47813 = ~decrypt_pad & ~\u1_uk_K_r0_reg[43]/NET0131  ;
  assign n47814 = ~n47812 & ~n47813 ;
  assign n47815 = \u1_R0_reg[24]/NET0131  & ~n47814 ;
  assign n47816 = ~\u1_R0_reg[24]/NET0131  & n47814 ;
  assign n47817 = ~n47815 & ~n47816 ;
  assign n47799 = decrypt_pad & ~\u1_uk_K_r0_reg[45]/NET0131  ;
  assign n47800 = ~decrypt_pad & ~\u1_uk_K_r0_reg[51]/NET0131  ;
  assign n47801 = ~n47799 & ~n47800 ;
  assign n47802 = \u1_R0_reg[29]/NET0131  & ~n47801 ;
  assign n47803 = ~\u1_R0_reg[29]/NET0131  & n47801 ;
  assign n47804 = ~n47802 & ~n47803 ;
  assign n47805 = decrypt_pad & ~\u1_uk_K_r0_reg[44]/NET0131  ;
  assign n47806 = ~decrypt_pad & ~\u1_uk_K_r0_reg[23]/NET0131  ;
  assign n47807 = ~n47805 & ~n47806 ;
  assign n47808 = \u1_R0_reg[25]/NET0131  & ~n47807 ;
  assign n47809 = ~\u1_R0_reg[25]/NET0131  & n47807 ;
  assign n47810 = ~n47808 & ~n47809 ;
  assign n47871 = ~n47804 & ~n47810 ;
  assign n47793 = decrypt_pad & ~\u1_uk_K_r0_reg[49]/NET0131  ;
  assign n47794 = ~decrypt_pad & ~\u1_uk_K_r0_reg[28]/NET0131  ;
  assign n47795 = ~n47793 & ~n47794 ;
  assign n47796 = \u1_R0_reg[28]/NET0131  & ~n47795 ;
  assign n47797 = ~\u1_R0_reg[28]/NET0131  & n47795 ;
  assign n47798 = ~n47796 & ~n47797 ;
  assign n47818 = decrypt_pad & ~\u1_uk_K_r0_reg[29]/NET0131  ;
  assign n47819 = ~decrypt_pad & ~\u1_uk_K_r0_reg[8]/NET0131  ;
  assign n47820 = ~n47818 & ~n47819 ;
  assign n47821 = \u1_R0_reg[26]/NET0131  & ~n47820 ;
  assign n47822 = ~\u1_R0_reg[26]/NET0131  & n47820 ;
  assign n47823 = ~n47821 & ~n47822 ;
  assign n47843 = ~n47810 & n47823 ;
  assign n47811 = n47804 & n47810 ;
  assign n47872 = n47811 & ~n47823 ;
  assign n47873 = ~n47843 & ~n47872 ;
  assign n47874 = n47798 & ~n47873 ;
  assign n47875 = ~n47871 & ~n47874 ;
  assign n47876 = n47817 & ~n47875 ;
  assign n47828 = n47804 & ~n47817 ;
  assign n47862 = n47828 & n47843 ;
  assign n47844 = ~n47804 & ~n47817 ;
  assign n47868 = n47810 & n47823 ;
  assign n47869 = n47844 & n47868 ;
  assign n47870 = ~n47862 & ~n47869 ;
  assign n47877 = ~n47823 & n47871 ;
  assign n47878 = n47870 & ~n47877 ;
  assign n47879 = ~n47876 & n47878 ;
  assign n47880 = n47834 & ~n47879 ;
  assign n47846 = n47810 & n47817 ;
  assign n47847 = ~n47804 & n47846 ;
  assign n47824 = n47817 & n47823 ;
  assign n47842 = n47804 & n47824 ;
  assign n47845 = n47843 & n47844 ;
  assign n47848 = ~n47842 & ~n47845 ;
  assign n47849 = ~n47847 & n47848 ;
  assign n47850 = ~n47834 & ~n47849 ;
  assign n47825 = ~n47817 & ~n47823 ;
  assign n47826 = ~n47824 & ~n47825 ;
  assign n47827 = n47811 & ~n47826 ;
  assign n47835 = n47828 & ~n47834 ;
  assign n47836 = ~n47804 & n47817 ;
  assign n47837 = n47817 & n47834 ;
  assign n47838 = ~n47836 & ~n47837 ;
  assign n47839 = ~n47810 & ~n47838 ;
  assign n47840 = ~n47835 & ~n47839 ;
  assign n47841 = ~n47823 & ~n47840 ;
  assign n47851 = ~n47827 & ~n47841 ;
  assign n47852 = ~n47850 & n47851 ;
  assign n47853 = ~n47798 & ~n47852 ;
  assign n47854 = n47810 & ~n47834 ;
  assign n47855 = ~n47826 & n47854 ;
  assign n47856 = n47804 & ~n47810 ;
  assign n47857 = n47817 & n47856 ;
  assign n47858 = ~n47823 & n47857 ;
  assign n47859 = n47810 & n47828 ;
  assign n47860 = ~n47858 & ~n47859 ;
  assign n47861 = ~n47834 & ~n47860 ;
  assign n47863 = ~n47810 & ~n47823 ;
  assign n47864 = n47844 & n47863 ;
  assign n47865 = ~n47862 & ~n47864 ;
  assign n47866 = ~n47861 & n47865 ;
  assign n47867 = n47798 & ~n47866 ;
  assign n47881 = ~n47855 & ~n47867 ;
  assign n47882 = ~n47853 & n47881 ;
  assign n47883 = ~n47880 & n47882 ;
  assign n47884 = ~\u1_L0_reg[22]/NET0131  & ~n47883 ;
  assign n47885 = \u1_L0_reg[22]/NET0131  & n47883 ;
  assign n47886 = ~n47884 & ~n47885 ;
  assign n47921 = decrypt_pad & ~\u1_uk_K_r0_reg[42]/NET0131  ;
  assign n47922 = ~decrypt_pad & ~\u1_uk_K_r0_reg[21]/NET0131  ;
  assign n47923 = ~n47921 & ~n47922 ;
  assign n47924 = \u1_R0_reg[24]/NET0131  & ~n47923 ;
  assign n47925 = ~\u1_R0_reg[24]/NET0131  & n47923 ;
  assign n47926 = ~n47924 & ~n47925 ;
  assign n47887 = decrypt_pad & ~\u1_uk_K_r0_reg[31]/NET0131  ;
  assign n47888 = ~decrypt_pad & ~\u1_uk_K_r0_reg[37]/NET0131  ;
  assign n47889 = ~n47887 & ~n47888 ;
  assign n47890 = \u1_R0_reg[22]/NET0131  & ~n47889 ;
  assign n47891 = ~\u1_R0_reg[22]/NET0131  & n47889 ;
  assign n47892 = ~n47890 & ~n47891 ;
  assign n47900 = decrypt_pad & ~\u1_uk_K_r0_reg[21]/NET0131  ;
  assign n47901 = ~decrypt_pad & ~\u1_uk_K_r0_reg[0]/NET0131  ;
  assign n47902 = ~n47900 & ~n47901 ;
  assign n47903 = \u1_R0_reg[20]/NET0131  & ~n47902 ;
  assign n47904 = ~\u1_R0_reg[20]/NET0131  & n47902 ;
  assign n47905 = ~n47903 & ~n47904 ;
  assign n47913 = decrypt_pad & ~\u1_uk_K_r0_reg[36]/NET0131  ;
  assign n47914 = ~decrypt_pad & ~\u1_uk_K_r0_reg[15]/NET0131  ;
  assign n47915 = ~n47913 & ~n47914 ;
  assign n47916 = \u1_R0_reg[21]/NET0131  & ~n47915 ;
  assign n47917 = ~\u1_R0_reg[21]/NET0131  & n47915 ;
  assign n47918 = ~n47916 & ~n47917 ;
  assign n47929 = ~n47905 & n47918 ;
  assign n47906 = decrypt_pad & ~\u1_uk_K_r0_reg[37]/NET0131  ;
  assign n47907 = ~decrypt_pad & ~\u1_uk_K_r0_reg[16]/NET0131  ;
  assign n47908 = ~n47906 & ~n47907 ;
  assign n47909 = \u1_R0_reg[25]/NET0131  & ~n47908 ;
  assign n47910 = ~\u1_R0_reg[25]/NET0131  & n47908 ;
  assign n47911 = ~n47909 & ~n47910 ;
  assign n47937 = n47905 & n47911 ;
  assign n47942 = ~n47929 & ~n47937 ;
  assign n47943 = n47892 & ~n47942 ;
  assign n47893 = decrypt_pad & ~\u1_uk_K_r0_reg[16]/NET0131  ;
  assign n47894 = ~decrypt_pad & ~\u1_uk_K_r0_reg[50]/NET0131  ;
  assign n47895 = ~n47893 & ~n47894 ;
  assign n47896 = \u1_R0_reg[23]/NET0131  & ~n47895 ;
  assign n47897 = ~\u1_R0_reg[23]/NET0131  & n47895 ;
  assign n47898 = ~n47896 & ~n47897 ;
  assign n47927 = n47911 & n47918 ;
  assign n47940 = ~n47905 & n47927 ;
  assign n47941 = ~n47892 & ~n47940 ;
  assign n47944 = ~n47898 & ~n47941 ;
  assign n47945 = ~n47943 & n47944 ;
  assign n47931 = n47905 & ~n47911 ;
  assign n47932 = ~n47892 & ~n47918 ;
  assign n47933 = n47931 & n47932 ;
  assign n47928 = n47905 & n47927 ;
  assign n47930 = n47892 & n47929 ;
  assign n47934 = ~n47928 & ~n47930 ;
  assign n47935 = ~n47933 & n47934 ;
  assign n47936 = n47898 & ~n47935 ;
  assign n47899 = ~n47892 & ~n47898 ;
  assign n47938 = n47899 & n47937 ;
  assign n47939 = ~n47918 & n47938 ;
  assign n47946 = ~n47936 & ~n47939 ;
  assign n47947 = ~n47945 & n47946 ;
  assign n47948 = n47926 & ~n47947 ;
  assign n47955 = ~n47911 & n47918 ;
  assign n47956 = n47905 & ~n47955 ;
  assign n47957 = ~n47898 & ~n47905 ;
  assign n47958 = ~n47892 & ~n47957 ;
  assign n47959 = ~n47956 & n47958 ;
  assign n47949 = ~n47905 & n47911 ;
  assign n47950 = ~n47918 & n47949 ;
  assign n47951 = n47898 & n47950 ;
  assign n47952 = n47905 & ~n47918 ;
  assign n47953 = n47892 & n47898 ;
  assign n47954 = n47952 & n47953 ;
  assign n47968 = ~n47951 & ~n47954 ;
  assign n47969 = ~n47959 & n47968 ;
  assign n47960 = n47892 & n47937 ;
  assign n47961 = ~n47918 & n47960 ;
  assign n47962 = n47899 & n47931 ;
  assign n47963 = ~n47961 & ~n47962 ;
  assign n47964 = ~n47892 & n47918 ;
  assign n47965 = n47905 & n47964 ;
  assign n47966 = ~n47930 & ~n47965 ;
  assign n47967 = ~n47898 & ~n47966 ;
  assign n47970 = n47963 & ~n47967 ;
  assign n47971 = n47969 & n47970 ;
  assign n47972 = ~n47926 & ~n47971 ;
  assign n47973 = n47918 & n47931 ;
  assign n47974 = ~n47898 & n47973 ;
  assign n47975 = ~n47951 & ~n47974 ;
  assign n47976 = ~n47892 & ~n47975 ;
  assign n47912 = ~n47905 & ~n47911 ;
  assign n47919 = n47912 & ~n47918 ;
  assign n47920 = n47899 & n47919 ;
  assign n47977 = n47912 & n47964 ;
  assign n47978 = ~n47960 & ~n47977 ;
  assign n47979 = n47898 & ~n47978 ;
  assign n47980 = ~n47920 & ~n47979 ;
  assign n47981 = ~n47976 & n47980 ;
  assign n47982 = ~n47972 & n47981 ;
  assign n47983 = ~n47948 & n47982 ;
  assign n47984 = \u1_L0_reg[11]/NET0131  & ~n47983 ;
  assign n47985 = ~\u1_L0_reg[11]/NET0131  & n47983 ;
  assign n47986 = ~n47984 & ~n47985 ;
  assign n47987 = decrypt_pad & ~\u1_uk_K_r0_reg[39]/NET0131  ;
  assign n47988 = ~decrypt_pad & ~\u1_uk_K_r0_reg[18]/NET0131  ;
  assign n47989 = ~n47987 & ~n47988 ;
  assign n47990 = \u1_R0_reg[15]/NET0131  & ~n47989 ;
  assign n47991 = ~\u1_R0_reg[15]/NET0131  & n47989 ;
  assign n47992 = ~n47990 & ~n47991 ;
  assign n47993 = decrypt_pad & ~\u1_uk_K_r0_reg[5]/NET0131  ;
  assign n47994 = ~decrypt_pad & ~\u1_uk_K_r0_reg[41]/NET0131  ;
  assign n47995 = ~n47993 & ~n47994 ;
  assign n47996 = \u1_R0_reg[13]/NET0131  & ~n47995 ;
  assign n47997 = ~\u1_R0_reg[13]/NET0131  & n47995 ;
  assign n47998 = ~n47996 & ~n47997 ;
  assign n47999 = decrypt_pad & ~\u1_uk_K_r0_reg[11]/NET0131  ;
  assign n48000 = ~decrypt_pad & ~\u1_uk_K_r0_reg[47]/NET0131  ;
  assign n48001 = ~n47999 & ~n48000 ;
  assign n48002 = \u1_R0_reg[12]/NET0131  & ~n48001 ;
  assign n48003 = ~\u1_R0_reg[12]/NET0131  & n48001 ;
  assign n48004 = ~n48002 & ~n48003 ;
  assign n48005 = n47998 & ~n48004 ;
  assign n48006 = decrypt_pad & ~\u1_uk_K_r0_reg[6]/NET0131  ;
  assign n48007 = ~decrypt_pad & ~\u1_uk_K_r0_reg[10]/NET0131  ;
  assign n48008 = ~n48006 & ~n48007 ;
  assign n48009 = \u1_R0_reg[14]/NET0131  & ~n48008 ;
  assign n48010 = ~\u1_R0_reg[14]/NET0131  & n48008 ;
  assign n48011 = ~n48009 & ~n48010 ;
  assign n48012 = decrypt_pad & ~\u1_uk_K_r0_reg[27]/NET0131  ;
  assign n48013 = ~decrypt_pad & ~\u1_uk_K_r0_reg[6]/NET0131  ;
  assign n48014 = ~n48012 & ~n48013 ;
  assign n48015 = \u1_R0_reg[17]/NET0131  & ~n48014 ;
  assign n48016 = ~\u1_R0_reg[17]/NET0131  & n48014 ;
  assign n48017 = ~n48015 & ~n48016 ;
  assign n48018 = ~n48011 & n48017 ;
  assign n48019 = n48005 & n48018 ;
  assign n48020 = ~n47992 & ~n48019 ;
  assign n48027 = ~n47998 & ~n48017 ;
  assign n48028 = ~n48004 & n48027 ;
  assign n48029 = ~n48011 & n48028 ;
  assign n48021 = n48004 & ~n48017 ;
  assign n48022 = ~n47998 & n48011 ;
  assign n48023 = n48021 & n48022 ;
  assign n48024 = n47992 & ~n48023 ;
  assign n48025 = n47998 & ~n48011 ;
  assign n48026 = n48021 & n48025 ;
  assign n48030 = n48024 & ~n48026 ;
  assign n48031 = ~n48029 & n48030 ;
  assign n48032 = ~n48020 & ~n48031 ;
  assign n48051 = ~n48004 & n48022 ;
  assign n48052 = ~n47992 & ~n48017 ;
  assign n48053 = n48051 & n48052 ;
  assign n48043 = decrypt_pad & ~\u1_uk_K_r0_reg[47]/NET0131  ;
  assign n48044 = ~decrypt_pad & ~\u1_uk_K_r0_reg[26]/NET0131  ;
  assign n48045 = ~n48043 & ~n48044 ;
  assign n48046 = \u1_R0_reg[16]/NET0131  & ~n48045 ;
  assign n48047 = ~\u1_R0_reg[16]/NET0131  & n48045 ;
  assign n48048 = ~n48046 & ~n48047 ;
  assign n48037 = ~n47998 & n48004 ;
  assign n48038 = ~n48005 & ~n48037 ;
  assign n48049 = ~n47992 & ~n48011 ;
  assign n48050 = ~n48038 & n48049 ;
  assign n48054 = n48048 & ~n48050 ;
  assign n48055 = ~n48053 & n48054 ;
  assign n48033 = n48004 & n48017 ;
  assign n48034 = n47998 & n48033 ;
  assign n48035 = n48011 & n48034 ;
  assign n48036 = ~n48019 & ~n48035 ;
  assign n48039 = ~n48004 & n48017 ;
  assign n48040 = ~n48021 & ~n48039 ;
  assign n48041 = n47992 & n48038 ;
  assign n48042 = ~n48040 & n48041 ;
  assign n48056 = n48036 & ~n48042 ;
  assign n48057 = n48055 & n48056 ;
  assign n48064 = n47992 & ~n48028 ;
  assign n48065 = ~n48034 & n48064 ;
  assign n48066 = n48011 & n48021 ;
  assign n48061 = ~n47998 & n48017 ;
  assign n48067 = ~n47992 & ~n48061 ;
  assign n48068 = ~n48066 & n48067 ;
  assign n48069 = ~n48065 & ~n48068 ;
  assign n48058 = n48005 & ~n48017 ;
  assign n48059 = n48011 & n48058 ;
  assign n48060 = ~n48029 & ~n48059 ;
  assign n48070 = n47992 & n48011 ;
  assign n48071 = n48005 & n48070 ;
  assign n48062 = n48004 & ~n48011 ;
  assign n48063 = n48061 & n48062 ;
  assign n48072 = ~n48048 & ~n48063 ;
  assign n48073 = ~n48071 & n48072 ;
  assign n48074 = n48060 & n48073 ;
  assign n48075 = ~n48069 & n48074 ;
  assign n48076 = ~n48057 & ~n48075 ;
  assign n48077 = ~n48032 & ~n48076 ;
  assign n48078 = ~\u1_L0_reg[20]/NET0131  & ~n48077 ;
  assign n48079 = \u1_L0_reg[20]/NET0131  & n48077 ;
  assign n48080 = ~n48078 & ~n48079 ;
  assign n48081 = decrypt_pad & ~\u1_uk_K_r0_reg[14]/NET0131  ;
  assign n48082 = ~decrypt_pad & ~\u1_uk_K_r0_reg[52]/P0001  ;
  assign n48083 = ~n48081 & ~n48082 ;
  assign n48084 = \u1_R0_reg[32]/NET0131  & ~n48083 ;
  assign n48085 = ~\u1_R0_reg[32]/NET0131  & n48083 ;
  assign n48086 = ~n48084 & ~n48085 ;
  assign n48112 = decrypt_pad & ~\u1_uk_K_r0_reg[51]/NET0131  ;
  assign n48113 = ~decrypt_pad & ~\u1_uk_K_r0_reg[30]/NET0131  ;
  assign n48114 = ~n48112 & ~n48113 ;
  assign n48115 = \u1_R0_reg[30]/NET0131  & ~n48114 ;
  assign n48116 = ~\u1_R0_reg[30]/NET0131  & n48114 ;
  assign n48117 = ~n48115 & ~n48116 ;
  assign n48105 = decrypt_pad & ~\u1_uk_K_r0_reg[23]/NET0131  ;
  assign n48106 = ~decrypt_pad & ~\u1_uk_K_r0_reg[2]/NET0131  ;
  assign n48107 = ~n48105 & ~n48106 ;
  assign n48108 = \u1_R0_reg[28]/NET0131  & ~n48107 ;
  assign n48109 = ~\u1_R0_reg[28]/NET0131  & n48107 ;
  assign n48110 = ~n48108 & ~n48109 ;
  assign n48093 = decrypt_pad & ~\u1_uk_K_r0_reg[35]/NET0131  ;
  assign n48094 = ~decrypt_pad & ~\u1_uk_K_r0_reg[14]/NET0131  ;
  assign n48095 = ~n48093 & ~n48094 ;
  assign n48096 = \u1_R0_reg[1]/NET0131  & ~n48095 ;
  assign n48097 = ~\u1_R0_reg[1]/NET0131  & n48095 ;
  assign n48098 = ~n48096 & ~n48097 ;
  assign n48099 = decrypt_pad & ~\u1_uk_K_r0_reg[50]/NET0131  ;
  assign n48100 = ~decrypt_pad & ~\u1_uk_K_r0_reg[29]/NET0131  ;
  assign n48101 = ~n48099 & ~n48100 ;
  assign n48102 = \u1_R0_reg[29]/NET0131  & ~n48101 ;
  assign n48103 = ~\u1_R0_reg[29]/NET0131  & n48101 ;
  assign n48104 = ~n48102 & ~n48103 ;
  assign n48124 = n48098 & n48104 ;
  assign n48153 = ~n48110 & n48124 ;
  assign n48154 = n48117 & n48153 ;
  assign n48147 = ~n48104 & ~n48117 ;
  assign n48148 = ~n48110 & n48147 ;
  assign n48087 = decrypt_pad & ~\u1_uk_K_r0_reg[8]/NET0131  ;
  assign n48088 = ~decrypt_pad & ~\u1_uk_K_r0_reg[42]/NET0131  ;
  assign n48089 = ~n48087 & ~n48088 ;
  assign n48090 = \u1_R0_reg[31]/P0001  & ~n48089 ;
  assign n48091 = ~\u1_R0_reg[31]/P0001  & n48089 ;
  assign n48092 = ~n48090 & ~n48091 ;
  assign n48111 = ~n48104 & n48110 ;
  assign n48118 = n48111 & n48117 ;
  assign n48155 = ~n48092 & ~n48118 ;
  assign n48156 = ~n48148 & n48155 ;
  assign n48130 = n48110 & ~n48117 ;
  assign n48157 = ~n48098 & n48104 ;
  assign n48159 = ~n48130 & n48157 ;
  assign n48158 = n48130 & ~n48157 ;
  assign n48160 = n48092 & ~n48158 ;
  assign n48161 = ~n48159 & n48160 ;
  assign n48162 = ~n48156 & ~n48161 ;
  assign n48163 = ~n48154 & ~n48162 ;
  assign n48164 = n48086 & ~n48163 ;
  assign n48119 = ~n48098 & n48118 ;
  assign n48120 = n48098 & ~n48110 ;
  assign n48121 = ~n48104 & n48120 ;
  assign n48122 = n48092 & ~n48121 ;
  assign n48123 = ~n48119 & n48122 ;
  assign n48125 = ~n48098 & ~n48110 ;
  assign n48126 = n48117 & n48125 ;
  assign n48127 = ~n48092 & ~n48124 ;
  assign n48128 = ~n48126 & n48127 ;
  assign n48129 = ~n48123 & ~n48128 ;
  assign n48131 = ~n48092 & n48130 ;
  assign n48134 = ~n48098 & ~n48130 ;
  assign n48132 = n48110 & n48117 ;
  assign n48133 = n48098 & ~n48132 ;
  assign n48135 = n48104 & ~n48133 ;
  assign n48136 = ~n48134 & n48135 ;
  assign n48137 = ~n48131 & ~n48136 ;
  assign n48138 = ~n48129 & n48137 ;
  assign n48139 = ~n48086 & ~n48138 ;
  assign n48141 = n48104 & ~n48117 ;
  assign n48142 = n48104 & ~n48110 ;
  assign n48143 = ~n48098 & ~n48142 ;
  assign n48144 = ~n48141 & ~n48143 ;
  assign n48145 = n48098 & ~n48130 ;
  assign n48146 = n48144 & ~n48145 ;
  assign n48140 = n48117 & n48121 ;
  assign n48149 = ~n48098 & n48148 ;
  assign n48150 = ~n48140 & ~n48149 ;
  assign n48151 = ~n48146 & n48150 ;
  assign n48152 = n48092 & ~n48151 ;
  assign n48165 = n48131 & n48157 ;
  assign n48166 = ~n48152 & ~n48165 ;
  assign n48167 = ~n48139 & n48166 ;
  assign n48168 = ~n48164 & n48167 ;
  assign n48169 = \u1_L0_reg[5]/NET0131  & ~n48168 ;
  assign n48170 = ~\u1_L0_reg[5]/NET0131  & n48168 ;
  assign n48171 = ~n48169 & ~n48170 ;
  assign n48199 = decrypt_pad & ~\u1_uk_K_r0_reg[20]/NET0131  ;
  assign n48200 = ~decrypt_pad & ~\u1_uk_K_r0_reg[24]/NET0131  ;
  assign n48201 = ~n48199 & ~n48200 ;
  assign n48202 = \u1_R0_reg[4]/NET0131  & ~n48201 ;
  assign n48203 = ~\u1_R0_reg[4]/NET0131  & n48201 ;
  assign n48204 = ~n48202 & ~n48203 ;
  assign n48172 = decrypt_pad & ~\u1_uk_K_r0_reg[10]/NET0131  ;
  assign n48173 = ~decrypt_pad & ~\u1_uk_K_r0_reg[46]/NET0131  ;
  assign n48174 = ~n48172 & ~n48173 ;
  assign n48175 = \u1_R0_reg[3]/NET0131  & ~n48174 ;
  assign n48176 = ~\u1_R0_reg[3]/NET0131  & n48174 ;
  assign n48177 = ~n48175 & ~n48176 ;
  assign n48191 = decrypt_pad & ~\u1_uk_K_r0_reg[18]/NET0131  ;
  assign n48192 = ~decrypt_pad & ~\u1_uk_K_r0_reg[54]/NET0131  ;
  assign n48193 = ~n48191 & ~n48192 ;
  assign n48194 = \u1_R0_reg[1]/NET0131  & ~n48193 ;
  assign n48195 = ~\u1_R0_reg[1]/NET0131  & n48193 ;
  assign n48196 = ~n48194 & ~n48195 ;
  assign n48206 = decrypt_pad & ~\u1_uk_K_r0_reg[48]/NET0131  ;
  assign n48207 = ~decrypt_pad & ~\u1_uk_K_r0_reg[27]/NET0131  ;
  assign n48208 = ~n48206 & ~n48207 ;
  assign n48209 = \u1_R0_reg[5]/NET0131  & ~n48208 ;
  assign n48210 = ~\u1_R0_reg[5]/NET0131  & n48208 ;
  assign n48211 = ~n48209 & ~n48210 ;
  assign n48219 = ~n48196 & n48211 ;
  assign n48178 = decrypt_pad & ~\u1_uk_K_r0_reg[33]/NET0131  ;
  assign n48179 = ~decrypt_pad & ~\u1_uk_K_r0_reg[12]/NET0131  ;
  assign n48180 = ~n48178 & ~n48179 ;
  assign n48181 = \u1_R0_reg[2]/NET0131  & ~n48180 ;
  assign n48182 = ~\u1_R0_reg[2]/NET0131  & n48180 ;
  assign n48183 = ~n48181 & ~n48182 ;
  assign n48185 = decrypt_pad & ~\u1_uk_K_r0_reg[54]/NET0131  ;
  assign n48186 = ~decrypt_pad & ~\u1_uk_K_r0_reg[33]/NET0131  ;
  assign n48187 = ~n48185 & ~n48186 ;
  assign n48188 = \u1_R0_reg[32]/NET0131  & ~n48187 ;
  assign n48189 = ~\u1_R0_reg[32]/NET0131  & n48187 ;
  assign n48190 = ~n48188 & ~n48189 ;
  assign n48237 = n48183 & ~n48190 ;
  assign n48238 = ~n48211 & n48237 ;
  assign n48239 = ~n48219 & ~n48238 ;
  assign n48240 = n48177 & ~n48239 ;
  assign n48224 = ~n48177 & n48196 ;
  assign n48233 = ~n48196 & ~n48211 ;
  assign n48234 = ~n48183 & n48233 ;
  assign n48235 = ~n48224 & ~n48234 ;
  assign n48236 = n48190 & ~n48235 ;
  assign n48184 = n48177 & ~n48183 ;
  assign n48242 = ~n48184 & n48196 ;
  assign n48241 = ~n48183 & ~n48211 ;
  assign n48243 = ~n48190 & ~n48241 ;
  assign n48244 = ~n48242 & n48243 ;
  assign n48245 = ~n48236 & ~n48244 ;
  assign n48246 = ~n48240 & n48245 ;
  assign n48247 = n48204 & ~n48246 ;
  assign n48197 = n48190 & ~n48196 ;
  assign n48217 = n48197 & ~n48211 ;
  assign n48218 = n48183 & n48217 ;
  assign n48220 = ~n48183 & ~n48190 ;
  assign n48221 = ~n48219 & n48220 ;
  assign n48222 = ~n48218 & ~n48221 ;
  assign n48223 = ~n48177 & ~n48222 ;
  assign n48205 = n48177 & n48183 ;
  assign n48212 = ~n48190 & ~n48211 ;
  assign n48213 = n48190 & n48211 ;
  assign n48214 = ~n48212 & ~n48213 ;
  assign n48215 = n48196 & n48214 ;
  assign n48216 = n48205 & n48215 ;
  assign n48225 = n48213 & ~n48224 ;
  assign n48226 = ~n48190 & n48196 ;
  assign n48227 = ~n48211 & n48226 ;
  assign n48228 = ~n48225 & ~n48227 ;
  assign n48229 = ~n48183 & ~n48228 ;
  assign n48230 = ~n48216 & ~n48229 ;
  assign n48231 = ~n48223 & n48230 ;
  assign n48232 = ~n48204 & ~n48231 ;
  assign n48248 = n48183 & n48213 ;
  assign n48249 = ~n48241 & ~n48248 ;
  assign n48250 = n48196 & ~n48249 ;
  assign n48251 = n48219 & n48237 ;
  assign n48252 = ~n48250 & ~n48251 ;
  assign n48253 = ~n48177 & ~n48252 ;
  assign n48198 = n48184 & n48197 ;
  assign n48254 = ~n48196 & n48205 ;
  assign n48255 = n48212 & n48254 ;
  assign n48256 = ~n48198 & ~n48255 ;
  assign n48257 = ~n48253 & n48256 ;
  assign n48258 = ~n48232 & n48257 ;
  assign n48259 = ~n48247 & n48258 ;
  assign n48260 = ~\u1_L0_reg[31]/NET0131  & ~n48259 ;
  assign n48261 = \u1_L0_reg[31]/NET0131  & n48259 ;
  assign n48262 = ~n48260 & ~n48261 ;
  assign n48280 = n48004 & n48025 ;
  assign n48281 = n48060 & ~n48280 ;
  assign n48274 = n48017 & n48062 ;
  assign n48275 = ~n48028 & ~n48274 ;
  assign n48276 = ~n47992 & ~n48275 ;
  assign n48277 = ~n48018 & ~n48037 ;
  assign n48278 = n47992 & ~n48274 ;
  assign n48279 = ~n48277 & n48278 ;
  assign n48282 = ~n48276 & ~n48279 ;
  assign n48283 = n48281 & n48282 ;
  assign n48284 = ~n48048 & ~n48283 ;
  assign n48268 = n48021 & ~n48025 ;
  assign n48269 = ~n48019 & ~n48268 ;
  assign n48270 = ~n47992 & ~n48269 ;
  assign n48264 = n48011 & n48038 ;
  assign n48265 = n48017 & n48264 ;
  assign n48266 = ~n48058 & ~n48063 ;
  assign n48267 = n47992 & ~n48266 ;
  assign n48271 = ~n48265 & ~n48267 ;
  assign n48272 = ~n48270 & n48271 ;
  assign n48273 = n48048 & ~n48272 ;
  assign n48285 = ~n48029 & ~n48265 ;
  assign n48286 = ~n47992 & ~n48285 ;
  assign n48263 = n47992 & n48026 ;
  assign n48287 = ~n48071 & ~n48263 ;
  assign n48288 = ~n48286 & n48287 ;
  assign n48289 = ~n48273 & n48288 ;
  assign n48290 = ~n48284 & n48289 ;
  assign n48291 = ~\u1_L0_reg[10]/NET0131  & ~n48290 ;
  assign n48292 = \u1_L0_reg[10]/NET0131  & n48290 ;
  assign n48293 = ~n48291 & ~n48292 ;
  assign n48304 = ~n47811 & ~n47817 ;
  assign n48305 = n47823 & ~n47837 ;
  assign n48306 = ~n48304 & n48305 ;
  assign n48298 = ~n47811 & ~n47871 ;
  assign n48299 = ~n47834 & ~n48298 ;
  assign n48307 = ~n47798 & ~n48299 ;
  assign n48308 = ~n48306 & n48307 ;
  assign n48295 = ~n47863 & ~n47868 ;
  assign n48294 = ~n47828 & ~n47836 ;
  assign n48296 = ~n47846 & n48294 ;
  assign n48297 = n48295 & n48296 ;
  assign n48300 = ~n47823 & n47836 ;
  assign n48301 = n47828 & n47834 ;
  assign n48302 = ~n48300 & ~n48301 ;
  assign n48303 = ~n47810 & ~n48302 ;
  assign n48309 = ~n48297 & ~n48303 ;
  assign n48310 = n48308 & n48309 ;
  assign n48311 = n47811 & n47825 ;
  assign n48316 = n47798 & ~n47869 ;
  assign n48317 = ~n48311 & n48316 ;
  assign n48318 = ~n47858 & n48317 ;
  assign n48312 = ~n47835 & ~n47836 ;
  assign n48313 = n47843 & ~n48312 ;
  assign n48314 = ~n47846 & ~n47864 ;
  assign n48315 = n47834 & ~n48314 ;
  assign n48319 = ~n48313 & ~n48315 ;
  assign n48320 = n48318 & n48319 ;
  assign n48321 = ~n48310 & ~n48320 ;
  assign n48322 = \u1_L0_reg[12]/NET0131  & n48321 ;
  assign n48323 = ~\u1_L0_reg[12]/NET0131  & ~n48321 ;
  assign n48324 = ~n48322 & ~n48323 ;
  assign n48385 = decrypt_pad & ~\u1_uk_K_r0_reg[30]/NET0131  ;
  assign n48386 = ~decrypt_pad & ~\u1_uk_K_r0_reg[9]/NET0131  ;
  assign n48387 = ~n48385 & ~n48386 ;
  assign n48388 = \u1_R0_reg[20]/NET0131  & ~n48387 ;
  assign n48389 = ~\u1_R0_reg[20]/NET0131  & n48387 ;
  assign n48390 = ~n48388 & ~n48389 ;
  assign n48365 = decrypt_pad & ~\u1_uk_K_r0_reg[15]/NET0131  ;
  assign n48366 = ~decrypt_pad & ~\u1_uk_K_r0_reg[49]/NET0131  ;
  assign n48367 = ~n48365 & ~n48366 ;
  assign n48368 = \u1_R0_reg[19]/NET0131  & ~n48367 ;
  assign n48369 = ~\u1_R0_reg[19]/NET0131  & n48367 ;
  assign n48370 = ~n48368 & ~n48369 ;
  assign n48325 = decrypt_pad & ~\u1_uk_K_r0_reg[0]/NET0131  ;
  assign n48326 = ~decrypt_pad & ~\u1_uk_K_r0_reg[38]/NET0131  ;
  assign n48327 = ~n48325 & ~n48326 ;
  assign n48328 = \u1_R0_reg[21]/NET0131  & ~n48327 ;
  assign n48329 = ~\u1_R0_reg[21]/NET0131  & n48327 ;
  assign n48330 = ~n48328 & ~n48329 ;
  assign n48338 = decrypt_pad & ~\u1_uk_K_r0_reg[38]/NET0131  ;
  assign n48339 = ~decrypt_pad & ~\u1_uk_K_r0_reg[44]/NET0131  ;
  assign n48340 = ~n48338 & ~n48339 ;
  assign n48341 = \u1_R0_reg[17]/NET0131  & ~n48340 ;
  assign n48342 = ~\u1_R0_reg[17]/NET0131  & n48340 ;
  assign n48343 = ~n48341 & ~n48342 ;
  assign n48344 = decrypt_pad & ~\u1_uk_K_r0_reg[43]/NET0131  ;
  assign n48345 = ~decrypt_pad & ~\u1_uk_K_r0_reg[22]/NET0131  ;
  assign n48346 = ~n48344 & ~n48345 ;
  assign n48347 = \u1_R0_reg[16]/NET0131  & ~n48346 ;
  assign n48348 = ~\u1_R0_reg[16]/NET0131  & n48346 ;
  assign n48349 = ~n48347 & ~n48348 ;
  assign n48356 = ~n48343 & ~n48349 ;
  assign n48357 = n48330 & n48356 ;
  assign n48392 = n48343 & n48349 ;
  assign n48393 = ~n48330 & n48392 ;
  assign n48396 = ~n48357 & ~n48393 ;
  assign n48331 = decrypt_pad & ~\u1_uk_K_r0_reg[28]/NET0131  ;
  assign n48332 = ~decrypt_pad & ~\u1_uk_K_r0_reg[7]/NET0131  ;
  assign n48333 = ~n48331 & ~n48332 ;
  assign n48334 = \u1_R0_reg[18]/NET0131  & ~n48333 ;
  assign n48335 = ~\u1_R0_reg[18]/NET0131  & n48333 ;
  assign n48336 = ~n48334 & ~n48335 ;
  assign n48337 = n48330 & ~n48336 ;
  assign n48394 = n48337 & n48349 ;
  assign n48375 = n48336 & ~n48349 ;
  assign n48395 = n48330 & n48375 ;
  assign n48397 = ~n48394 & ~n48395 ;
  assign n48398 = n48396 & n48397 ;
  assign n48399 = n48370 & ~n48398 ;
  assign n48407 = ~n48336 & ~n48370 ;
  assign n48379 = ~n48330 & ~n48349 ;
  assign n48380 = ~n48343 & n48379 ;
  assign n48352 = n48343 & ~n48349 ;
  assign n48408 = n48330 & n48352 ;
  assign n48409 = ~n48380 & ~n48408 ;
  assign n48410 = n48407 & ~n48409 ;
  assign n48358 = ~n48330 & n48349 ;
  assign n48400 = n48336 & ~n48343 ;
  assign n48401 = n48358 & n48400 ;
  assign n48402 = n48336 & ~n48370 ;
  assign n48403 = n48330 & n48392 ;
  assign n48404 = n48402 & n48403 ;
  assign n48411 = ~n48401 & ~n48404 ;
  assign n48405 = ~n48343 & n48394 ;
  assign n48406 = ~n48336 & n48393 ;
  assign n48412 = ~n48405 & ~n48406 ;
  assign n48413 = n48411 & n48412 ;
  assign n48414 = ~n48410 & n48413 ;
  assign n48415 = ~n48399 & n48414 ;
  assign n48416 = n48390 & ~n48415 ;
  assign n48350 = ~n48343 & n48349 ;
  assign n48351 = n48330 & n48350 ;
  assign n48353 = ~n48336 & n48352 ;
  assign n48354 = ~n48351 & ~n48353 ;
  assign n48355 = ~n48337 & ~n48354 ;
  assign n48361 = n48337 & n48343 ;
  assign n48362 = n48349 & n48361 ;
  assign n48371 = ~n48357 & ~n48370 ;
  assign n48359 = ~n48336 & ~n48343 ;
  assign n48360 = n48358 & n48359 ;
  assign n48363 = ~n48330 & n48343 ;
  assign n48364 = n48336 & n48363 ;
  assign n48372 = ~n48360 & ~n48364 ;
  assign n48373 = n48371 & n48372 ;
  assign n48374 = ~n48362 & n48373 ;
  assign n48376 = n48330 & n48336 ;
  assign n48377 = ~n48352 & ~n48376 ;
  assign n48378 = ~n48375 & ~n48377 ;
  assign n48381 = n48370 & ~n48380 ;
  assign n48382 = ~n48378 & n48381 ;
  assign n48383 = ~n48374 & ~n48382 ;
  assign n48384 = ~n48355 & ~n48383 ;
  assign n48391 = ~n48384 & ~n48390 ;
  assign n48417 = n48336 & n48357 ;
  assign n48418 = ~n48364 & ~n48417 ;
  assign n48419 = ~n48349 & ~n48418 ;
  assign n48420 = ~n48370 & n48419 ;
  assign n48421 = n48336 & n48380 ;
  assign n48422 = ~n48406 & ~n48421 ;
  assign n48423 = n48370 & ~n48422 ;
  assign n48424 = ~n48420 & ~n48423 ;
  assign n48425 = ~n48391 & n48424 ;
  assign n48426 = ~n48416 & n48425 ;
  assign n48427 = ~\u1_L0_reg[14]/NET0131  & ~n48426 ;
  assign n48428 = \u1_L0_reg[14]/NET0131  & n48426 ;
  assign n48429 = ~n48427 & ~n48428 ;
  assign n48441 = ~n48104 & n48117 ;
  assign n48442 = ~n48092 & n48098 ;
  assign n48443 = n48441 & n48442 ;
  assign n48449 = n48086 & ~n48443 ;
  assign n48445 = n48104 & n48110 ;
  assign n48446 = ~n48117 & n48445 ;
  assign n48447 = n48092 & ~n48104 ;
  assign n48448 = n48125 & n48447 ;
  assign n48450 = ~n48446 & ~n48448 ;
  assign n48451 = n48449 & n48450 ;
  assign n48431 = n48104 & n48126 ;
  assign n48444 = n48098 & n48118 ;
  assign n48452 = ~n48431 & ~n48444 ;
  assign n48453 = n48451 & n48452 ;
  assign n48454 = ~n48117 & n48157 ;
  assign n48455 = ~n48121 & ~n48445 ;
  assign n48456 = ~n48454 & n48455 ;
  assign n48457 = n48092 & ~n48456 ;
  assign n48458 = ~n48098 & n48130 ;
  assign n48459 = ~n48104 & n48458 ;
  assign n48460 = ~n48086 & ~n48459 ;
  assign n48461 = ~n48457 & n48460 ;
  assign n48462 = ~n48453 & ~n48461 ;
  assign n48430 = n48120 & n48141 ;
  assign n48432 = ~n48149 & ~n48430 ;
  assign n48433 = n48155 & ~n48431 ;
  assign n48434 = n48432 & n48433 ;
  assign n48435 = ~n48117 & n48121 ;
  assign n48436 = n48092 & ~n48154 ;
  assign n48437 = ~n48435 & n48436 ;
  assign n48438 = ~n48434 & ~n48437 ;
  assign n48439 = ~n48086 & ~n48092 ;
  assign n48440 = n48111 & n48439 ;
  assign n48463 = ~n48438 & ~n48440 ;
  assign n48464 = ~n48462 & n48463 ;
  assign n48465 = \u1_L0_reg[15]/P0001  & n48464 ;
  assign n48466 = ~\u1_L0_reg[15]/P0001  & ~n48464 ;
  assign n48467 = ~n48465 & ~n48466 ;
  assign n48479 = ~n47998 & n48018 ;
  assign n48480 = ~n48033 & ~n48479 ;
  assign n48481 = ~n47992 & ~n48062 ;
  assign n48482 = ~n48480 & n48481 ;
  assign n48484 = ~n48011 & ~n48017 ;
  assign n48485 = n48005 & n48484 ;
  assign n48483 = n48039 & n48070 ;
  assign n48486 = n48048 & ~n48483 ;
  assign n48487 = ~n48485 & n48486 ;
  assign n48476 = n47998 & n48011 ;
  assign n48477 = ~n48040 & n48476 ;
  assign n48478 = n47992 & n48028 ;
  assign n48488 = ~n48477 & ~n48478 ;
  assign n48489 = n48487 & n48488 ;
  assign n48490 = ~n48482 & n48489 ;
  assign n48491 = n48011 & ~n48039 ;
  assign n48492 = ~n48021 & ~n48491 ;
  assign n48493 = n47992 & n47998 ;
  assign n48494 = ~n48492 & n48493 ;
  assign n48495 = ~n48011 & n48037 ;
  assign n48496 = ~n48019 & ~n48048 ;
  assign n48497 = ~n48495 & n48496 ;
  assign n48498 = ~n48494 & n48497 ;
  assign n48499 = ~n48490 & ~n48498 ;
  assign n48468 = ~n48017 & ~n48038 ;
  assign n48469 = ~n48034 & ~n48468 ;
  assign n48470 = n48049 & ~n48469 ;
  assign n48471 = n47992 & n48018 ;
  assign n48472 = ~n48038 & n48471 ;
  assign n48473 = ~n48027 & ~n48051 ;
  assign n48474 = ~n47992 & ~n48048 ;
  assign n48475 = ~n48473 & n48474 ;
  assign n48500 = ~n48472 & ~n48475 ;
  assign n48501 = ~n48470 & n48500 ;
  assign n48502 = ~n48499 & n48501 ;
  assign n48503 = ~\u1_L0_reg[26]/NET0131  & ~n48502 ;
  assign n48504 = \u1_L0_reg[26]/NET0131  & n48502 ;
  assign n48505 = ~n48503 & ~n48504 ;
  assign n48514 = ~n48061 & ~n48484 ;
  assign n48515 = n48004 & ~n48514 ;
  assign n48516 = ~n47992 & ~n48515 ;
  assign n48517 = ~n48004 & n48484 ;
  assign n48518 = n48024 & ~n48517 ;
  assign n48519 = ~n48516 & ~n48518 ;
  assign n48520 = ~n48026 & n48036 ;
  assign n48521 = ~n48519 & n48520 ;
  assign n48522 = ~n48048 & ~n48521 ;
  assign n48509 = ~n47992 & n47998 ;
  assign n48510 = n48492 & n48509 ;
  assign n48506 = ~n48033 & n48264 ;
  assign n48507 = ~n48061 & ~n48495 ;
  assign n48508 = n47992 & ~n48507 ;
  assign n48511 = ~n48506 & ~n48508 ;
  assign n48512 = ~n48510 & n48511 ;
  assign n48513 = n48048 & ~n48512 ;
  assign n48524 = ~n48059 & ~n48265 ;
  assign n48525 = n47992 & ~n48524 ;
  assign n48523 = n48066 & n48509 ;
  assign n48526 = ~n48053 & ~n48523 ;
  assign n48527 = ~n48525 & n48526 ;
  assign n48528 = ~n48513 & n48527 ;
  assign n48529 = ~n48522 & n48528 ;
  assign n48530 = ~\u1_L0_reg[1]/NET0131  & ~n48529 ;
  assign n48531 = \u1_L0_reg[1]/NET0131  & n48529 ;
  assign n48532 = ~n48530 & ~n48531 ;
  assign n48537 = n48092 & ~n48153 ;
  assign n48535 = n48117 & n48445 ;
  assign n48536 = n48098 & n48147 ;
  assign n48538 = ~n48535 & ~n48536 ;
  assign n48539 = n48537 & n48538 ;
  assign n48540 = ~n48092 & ~n48458 ;
  assign n48541 = ~n48444 & n48540 ;
  assign n48542 = ~n48539 & ~n48541 ;
  assign n48543 = ~n48111 & n48117 ;
  assign n48544 = n48143 & n48543 ;
  assign n48545 = n48086 & ~n48435 ;
  assign n48546 = ~n48544 & n48545 ;
  assign n48547 = ~n48542 & n48546 ;
  assign n48548 = n48092 & ~n48098 ;
  assign n48549 = ~n48120 & ~n48548 ;
  assign n48550 = ~n48117 & ~n48549 ;
  assign n48551 = ~n48132 & ~n48447 ;
  assign n48552 = ~n48143 & n48551 ;
  assign n48553 = ~n48550 & n48552 ;
  assign n48557 = ~n48086 & ~n48119 ;
  assign n48554 = n48110 & ~n48124 ;
  assign n48555 = n48092 & ~n48147 ;
  assign n48556 = n48554 & n48555 ;
  assign n48558 = ~n48149 & ~n48556 ;
  assign n48559 = n48557 & n48558 ;
  assign n48560 = ~n48553 & n48559 ;
  assign n48561 = ~n48547 & ~n48560 ;
  assign n48533 = n48092 & n48148 ;
  assign n48534 = n48442 & n48446 ;
  assign n48562 = ~n48533 & ~n48534 ;
  assign n48563 = ~n48561 & n48562 ;
  assign n48564 = ~\u1_L0_reg[21]/NET0131  & ~n48563 ;
  assign n48565 = \u1_L0_reg[21]/NET0131  & n48563 ;
  assign n48566 = ~n48564 & ~n48565 ;
  assign n48567 = ~n48359 & ~n48375 ;
  assign n48568 = ~n48330 & ~n48567 ;
  assign n48569 = ~n48356 & ~n48403 ;
  assign n48570 = ~n48568 & n48569 ;
  assign n48571 = n48370 & ~n48570 ;
  assign n48572 = ~n48354 & ~n48370 ;
  assign n48573 = n48336 & n48393 ;
  assign n48574 = ~n48361 & ~n48573 ;
  assign n48575 = ~n48572 & n48574 ;
  assign n48576 = ~n48571 & n48575 ;
  assign n48577 = n48390 & ~n48576 ;
  assign n48589 = ~n48421 & ~n48573 ;
  assign n48590 = n48337 & n48356 ;
  assign n48591 = n48589 & ~n48590 ;
  assign n48592 = n48370 & ~n48591 ;
  assign n48578 = ~n48330 & n48370 ;
  assign n48579 = ~n48330 & n48350 ;
  assign n48580 = n48343 & n48375 ;
  assign n48581 = ~n48579 & ~n48580 ;
  assign n48582 = ~n48578 & ~n48581 ;
  assign n48584 = ~n48363 & n48370 ;
  assign n48583 = ~n48356 & ~n48370 ;
  assign n48585 = ~n48336 & ~n48583 ;
  assign n48586 = ~n48584 & n48585 ;
  assign n48587 = ~n48582 & ~n48586 ;
  assign n48588 = ~n48390 & ~n48587 ;
  assign n48593 = n48350 & n48402 ;
  assign n48594 = ~n48362 & ~n48593 ;
  assign n48595 = ~n48588 & n48594 ;
  assign n48596 = ~n48592 & n48595 ;
  assign n48597 = ~n48577 & n48596 ;
  assign n48598 = ~\u1_L0_reg[25]/NET0131  & ~n48597 ;
  assign n48599 = \u1_L0_reg[25]/NET0131  & n48597 ;
  assign n48600 = ~n48598 & ~n48599 ;
  assign n48613 = decrypt_pad & ~\u1_uk_K_r0_reg[26]/NET0131  ;
  assign n48614 = ~decrypt_pad & ~\u1_uk_K_r0_reg[5]/NET0131  ;
  assign n48615 = ~n48613 & ~n48614 ;
  assign n48616 = \u1_R0_reg[9]/NET0131  & ~n48615 ;
  assign n48617 = ~\u1_R0_reg[9]/NET0131  & n48615 ;
  assign n48618 = ~n48616 & ~n48617 ;
  assign n48619 = decrypt_pad & ~\u1_uk_K_r0_reg[13]/NET0131  ;
  assign n48620 = ~decrypt_pad & ~\u1_uk_K_r0_reg[17]/NET0131  ;
  assign n48621 = ~n48619 & ~n48620 ;
  assign n48622 = \u1_R0_reg[5]/NET0131  & ~n48621 ;
  assign n48623 = ~\u1_R0_reg[5]/NET0131  & n48621 ;
  assign n48624 = ~n48622 & ~n48623 ;
  assign n48625 = n48618 & ~n48624 ;
  assign n48607 = decrypt_pad & ~\u1_uk_K_r0_reg[34]/NET0131  ;
  assign n48608 = ~decrypt_pad & ~\u1_uk_K_r0_reg[13]/NET0131  ;
  assign n48609 = ~n48607 & ~n48608 ;
  assign n48610 = \u1_R0_reg[4]/NET0131  & ~n48609 ;
  assign n48611 = ~\u1_R0_reg[4]/NET0131  & n48609 ;
  assign n48612 = ~n48610 & ~n48611 ;
  assign n48641 = ~n48618 & n48624 ;
  assign n48644 = n48612 & ~n48641 ;
  assign n48645 = ~n48625 & n48644 ;
  assign n48626 = decrypt_pad & ~\u1_uk_K_r0_reg[55]/NET0131  ;
  assign n48627 = ~decrypt_pad & ~\u1_uk_K_r0_reg[34]/NET0131  ;
  assign n48628 = ~n48626 & ~n48627 ;
  assign n48629 = \u1_R0_reg[7]/NET0131  & ~n48628 ;
  assign n48630 = ~\u1_R0_reg[7]/NET0131  & n48628 ;
  assign n48631 = ~n48629 & ~n48630 ;
  assign n48633 = decrypt_pad & ~\u1_uk_K_r0_reg[4]/NET0131  ;
  assign n48634 = ~decrypt_pad & ~\u1_uk_K_r0_reg[40]/NET0131  ;
  assign n48635 = ~n48633 & ~n48634 ;
  assign n48636 = \u1_R0_reg[6]/NET0131  & ~n48635 ;
  assign n48637 = ~\u1_R0_reg[6]/NET0131  & n48635 ;
  assign n48638 = ~n48636 & ~n48637 ;
  assign n48642 = ~n48612 & n48641 ;
  assign n48643 = n48638 & n48642 ;
  assign n48646 = n48631 & ~n48643 ;
  assign n48647 = ~n48645 & n48646 ;
  assign n48655 = ~n48624 & n48638 ;
  assign n48656 = ~n48612 & n48655 ;
  assign n48657 = ~n48631 & ~n48656 ;
  assign n48648 = ~n48612 & n48618 ;
  assign n48649 = n48624 & n48648 ;
  assign n48650 = ~n48618 & ~n48638 ;
  assign n48651 = ~n48612 & n48650 ;
  assign n48652 = ~n48649 & ~n48651 ;
  assign n48653 = n48612 & n48638 ;
  assign n48654 = n48641 & n48653 ;
  assign n48658 = n48652 & ~n48654 ;
  assign n48659 = n48657 & n48658 ;
  assign n48660 = ~n48647 & ~n48659 ;
  assign n48632 = ~n48625 & ~n48631 ;
  assign n48639 = n48612 & ~n48638 ;
  assign n48640 = ~n48632 & n48639 ;
  assign n48601 = decrypt_pad & ~\u1_uk_K_r0_reg[46]/NET0131  ;
  assign n48602 = ~decrypt_pad & ~\u1_uk_K_r0_reg[25]/P0001  ;
  assign n48603 = ~n48601 & ~n48602 ;
  assign n48604 = \u1_R0_reg[8]/NET0131  & ~n48603 ;
  assign n48605 = ~\u1_R0_reg[8]/NET0131  & n48603 ;
  assign n48606 = ~n48604 & ~n48605 ;
  assign n48661 = ~n48612 & n48638 ;
  assign n48662 = n48625 & n48661 ;
  assign n48663 = n48606 & ~n48662 ;
  assign n48664 = ~n48640 & n48663 ;
  assign n48665 = ~n48660 & n48664 ;
  assign n48670 = n48631 & n48652 ;
  assign n48671 = ~n48612 & ~n48625 ;
  assign n48672 = ~n48624 & ~n48648 ;
  assign n48673 = ~n48650 & n48672 ;
  assign n48674 = ~n48671 & ~n48673 ;
  assign n48675 = n48657 & ~n48674 ;
  assign n48676 = ~n48670 & ~n48675 ;
  assign n48666 = n48612 & n48618 ;
  assign n48667 = ~n48612 & ~n48618 ;
  assign n48668 = ~n48666 & ~n48667 ;
  assign n48669 = n48655 & ~n48668 ;
  assign n48677 = ~n48606 & ~n48654 ;
  assign n48678 = ~n48669 & n48677 ;
  assign n48679 = ~n48676 & n48678 ;
  assign n48680 = ~n48665 & ~n48679 ;
  assign n48681 = ~\u1_L0_reg[28]/NET0131  & n48680 ;
  assign n48682 = \u1_L0_reg[28]/NET0131  & ~n48680 ;
  assign n48683 = ~n48681 & ~n48682 ;
  assign n48708 = n47892 & ~n47931 ;
  assign n48709 = ~n47949 & n48708 ;
  assign n48710 = ~n47919 & ~n48709 ;
  assign n48711 = ~n47898 & ~n48710 ;
  assign n48690 = n47892 & n47973 ;
  assign n48701 = n47892 & ~n47911 ;
  assign n48705 = n47929 & ~n48701 ;
  assign n48706 = ~n48690 & ~n48705 ;
  assign n48707 = n47898 & ~n48706 ;
  assign n48700 = ~n47892 & n47949 ;
  assign n48702 = ~n47905 & n48701 ;
  assign n48703 = ~n48700 & ~n48702 ;
  assign n48704 = ~n47918 & ~n48703 ;
  assign n48712 = n47963 & ~n48704 ;
  assign n48713 = ~n48707 & n48712 ;
  assign n48714 = ~n48711 & n48713 ;
  assign n48715 = n47926 & ~n48714 ;
  assign n48684 = ~n47918 & n47931 ;
  assign n48685 = ~n47928 & ~n48684 ;
  assign n48686 = ~n47930 & ~n47932 ;
  assign n48687 = ~n47911 & ~n48686 ;
  assign n48688 = n48685 & ~n48687 ;
  assign n48689 = n47898 & ~n48688 ;
  assign n48691 = ~n47892 & ~n47942 ;
  assign n48692 = ~n48690 & ~n48691 ;
  assign n48693 = ~n47898 & ~n48692 ;
  assign n48694 = n47892 & n47950 ;
  assign n48695 = ~n48693 & ~n48694 ;
  assign n48696 = ~n48689 & n48695 ;
  assign n48697 = ~n47926 & ~n48696 ;
  assign n48698 = ~n47892 & n47898 ;
  assign n48699 = n47927 & n48698 ;
  assign n48716 = ~n47933 & ~n48699 ;
  assign n48717 = ~n48697 & n48716 ;
  assign n48718 = ~n48715 & n48717 ;
  assign n48719 = \u1_L0_reg[29]/NET0131  & ~n48718 ;
  assign n48720 = ~\u1_L0_reg[29]/NET0131  & n48718 ;
  assign n48721 = ~n48719 & ~n48720 ;
  assign n48733 = n48625 & n48653 ;
  assign n48734 = n48631 & n48733 ;
  assign n48722 = ~n48624 & ~n48631 ;
  assign n48723 = ~n48661 & ~n48722 ;
  assign n48724 = n48618 & ~n48655 ;
  assign n48725 = ~n48723 & n48724 ;
  assign n48735 = ~n48606 & ~n48725 ;
  assign n48736 = ~n48734 & n48735 ;
  assign n48726 = ~n48625 & ~n48641 ;
  assign n48727 = ~n48666 & ~n48726 ;
  assign n48728 = ~n48638 & n48727 ;
  assign n48730 = ~n48624 & n48666 ;
  assign n48729 = ~n48625 & ~n48653 ;
  assign n48731 = ~n48631 & ~n48729 ;
  assign n48732 = ~n48730 & n48731 ;
  assign n48737 = ~n48728 & ~n48732 ;
  assign n48738 = n48736 & n48737 ;
  assign n48743 = ~n48624 & n48650 ;
  assign n48744 = n48612 & n48743 ;
  assign n48741 = n48624 & ~n48638 ;
  assign n48742 = n48666 & n48741 ;
  assign n48739 = n48624 & n48631 ;
  assign n48740 = ~n48661 & n48739 ;
  assign n48745 = n48606 & ~n48740 ;
  assign n48746 = ~n48742 & n48745 ;
  assign n48747 = ~n48744 & n48746 ;
  assign n48748 = ~n48738 & ~n48747 ;
  assign n48750 = ~n48618 & n48656 ;
  assign n48749 = n48612 & n48741 ;
  assign n48751 = n48631 & ~n48749 ;
  assign n48752 = ~n48750 & n48751 ;
  assign n48755 = n48667 & ~n48741 ;
  assign n48756 = ~n48733 & ~n48755 ;
  assign n48757 = n48606 & ~n48756 ;
  assign n48753 = ~n48655 & ~n48741 ;
  assign n48754 = n48648 & n48753 ;
  assign n48758 = ~n48631 & ~n48754 ;
  assign n48759 = ~n48757 & n48758 ;
  assign n48760 = ~n48752 & ~n48759 ;
  assign n48761 = ~n48748 & ~n48760 ;
  assign n48762 = \u1_L0_reg[2]/NET0131  & n48761 ;
  assign n48763 = ~\u1_L0_reg[2]/NET0131  & ~n48761 ;
  assign n48764 = ~n48762 & ~n48763 ;
  assign n48782 = ~n47905 & n47955 ;
  assign n48783 = ~n48694 & ~n48782 ;
  assign n48784 = ~n47898 & ~n48783 ;
  assign n48779 = ~n47973 & ~n48700 ;
  assign n48780 = ~n47961 & n48779 ;
  assign n48781 = n47898 & ~n48780 ;
  assign n48785 = ~n47933 & ~n47938 ;
  assign n48786 = ~n48781 & n48785 ;
  assign n48787 = ~n48784 & n48786 ;
  assign n48788 = ~n47926 & ~n48787 ;
  assign n48766 = n47899 & ~n47956 ;
  assign n48767 = n47937 & n48698 ;
  assign n48765 = n47892 & n47927 ;
  assign n48768 = ~n47977 & ~n48765 ;
  assign n48769 = ~n48767 & n48768 ;
  assign n48770 = ~n48766 & n48769 ;
  assign n48771 = n47926 & ~n48770 ;
  assign n48772 = ~n47919 & ~n47940 ;
  assign n48773 = ~n47973 & n48772 ;
  assign n48774 = n47953 & ~n48773 ;
  assign n48775 = n47892 & n48685 ;
  assign n48776 = ~n47892 & ~n47912 ;
  assign n48777 = ~n47898 & ~n48776 ;
  assign n48778 = ~n48775 & n48777 ;
  assign n48789 = ~n48774 & ~n48778 ;
  assign n48790 = ~n48771 & n48789 ;
  assign n48791 = ~n48788 & n48790 ;
  assign n48792 = ~\u1_L0_reg[4]/NET0131  & ~n48791 ;
  assign n48793 = \u1_L0_reg[4]/NET0131  & n48791 ;
  assign n48794 = ~n48792 & ~n48793 ;
  assign n48795 = ~n48654 & ~n48742 ;
  assign n48796 = ~n48642 & ~n48662 ;
  assign n48797 = ~n48744 & n48796 ;
  assign n48798 = ~n48606 & ~n48797 ;
  assign n48799 = n48795 & ~n48798 ;
  assign n48800 = ~n48631 & ~n48799 ;
  assign n48805 = ~n48618 & n48749 ;
  assign n48803 = ~n48641 & n48653 ;
  assign n48804 = ~n48624 & ~n48668 ;
  assign n48806 = ~n48803 & ~n48804 ;
  assign n48807 = ~n48805 & n48806 ;
  assign n48808 = n48631 & ~n48807 ;
  assign n48801 = ~n48638 & n48648 ;
  assign n48802 = ~n48722 & n48801 ;
  assign n48809 = ~n48606 & ~n48802 ;
  assign n48810 = ~n48808 & n48809 ;
  assign n48812 = ~n48631 & ~n48673 ;
  assign n48813 = n48618 & n48661 ;
  assign n48814 = n48631 & ~n48743 ;
  assign n48815 = ~n48813 & n48814 ;
  assign n48816 = ~n48812 & ~n48815 ;
  assign n48817 = n48606 & ~n48725 ;
  assign n48811 = ~n48638 & n48642 ;
  assign n48818 = n48795 & ~n48811 ;
  assign n48819 = n48817 & n48818 ;
  assign n48820 = ~n48816 & n48819 ;
  assign n48821 = ~n48810 & ~n48820 ;
  assign n48822 = ~n48800 & ~n48821 ;
  assign n48823 = ~\u1_L0_reg[13]/NET0131  & n48822 ;
  assign n48824 = \u1_L0_reg[13]/NET0131  & ~n48822 ;
  assign n48825 = ~n48823 & ~n48824 ;
  assign n48829 = ~n48196 & ~n48214 ;
  assign n48830 = ~n48190 & n48241 ;
  assign n48831 = ~n48829 & ~n48830 ;
  assign n48832 = ~n48177 & ~n48831 ;
  assign n48833 = n48190 & n48196 ;
  assign n48834 = n48211 & n48833 ;
  assign n48835 = ~n48217 & ~n48834 ;
  assign n48836 = n48177 & ~n48835 ;
  assign n48826 = n48183 & n48196 ;
  assign n48827 = ~n48211 & n48826 ;
  assign n48828 = n48190 & n48827 ;
  assign n48837 = ~n48251 & ~n48828 ;
  assign n48838 = ~n48836 & n48837 ;
  assign n48839 = ~n48832 & n48838 ;
  assign n48840 = ~n48204 & ~n48839 ;
  assign n48842 = ~n48190 & n48211 ;
  assign n48843 = n48196 & n48842 ;
  assign n48844 = ~n48183 & ~n48843 ;
  assign n48841 = n48183 & ~n48227 ;
  assign n48845 = n48177 & ~n48841 ;
  assign n48846 = ~n48844 & n48845 ;
  assign n48849 = ~n48226 & ~n48237 ;
  assign n48850 = ~n48183 & n48190 ;
  assign n48851 = n48219 & n48850 ;
  assign n48852 = n48849 & ~n48851 ;
  assign n48853 = n48177 & ~n48852 ;
  assign n48854 = ~n48177 & ~n48850 ;
  assign n48855 = n48849 & n48854 ;
  assign n48847 = n48241 & n48833 ;
  assign n48848 = n48211 & n48826 ;
  assign n48856 = ~n48847 & ~n48848 ;
  assign n48857 = ~n48855 & n48856 ;
  assign n48858 = ~n48853 & n48857 ;
  assign n48859 = n48204 & ~n48858 ;
  assign n48860 = ~n48846 & ~n48859 ;
  assign n48861 = ~n48840 & n48860 ;
  assign n48862 = ~\u1_L0_reg[17]/NET0131  & ~n48861 ;
  assign n48863 = \u1_L0_reg[17]/NET0131  & n48861 ;
  assign n48864 = ~n48862 & ~n48863 ;
  assign n48868 = ~n47898 & ~n48772 ;
  assign n48869 = n47898 & n48782 ;
  assign n48865 = ~n47898 & ~n47927 ;
  assign n48866 = n47905 & ~n47964 ;
  assign n48867 = ~n48865 & n48866 ;
  assign n48870 = ~n47926 & ~n48867 ;
  assign n48871 = ~n48869 & n48870 ;
  assign n48872 = ~n48868 & n48871 ;
  assign n48877 = ~n47905 & n48765 ;
  assign n48876 = ~n47898 & n47952 ;
  assign n48873 = ~n47892 & n47955 ;
  assign n48878 = n47926 & ~n48873 ;
  assign n48879 = ~n48876 & n48878 ;
  assign n48880 = ~n48877 & n48879 ;
  assign n48874 = ~n47950 & ~n47965 ;
  assign n48875 = n47898 & ~n48874 ;
  assign n48881 = ~n48704 & ~n48875 ;
  assign n48882 = n48880 & n48881 ;
  assign n48883 = ~n48872 & ~n48882 ;
  assign n48884 = ~n47939 & ~n47976 ;
  assign n48885 = ~n48883 & n48884 ;
  assign n48886 = ~\u1_L0_reg[19]/NET0131  & ~n48885 ;
  assign n48887 = \u1_L0_reg[19]/NET0131  & n48885 ;
  assign n48888 = ~n48886 & ~n48887 ;
  assign n48889 = n48110 & n48157 ;
  assign n48890 = ~n48148 & ~n48153 ;
  assign n48891 = ~n48889 & n48890 ;
  assign n48892 = ~n48092 & ~n48891 ;
  assign n48893 = ~n48110 & ~n48454 ;
  assign n48894 = n48092 & ~n48554 ;
  assign n48895 = ~n48893 & n48894 ;
  assign n48896 = ~n48119 & ~n48536 ;
  assign n48897 = ~n48154 & n48896 ;
  assign n48898 = ~n48895 & n48897 ;
  assign n48899 = ~n48892 & n48898 ;
  assign n48900 = n48086 & ~n48899 ;
  assign n48901 = n48092 & ~n48454 ;
  assign n48902 = ~n48144 & n48901 ;
  assign n48903 = ~n48140 & ~n48902 ;
  assign n48904 = ~n48086 & ~n48903 ;
  assign n48907 = ~n48092 & n48146 ;
  assign n48905 = ~n48133 & n48439 ;
  assign n48906 = ~n48143 & n48905 ;
  assign n48908 = n48441 & n48548 ;
  assign n48909 = ~n48165 & ~n48908 ;
  assign n48910 = ~n48906 & n48909 ;
  assign n48911 = ~n48907 & n48910 ;
  assign n48912 = ~n48904 & n48911 ;
  assign n48913 = ~n48900 & n48912 ;
  assign n48914 = ~\u1_L0_reg[27]/NET0131  & ~n48913 ;
  assign n48915 = \u1_L0_reg[27]/NET0131  & n48913 ;
  assign n48916 = ~n48914 & ~n48915 ;
  assign n48919 = ~n47810 & n47842 ;
  assign n48920 = ~n47810 & n48294 ;
  assign n48921 = ~n47844 & ~n47863 ;
  assign n48922 = ~n48920 & ~n48921 ;
  assign n48923 = ~n48919 & ~n48922 ;
  assign n48924 = ~n47834 & ~n48923 ;
  assign n48917 = n47823 & n47836 ;
  assign n48918 = n47810 & n48917 ;
  assign n48925 = ~n47817 & n47871 ;
  assign n48926 = ~n47872 & ~n48917 ;
  assign n48927 = ~n48925 & n48926 ;
  assign n48928 = n47834 & ~n48927 ;
  assign n48929 = ~n48918 & ~n48928 ;
  assign n48930 = ~n48924 & n48929 ;
  assign n48931 = n47798 & ~n48930 ;
  assign n48933 = ~n47842 & ~n48300 ;
  assign n48934 = n47810 & ~n48933 ;
  assign n48938 = n47870 & ~n48934 ;
  assign n48935 = ~n47857 & ~n48300 ;
  assign n48936 = n47834 & ~n48935 ;
  assign n48937 = n48299 & ~n48300 ;
  assign n48939 = ~n48936 & ~n48937 ;
  assign n48940 = n48938 & n48939 ;
  assign n48941 = ~n47798 & ~n48940 ;
  assign n48932 = n47843 & n48301 ;
  assign n48942 = ~n47836 & n47854 ;
  assign n48943 = n47826 & n48942 ;
  assign n48944 = ~n48932 & ~n48943 ;
  assign n48945 = ~n48941 & n48944 ;
  assign n48946 = ~n48931 & n48945 ;
  assign n48947 = \u1_L0_reg[32]/NET0131  & n48946 ;
  assign n48948 = ~\u1_L0_reg[32]/NET0131  & ~n48946 ;
  assign n48949 = ~n48947 & ~n48948 ;
  assign n48984 = decrypt_pad & ~\u1_uk_K_r0_reg[41]/NET0131  ;
  assign n48985 = ~decrypt_pad & ~\u1_uk_K_r0_reg[20]/NET0131  ;
  assign n48986 = ~n48984 & ~n48985 ;
  assign n48987 = \u1_R0_reg[11]/NET0131  & ~n48986 ;
  assign n48988 = ~\u1_R0_reg[11]/NET0131  & n48986 ;
  assign n48989 = ~n48987 & ~n48988 ;
  assign n48950 = decrypt_pad & ~\u1_uk_K_r0_reg[24]/NET0131  ;
  assign n48951 = ~decrypt_pad & ~\u1_uk_K_r0_reg[3]/NET0131  ;
  assign n48952 = ~n48950 & ~n48951 ;
  assign n48953 = \u1_R0_reg[12]/NET0131  & ~n48952 ;
  assign n48954 = ~\u1_R0_reg[12]/NET0131  & n48952 ;
  assign n48955 = ~n48953 & ~n48954 ;
  assign n48963 = decrypt_pad & ~\u1_uk_K_r0_reg[12]/NET0131  ;
  assign n48964 = ~decrypt_pad & ~\u1_uk_K_r0_reg[48]/NET0131  ;
  assign n48965 = ~n48963 & ~n48964 ;
  assign n48966 = \u1_R0_reg[13]/NET0131  & ~n48965 ;
  assign n48967 = ~\u1_R0_reg[13]/NET0131  & n48965 ;
  assign n48968 = ~n48966 & ~n48967 ;
  assign n48976 = decrypt_pad & ~\u1_uk_K_r0_reg[32]/NET0131  ;
  assign n48977 = ~decrypt_pad & ~\u1_uk_K_r0_reg[11]/NET0131  ;
  assign n48978 = ~n48976 & ~n48977 ;
  assign n48979 = \u1_R0_reg[9]/NET0131  & ~n48978 ;
  assign n48980 = ~\u1_R0_reg[9]/NET0131  & n48978 ;
  assign n48981 = ~n48979 & ~n48980 ;
  assign n48992 = n48968 & ~n48981 ;
  assign n48956 = decrypt_pad & ~\u1_uk_K_r0_reg[40]/NET0131  ;
  assign n48957 = ~decrypt_pad & ~\u1_uk_K_r0_reg[19]/NET0131  ;
  assign n48958 = ~n48956 & ~n48957 ;
  assign n48959 = \u1_R0_reg[10]/NET0131  & ~n48958 ;
  assign n48960 = ~\u1_R0_reg[10]/NET0131  & n48958 ;
  assign n48961 = ~n48959 & ~n48960 ;
  assign n48969 = decrypt_pad & ~\u1_uk_K_r0_reg[3]/NET0131  ;
  assign n48970 = ~decrypt_pad & ~\u1_uk_K_r0_reg[39]/NET0131  ;
  assign n48971 = ~n48969 & ~n48970 ;
  assign n48972 = \u1_R0_reg[8]/NET0131  & ~n48971 ;
  assign n48973 = ~\u1_R0_reg[8]/NET0131  & n48971 ;
  assign n48974 = ~n48972 & ~n48973 ;
  assign n48993 = n48968 & ~n48974 ;
  assign n48994 = n48961 & n48993 ;
  assign n48995 = ~n48968 & n48974 ;
  assign n48996 = n48981 & n48995 ;
  assign n48997 = ~n48994 & ~n48996 ;
  assign n48998 = ~n48992 & n48997 ;
  assign n48999 = n48955 & ~n48998 ;
  assign n48975 = ~n48968 & ~n48974 ;
  assign n48990 = ~n48961 & ~n48981 ;
  assign n48991 = n48975 & n48990 ;
  assign n49000 = n48961 & ~n48981 ;
  assign n49001 = n48968 & n49000 ;
  assign n49002 = ~n48991 & ~n49001 ;
  assign n49003 = ~n48999 & n49002 ;
  assign n49004 = n48989 & ~n49003 ;
  assign n49007 = ~n48961 & n48981 ;
  assign n49008 = ~n49000 & ~n49007 ;
  assign n49005 = n48968 & n48974 ;
  assign n49006 = ~n48975 & ~n49005 ;
  assign n49009 = ~n48974 & n48989 ;
  assign n49013 = n49006 & ~n49009 ;
  assign n49014 = n49008 & ~n49013 ;
  assign n49010 = ~n48961 & n49009 ;
  assign n49011 = n49006 & ~n49008 ;
  assign n49012 = ~n49010 & n49011 ;
  assign n49015 = ~n48955 & ~n49012 ;
  assign n49016 = ~n49014 & n49015 ;
  assign n48962 = n48955 & n48961 ;
  assign n48982 = n48975 & n48981 ;
  assign n48983 = n48962 & n48982 ;
  assign n49017 = n48974 & ~n48992 ;
  assign n49018 = ~n49007 & ~n49017 ;
  assign n49019 = ~n48968 & n48981 ;
  assign n49020 = n48955 & ~n48989 ;
  assign n49021 = ~n49019 & n49020 ;
  assign n49022 = ~n49018 & n49021 ;
  assign n49023 = ~n48983 & ~n49022 ;
  assign n49024 = ~n49016 & n49023 ;
  assign n49025 = ~n49004 & n49024 ;
  assign n49026 = ~\u1_L0_reg[6]/NET0131  & ~n49025 ;
  assign n49027 = \u1_L0_reg[6]/NET0131  & n49025 ;
  assign n49028 = ~n49026 & ~n49027 ;
  assign n49030 = ~n47817 & ~n48295 ;
  assign n49029 = n47810 & ~n48294 ;
  assign n49031 = ~n48917 & ~n49029 ;
  assign n49032 = ~n49030 & n49031 ;
  assign n49033 = ~n47834 & ~n49032 ;
  assign n49037 = ~n47857 & ~n49029 ;
  assign n49038 = n47823 & ~n49037 ;
  assign n49034 = ~n47823 & n48294 ;
  assign n49035 = ~n47871 & n49034 ;
  assign n49036 = n47834 & n49035 ;
  assign n49039 = n47798 & ~n49036 ;
  assign n49040 = ~n49038 & n49039 ;
  assign n49041 = ~n49033 & n49040 ;
  assign n49042 = n47868 & ~n48294 ;
  assign n49043 = n47834 & ~n47857 ;
  assign n49044 = ~n49034 & n49043 ;
  assign n49045 = ~n49042 & n49044 ;
  assign n49046 = ~n47798 & ~n49045 ;
  assign n49047 = ~n49041 & ~n49046 ;
  assign n49048 = ~n47834 & n49038 ;
  assign n49049 = ~n47834 & n49035 ;
  assign n49050 = ~n47845 & ~n49049 ;
  assign n49051 = n47798 & ~n47834 ;
  assign n49052 = ~n49050 & ~n49051 ;
  assign n49053 = ~n49048 & ~n49052 ;
  assign n49054 = ~n49047 & n49053 ;
  assign n49055 = ~\u1_L0_reg[7]/NET0131  & ~n49054 ;
  assign n49056 = \u1_L0_reg[7]/NET0131  & n49054 ;
  assign n49057 = ~n49055 & ~n49056 ;
  assign n49058 = n48337 & ~n48349 ;
  assign n49059 = ~n48351 & ~n48408 ;
  assign n49060 = ~n49058 & n49059 ;
  assign n49061 = ~n48370 & ~n49060 ;
  assign n49062 = ~n48360 & ~n48403 ;
  assign n49063 = n48370 & ~n49062 ;
  assign n49064 = ~n48353 & n48589 ;
  assign n49065 = ~n49063 & n49064 ;
  assign n49066 = ~n49061 & n49065 ;
  assign n49067 = ~n48390 & ~n49066 ;
  assign n49068 = n48359 & n48379 ;
  assign n49069 = ~n48351 & ~n49068 ;
  assign n49070 = n48370 & ~n49069 ;
  assign n49071 = n48349 & n48407 ;
  assign n49072 = ~n49070 & ~n49071 ;
  assign n49073 = ~n48419 & n49072 ;
  assign n49074 = n48390 & ~n49073 ;
  assign n49075 = ~n48370 & n48401 ;
  assign n49076 = n48343 & n49058 ;
  assign n49077 = n48418 & ~n49076 ;
  assign n49078 = n48370 & ~n49077 ;
  assign n49079 = ~n49075 & ~n49078 ;
  assign n49080 = ~n49074 & n49079 ;
  assign n49081 = ~n49067 & n49080 ;
  assign n49082 = ~\u1_L0_reg[8]/NET0131  & ~n49081 ;
  assign n49083 = \u1_L0_reg[8]/NET0131  & n49081 ;
  assign n49084 = ~n49082 & ~n49083 ;
  assign n49095 = n48981 & n49005 ;
  assign n49096 = ~n48981 & n48993 ;
  assign n49097 = ~n49095 & ~n49096 ;
  assign n49110 = ~n48961 & n48975 ;
  assign n49111 = n49097 & ~n49110 ;
  assign n49112 = ~n48989 & ~n49111 ;
  assign n49113 = ~n48981 & ~n49005 ;
  assign n49114 = ~n48975 & n48989 ;
  assign n49115 = ~n49095 & n49114 ;
  assign n49116 = ~n49113 & n49115 ;
  assign n49117 = ~n48991 & ~n49116 ;
  assign n49118 = ~n49112 & n49117 ;
  assign n49119 = ~n48955 & ~n49118 ;
  assign n49098 = ~n48981 & n48995 ;
  assign n49099 = n49009 & n49019 ;
  assign n49100 = ~n49098 & ~n49099 ;
  assign n49101 = n49097 & n49100 ;
  assign n49102 = ~n48961 & ~n49101 ;
  assign n49088 = n48981 & n48993 ;
  assign n49089 = n48961 & n49088 ;
  assign n49090 = n48961 & n48975 ;
  assign n49091 = ~n48961 & n48974 ;
  assign n49092 = ~n48968 & n49091 ;
  assign n49093 = ~n49090 & ~n49092 ;
  assign n49094 = ~n48989 & ~n49093 ;
  assign n49103 = ~n49089 & ~n49094 ;
  assign n49104 = ~n49102 & n49103 ;
  assign n49105 = n48955 & ~n49104 ;
  assign n49085 = n48961 & n48974 ;
  assign n49086 = ~n48981 & n49085 ;
  assign n49087 = ~n48989 & n49086 ;
  assign n49106 = n49019 & n49085 ;
  assign n49107 = ~n48981 & n49090 ;
  assign n49108 = ~n49106 & ~n49107 ;
  assign n49109 = n48989 & ~n49108 ;
  assign n49120 = ~n49087 & ~n49109 ;
  assign n49121 = ~n49105 & n49120 ;
  assign n49122 = ~n49119 & n49121 ;
  assign n49123 = ~\u1_L0_reg[16]/NET0131  & ~n49122 ;
  assign n49124 = \u1_L0_reg[16]/NET0131  & n49122 ;
  assign n49125 = ~n49123 & ~n49124 ;
  assign n49142 = ~n48219 & ~n48227 ;
  assign n49143 = ~n48190 & ~n49142 ;
  assign n49144 = ~n48218 & ~n49143 ;
  assign n49145 = ~n48177 & ~n49144 ;
  assign n49146 = n48177 & ~n48241 ;
  assign n49147 = n48215 & n49146 ;
  assign n49148 = ~n48255 & ~n48851 ;
  assign n49149 = ~n49147 & n49148 ;
  assign n49150 = ~n49145 & n49149 ;
  assign n49151 = n48204 & ~n49150 ;
  assign n49133 = ~n48248 & ~n48833 ;
  assign n49134 = ~n48177 & ~n49133 ;
  assign n49135 = n48177 & n48227 ;
  assign n49136 = n48205 & n48842 ;
  assign n49137 = ~n48234 & ~n48848 ;
  assign n49138 = ~n49136 & n49137 ;
  assign n49139 = ~n49135 & n49138 ;
  assign n49140 = ~n49134 & n49139 ;
  assign n49141 = ~n48204 & ~n49140 ;
  assign n49126 = ~n48197 & ~n48227 ;
  assign n49127 = n48184 & ~n49126 ;
  assign n49129 = n48213 & n48826 ;
  assign n49128 = n48219 & n48220 ;
  assign n49130 = ~n48847 & ~n49128 ;
  assign n49131 = ~n49129 & n49130 ;
  assign n49132 = ~n48177 & ~n49131 ;
  assign n49152 = ~n49127 & ~n49132 ;
  assign n49153 = ~n49141 & n49152 ;
  assign n49154 = ~n49151 & n49153 ;
  assign n49155 = \u1_L0_reg[23]/NET0131  & ~n49154 ;
  assign n49156 = ~\u1_L0_reg[23]/NET0131  & n49154 ;
  assign n49157 = ~n49155 & ~n49156 ;
  assign n49173 = ~n48961 & n48993 ;
  assign n49174 = ~n49090 & ~n49173 ;
  assign n49175 = ~n48982 & ~n49086 ;
  assign n49176 = n49174 & n49175 ;
  assign n49177 = n48989 & ~n49176 ;
  assign n49178 = n48961 & n49098 ;
  assign n49179 = ~n49177 & ~n49178 ;
  assign n49180 = ~n48955 & ~n49179 ;
  assign n49160 = ~n48989 & ~n48990 ;
  assign n49161 = ~n48995 & n49160 ;
  assign n49162 = ~n48961 & n48989 ;
  assign n49163 = ~n48981 & n49162 ;
  assign n49164 = ~n49161 & ~n49163 ;
  assign n49165 = ~n48993 & ~n49164 ;
  assign n49166 = n48990 & n49013 ;
  assign n49167 = n48981 & n49085 ;
  assign n49168 = ~n48994 & ~n49167 ;
  assign n49169 = n48989 & ~n49168 ;
  assign n49170 = ~n49166 & ~n49169 ;
  assign n49171 = ~n49165 & n49170 ;
  assign n49172 = n48955 & ~n49171 ;
  assign n49183 = n48990 & ~n49006 ;
  assign n49184 = n48997 & ~n49183 ;
  assign n49185 = ~n48955 & ~n48989 ;
  assign n49186 = ~n49184 & n49185 ;
  assign n49158 = n48961 & ~n48989 ;
  assign n49159 = n49095 & n49158 ;
  assign n49181 = ~n49088 & ~n49098 ;
  assign n49182 = n49162 & ~n49181 ;
  assign n49187 = ~n49159 & ~n49182 ;
  assign n49188 = ~n49186 & n49187 ;
  assign n49189 = ~n49172 & n49188 ;
  assign n49190 = ~n49180 & n49189 ;
  assign n49191 = ~\u1_L0_reg[24]/NET0131  & ~n49190 ;
  assign n49192 = \u1_L0_reg[24]/NET0131  & n49190 ;
  assign n49193 = ~n49191 & ~n49192 ;
  assign n49194 = ~n48961 & n49098 ;
  assign n49195 = n48989 & n49174 ;
  assign n49196 = ~n49194 & n49195 ;
  assign n49197 = ~n48989 & ~n49085 ;
  assign n49198 = ~n48982 & n49197 ;
  assign n49199 = ~n49196 & ~n49198 ;
  assign n49200 = n48955 & ~n49199 ;
  assign n49203 = ~n48968 & n49007 ;
  assign n49202 = ~n49019 & n49085 ;
  assign n49204 = n48989 & ~n49202 ;
  assign n49205 = ~n49203 & n49204 ;
  assign n49206 = ~n49019 & n49091 ;
  assign n49207 = ~n48989 & ~n49088 ;
  assign n49208 = ~n49206 & n49207 ;
  assign n49209 = ~n49205 & ~n49208 ;
  assign n49201 = n48993 & n49000 ;
  assign n49210 = ~n48955 & ~n49201 ;
  assign n49211 = ~n49183 & n49210 ;
  assign n49212 = ~n49209 & n49211 ;
  assign n49213 = ~n49200 & ~n49212 ;
  assign n49217 = n48962 & n48981 ;
  assign n49218 = ~n49005 & n49217 ;
  assign n49214 = n49019 & n49158 ;
  assign n49215 = n48989 & n49000 ;
  assign n49216 = n49005 & n49215 ;
  assign n49219 = ~n49214 & ~n49216 ;
  assign n49220 = ~n49218 & n49219 ;
  assign n49221 = ~n49213 & n49220 ;
  assign n49222 = \u1_L0_reg[30]/NET0131  & ~n49221 ;
  assign n49223 = ~\u1_L0_reg[30]/NET0131  & n49221 ;
  assign n49224 = ~n49222 & ~n49223 ;
  assign n49225 = n48390 & ~n48401 ;
  assign n49226 = ~n48362 & n49225 ;
  assign n49227 = ~n48408 & n49226 ;
  assign n49228 = ~n48358 & n48400 ;
  assign n49229 = ~n48390 & ~n49228 ;
  assign n49230 = ~n48376 & ~n48379 ;
  assign n49231 = ~n48351 & n49230 ;
  assign n49232 = n49229 & n49231 ;
  assign n49233 = ~n49227 & ~n49232 ;
  assign n49234 = n48350 & n48376 ;
  assign n49235 = ~n48370 & ~n49068 ;
  assign n49236 = ~n49234 & n49235 ;
  assign n49237 = ~n48406 & n49236 ;
  assign n49238 = ~n49233 & n49237 ;
  assign n49239 = n48343 & n48379 ;
  assign n49240 = ~n48394 & ~n49239 ;
  assign n49241 = n49226 & n49240 ;
  assign n49242 = ~n48393 & ~n49058 ;
  assign n49243 = n49229 & n49242 ;
  assign n49244 = ~n49241 & ~n49243 ;
  assign n49245 = ~n48360 & n48370 ;
  assign n49246 = ~n48417 & n49245 ;
  assign n49247 = ~n49244 & n49246 ;
  assign n49248 = ~n49238 & ~n49247 ;
  assign n49249 = ~\u1_L0_reg[3]/NET0131  & n49248 ;
  assign n49250 = \u1_L0_reg[3]/NET0131  & ~n49248 ;
  assign n49251 = ~n49249 & ~n49250 ;
  assign n49253 = ~n48827 & n49142 ;
  assign n49254 = n48177 & ~n49253 ;
  assign n49255 = ~n48233 & ~n48843 ;
  assign n49256 = ~n48177 & ~n49255 ;
  assign n49252 = n48183 & n48829 ;
  assign n49257 = ~n48183 & n48834 ;
  assign n49258 = ~n49252 & ~n49257 ;
  assign n49259 = ~n49256 & n49258 ;
  assign n49260 = ~n49254 & n49259 ;
  assign n49261 = ~n48204 & ~n49260 ;
  assign n49262 = ~n48190 & n48848 ;
  assign n49263 = ~n49257 & ~n49262 ;
  assign n49264 = ~n48177 & ~n49263 ;
  assign n49266 = n48183 & ~n48215 ;
  assign n49267 = ~n48829 & n49266 ;
  assign n49265 = n48184 & ~n49255 ;
  assign n49268 = ~n48847 & ~n49265 ;
  assign n49269 = ~n49267 & n49268 ;
  assign n49270 = n48204 & ~n49269 ;
  assign n49271 = ~n49264 & ~n49270 ;
  assign n49272 = ~n49261 & n49271 ;
  assign n49273 = ~\u1_L0_reg[9]/NET0131  & ~n49272 ;
  assign n49274 = \u1_L0_reg[9]/NET0131  & n49272 ;
  assign n49275 = ~n49273 & ~n49274 ;
  assign n49285 = n48631 & n48727 ;
  assign n49286 = n48618 & n48638 ;
  assign n49287 = ~n48631 & ~n49286 ;
  assign n49288 = n48644 & n49287 ;
  assign n49289 = ~n48750 & ~n49288 ;
  assign n49290 = ~n49285 & n49289 ;
  assign n49291 = n48606 & ~n49290 ;
  assign n49279 = n48653 & ~n48726 ;
  assign n49277 = ~n48612 & ~n48739 ;
  assign n49278 = n48753 & n49277 ;
  assign n49280 = n48666 & n48739 ;
  assign n49281 = ~n48743 & ~n49280 ;
  assign n49282 = ~n49278 & n49281 ;
  assign n49283 = ~n49279 & n49282 ;
  assign n49284 = ~n48606 & ~n49283 ;
  assign n49276 = ~n48631 & n48649 ;
  assign n49292 = n48638 & n48666 ;
  assign n49293 = ~n48811 & ~n49292 ;
  assign n49294 = n48631 & ~n49293 ;
  assign n49295 = ~n49276 & ~n49294 ;
  assign n49296 = ~n49284 & n49295 ;
  assign n49297 = ~n49291 & n49296 ;
  assign n49298 = \u1_L0_reg[18]/NET0131  & n49297 ;
  assign n49299 = ~\u1_L0_reg[18]/NET0131  & ~n49297 ;
  assign n49300 = ~n49298 & ~n49299 ;
  assign n49301 = decrypt_pad & ~\u1_key_r_reg[13]/NET0131  ;
  assign n49302 = ~decrypt_pad & ~\u1_key_r_reg[6]/NET0131  ;
  assign n49303 = ~n49301 & ~n49302 ;
  assign n49304 = \u1_desIn_r_reg[31]/NET0131  & ~n49303 ;
  assign n49305 = ~\u1_desIn_r_reg[31]/NET0131  & n49303 ;
  assign n49306 = ~n49304 & ~n49305 ;
  assign n49326 = decrypt_pad & ~\u1_key_r_reg[47]/NET0131  ;
  assign n49327 = ~decrypt_pad & ~\u1_key_r_reg[40]/NET0131  ;
  assign n49328 = ~n49326 & ~n49327 ;
  assign n49329 = \u1_desIn_r_reg[57]/NET0131  & ~n49328 ;
  assign n49330 = ~\u1_desIn_r_reg[57]/NET0131  & n49328 ;
  assign n49331 = ~n49329 & ~n49330 ;
  assign n49335 = decrypt_pad & ~\u1_key_r_reg[11]/NET0131  ;
  assign n49336 = ~decrypt_pad & ~\u1_key_r_reg[4]/NET0131  ;
  assign n49337 = ~n49335 & ~n49336 ;
  assign n49338 = \u1_desIn_r_reg[7]/NET0131  & ~n49337 ;
  assign n49339 = ~\u1_desIn_r_reg[7]/NET0131  & n49337 ;
  assign n49340 = ~n49338 & ~n49339 ;
  assign n49307 = decrypt_pad & ~\u1_key_r_reg[26]/NET0131  ;
  assign n49308 = ~decrypt_pad & ~\u1_key_r_reg[19]/NET0131  ;
  assign n49309 = ~n49307 & ~n49308 ;
  assign n49310 = \u1_desIn_r_reg[15]/NET0131  & ~n49309 ;
  assign n49311 = ~\u1_desIn_r_reg[15]/NET0131  & n49309 ;
  assign n49312 = ~n49310 & ~n49311 ;
  assign n49320 = decrypt_pad & ~\u1_key_r_reg[41]/NET0131  ;
  assign n49321 = ~decrypt_pad & ~\u1_key_r_reg[34]/NET0131  ;
  assign n49322 = ~n49320 & ~n49321 ;
  assign n49323 = \u1_desIn_r_reg[39]/NET0131  & ~n49322 ;
  assign n49324 = ~\u1_desIn_r_reg[39]/NET0131  & n49322 ;
  assign n49325 = ~n49323 & ~n49324 ;
  assign n49368 = ~n49312 & ~n49325 ;
  assign n49369 = ~n49340 & n49368 ;
  assign n49370 = n49331 & ~n49369 ;
  assign n49333 = ~n49325 & ~n49331 ;
  assign n49313 = decrypt_pad & ~\u1_key_r_reg[3]/NET0131  ;
  assign n49314 = ~decrypt_pad & ~\u1_key_r_reg[53]/NET0131  ;
  assign n49315 = ~n49313 & ~n49314 ;
  assign n49316 = \u1_desIn_r_reg[23]/NET0131  & ~n49315 ;
  assign n49317 = ~\u1_desIn_r_reg[23]/NET0131  & n49315 ;
  assign n49318 = ~n49316 & ~n49317 ;
  assign n49366 = ~n49312 & n49318 ;
  assign n49367 = n49340 & ~n49366 ;
  assign n49371 = ~n49333 & ~n49367 ;
  assign n49372 = ~n49370 & n49371 ;
  assign n49349 = n49325 & ~n49340 ;
  assign n49359 = n49312 & ~n49331 ;
  assign n49360 = ~n49325 & n49359 ;
  assign n49361 = ~n49349 & ~n49360 ;
  assign n49362 = n49318 & ~n49361 ;
  assign n49363 = ~n49331 & n49340 ;
  assign n49343 = ~n49318 & n49340 ;
  assign n49364 = ~n49343 & ~n49359 ;
  assign n49365 = ~n49363 & ~n49364 ;
  assign n49373 = ~n49362 & ~n49365 ;
  assign n49374 = ~n49372 & n49373 ;
  assign n49375 = n49306 & ~n49374 ;
  assign n49350 = ~n49312 & ~n49331 ;
  assign n49351 = n49331 & ~n49340 ;
  assign n49352 = n49312 & n49351 ;
  assign n49353 = ~n49350 & ~n49352 ;
  assign n49354 = ~n49318 & ~n49349 ;
  assign n49355 = ~n49353 & n49354 ;
  assign n49319 = n49312 & n49318 ;
  assign n49332 = n49325 & n49331 ;
  assign n49334 = ~n49332 & ~n49333 ;
  assign n49341 = n49334 & n49340 ;
  assign n49342 = n49319 & n49341 ;
  assign n49344 = n49332 & ~n49343 ;
  assign n49345 = ~n49325 & n49340 ;
  assign n49346 = ~n49331 & n49345 ;
  assign n49347 = ~n49344 & ~n49346 ;
  assign n49348 = ~n49312 & ~n49347 ;
  assign n49356 = ~n49342 & ~n49348 ;
  assign n49357 = ~n49355 & n49356 ;
  assign n49358 = ~n49306 & ~n49357 ;
  assign n49376 = n49318 & ~n49340 ;
  assign n49377 = ~n49312 & n49331 ;
  assign n49378 = ~n49360 & ~n49377 ;
  assign n49379 = n49376 & ~n49378 ;
  assign n49381 = n49312 & n49325 ;
  assign n49382 = n49340 & n49381 ;
  assign n49383 = n49331 & n49382 ;
  assign n49380 = n49349 & n49359 ;
  assign n49384 = n49340 & n49368 ;
  assign n49385 = ~n49380 & ~n49384 ;
  assign n49386 = ~n49383 & n49385 ;
  assign n49387 = ~n49318 & ~n49386 ;
  assign n49388 = ~n49379 & ~n49387 ;
  assign n49389 = ~n49358 & n49388 ;
  assign n49390 = ~n49375 & n49389 ;
  assign n49391 = ~\u1_desIn_r_reg[48]/NET0131  & ~n49390 ;
  assign n49392 = \u1_desIn_r_reg[48]/NET0131  & n49390 ;
  assign n49393 = ~n49391 & ~n49392 ;
  assign n49416 = decrypt_pad & ~\u1_key_r_reg[9]/NET0131  ;
  assign n49417 = ~decrypt_pad & ~\u1_key_r_reg[2]/NET0131  ;
  assign n49418 = ~n49416 & ~n49417 ;
  assign n49419 = \u1_desIn_r_reg[51]/NET0131  & ~n49418 ;
  assign n49420 = ~\u1_desIn_r_reg[51]/NET0131  & n49418 ;
  assign n49421 = ~n49419 & ~n49420 ;
  assign n49448 = decrypt_pad & ~\u1_key_r_reg[35]/P0001  ;
  assign n49449 = ~decrypt_pad & ~\u1_key_r_reg[28]/NET0131  ;
  assign n49450 = ~n49448 & ~n49449 ;
  assign n49451 = \u1_desIn_r_reg[59]/NET0131  & ~n49450 ;
  assign n49452 = ~\u1_desIn_r_reg[59]/NET0131  & n49450 ;
  assign n49453 = ~n49451 & ~n49452 ;
  assign n49394 = decrypt_pad & ~\u1_key_r_reg[29]/NET0131  ;
  assign n49395 = ~decrypt_pad & ~\u1_key_r_reg[22]/NET0131  ;
  assign n49396 = ~n49394 & ~n49395 ;
  assign n49397 = \u1_desIn_r_reg[35]/NET0131  & ~n49396 ;
  assign n49398 = ~\u1_desIn_r_reg[35]/NET0131  & n49396 ;
  assign n49399 = ~n49397 & ~n49398 ;
  assign n49400 = decrypt_pad & ~\u1_key_r_reg[51]/NET0131  ;
  assign n49401 = ~decrypt_pad & ~\u1_key_r_reg[44]/NET0131  ;
  assign n49402 = ~n49400 & ~n49401 ;
  assign n49403 = \u1_desIn_r_reg[43]/NET0131  & ~n49402 ;
  assign n49404 = ~\u1_desIn_r_reg[43]/NET0131  & n49402 ;
  assign n49405 = ~n49403 & ~n49404 ;
  assign n49407 = decrypt_pad & ~\u1_key_r_reg[14]/NET0131  ;
  assign n49408 = ~decrypt_pad & ~\u1_key_r_reg[7]/NET0131  ;
  assign n49409 = ~n49407 & ~n49408 ;
  assign n49410 = \u1_desIn_r_reg[27]/NET0131  & ~n49409 ;
  assign n49411 = ~\u1_desIn_r_reg[27]/NET0131  & n49409 ;
  assign n49412 = ~n49410 & ~n49411 ;
  assign n49414 = n49405 & ~n49412 ;
  assign n49415 = n49399 & n49414 ;
  assign n49425 = decrypt_pad & ~\u1_key_r_reg[30]/NET0131  ;
  assign n49426 = ~decrypt_pad & ~\u1_key_r_reg[23]/NET0131  ;
  assign n49427 = ~n49425 & ~n49426 ;
  assign n49428 = \u1_desIn_r_reg[1]/NET0131  & ~n49427 ;
  assign n49429 = ~\u1_desIn_r_reg[1]/NET0131  & n49427 ;
  assign n49430 = ~n49428 & ~n49429 ;
  assign n49457 = n49399 & n49430 ;
  assign n49468 = ~n49399 & ~n49430 ;
  assign n49469 = ~n49405 & n49468 ;
  assign n49470 = ~n49457 & ~n49469 ;
  assign n49471 = n49412 & ~n49470 ;
  assign n49472 = ~n49415 & ~n49471 ;
  assign n49473 = n49453 & ~n49472 ;
  assign n49474 = ~n49399 & n49430 ;
  assign n49475 = ~n49412 & n49474 ;
  assign n49476 = ~n49405 & n49475 ;
  assign n49437 = n49412 & n49430 ;
  assign n49438 = n49405 & n49437 ;
  assign n49406 = n49399 & ~n49405 ;
  assign n49444 = n49406 & ~n49430 ;
  assign n49467 = ~n49412 & n49444 ;
  assign n49477 = ~n49438 & ~n49467 ;
  assign n49478 = ~n49476 & n49477 ;
  assign n49479 = ~n49473 & n49478 ;
  assign n49480 = n49421 & ~n49479 ;
  assign n49413 = n49406 & n49412 ;
  assign n49422 = ~n49415 & ~n49421 ;
  assign n49423 = ~n49413 & n49422 ;
  assign n49431 = ~n49412 & ~n49430 ;
  assign n49432 = ~n49399 & ~n49431 ;
  assign n49433 = n49405 & n49432 ;
  assign n49424 = ~n49405 & ~n49412 ;
  assign n49434 = n49421 & ~n49424 ;
  assign n49435 = ~n49433 & n49434 ;
  assign n49436 = ~n49423 & ~n49435 ;
  assign n49439 = ~n49399 & n49438 ;
  assign n49440 = ~n49405 & ~n49421 ;
  assign n49441 = n49412 & ~n49430 ;
  assign n49442 = n49440 & n49441 ;
  assign n49443 = ~n49439 & ~n49442 ;
  assign n49445 = n49412 & n49444 ;
  assign n49446 = n49443 & ~n49445 ;
  assign n49447 = ~n49436 & n49446 ;
  assign n49454 = ~n49447 & ~n49453 ;
  assign n49458 = ~n49412 & n49457 ;
  assign n49455 = ~n49399 & n49412 ;
  assign n49456 = n49430 & n49455 ;
  assign n49459 = ~n49405 & ~n49456 ;
  assign n49460 = ~n49458 & n49459 ;
  assign n49461 = ~n49438 & n49453 ;
  assign n49462 = n49422 & n49461 ;
  assign n49463 = ~n49460 & n49462 ;
  assign n49464 = n49399 & ~n49441 ;
  assign n49465 = ~n49432 & n49440 ;
  assign n49466 = ~n49464 & n49465 ;
  assign n49481 = ~n49463 & ~n49466 ;
  assign n49482 = ~n49454 & n49481 ;
  assign n49483 = ~n49480 & n49482 ;
  assign n49484 = \u1_desIn_r_reg[20]/NET0131  & ~n49483 ;
  assign n49485 = ~\u1_desIn_r_reg[20]/NET0131  & n49483 ;
  assign n49486 = ~n49484 & ~n49485 ;
  assign n49487 = decrypt_pad & ~\u1_key_r_reg[22]/NET0131  ;
  assign n49488 = ~decrypt_pad & ~\u1_key_r_reg[15]/NET0131  ;
  assign n49489 = ~n49487 & ~n49488 ;
  assign n49490 = \u1_desIn_r_reg[9]/NET0131  & ~n49489 ;
  assign n49491 = ~\u1_desIn_r_reg[9]/NET0131  & n49489 ;
  assign n49492 = ~n49490 & ~n49491 ;
  assign n49493 = decrypt_pad & ~\u1_key_r_reg[37]/NET0131  ;
  assign n49494 = ~decrypt_pad & ~\u1_key_r_reg[30]/NET0131  ;
  assign n49495 = ~n49493 & ~n49494 ;
  assign n49496 = \u1_desIn_r_reg[1]/NET0131  & ~n49495 ;
  assign n49497 = ~\u1_desIn_r_reg[1]/NET0131  & n49495 ;
  assign n49498 = ~n49496 & ~n49497 ;
  assign n49499 = n49492 & ~n49498 ;
  assign n49500 = decrypt_pad & ~\u1_key_r_reg[2]/NET0131  ;
  assign n49501 = ~decrypt_pad & ~\u1_key_r_reg[50]/NET0131  ;
  assign n49502 = ~n49500 & ~n49501 ;
  assign n49503 = \u1_desIn_r_reg[59]/NET0131  & ~n49502 ;
  assign n49504 = ~\u1_desIn_r_reg[59]/NET0131  & n49502 ;
  assign n49505 = ~n49503 & ~n49504 ;
  assign n49506 = decrypt_pad & ~\u1_key_r_reg[38]/NET0131  ;
  assign n49507 = ~decrypt_pad & ~\u1_key_r_reg[31]/NET0131  ;
  assign n49508 = ~n49506 & ~n49507 ;
  assign n49509 = \u1_desIn_r_reg[33]/NET0131  & ~n49508 ;
  assign n49510 = ~\u1_desIn_r_reg[33]/NET0131  & n49508 ;
  assign n49511 = ~n49509 & ~n49510 ;
  assign n49512 = ~n49505 & n49511 ;
  assign n49513 = n49499 & n49512 ;
  assign n49514 = ~n49505 & ~n49511 ;
  assign n49515 = n49492 & n49498 ;
  assign n49516 = n49514 & n49515 ;
  assign n49517 = ~n49513 & ~n49516 ;
  assign n49518 = ~n49498 & ~n49511 ;
  assign n49519 = n49498 & n49511 ;
  assign n49520 = ~n49492 & n49519 ;
  assign n49521 = ~n49499 & ~n49520 ;
  assign n49522 = decrypt_pad & ~\u1_key_r_reg[42]/P0001  ;
  assign n49523 = ~decrypt_pad & ~\u1_key_r_reg[35]/P0001  ;
  assign n49524 = ~n49522 & ~n49523 ;
  assign n49525 = \u1_desIn_r_reg[25]/NET0131  & ~n49524 ;
  assign n49526 = ~\u1_desIn_r_reg[25]/NET0131  & n49524 ;
  assign n49527 = ~n49525 & ~n49526 ;
  assign n49528 = ~n49521 & n49527 ;
  assign n49529 = ~n49518 & ~n49528 ;
  assign n49530 = n49505 & ~n49529 ;
  assign n49531 = n49517 & ~n49530 ;
  assign n49532 = decrypt_pad & ~\u1_key_r_reg[0]/NET0131  ;
  assign n49533 = ~decrypt_pad & ~\u1_key_r_reg[52]/NET0131  ;
  assign n49534 = ~n49532 & ~n49533 ;
  assign n49535 = \u1_desIn_r_reg[17]/NET0131  & ~n49534 ;
  assign n49536 = ~\u1_desIn_r_reg[17]/NET0131  & n49534 ;
  assign n49537 = ~n49535 & ~n49536 ;
  assign n49538 = ~n49531 & n49537 ;
  assign n49539 = ~n49498 & n49537 ;
  assign n49540 = ~n49492 & n49539 ;
  assign n49541 = ~n49492 & n49511 ;
  assign n49542 = ~n49499 & ~n49537 ;
  assign n49543 = ~n49541 & n49542 ;
  assign n49544 = ~n49540 & ~n49543 ;
  assign n49545 = n49505 & ~n49544 ;
  assign n49546 = ~n49505 & n49518 ;
  assign n49547 = n49492 & n49546 ;
  assign n49548 = ~n49537 & n49547 ;
  assign n49549 = ~n49492 & ~n49505 ;
  assign n49550 = n49492 & n49505 ;
  assign n49551 = ~n49549 & ~n49550 ;
  assign n49552 = n49511 & ~n49539 ;
  assign n49553 = ~n49551 & n49552 ;
  assign n49554 = ~n49548 & ~n49553 ;
  assign n49555 = ~n49545 & n49554 ;
  assign n49556 = ~n49527 & ~n49555 ;
  assign n49560 = n49505 & n49511 ;
  assign n49561 = ~n49492 & ~n49498 ;
  assign n49562 = n49560 & n49561 ;
  assign n49563 = n49498 & n49512 ;
  assign n49564 = ~n49562 & ~n49563 ;
  assign n49565 = ~n49537 & ~n49564 ;
  assign n49566 = n49518 & n49549 ;
  assign n49567 = ~n49513 & ~n49566 ;
  assign n49568 = ~n49565 & n49567 ;
  assign n49569 = n49527 & ~n49568 ;
  assign n49557 = n49498 & ~n49537 ;
  assign n49558 = ~n49551 & n49557 ;
  assign n49559 = ~n49511 & n49540 ;
  assign n49570 = ~n49558 & ~n49559 ;
  assign n49571 = ~n49569 & n49570 ;
  assign n49572 = ~n49556 & n49571 ;
  assign n49573 = ~n49538 & n49572 ;
  assign n49574 = ~\u1_desIn_r_reg[42]/NET0131  & ~n49573 ;
  assign n49575 = \u1_desIn_r_reg[42]/NET0131  & n49573 ;
  assign n49576 = ~n49574 & ~n49575 ;
  assign n49582 = ~n49334 & ~n49340 ;
  assign n49583 = ~n49325 & n49350 ;
  assign n49584 = ~n49582 & ~n49583 ;
  assign n49585 = ~n49318 & ~n49584 ;
  assign n49577 = ~n49345 & ~n49349 ;
  assign n49578 = n49318 & n49577 ;
  assign n49579 = n49312 & n49345 ;
  assign n49580 = ~n49578 & ~n49579 ;
  assign n49581 = n49331 & ~n49580 ;
  assign n49586 = ~n49306 & ~n49380 ;
  assign n49587 = ~n49581 & n49586 ;
  assign n49588 = ~n49585 & n49587 ;
  assign n49589 = ~n49359 & ~n49363 ;
  assign n49592 = n49349 & n49377 ;
  assign n49593 = n49589 & ~n49592 ;
  assign n49594 = n49318 & ~n49593 ;
  assign n49595 = n49331 & n49384 ;
  assign n49590 = ~n49318 & ~n49377 ;
  assign n49591 = n49589 & n49590 ;
  assign n49596 = n49306 & ~n49382 ;
  assign n49597 = ~n49591 & n49596 ;
  assign n49598 = ~n49595 & n49597 ;
  assign n49599 = ~n49594 & n49598 ;
  assign n49600 = ~n49588 & ~n49599 ;
  assign n49602 = n49340 & ~n49368 ;
  assign n49601 = n49318 & ~n49331 ;
  assign n49603 = ~n49381 & n49601 ;
  assign n49604 = n49602 & n49603 ;
  assign n49605 = ~n49600 & ~n49604 ;
  assign n49606 = ~\u1_desIn_r_reg[2]/NET0131  & ~n49605 ;
  assign n49607 = \u1_desIn_r_reg[2]/NET0131  & n49605 ;
  assign n49608 = ~n49606 & ~n49607 ;
  assign n49609 = n49399 & n49431 ;
  assign n49610 = ~n49406 & n49412 ;
  assign n49611 = ~n49609 & ~n49610 ;
  assign n49612 = ~n49476 & n49611 ;
  assign n49613 = n49421 & ~n49612 ;
  assign n49615 = ~n49457 & ~n49468 ;
  assign n49616 = ~n49412 & ~n49421 ;
  assign n49617 = ~n49615 & n49616 ;
  assign n49614 = n49399 & n49438 ;
  assign n49618 = ~n49453 & ~n49614 ;
  assign n49619 = ~n49617 & n49618 ;
  assign n49620 = ~n49613 & n49619 ;
  assign n49623 = ~n49413 & ~n49475 ;
  assign n49624 = n49421 & ~n49623 ;
  assign n49621 = ~n49421 & n49455 ;
  assign n49625 = ~n49444 & n49453 ;
  assign n49626 = ~n49621 & n49625 ;
  assign n49622 = n49414 & ~n49615 ;
  assign n49627 = ~n49476 & ~n49622 ;
  assign n49628 = n49626 & n49627 ;
  assign n49629 = ~n49624 & n49628 ;
  assign n49630 = ~n49620 & ~n49629 ;
  assign n49631 = n49412 & n49440 ;
  assign n49632 = n49615 & n49631 ;
  assign n49633 = ~n49630 & ~n49632 ;
  assign n49634 = ~\u1_desIn_r_reg[18]/P0001  & ~n49633 ;
  assign n49635 = \u1_desIn_r_reg[18]/P0001  & n49633 ;
  assign n49636 = ~n49634 & ~n49635 ;
  assign n49637 = decrypt_pad & ~\u1_key_r_reg[55]/NET0131  ;
  assign n49638 = ~decrypt_pad & ~\u1_key_r_reg[48]/NET0131  ;
  assign n49639 = ~n49637 & ~n49638 ;
  assign n49640 = \u1_desIn_r_reg[37]/NET0131  & ~n49639 ;
  assign n49641 = ~\u1_desIn_r_reg[37]/NET0131  & n49639 ;
  assign n49642 = ~n49640 & ~n49641 ;
  assign n49650 = decrypt_pad & ~\u1_key_r_reg[4]/NET0131  ;
  assign n49651 = ~decrypt_pad & ~\u1_key_r_reg[54]/NET0131  ;
  assign n49652 = ~n49650 & ~n49651 ;
  assign n49653 = \u1_desIn_r_reg[29]/NET0131  & ~n49652 ;
  assign n49654 = ~\u1_desIn_r_reg[29]/NET0131  & n49652 ;
  assign n49655 = ~n49653 & ~n49654 ;
  assign n49689 = n49642 & ~n49655 ;
  assign n49690 = ~n49642 & n49655 ;
  assign n49691 = ~n49689 & ~n49690 ;
  assign n49643 = decrypt_pad & ~\u1_key_r_reg[32]/NET0131  ;
  assign n49644 = ~decrypt_pad & ~\u1_key_r_reg[25]/NET0131  ;
  assign n49645 = ~n49643 & ~n49644 ;
  assign n49646 = \u1_desIn_r_reg[53]/NET0131  & ~n49645 ;
  assign n49647 = ~\u1_desIn_r_reg[53]/NET0131  & n49645 ;
  assign n49648 = ~n49646 & ~n49647 ;
  assign n49667 = decrypt_pad & ~\u1_key_r_reg[24]/NET0131  ;
  assign n49668 = ~decrypt_pad & ~\u1_key_r_reg[17]/NET0131  ;
  assign n49669 = ~n49667 & ~n49668 ;
  assign n49670 = \u1_desIn_r_reg[45]/NET0131  & ~n49669 ;
  assign n49671 = ~\u1_desIn_r_reg[45]/NET0131  & n49669 ;
  assign n49672 = ~n49670 & ~n49671 ;
  assign n49692 = ~n49648 & ~n49672 ;
  assign n49693 = ~n49691 & n49692 ;
  assign n49656 = decrypt_pad & ~\u1_key_r_reg[20]/NET0131  ;
  assign n49657 = ~decrypt_pad & ~\u1_key_r_reg[13]/NET0131  ;
  assign n49658 = ~n49656 & ~n49657 ;
  assign n49659 = \u1_desIn_r_reg[3]/NET0131  & ~n49658 ;
  assign n49660 = ~\u1_desIn_r_reg[3]/NET0131  & n49658 ;
  assign n49661 = ~n49659 & ~n49660 ;
  assign n49680 = n49655 & ~n49661 ;
  assign n49681 = n49642 & n49648 ;
  assign n49682 = n49680 & n49681 ;
  assign n49649 = ~n49642 & n49648 ;
  assign n49662 = ~n49655 & n49661 ;
  assign n49663 = n49649 & n49662 ;
  assign n49683 = decrypt_pad & ~\u1_key_r_reg[40]/NET0131  ;
  assign n49684 = ~decrypt_pad & ~\u1_key_r_reg[33]/NET0131  ;
  assign n49685 = ~n49683 & ~n49684 ;
  assign n49686 = \u1_desIn_r_reg[61]/NET0131  & ~n49685 ;
  assign n49687 = ~\u1_desIn_r_reg[61]/NET0131  & n49685 ;
  assign n49688 = ~n49686 & ~n49687 ;
  assign n49694 = ~n49663 & n49688 ;
  assign n49695 = ~n49682 & n49694 ;
  assign n49696 = ~n49693 & n49695 ;
  assign n49664 = ~n49642 & ~n49661 ;
  assign n49665 = ~n49655 & n49664 ;
  assign n49666 = ~n49648 & n49665 ;
  assign n49673 = n49666 & n49672 ;
  assign n49674 = n49642 & ~n49672 ;
  assign n49675 = n49662 & n49674 ;
  assign n49676 = n49655 & n49661 ;
  assign n49677 = n49642 & n49676 ;
  assign n49678 = n49672 & n49677 ;
  assign n49679 = ~n49675 & ~n49678 ;
  assign n49697 = ~n49673 & n49679 ;
  assign n49698 = n49696 & n49697 ;
  assign n49709 = ~n49672 & n49690 ;
  assign n49710 = n49661 & n49709 ;
  assign n49714 = n49676 & n49681 ;
  assign n49715 = ~n49688 & ~n49714 ;
  assign n49716 = ~n49710 & n49715 ;
  assign n49711 = n49648 & n49665 ;
  assign n49712 = n49672 & n49681 ;
  assign n49713 = ~n49655 & n49712 ;
  assign n49717 = ~n49711 & ~n49713 ;
  assign n49718 = n49716 & n49717 ;
  assign n49699 = ~n49661 & n49689 ;
  assign n49700 = n49672 & n49699 ;
  assign n49701 = ~n49655 & ~n49672 ;
  assign n49702 = ~n49661 & n49701 ;
  assign n49703 = ~n49642 & n49702 ;
  assign n49704 = ~n49700 & ~n49703 ;
  assign n49705 = n49672 & n49680 ;
  assign n49706 = ~n49642 & n49661 ;
  assign n49707 = ~n49705 & ~n49706 ;
  assign n49708 = ~n49648 & ~n49707 ;
  assign n49719 = n49704 & ~n49708 ;
  assign n49720 = n49718 & n49719 ;
  assign n49721 = ~n49698 & ~n49720 ;
  assign n49722 = ~n49702 & ~n49705 ;
  assign n49723 = n49649 & ~n49722 ;
  assign n49724 = n49661 & ~n49672 ;
  assign n49725 = ~n49648 & n49724 ;
  assign n49726 = n49689 & n49725 ;
  assign n49727 = ~n49672 & n49680 ;
  assign n49728 = n49681 & n49727 ;
  assign n49729 = ~n49726 & ~n49728 ;
  assign n49730 = ~n49723 & n49729 ;
  assign n49731 = ~n49721 & n49730 ;
  assign n49732 = ~\u1_desIn_r_reg[26]/NET0131  & ~n49731 ;
  assign n49733 = \u1_desIn_r_reg[26]/NET0131  & n49731 ;
  assign n49734 = ~n49732 & ~n49733 ;
  assign n49735 = n49405 & n49441 ;
  assign n49736 = ~n49424 & ~n49735 ;
  assign n49737 = n49399 & ~n49736 ;
  assign n49758 = ~n49405 & n49437 ;
  assign n49759 = ~n49737 & ~n49758 ;
  assign n49760 = ~n49421 & ~n49759 ;
  assign n49754 = n49412 & ~n49615 ;
  assign n49753 = n49415 & ~n49430 ;
  assign n49755 = ~n49469 & ~n49753 ;
  assign n49756 = ~n49754 & n49755 ;
  assign n49757 = n49421 & ~n49756 ;
  assign n49761 = n49414 & n49474 ;
  assign n49762 = ~n49757 & ~n49761 ;
  assign n49763 = ~n49760 & n49762 ;
  assign n49764 = ~n49453 & ~n49763 ;
  assign n49738 = ~n49458 & ~n49737 ;
  assign n49739 = n49421 & ~n49738 ;
  assign n49742 = ~n49431 & ~n49437 ;
  assign n49741 = ~n49405 & ~n49468 ;
  assign n49743 = ~n49421 & ~n49741 ;
  assign n49744 = ~n49742 & n49743 ;
  assign n49740 = n49414 & n49468 ;
  assign n49745 = ~n49476 & ~n49740 ;
  assign n49746 = n49443 & n49745 ;
  assign n49747 = ~n49744 & n49746 ;
  assign n49748 = ~n49739 & n49747 ;
  assign n49749 = n49453 & ~n49748 ;
  assign n49750 = n49412 & n49469 ;
  assign n49751 = ~n49405 & n49421 ;
  assign n49752 = n49457 & n49751 ;
  assign n49765 = ~n49750 & ~n49752 ;
  assign n49766 = ~n49749 & n49765 ;
  assign n49767 = ~n49764 & n49766 ;
  assign n49768 = \u1_desIn_r_reg[32]/NET0131  & ~n49767 ;
  assign n49769 = ~\u1_desIn_r_reg[32]/NET0131  & n49767 ;
  assign n49770 = ~n49768 & ~n49769 ;
  assign n49771 = decrypt_pad & ~\u1_key_r_reg[39]/P0001  ;
  assign n49772 = ~decrypt_pad & ~\u1_key_r_reg[32]/NET0131  ;
  assign n49773 = ~n49771 & ~n49772 ;
  assign n49774 = \u1_desIn_r_reg[63]/NET0131  & ~n49773 ;
  assign n49775 = ~\u1_desIn_r_reg[63]/NET0131  & n49773 ;
  assign n49776 = ~n49774 & ~n49775 ;
  assign n49777 = decrypt_pad & ~\u1_key_r_reg[48]/NET0131  ;
  assign n49778 = ~decrypt_pad & ~\u1_key_r_reg[41]/NET0131  ;
  assign n49779 = ~n49777 & ~n49778 ;
  assign n49780 = \u1_desIn_r_reg[55]/NET0131  & ~n49779 ;
  assign n49781 = ~\u1_desIn_r_reg[55]/NET0131  & n49779 ;
  assign n49782 = ~n49780 & ~n49781 ;
  assign n49796 = decrypt_pad & ~\u1_key_r_reg[6]/NET0131  ;
  assign n49797 = ~decrypt_pad & ~\u1_key_r_reg[24]/NET0131  ;
  assign n49798 = ~n49796 & ~n49797 ;
  assign n49799 = \u1_desIn_r_reg[39]/NET0131  & ~n49798 ;
  assign n49800 = ~\u1_desIn_r_reg[39]/NET0131  & n49798 ;
  assign n49801 = ~n49799 & ~n49800 ;
  assign n49783 = decrypt_pad & ~\u1_key_r_reg[27]/NET0131  ;
  assign n49784 = ~decrypt_pad & ~\u1_key_r_reg[20]/NET0131  ;
  assign n49785 = ~n49783 & ~n49784 ;
  assign n49786 = \u1_desIn_r_reg[31]/NET0131  & ~n49785 ;
  assign n49787 = ~\u1_desIn_r_reg[31]/NET0131  & n49785 ;
  assign n49788 = ~n49786 & ~n49787 ;
  assign n49789 = decrypt_pad & ~\u1_key_r_reg[19]/NET0131  ;
  assign n49790 = ~decrypt_pad & ~\u1_key_r_reg[12]/NET0131  ;
  assign n49791 = ~n49789 & ~n49790 ;
  assign n49792 = \u1_desIn_r_reg[5]/NET0131  & ~n49791 ;
  assign n49793 = ~\u1_desIn_r_reg[5]/NET0131  & n49791 ;
  assign n49794 = ~n49792 & ~n49793 ;
  assign n49811 = ~n49788 & n49794 ;
  assign n49812 = ~n49801 & n49811 ;
  assign n49803 = decrypt_pad & ~\u1_key_r_reg[54]/NET0131  ;
  assign n49804 = ~decrypt_pad & ~\u1_key_r_reg[47]/NET0131  ;
  assign n49805 = ~n49803 & ~n49804 ;
  assign n49806 = \u1_desIn_r_reg[47]/NET0131  & ~n49805 ;
  assign n49807 = ~\u1_desIn_r_reg[47]/NET0131  & n49805 ;
  assign n49808 = ~n49806 & ~n49807 ;
  assign n49813 = n49788 & n49801 ;
  assign n49814 = n49788 & ~n49794 ;
  assign n49815 = ~n49813 & ~n49814 ;
  assign n49816 = n49808 & ~n49815 ;
  assign n49817 = ~n49812 & ~n49816 ;
  assign n49818 = ~n49782 & ~n49817 ;
  assign n49819 = ~n49794 & n49801 ;
  assign n49820 = ~n49812 & ~n49819 ;
  assign n49821 = ~n49808 & ~n49820 ;
  assign n49795 = n49788 & n49794 ;
  assign n49802 = n49795 & ~n49801 ;
  assign n49809 = n49802 & n49808 ;
  assign n49810 = n49782 & n49809 ;
  assign n49822 = ~n49782 & ~n49801 ;
  assign n49823 = n49794 & ~n49808 ;
  assign n49824 = n49822 & n49823 ;
  assign n49825 = n49801 & n49808 ;
  assign n49826 = n49811 & n49825 ;
  assign n49827 = ~n49824 & ~n49826 ;
  assign n49828 = ~n49810 & n49827 ;
  assign n49829 = ~n49821 & n49828 ;
  assign n49830 = ~n49818 & n49829 ;
  assign n49831 = ~n49776 & ~n49830 ;
  assign n49848 = ~n49788 & ~n49794 ;
  assign n49849 = ~n49809 & ~n49848 ;
  assign n49850 = n49776 & ~n49849 ;
  assign n49832 = ~n49801 & n49808 ;
  assign n49851 = n49811 & ~n49832 ;
  assign n49852 = ~n49850 & ~n49851 ;
  assign n49847 = n49801 & ~n49808 ;
  assign n49853 = ~n49782 & ~n49847 ;
  assign n49854 = ~n49852 & n49853 ;
  assign n49833 = ~n49794 & n49832 ;
  assign n49834 = ~n49788 & n49833 ;
  assign n49835 = ~n49808 & n49813 ;
  assign n49836 = ~n49834 & ~n49835 ;
  assign n49837 = n49782 & ~n49836 ;
  assign n49838 = ~n49801 & n49814 ;
  assign n49839 = n49795 & n49801 ;
  assign n49840 = ~n49838 & ~n49839 ;
  assign n49841 = ~n49808 & ~n49840 ;
  assign n49842 = ~n49788 & n49808 ;
  assign n49843 = n49782 & n49801 ;
  assign n49844 = ~n49842 & n49843 ;
  assign n49845 = ~n49841 & ~n49844 ;
  assign n49846 = n49776 & ~n49845 ;
  assign n49855 = ~n49837 & ~n49846 ;
  assign n49856 = ~n49854 & n49855 ;
  assign n49857 = ~n49831 & n49856 ;
  assign n49858 = \u1_desIn_r_reg[14]/NET0131  & n49857 ;
  assign n49859 = ~\u1_desIn_r_reg[14]/NET0131  & ~n49857 ;
  assign n49860 = ~n49858 & ~n49859 ;
  assign n49863 = n49421 & ~n49437 ;
  assign n49864 = ~n49432 & n49863 ;
  assign n49865 = ~n49609 & n49864 ;
  assign n49861 = ~n49421 & n49754 ;
  assign n49862 = n49453 & n49457 ;
  assign n49866 = ~n49861 & ~n49862 ;
  assign n49867 = ~n49865 & n49866 ;
  assign n49868 = n49405 & ~n49867 ;
  assign n49870 = ~n49424 & ~n49444 ;
  assign n49871 = n49421 & ~n49467 ;
  assign n49872 = ~n49870 & ~n49871 ;
  assign n49869 = n49437 & n49751 ;
  assign n49873 = n49453 & ~n49869 ;
  assign n49874 = ~n49872 & n49873 ;
  assign n49875 = ~n49405 & ~n49742 ;
  assign n49876 = ~n49421 & ~n49609 ;
  assign n49877 = ~n49761 & n49876 ;
  assign n49878 = ~n49875 & n49877 ;
  assign n49879 = ~n49414 & ~n49455 ;
  assign n49880 = n49742 & n49879 ;
  assign n49881 = n49421 & ~n49439 ;
  assign n49882 = ~n49880 & n49881 ;
  assign n49883 = ~n49878 & ~n49882 ;
  assign n49884 = ~n49453 & ~n49750 ;
  assign n49885 = ~n49883 & n49884 ;
  assign n49886 = ~n49874 & ~n49885 ;
  assign n49887 = ~n49868 & ~n49886 ;
  assign n49888 = ~\u1_desIn_r_reg[30]/NET0131  & ~n49887 ;
  assign n49889 = \u1_desIn_r_reg[30]/NET0131  & n49887 ;
  assign n49890 = ~n49888 & ~n49889 ;
  assign n49901 = ~n49518 & ~n49519 ;
  assign n49902 = ~n49537 & ~n49901 ;
  assign n49891 = n49498 & n49514 ;
  assign n49892 = ~n49492 & n49891 ;
  assign n49893 = ~n49515 & ~n49539 ;
  assign n49894 = n49512 & ~n49893 ;
  assign n49905 = ~n49892 & ~n49894 ;
  assign n49906 = ~n49902 & n49905 ;
  assign n49896 = n49505 & ~n49511 ;
  assign n49897 = ~n49492 & n49896 ;
  assign n49898 = n49511 & n49550 ;
  assign n49899 = ~n49897 & ~n49898 ;
  assign n49900 = ~n49498 & ~n49899 ;
  assign n49895 = ~n49537 & n49550 ;
  assign n49903 = ~n49527 & ~n49895 ;
  assign n49904 = ~n49547 & n49903 ;
  assign n49907 = ~n49900 & n49904 ;
  assign n49908 = n49906 & n49907 ;
  assign n49909 = n49498 & n49505 ;
  assign n49910 = ~n49566 & ~n49909 ;
  assign n49911 = n49537 & ~n49910 ;
  assign n49917 = ~n49516 & n49527 ;
  assign n49918 = ~n49562 & n49917 ;
  assign n49912 = ~n49505 & n49520 ;
  assign n49913 = ~n49514 & ~n49560 ;
  assign n49914 = ~n49505 & n49537 ;
  assign n49915 = n49499 & ~n49914 ;
  assign n49916 = n49913 & n49915 ;
  assign n49919 = ~n49912 & ~n49916 ;
  assign n49920 = n49918 & n49919 ;
  assign n49921 = ~n49911 & n49920 ;
  assign n49922 = ~n49908 & ~n49921 ;
  assign n49923 = \u1_desIn_r_reg[28]/NET0131  & n49922 ;
  assign n49924 = ~\u1_desIn_r_reg[28]/NET0131  & ~n49922 ;
  assign n49925 = ~n49923 & ~n49924 ;
  assign n49930 = ~n49782 & ~n49802 ;
  assign n49931 = ~n49833 & n49930 ;
  assign n49934 = n49794 & n49842 ;
  assign n49932 = ~n49801 & ~n49808 ;
  assign n49933 = ~n49794 & n49932 ;
  assign n49935 = n49782 & ~n49933 ;
  assign n49936 = ~n49934 & n49935 ;
  assign n49937 = ~n49931 & ~n49936 ;
  assign n49928 = n49801 & n49848 ;
  assign n49929 = ~n49808 & n49928 ;
  assign n49938 = n49776 & n49827 ;
  assign n49939 = ~n49929 & n49938 ;
  assign n49940 = ~n49937 & n49939 ;
  assign n49944 = ~n49788 & ~n49822 ;
  assign n49945 = n49823 & n49944 ;
  assign n49941 = n49782 & n49788 ;
  assign n49942 = n49808 & ~n49819 ;
  assign n49943 = n49941 & n49942 ;
  assign n49946 = ~n49776 & ~n49943 ;
  assign n49947 = ~n49945 & n49946 ;
  assign n49950 = ~n49782 & ~n49928 ;
  assign n49948 = n49811 & n49832 ;
  assign n49949 = n49814 & n49932 ;
  assign n49951 = ~n49948 & ~n49949 ;
  assign n49952 = n49950 & n49951 ;
  assign n49953 = n49947 & n49952 ;
  assign n49954 = ~n49940 & ~n49953 ;
  assign n49926 = n49814 & n49825 ;
  assign n49927 = n49794 & n49835 ;
  assign n49955 = ~n49926 & ~n49927 ;
  assign n49956 = ~n49954 & n49955 ;
  assign n49959 = ~n49795 & ~n49848 ;
  assign n49960 = ~n49801 & ~n49959 ;
  assign n49957 = ~n49808 & n49814 ;
  assign n49958 = n49801 & n49957 ;
  assign n49961 = n49782 & ~n49958 ;
  assign n49962 = ~n49960 & n49961 ;
  assign n49963 = n49947 & n49962 ;
  assign n49964 = ~n49956 & ~n49963 ;
  assign n49965 = ~\u1_desIn_r_reg[36]/NET0131  & ~n49964 ;
  assign n49966 = \u1_desIn_r_reg[36]/NET0131  & n49964 ;
  assign n49967 = ~n49965 & ~n49966 ;
  assign n50001 = decrypt_pad & ~\u1_key_r_reg[44]/NET0131  ;
  assign n50002 = ~decrypt_pad & ~\u1_key_r_reg[37]/NET0131  ;
  assign n50003 = ~n50001 & ~n50002 ;
  assign n50004 = \u1_desIn_r_reg[41]/NET0131  & ~n50003 ;
  assign n50005 = ~\u1_desIn_r_reg[41]/NET0131  & n50003 ;
  assign n50006 = ~n50004 & ~n50005 ;
  assign n49980 = decrypt_pad & ~\u1_key_r_reg[16]/NET0131  ;
  assign n49981 = ~decrypt_pad & ~\u1_key_r_reg[9]/NET0131  ;
  assign n49982 = ~n49980 & ~n49981 ;
  assign n49983 = \u1_desIn_r_reg[25]/NET0131  & ~n49982 ;
  assign n49984 = ~\u1_desIn_r_reg[25]/NET0131  & n49982 ;
  assign n49985 = ~n49983 & ~n49984 ;
  assign n49986 = decrypt_pad & ~\u1_key_r_reg[43]/NET0131  ;
  assign n49987 = ~decrypt_pad & ~\u1_key_r_reg[36]/NET0131  ;
  assign n49988 = ~n49986 & ~n49987 ;
  assign n49989 = \u1_desIn_r_reg[33]/NET0131  & ~n49988 ;
  assign n49990 = ~\u1_desIn_r_reg[33]/NET0131  & n49988 ;
  assign n49991 = ~n49989 & ~n49990 ;
  assign n49993 = decrypt_pad & ~\u1_key_r_reg[28]/NET0131  ;
  assign n49994 = ~decrypt_pad & ~\u1_key_r_reg[21]/NET0131  ;
  assign n49995 = ~n49993 & ~n49994 ;
  assign n49996 = \u1_desIn_r_reg[7]/NET0131  & ~n49995 ;
  assign n49997 = ~\u1_desIn_r_reg[7]/NET0131  & n49995 ;
  assign n49998 = ~n49996 & ~n49997 ;
  assign n50017 = ~n49991 & ~n49998 ;
  assign n50018 = ~n49985 & n50017 ;
  assign n50038 = ~n50006 & n50018 ;
  assign n50039 = n49991 & ~n49998 ;
  assign n50040 = ~n49985 & n50039 ;
  assign n50041 = n50006 & n50040 ;
  assign n50042 = ~n50038 & ~n50041 ;
  assign n49974 = decrypt_pad & ~\u1_key_r_reg[1]/NET0131  ;
  assign n49975 = ~decrypt_pad & ~\u1_key_r_reg[49]/NET0131  ;
  assign n49976 = ~n49974 & ~n49975 ;
  assign n49977 = \u1_desIn_r_reg[49]/NET0131  & ~n49976 ;
  assign n49978 = ~\u1_desIn_r_reg[49]/NET0131  & n49976 ;
  assign n49979 = ~n49977 & ~n49978 ;
  assign n50020 = ~n49985 & n50006 ;
  assign n50024 = ~n49991 & n50006 ;
  assign n49999 = ~n49985 & n49998 ;
  assign n50035 = n49991 & n49999 ;
  assign n50036 = ~n50024 & ~n50035 ;
  assign n50037 = ~n50020 & ~n50036 ;
  assign n50043 = ~n49979 & ~n50037 ;
  assign n50044 = n50042 & n50043 ;
  assign n50047 = ~n49991 & ~n50006 ;
  assign n50048 = n49998 & n50047 ;
  assign n50049 = ~n49985 & n50048 ;
  assign n50045 = n49991 & n50020 ;
  assign n50046 = n49998 & n50045 ;
  assign n50050 = n49979 & ~n50046 ;
  assign n50051 = ~n50049 & n50050 ;
  assign n50052 = ~n50044 & ~n50051 ;
  assign n49968 = decrypt_pad & ~\u1_key_r_reg[7]/NET0131  ;
  assign n49969 = ~decrypt_pad & ~\u1_key_r_reg[0]/NET0131  ;
  assign n49970 = ~n49968 & ~n49969 ;
  assign n49971 = \u1_desIn_r_reg[57]/NET0131  & ~n49970 ;
  assign n49972 = ~\u1_desIn_r_reg[57]/NET0131  & n49970 ;
  assign n49973 = ~n49971 & ~n49972 ;
  assign n50007 = n49991 & ~n50006 ;
  assign n50008 = ~n49998 & n50007 ;
  assign n49992 = n49985 & n49991 ;
  assign n50000 = ~n49991 & n49999 ;
  assign n50009 = ~n49992 & ~n50000 ;
  assign n50010 = ~n50008 & n50009 ;
  assign n50011 = n49979 & ~n50010 ;
  assign n50012 = n49985 & ~n50006 ;
  assign n50013 = ~n49998 & n50012 ;
  assign n50014 = ~n49991 & n50013 ;
  assign n50015 = ~n50011 & ~n50014 ;
  assign n50016 = ~n49973 & ~n50015 ;
  assign n50021 = ~n50012 & ~n50020 ;
  assign n50022 = ~n49999 & ~n50021 ;
  assign n50023 = n49991 & n50022 ;
  assign n50019 = n49979 & n50018 ;
  assign n50025 = ~n49979 & n49998 ;
  assign n50026 = n49985 & n49998 ;
  assign n50027 = ~n50025 & ~n50026 ;
  assign n50028 = n50024 & ~n50027 ;
  assign n50029 = ~n50019 & ~n50028 ;
  assign n50030 = ~n50023 & n50029 ;
  assign n50031 = n49973 & ~n50030 ;
  assign n50032 = ~n49979 & ~n49991 ;
  assign n50033 = ~n49973 & n49985 ;
  assign n50034 = n50032 & n50033 ;
  assign n50053 = ~n50031 & ~n50034 ;
  assign n50054 = ~n50016 & n50053 ;
  assign n50055 = ~n50052 & n50054 ;
  assign n50056 = \u1_desIn_r_reg[52]/P0001  & n50055 ;
  assign n50057 = ~\u1_desIn_r_reg[52]/P0001  & ~n50055 ;
  assign n50058 = ~n50056 & ~n50057 ;
  assign n50059 = decrypt_pad & ~\u1_key_r_reg[23]/NET0131  ;
  assign n50060 = ~decrypt_pad & ~\u1_key_r_reg[16]/NET0131  ;
  assign n50061 = ~n50059 & ~n50060 ;
  assign n50062 = \u1_desIn_r_reg[27]/NET0131  & ~n50061 ;
  assign n50063 = ~\u1_desIn_r_reg[27]/NET0131  & n50061 ;
  assign n50064 = ~n50062 & ~n50063 ;
  assign n50092 = decrypt_pad & ~\u1_key_r_reg[8]/NET0131  ;
  assign n50093 = ~decrypt_pad & ~\u1_key_r_reg[1]/NET0131  ;
  assign n50094 = ~n50092 & ~n50093 ;
  assign n50095 = \u1_desIn_r_reg[19]/NET0131  & ~n50094 ;
  assign n50096 = ~\u1_desIn_r_reg[19]/NET0131  & n50094 ;
  assign n50097 = ~n50095 & ~n50096 ;
  assign n50065 = decrypt_pad & ~\u1_key_r_reg[31]/NET0131  ;
  assign n50066 = ~decrypt_pad & ~\u1_key_r_reg[51]/NET0131  ;
  assign n50067 = ~n50065 & ~n50066 ;
  assign n50068 = \u1_desIn_r_reg[3]/NET0131  & ~n50067 ;
  assign n50069 = ~\u1_desIn_r_reg[3]/NET0131  & n50067 ;
  assign n50070 = ~n50068 & ~n50069 ;
  assign n50078 = decrypt_pad & ~\u1_key_r_reg[36]/NET0131  ;
  assign n50079 = ~decrypt_pad & ~\u1_key_r_reg[29]/NET0131  ;
  assign n50080 = ~n50078 & ~n50079 ;
  assign n50081 = \u1_desIn_r_reg[61]/NET0131  & ~n50080 ;
  assign n50082 = ~\u1_desIn_r_reg[61]/NET0131  & n50080 ;
  assign n50083 = ~n50081 & ~n50082 ;
  assign n50085 = decrypt_pad & ~\u1_key_r_reg[52]/NET0131  ;
  assign n50086 = ~decrypt_pad & ~\u1_key_r_reg[45]/NET0131  ;
  assign n50087 = ~n50085 & ~n50086 ;
  assign n50088 = \u1_desIn_r_reg[35]/NET0131  & ~n50087 ;
  assign n50089 = ~\u1_desIn_r_reg[35]/NET0131  & n50087 ;
  assign n50090 = ~n50088 & ~n50089 ;
  assign n50101 = ~n50083 & n50090 ;
  assign n50102 = ~n50070 & n50101 ;
  assign n50103 = n50070 & ~n50090 ;
  assign n50125 = n50083 & n50103 ;
  assign n50138 = ~n50102 & ~n50125 ;
  assign n50071 = decrypt_pad & ~\u1_key_r_reg[21]/NET0131  ;
  assign n50072 = ~decrypt_pad & ~\u1_key_r_reg[14]/NET0131  ;
  assign n50073 = ~n50071 & ~n50072 ;
  assign n50074 = \u1_desIn_r_reg[11]/NET0131  & ~n50073 ;
  assign n50075 = ~\u1_desIn_r_reg[11]/NET0131  & n50073 ;
  assign n50076 = ~n50074 & ~n50075 ;
  assign n50105 = n50083 & n50090 ;
  assign n50136 = ~n50076 & n50105 ;
  assign n50137 = n50076 & n50101 ;
  assign n50139 = ~n50136 & ~n50137 ;
  assign n50140 = n50138 & n50139 ;
  assign n50141 = n50097 & ~n50140 ;
  assign n50127 = ~n50076 & ~n50097 ;
  assign n50112 = ~n50083 & ~n50090 ;
  assign n50113 = ~n50070 & n50112 ;
  assign n50128 = n50070 & n50101 ;
  assign n50129 = ~n50113 & ~n50128 ;
  assign n50130 = n50127 & ~n50129 ;
  assign n50131 = n50070 & ~n50097 ;
  assign n50132 = n50076 & ~n50131 ;
  assign n50077 = n50070 & ~n50076 ;
  assign n50133 = ~n50077 & n50105 ;
  assign n50134 = ~n50132 & n50133 ;
  assign n50126 = ~n50076 & n50125 ;
  assign n50098 = n50083 & ~n50090 ;
  assign n50119 = ~n50070 & n50076 ;
  assign n50135 = n50098 & n50119 ;
  assign n50142 = ~n50126 & ~n50135 ;
  assign n50143 = ~n50134 & n50142 ;
  assign n50144 = ~n50130 & n50143 ;
  assign n50145 = ~n50141 & n50144 ;
  assign n50146 = n50064 & ~n50145 ;
  assign n50106 = n50070 & n50105 ;
  assign n50107 = ~n50076 & n50106 ;
  assign n50104 = n50076 & n50103 ;
  assign n50099 = ~n50070 & ~n50076 ;
  assign n50100 = n50098 & n50099 ;
  assign n50108 = ~n50100 & ~n50102 ;
  assign n50109 = ~n50104 & n50108 ;
  assign n50110 = ~n50107 & n50109 ;
  assign n50111 = ~n50097 & ~n50110 ;
  assign n50114 = n50076 & n50090 ;
  assign n50115 = n50083 & n50114 ;
  assign n50084 = n50077 & ~n50083 ;
  assign n50116 = ~n50084 & ~n50113 ;
  assign n50117 = ~n50115 & n50116 ;
  assign n50118 = n50097 & ~n50117 ;
  assign n50091 = n50084 & ~n50090 ;
  assign n50120 = n50105 & n50119 ;
  assign n50121 = ~n50091 & ~n50120 ;
  assign n50122 = ~n50118 & n50121 ;
  assign n50123 = ~n50111 & n50122 ;
  assign n50124 = ~n50064 & ~n50123 ;
  assign n50147 = n50076 & n50113 ;
  assign n50148 = ~n50126 & ~n50147 ;
  assign n50149 = n50097 & ~n50148 ;
  assign n50150 = n50076 & n50102 ;
  assign n50151 = n50076 & ~n50083 ;
  assign n50152 = n50103 & n50151 ;
  assign n50153 = ~n50150 & ~n50152 ;
  assign n50154 = ~n50097 & ~n50153 ;
  assign n50155 = ~n50149 & ~n50154 ;
  assign n50156 = ~n50124 & n50155 ;
  assign n50157 = ~n50146 & n50156 ;
  assign n50158 = ~\u1_desIn_r_reg[44]/NET0131  & ~n50157 ;
  assign n50159 = \u1_desIn_r_reg[44]/NET0131  & n50157 ;
  assign n50160 = ~n50158 & ~n50159 ;
  assign n50161 = ~n49642 & n49672 ;
  assign n50179 = n49680 & n50161 ;
  assign n50180 = n49648 & ~n49702 ;
  assign n50181 = ~n50179 & n50180 ;
  assign n50182 = n49655 & n49706 ;
  assign n50183 = ~n49648 & ~n49727 ;
  assign n50184 = ~n50182 & n50183 ;
  assign n50185 = ~n50181 & ~n50184 ;
  assign n50186 = n49642 & n49727 ;
  assign n50187 = n49679 & ~n50186 ;
  assign n50188 = ~n50185 & n50187 ;
  assign n50189 = ~n49688 & ~n50188 ;
  assign n50171 = n49674 & ~n49680 ;
  assign n50172 = n49642 & n49662 ;
  assign n50173 = ~n50171 & ~n50172 ;
  assign n50174 = ~n49648 & ~n50173 ;
  assign n50169 = n49642 & n49705 ;
  assign n50175 = ~n49655 & n50161 ;
  assign n50176 = ~n50169 & ~n50175 ;
  assign n50177 = ~n50174 & n50176 ;
  assign n50178 = n49688 & ~n50177 ;
  assign n50162 = n49662 & n50161 ;
  assign n50163 = ~n49678 & ~n50162 ;
  assign n50164 = ~n49700 & n50163 ;
  assign n50165 = n49648 & ~n50164 ;
  assign n50170 = ~n49648 & n50169 ;
  assign n50166 = ~n49706 & ~n49709 ;
  assign n50167 = n49648 & n49688 ;
  assign n50168 = ~n50166 & n50167 ;
  assign n50190 = ~n49673 & ~n50168 ;
  assign n50191 = ~n50170 & n50190 ;
  assign n50192 = ~n50165 & n50191 ;
  assign n50193 = ~n50178 & n50192 ;
  assign n50194 = ~n50189 & n50193 ;
  assign n50195 = ~\u1_desIn_r_reg[6]/NET0131  & ~n50194 ;
  assign n50196 = \u1_desIn_r_reg[6]/NET0131  & n50194 ;
  assign n50197 = ~n50195 & ~n50196 ;
  assign n50218 = n49998 & ~n50021 ;
  assign n50219 = ~n50040 & ~n50218 ;
  assign n50220 = ~n49979 & ~n50219 ;
  assign n50213 = n49991 & n49998 ;
  assign n50214 = n50012 & n50213 ;
  assign n50223 = ~n50045 & ~n50214 ;
  assign n50224 = ~n50038 & n50223 ;
  assign n50215 = n49985 & ~n50213 ;
  assign n50216 = n49979 & ~n50047 ;
  assign n50217 = n50215 & n50216 ;
  assign n50221 = ~n49998 & n50024 ;
  assign n50222 = n49985 & n50221 ;
  assign n50225 = ~n50217 & ~n50222 ;
  assign n50226 = n50224 & n50225 ;
  assign n50227 = ~n50220 & n50226 ;
  assign n50228 = ~n49973 & ~n50227 ;
  assign n50199 = n49979 & ~n50035 ;
  assign n50198 = n49992 & n50006 ;
  assign n50200 = ~n50048 & ~n50198 ;
  assign n50201 = n50199 & n50200 ;
  assign n50202 = n50006 & n50026 ;
  assign n50203 = ~n49991 & n50202 ;
  assign n50204 = ~n49979 & ~n50013 ;
  assign n50205 = ~n50203 & n50204 ;
  assign n50206 = ~n50201 & ~n50205 ;
  assign n50207 = n49992 & ~n49998 ;
  assign n50208 = ~n50018 & ~n50207 ;
  assign n50209 = n50006 & ~n50208 ;
  assign n50210 = ~n50049 & ~n50209 ;
  assign n50211 = ~n50206 & n50210 ;
  assign n50212 = n49973 & ~n50211 ;
  assign n50229 = ~n49985 & n50047 ;
  assign n50230 = n49979 & n50229 ;
  assign n50231 = ~n49979 & n50214 ;
  assign n50232 = ~n50230 & ~n50231 ;
  assign n50233 = ~n50212 & n50232 ;
  assign n50234 = ~n50228 & n50233 ;
  assign n50235 = ~\u1_desIn_r_reg[34]/NET0131  & ~n50234 ;
  assign n50236 = \u1_desIn_r_reg[34]/NET0131  & n50234 ;
  assign n50237 = ~n50235 & ~n50236 ;
  assign n50259 = ~n49331 & ~n49577 ;
  assign n50260 = ~n49325 & n49352 ;
  assign n50261 = ~n50259 & ~n50260 ;
  assign n50262 = n49306 & ~n50261 ;
  assign n50258 = n49349 & n49350 ;
  assign n50263 = ~n49595 & ~n50258 ;
  assign n50264 = ~n50262 & n50263 ;
  assign n50265 = ~n49318 & ~n50264 ;
  assign n50238 = ~n49346 & ~n49351 ;
  assign n50239 = n49318 & ~n50238 ;
  assign n50240 = ~n49383 & ~n50239 ;
  assign n50241 = ~n49319 & ~n50240 ;
  assign n50242 = n49318 & ~n49377 ;
  assign n50243 = n49341 & n50242 ;
  assign n50244 = n49360 & n49376 ;
  assign n50245 = n49306 & ~n49592 ;
  assign n50246 = ~n50244 & n50245 ;
  assign n50247 = ~n50243 & n50246 ;
  assign n50253 = ~n49306 & ~n49369 ;
  assign n50254 = ~n49382 & n50253 ;
  assign n50248 = ~n49345 & ~n49381 ;
  assign n50249 = n49601 & ~n50248 ;
  assign n50250 = ~n49340 & ~n49381 ;
  assign n50251 = ~n49318 & n49331 ;
  assign n50252 = ~n50250 & n50251 ;
  assign n50255 = ~n50249 & ~n50252 ;
  assign n50256 = n50254 & n50255 ;
  assign n50257 = ~n50247 & ~n50256 ;
  assign n50266 = ~n50241 & ~n50257 ;
  assign n50267 = ~n50265 & n50266 ;
  assign n50268 = \u1_desIn_r_reg[50]/NET0131  & ~n50267 ;
  assign n50269 = ~\u1_desIn_r_reg[50]/NET0131  & n50267 ;
  assign n50270 = ~n50268 & ~n50269 ;
  assign n50281 = ~n50070 & n50105 ;
  assign n50282 = ~n50097 & ~n50281 ;
  assign n50283 = ~n50084 & n50282 ;
  assign n50287 = n50097 & ~n50106 ;
  assign n50284 = ~n50099 & ~n50151 ;
  assign n50285 = ~n50090 & ~n50284 ;
  assign n50286 = ~n50070 & ~n50083 ;
  assign n50288 = ~n50285 & ~n50286 ;
  assign n50289 = n50287 & n50288 ;
  assign n50290 = ~n50283 & ~n50289 ;
  assign n50276 = n50083 & n50104 ;
  assign n50271 = n50077 & n50090 ;
  assign n50291 = n50064 & ~n50271 ;
  assign n50292 = ~n50276 & n50291 ;
  assign n50293 = ~n50290 & n50292 ;
  assign n50272 = ~n50070 & ~n50097 ;
  assign n50295 = ~n50083 & n50272 ;
  assign n50296 = n50097 & n50103 ;
  assign n50297 = ~n50295 & ~n50296 ;
  assign n50298 = ~n50076 & ~n50297 ;
  assign n50299 = ~n50090 & n50097 ;
  assign n50300 = n50070 & n50151 ;
  assign n50301 = ~n50299 & n50300 ;
  assign n50294 = n50098 & n50272 ;
  assign n50302 = ~n50064 & ~n50294 ;
  assign n50303 = ~n50301 & n50302 ;
  assign n50304 = ~n50298 & n50303 ;
  assign n50305 = ~n50293 & ~n50304 ;
  assign n50273 = n50076 & n50272 ;
  assign n50274 = ~n50271 & ~n50273 ;
  assign n50275 = n50083 & ~n50274 ;
  assign n50277 = ~n50147 & ~n50276 ;
  assign n50278 = n50099 & n50101 ;
  assign n50279 = n50277 & ~n50278 ;
  assign n50280 = n50097 & ~n50279 ;
  assign n50306 = ~n50275 & ~n50280 ;
  assign n50307 = ~n50305 & n50306 ;
  assign n50308 = ~\u1_desIn_r_reg[0]/NET0131  & ~n50307 ;
  assign n50309 = \u1_desIn_r_reg[0]/NET0131  & n50307 ;
  assign n50310 = ~n50308 & ~n50309 ;
  assign n50329 = n49808 & n49928 ;
  assign n50330 = n49840 & ~n50329 ;
  assign n50331 = n49782 & ~n50330 ;
  assign n50314 = ~n49808 & n49848 ;
  assign n50315 = n49801 & n49811 ;
  assign n50316 = ~n50314 & ~n50315 ;
  assign n50328 = ~n49782 & ~n50316 ;
  assign n50326 = ~n49802 & ~n49941 ;
  assign n50327 = ~n49808 & ~n50326 ;
  assign n50332 = ~n49948 & ~n50327 ;
  assign n50333 = ~n50328 & n50332 ;
  assign n50334 = ~n50331 & n50333 ;
  assign n50335 = n49776 & ~n50334 ;
  assign n50311 = ~n49801 & n49842 ;
  assign n50312 = ~n49926 & ~n50311 ;
  assign n50313 = ~n49782 & ~n50312 ;
  assign n50317 = n49782 & n50316 ;
  assign n50318 = ~n49782 & ~n49813 ;
  assign n50319 = ~n49812 & n50318 ;
  assign n50320 = ~n49957 & n50319 ;
  assign n50321 = ~n50317 & ~n50320 ;
  assign n50322 = n49832 & ~n49959 ;
  assign n50323 = ~n49926 & ~n50322 ;
  assign n50324 = ~n50321 & n50323 ;
  assign n50325 = ~n49776 & ~n50324 ;
  assign n50336 = ~n50313 & ~n50325 ;
  assign n50337 = ~n50335 & n50336 ;
  assign n50338 = ~\u1_desIn_r_reg[24]/NET0131  & ~n50337 ;
  assign n50339 = \u1_desIn_r_reg[24]/NET0131  & n50337 ;
  assign n50340 = ~n50338 & ~n50339 ;
  assign n50348 = n49648 & n49662 ;
  assign n50349 = ~n50172 & ~n50348 ;
  assign n50350 = n49672 & ~n50349 ;
  assign n50356 = ~n49711 & ~n50350 ;
  assign n50351 = n49642 & ~n49722 ;
  assign n50352 = n49672 & n49676 ;
  assign n50353 = n49701 & n49706 ;
  assign n50354 = ~n50352 & ~n50353 ;
  assign n50355 = ~n49648 & ~n50354 ;
  assign n50357 = ~n50351 & ~n50355 ;
  assign n50358 = n50356 & n50357 ;
  assign n50359 = n49688 & ~n50358 ;
  assign n50341 = ~n49664 & ~n50175 ;
  assign n50342 = ~n49688 & ~n50341 ;
  assign n50343 = ~n49661 & ~n49691 ;
  assign n50344 = ~n49677 & ~n50343 ;
  assign n50345 = ~n49672 & ~n50344 ;
  assign n50346 = ~n50342 & ~n50345 ;
  assign n50347 = ~n49648 & ~n50346 ;
  assign n50360 = ~n49662 & n49712 ;
  assign n50361 = ~n49675 & ~n49682 ;
  assign n50362 = ~n49709 & n50361 ;
  assign n50363 = ~n50360 & n50362 ;
  assign n50364 = ~n49688 & ~n50363 ;
  assign n50365 = n49648 & n49724 ;
  assign n50366 = ~n49691 & n50365 ;
  assign n50367 = ~n50364 & ~n50366 ;
  assign n50368 = ~n50347 & n50367 ;
  assign n50369 = ~n50359 & n50368 ;
  assign n50370 = ~\u1_desIn_r_reg[8]/NET0131  & ~n50369 ;
  assign n50371 = \u1_desIn_r_reg[8]/NET0131  & n50369 ;
  assign n50372 = ~n50370 & ~n50371 ;
  assign n50381 = ~n49979 & n50022 ;
  assign n50382 = ~n50013 & ~n50025 ;
  assign n50383 = ~n50202 & n50382 ;
  assign n50384 = n49991 & ~n50383 ;
  assign n50385 = ~n50381 & ~n50384 ;
  assign n50386 = ~n49973 & ~n50385 ;
  assign n50375 = ~n50000 & ~n50222 ;
  assign n50376 = ~n49973 & ~n50375 ;
  assign n50377 = ~n49991 & n50218 ;
  assign n50378 = n50042 & ~n50377 ;
  assign n50379 = ~n50376 & n50378 ;
  assign n50380 = n49979 & ~n50379 ;
  assign n50373 = n50012 & n50039 ;
  assign n50374 = ~n49979 & n50373 ;
  assign n50388 = ~n50012 & ~n50039 ;
  assign n50389 = n49979 & ~n50373 ;
  assign n50390 = ~n50388 & n50389 ;
  assign n50387 = n50021 & n50032 ;
  assign n50391 = ~n50046 & ~n50387 ;
  assign n50392 = ~n50390 & n50391 ;
  assign n50393 = n49973 & ~n50392 ;
  assign n50394 = ~n50374 & ~n50393 ;
  assign n50395 = ~n50380 & n50394 ;
  assign n50396 = ~n50386 & n50395 ;
  assign n50397 = \u1_desIn_r_reg[38]/NET0131  & ~n50396 ;
  assign n50398 = ~\u1_desIn_r_reg[38]/NET0131  & n50396 ;
  assign n50399 = ~n50397 & ~n50398 ;
  assign n50400 = ~n50097 & ~n50135 ;
  assign n50401 = n50097 & ~n50150 ;
  assign n50402 = ~n50076 & n50101 ;
  assign n50403 = n50070 & n50402 ;
  assign n50404 = ~n50104 & ~n50403 ;
  assign n50405 = n50401 & n50404 ;
  assign n50406 = ~n50400 & ~n50405 ;
  assign n50408 = ~n50076 & n50113 ;
  assign n50409 = ~n50281 & ~n50408 ;
  assign n50410 = n50097 & ~n50409 ;
  assign n50407 = n50083 & n50127 ;
  assign n50411 = n50064 & ~n50407 ;
  assign n50412 = n50153 & n50411 ;
  assign n50413 = ~n50410 & n50412 ;
  assign n50414 = n50101 & ~n50119 ;
  assign n50415 = n50282 & ~n50414 ;
  assign n50416 = ~n50100 & n50287 ;
  assign n50417 = ~n50415 & ~n50416 ;
  assign n50418 = ~n50064 & ~n50084 ;
  assign n50419 = n50277 & n50418 ;
  assign n50420 = ~n50417 & n50419 ;
  assign n50421 = ~n50413 & ~n50420 ;
  assign n50422 = ~n50406 & ~n50421 ;
  assign n50423 = ~\u1_desIn_r_reg[62]/NET0131  & ~n50422 ;
  assign n50424 = \u1_desIn_r_reg[62]/NET0131  & n50422 ;
  assign n50425 = ~n50423 & ~n50424 ;
  assign n50436 = ~n49672 & n50348 ;
  assign n50434 = n49649 & n49655 ;
  assign n50435 = ~n49724 & n50434 ;
  assign n50439 = ~n49666 & ~n50435 ;
  assign n50440 = ~n50436 & n50439 ;
  assign n50437 = ~n49674 & ~n49725 ;
  assign n50438 = n49655 & ~n50437 ;
  assign n50441 = n49704 & ~n50438 ;
  assign n50442 = n50440 & n50441 ;
  assign n50443 = ~n49688 & ~n50442 ;
  assign n50429 = ~n49699 & ~n49710 ;
  assign n50430 = n49648 & ~n50429 ;
  assign n50426 = ~n49674 & n49680 ;
  assign n50427 = ~n49675 & ~n50426 ;
  assign n50428 = ~n49648 & ~n50427 ;
  assign n50431 = n50163 & ~n50428 ;
  assign n50432 = ~n50430 & n50431 ;
  assign n50433 = n49688 & ~n50432 ;
  assign n50444 = ~n49703 & n50163 ;
  assign n50445 = ~n49648 & ~n50444 ;
  assign n50446 = ~n49713 & ~n49728 ;
  assign n50447 = ~n50445 & n50446 ;
  assign n50448 = ~n50433 & n50447 ;
  assign n50449 = ~n50443 & n50448 ;
  assign n50450 = ~\u1_desIn_r_reg[12]/NET0131  & ~n50449 ;
  assign n50451 = \u1_desIn_r_reg[12]/NET0131  & n50449 ;
  assign n50452 = ~n50450 & ~n50451 ;
  assign n50453 = ~n50035 & ~n50207 ;
  assign n50454 = ~n50229 & n50453 ;
  assign n50455 = ~n49979 & ~n50454 ;
  assign n50456 = ~n49985 & ~n50008 ;
  assign n50457 = n49979 & ~n50215 ;
  assign n50458 = ~n50456 & n50457 ;
  assign n50459 = ~n50046 & ~n50048 ;
  assign n50460 = ~n50222 & n50459 ;
  assign n50461 = ~n50458 & n50460 ;
  assign n50462 = ~n50455 & n50461 ;
  assign n50463 = n49973 & ~n50462 ;
  assign n50470 = ~n49973 & ~n50008 ;
  assign n50469 = n49998 & ~n50007 ;
  assign n50471 = ~n50045 & ~n50469 ;
  assign n50472 = n50470 & n50471 ;
  assign n50473 = ~n50221 & ~n50472 ;
  assign n50474 = n49979 & ~n50473 ;
  assign n50464 = ~n50040 & ~n50202 ;
  assign n50465 = ~n49979 & ~n50464 ;
  assign n50466 = n49999 & n50024 ;
  assign n50467 = ~n50465 & ~n50466 ;
  assign n50468 = ~n49973 & ~n50467 ;
  assign n50475 = ~n50017 & ~n50213 ;
  assign n50476 = n50381 & n50475 ;
  assign n50477 = ~n50468 & ~n50476 ;
  assign n50478 = ~n50474 & n50477 ;
  assign n50479 = ~n50463 & n50478 ;
  assign n50480 = ~\u1_desIn_r_reg[16]/NET0131  & ~n50479 ;
  assign n50481 = \u1_desIn_r_reg[16]/NET0131  & n50479 ;
  assign n50482 = ~n50480 & ~n50481 ;
  assign n50485 = ~n49492 & ~n49913 ;
  assign n50486 = ~n49498 & n49560 ;
  assign n50487 = ~n49561 & ~n50486 ;
  assign n50488 = ~n50485 & ~n50487 ;
  assign n50489 = ~n49891 & ~n50488 ;
  assign n50490 = ~n49537 & ~n50489 ;
  assign n50483 = n49492 & n49896 ;
  assign n50484 = n49498 & n50483 ;
  assign n50491 = ~n49520 & ~n49546 ;
  assign n50492 = ~n50483 & n50491 ;
  assign n50493 = n49537 & ~n50492 ;
  assign n50494 = ~n50484 & ~n50493 ;
  assign n50495 = ~n50490 & n50494 ;
  assign n50496 = n49527 & ~n50495 ;
  assign n50497 = n49498 & ~n49899 ;
  assign n50501 = n49517 & ~n50497 ;
  assign n50498 = ~n49897 & n49902 ;
  assign n50499 = ~n49897 & ~n50486 ;
  assign n50500 = n49537 & ~n50499 ;
  assign n50502 = ~n50498 & ~n50500 ;
  assign n50503 = n50501 & n50502 ;
  assign n50504 = ~n49527 & ~n50503 ;
  assign n50505 = n49513 & n49537 ;
  assign n50506 = n49557 & ~n49896 ;
  assign n50507 = n49551 & n50506 ;
  assign n50508 = ~n50505 & ~n50507 ;
  assign n50509 = ~n50504 & n50508 ;
  assign n50510 = ~n50496 & n50509 ;
  assign n50511 = \u1_desIn_r_reg[56]/NET0131  & n50510 ;
  assign n50512 = ~\u1_desIn_r_reg[56]/NET0131  & ~n50510 ;
  assign n50513 = ~n50511 & ~n50512 ;
  assign n50515 = ~n50083 & n50103 ;
  assign n50516 = ~n50136 & ~n50515 ;
  assign n50517 = n50097 & ~n50516 ;
  assign n50514 = ~n50097 & n50128 ;
  assign n50518 = ~n50107 & ~n50135 ;
  assign n50519 = ~n50514 & n50518 ;
  assign n50520 = ~n50517 & n50519 ;
  assign n50521 = n50064 & ~n50520 ;
  assign n50522 = ~n50098 & n50119 ;
  assign n50523 = ~n50125 & ~n50402 ;
  assign n50524 = ~n50522 & n50523 ;
  assign n50525 = ~n50064 & ~n50524 ;
  assign n50526 = ~n50100 & n50401 ;
  assign n50527 = ~n50525 & n50526 ;
  assign n50528 = n50064 & ~n50120 ;
  assign n50529 = ~n50112 & ~n50114 ;
  assign n50530 = ~n50281 & n50529 ;
  assign n50531 = ~n50528 & ~n50530 ;
  assign n50532 = ~n50097 & ~n50126 ;
  assign n50533 = ~n50408 & n50532 ;
  assign n50534 = ~n50531 & n50533 ;
  assign n50535 = ~n50527 & ~n50534 ;
  assign n50536 = ~n50521 & ~n50535 ;
  assign n50537 = ~\u1_desIn_r_reg[22]/NET0131  & ~n50536 ;
  assign n50538 = \u1_desIn_r_reg[22]/NET0131  & n50536 ;
  assign n50539 = ~n50537 & ~n50538 ;
  assign n50540 = decrypt_pad & ~\u1_key_r_reg[25]/NET0131  ;
  assign n50541 = ~decrypt_pad & ~\u1_key_r_reg[18]/NET0131  ;
  assign n50542 = ~n50540 & ~n50541 ;
  assign n50543 = \u1_desIn_r_reg[5]/NET0131  & ~n50542 ;
  assign n50544 = ~\u1_desIn_r_reg[5]/NET0131  & n50542 ;
  assign n50545 = ~n50543 & ~n50544 ;
  assign n50546 = decrypt_pad & ~\u1_key_r_reg[33]/NET0131  ;
  assign n50547 = ~decrypt_pad & ~\u1_key_r_reg[26]/NET0131  ;
  assign n50548 = ~n50546 & ~n50547 ;
  assign n50549 = \u1_desIn_r_reg[13]/NET0131  & ~n50548 ;
  assign n50550 = ~\u1_desIn_r_reg[13]/NET0131  & n50548 ;
  assign n50551 = ~n50549 & ~n50550 ;
  assign n50552 = n50545 & n50551 ;
  assign n50553 = ~n50545 & ~n50551 ;
  assign n50554 = decrypt_pad & ~\u1_key_r_reg[5]/NET0131  ;
  assign n50555 = ~decrypt_pad & ~\u1_key_r_reg[55]/NET0131  ;
  assign n50556 = ~n50554 & ~n50555 ;
  assign n50557 = \u1_desIn_r_reg[37]/NET0131  & ~n50556 ;
  assign n50558 = ~\u1_desIn_r_reg[37]/NET0131  & n50556 ;
  assign n50559 = ~n50557 & ~n50558 ;
  assign n50560 = decrypt_pad & ~\u1_key_r_reg[53]/NET0131  ;
  assign n50561 = ~decrypt_pad & ~\u1_key_r_reg[46]/NET0131  ;
  assign n50562 = ~n50560 & ~n50561 ;
  assign n50563 = \u1_desIn_r_reg[63]/NET0131  & ~n50562 ;
  assign n50564 = ~\u1_desIn_r_reg[63]/NET0131  & n50562 ;
  assign n50565 = ~n50563 & ~n50564 ;
  assign n50566 = ~n50559 & ~n50565 ;
  assign n50567 = n50559 & n50565 ;
  assign n50568 = ~n50566 & ~n50567 ;
  assign n50569 = ~n50553 & ~n50568 ;
  assign n50570 = n50559 & ~n50565 ;
  assign n50571 = ~n50551 & n50570 ;
  assign n50572 = decrypt_pad & ~\u1_key_r_reg[34]/NET0131  ;
  assign n50573 = ~decrypt_pad & ~\u1_key_r_reg[27]/NET0131  ;
  assign n50574 = ~n50572 & ~n50573 ;
  assign n50575 = \u1_desIn_r_reg[21]/NET0131  & ~n50574 ;
  assign n50576 = ~\u1_desIn_r_reg[21]/NET0131  & n50574 ;
  assign n50577 = ~n50575 & ~n50576 ;
  assign n50578 = n50571 & ~n50577 ;
  assign n50579 = ~n50559 & n50565 ;
  assign n50580 = ~n50551 & n50579 ;
  assign n50581 = ~n50578 & ~n50580 ;
  assign n50582 = ~n50545 & ~n50581 ;
  assign n50583 = ~n50569 & ~n50582 ;
  assign n50584 = ~n50552 & ~n50583 ;
  assign n50588 = n50552 & ~n50577 ;
  assign n50589 = n50570 & n50588 ;
  assign n50585 = ~n50551 & n50577 ;
  assign n50586 = n50545 & ~n50565 ;
  assign n50587 = n50585 & n50586 ;
  assign n50590 = n50552 & n50579 ;
  assign n50591 = ~n50587 & ~n50590 ;
  assign n50592 = ~n50589 & n50591 ;
  assign n50593 = ~n50584 & n50592 ;
  assign n50594 = decrypt_pad & ~\u1_key_r_reg[17]/NET0131  ;
  assign n50595 = ~decrypt_pad & ~\u1_key_r_reg[10]/NET0131  ;
  assign n50596 = ~n50594 & ~n50595 ;
  assign n50597 = \u1_desIn_r_reg[29]/NET0131  & ~n50596 ;
  assign n50598 = ~\u1_desIn_r_reg[29]/NET0131  & n50596 ;
  assign n50599 = ~n50597 & ~n50598 ;
  assign n50600 = ~n50593 & ~n50599 ;
  assign n50603 = ~n50545 & n50559 ;
  assign n50604 = n50551 & n50570 ;
  assign n50605 = n50545 & n50579 ;
  assign n50606 = ~n50604 & ~n50605 ;
  assign n50607 = ~n50603 & n50606 ;
  assign n50608 = n50577 & ~n50607 ;
  assign n50601 = n50551 & n50566 ;
  assign n50602 = n50545 & n50601 ;
  assign n50609 = n50545 & ~n50559 ;
  assign n50610 = ~n50545 & ~n50565 ;
  assign n50611 = ~n50609 & ~n50610 ;
  assign n50612 = ~n50577 & n50611 ;
  assign n50613 = n50545 & ~n50551 ;
  assign n50614 = n50565 & ~n50603 ;
  assign n50615 = ~n50613 & ~n50614 ;
  assign n50616 = n50612 & ~n50615 ;
  assign n50617 = ~n50602 & ~n50616 ;
  assign n50618 = ~n50608 & n50617 ;
  assign n50619 = n50599 & ~n50618 ;
  assign n50620 = ~n50551 & n50566 ;
  assign n50621 = ~n50545 & n50620 ;
  assign n50622 = ~n50545 & n50551 ;
  assign n50623 = n50559 & n50622 ;
  assign n50624 = ~n50621 & ~n50623 ;
  assign n50625 = n50577 & ~n50624 ;
  assign n50626 = ~n50619 & ~n50625 ;
  assign n50627 = ~n50600 & n50626 ;
  assign n50628 = ~\u1_desIn_r_reg[46]/NET0131  & ~n50627 ;
  assign n50629 = \u1_desIn_r_reg[46]/NET0131  & n50627 ;
  assign n50630 = ~n50628 & ~n50629 ;
  assign n50634 = ~n49518 & n50485 ;
  assign n50635 = n49537 & ~n50634 ;
  assign n50636 = ~n49515 & ~n49561 ;
  assign n50637 = ~n49505 & ~n50636 ;
  assign n50631 = n49498 & n49913 ;
  assign n50638 = ~n49537 & ~n50483 ;
  assign n50639 = ~n50631 & n50638 ;
  assign n50640 = ~n50637 & n50639 ;
  assign n50641 = ~n50635 & ~n50640 ;
  assign n50632 = ~n50486 & ~n50631 ;
  assign n50633 = n49492 & ~n50632 ;
  assign n50642 = n49527 & ~n50633 ;
  assign n50643 = ~n50641 & n50642 ;
  assign n50644 = n49515 & n49913 ;
  assign n50645 = n49537 & ~n50486 ;
  assign n50646 = ~n50485 & n50645 ;
  assign n50647 = ~n50644 & n50646 ;
  assign n50648 = ~n49527 & ~n50647 ;
  assign n50649 = ~n50643 & ~n50648 ;
  assign n50650 = ~n49537 & n50633 ;
  assign n50651 = ~n49537 & n50634 ;
  assign n50652 = ~n49547 & ~n50651 ;
  assign n50653 = n49527 & ~n49537 ;
  assign n50654 = ~n50652 & ~n50653 ;
  assign n50655 = ~n50650 & ~n50654 ;
  assign n50656 = ~n50649 & n50655 ;
  assign n50657 = ~\u1_desIn_r_reg[54]/NET0131  & ~n50656 ;
  assign n50658 = \u1_desIn_r_reg[54]/NET0131  & n50656 ;
  assign n50659 = ~n50657 & ~n50658 ;
  assign n50665 = ~n49346 & ~n49349 ;
  assign n50666 = ~n49579 & n50665 ;
  assign n50667 = n49318 & ~n50666 ;
  assign n50662 = n49312 & n49582 ;
  assign n50660 = ~n49332 & n49577 ;
  assign n50661 = ~n49318 & n50660 ;
  assign n50663 = ~n49312 & n49340 ;
  assign n50664 = n49332 & n50663 ;
  assign n50668 = ~n50661 & ~n50664 ;
  assign n50669 = ~n50662 & n50668 ;
  assign n50670 = ~n50667 & n50669 ;
  assign n50671 = ~n49306 & ~n50670 ;
  assign n50672 = n49363 & n49381 ;
  assign n50673 = ~n50664 & ~n50672 ;
  assign n50674 = ~n49318 & ~n50673 ;
  assign n50676 = n49312 & ~n49341 ;
  assign n50677 = ~n49582 & n50676 ;
  assign n50675 = n49366 & n50660 ;
  assign n50678 = ~n49595 & ~n50675 ;
  assign n50679 = ~n50677 & n50678 ;
  assign n50680 = n49306 & ~n50679 ;
  assign n50681 = ~n50674 & ~n50680 ;
  assign n50682 = ~n50671 & n50681 ;
  assign n50683 = ~\u1_desIn_r_reg[4]/NET0131  & ~n50682 ;
  assign n50684 = \u1_desIn_r_reg[4]/NET0131  & n50682 ;
  assign n50685 = ~n50683 & ~n50684 ;
  assign n50687 = n50545 & n50565 ;
  assign n50688 = ~n50610 & ~n50687 ;
  assign n50689 = n50559 & ~n50688 ;
  assign n50690 = ~n50559 & ~n50687 ;
  assign n50691 = ~n50689 & ~n50690 ;
  assign n50692 = n50545 & n50577 ;
  assign n50693 = n50566 & ~n50692 ;
  assign n50694 = ~n50551 & ~n50693 ;
  assign n50695 = ~n50691 & n50694 ;
  assign n50696 = ~n50580 & ~n50601 ;
  assign n50697 = ~n50577 & ~n50696 ;
  assign n50686 = n50552 & n50570 ;
  assign n50698 = n50599 & ~n50686 ;
  assign n50699 = ~n50697 & n50698 ;
  assign n50700 = ~n50695 & n50699 ;
  assign n50701 = n50577 & ~n50691 ;
  assign n50702 = ~n50577 & ~n50620 ;
  assign n50703 = ~n50689 & n50702 ;
  assign n50704 = ~n50701 & ~n50703 ;
  assign n50705 = ~n50599 & ~n50621 ;
  assign n50706 = ~n50704 & n50705 ;
  assign n50707 = ~n50700 & ~n50706 ;
  assign n50708 = n50551 & n50565 ;
  assign n50709 = ~n50545 & n50708 ;
  assign n50710 = ~n50577 & n50709 ;
  assign n50711 = ~n50545 & n50601 ;
  assign n50712 = ~n50590 & ~n50711 ;
  assign n50713 = n50577 & ~n50712 ;
  assign n50714 = ~n50710 & ~n50713 ;
  assign n50715 = ~n50707 & n50714 ;
  assign n50716 = ~\u1_desIn_r_reg[60]/NET0131  & ~n50715 ;
  assign n50717 = \u1_desIn_r_reg[60]/NET0131  & n50715 ;
  assign n50718 = ~n50716 & ~n50717 ;
  assign n50720 = n49788 & n49823 ;
  assign n50721 = ~n49838 & ~n50720 ;
  assign n50722 = ~n49782 & ~n50721 ;
  assign n50719 = n49782 & ~n49820 ;
  assign n50723 = n49776 & ~n49834 ;
  assign n50724 = ~n50719 & n50723 ;
  assign n50725 = ~n50722 & n50724 ;
  assign n50727 = ~n49782 & n49825 ;
  assign n50728 = ~n49932 & ~n50727 ;
  assign n50729 = ~n49788 & ~n50728 ;
  assign n50730 = ~n49776 & ~n49926 ;
  assign n50731 = ~n49933 & n50730 ;
  assign n50726 = n49782 & n49839 ;
  assign n50732 = ~n49809 & ~n50726 ;
  assign n50733 = n50731 & n50732 ;
  assign n50734 = ~n50729 & n50733 ;
  assign n50735 = ~n50725 & ~n50734 ;
  assign n50736 = ~n49782 & n50315 ;
  assign n50737 = n49795 & n49808 ;
  assign n50738 = ~n49929 & ~n50737 ;
  assign n50739 = n49782 & ~n50738 ;
  assign n50740 = ~n50736 & ~n50739 ;
  assign n50741 = ~n50735 & n50740 ;
  assign n50742 = \u1_desIn_r_reg[10]/NET0131  & n50741 ;
  assign n50743 = ~\u1_desIn_r_reg[10]/NET0131  & ~n50741 ;
  assign n50744 = ~n50742 & ~n50743 ;
  assign n50747 = ~n50571 & n50577 ;
  assign n50748 = ~n50601 & n50747 ;
  assign n50746 = n50545 & n50566 ;
  assign n50749 = ~n50709 & ~n50746 ;
  assign n50750 = n50748 & n50749 ;
  assign n50751 = n50553 & ~n50568 ;
  assign n50752 = ~n50577 & n50606 ;
  assign n50753 = ~n50751 & n50752 ;
  assign n50754 = ~n50750 & ~n50753 ;
  assign n50745 = n50579 & n50622 ;
  assign n50755 = ~n50599 & ~n50745 ;
  assign n50756 = ~n50754 & n50755 ;
  assign n50762 = n50569 & ~n50577 ;
  assign n50760 = ~n50545 & ~n50570 ;
  assign n50761 = n50585 & n50760 ;
  assign n50757 = ~n50570 & ~n50687 ;
  assign n50758 = n50551 & n50577 ;
  assign n50759 = ~n50757 & n50758 ;
  assign n50763 = n50599 & ~n50759 ;
  assign n50764 = ~n50761 & n50763 ;
  assign n50765 = ~n50762 & n50764 ;
  assign n50766 = ~n50582 & n50765 ;
  assign n50767 = ~n50756 & ~n50766 ;
  assign n50768 = n50567 & n50588 ;
  assign n50769 = ~n50567 & n50585 ;
  assign n50770 = n50611 & n50769 ;
  assign n50771 = ~n50768 & ~n50770 ;
  assign n50772 = ~n50767 & n50771 ;
  assign n50773 = ~\u1_desIn_r_reg[58]/NET0131  & ~n50772 ;
  assign n50774 = \u1_desIn_r_reg[58]/NET0131  & n50772 ;
  assign n50775 = ~n50773 & ~n50774 ;
  assign n50776 = n50553 & n50579 ;
  assign n50777 = n50748 & ~n50776 ;
  assign n50778 = ~n50577 & ~n50708 ;
  assign n50779 = ~n50746 & n50778 ;
  assign n50780 = ~n50777 & ~n50779 ;
  assign n50781 = n50599 & ~n50780 ;
  assign n50783 = ~n50545 & n50604 ;
  assign n50788 = ~n50599 & ~n50751 ;
  assign n50789 = ~n50783 & n50788 ;
  assign n50782 = n50612 & ~n50708 ;
  assign n50784 = ~n50609 & n50708 ;
  assign n50785 = ~n50559 & n50613 ;
  assign n50786 = ~n50784 & ~n50785 ;
  assign n50787 = n50577 & ~n50786 ;
  assign n50790 = ~n50782 & ~n50787 ;
  assign n50791 = n50789 & n50790 ;
  assign n50792 = ~n50781 & ~n50791 ;
  assign n50796 = n50567 & n50577 ;
  assign n50797 = n50622 & n50796 ;
  assign n50793 = ~n50559 & n50588 ;
  assign n50794 = n50552 & n50599 ;
  assign n50795 = ~n50567 & n50794 ;
  assign n50798 = ~n50793 & ~n50795 ;
  assign n50799 = ~n50797 & n50798 ;
  assign n50800 = ~n50792 & n50799 ;
  assign n50801 = ~\u1_desIn_r_reg[40]/NET0131  & n50800 ;
  assign n50802 = \u1_desIn_r_reg[40]/NET0131  & ~n50800 ;
  assign n50803 = ~n50801 & ~n50802 ;
  assign n50817 = decrypt_pad & ~\u0_uk_K_r14_reg[43]/NET0131  ;
  assign n50818 = ~decrypt_pad & ~\u0_uk_K_r14_reg[36]/NET0131  ;
  assign n50819 = ~n50817 & ~n50818 ;
  assign n50820 = \u0_R14_reg[29]/NET0131  & ~n50819 ;
  assign n50821 = ~\u0_R14_reg[29]/NET0131  & n50819 ;
  assign n50822 = ~n50820 & ~n50821 ;
  assign n50824 = decrypt_pad & ~\u0_uk_K_r14_reg[44]/NET0131  ;
  assign n50825 = ~decrypt_pad & ~\u0_uk_K_r14_reg[37]/NET0131  ;
  assign n50826 = ~n50824 & ~n50825 ;
  assign n50827 = \u0_R14_reg[30]/NET0131  & ~n50826 ;
  assign n50828 = ~\u0_R14_reg[30]/NET0131  & n50826 ;
  assign n50829 = ~n50827 & ~n50828 ;
  assign n50830 = ~n50822 & n50829 ;
  assign n50831 = n50822 & ~n50829 ;
  assign n50832 = ~n50830 & ~n50831 ;
  assign n50804 = decrypt_pad & ~\u0_uk_K_r14_reg[16]/NET0131  ;
  assign n50805 = ~decrypt_pad & ~\u0_uk_K_r14_reg[9]/NET0131  ;
  assign n50806 = ~n50804 & ~n50805 ;
  assign n50807 = \u0_R14_reg[28]/NET0131  & ~n50806 ;
  assign n50808 = ~\u0_R14_reg[28]/NET0131  & n50806 ;
  assign n50809 = ~n50807 & ~n50808 ;
  assign n50810 = decrypt_pad & ~\u0_uk_K_r14_reg[28]/NET0131  ;
  assign n50811 = ~decrypt_pad & ~\u0_uk_K_r14_reg[21]/NET0131  ;
  assign n50812 = ~n50810 & ~n50811 ;
  assign n50813 = \u0_R14_reg[1]/NET0131  & ~n50812 ;
  assign n50814 = ~\u0_R14_reg[1]/NET0131  & n50812 ;
  assign n50815 = ~n50813 & ~n50814 ;
  assign n50833 = ~n50809 & ~n50815 ;
  assign n50834 = n50832 & n50833 ;
  assign n50835 = n50815 & ~n50822 ;
  assign n50836 = n50809 & ~n50829 ;
  assign n50837 = n50835 & n50836 ;
  assign n50816 = ~n50809 & n50815 ;
  assign n50838 = n50816 & n50830 ;
  assign n50839 = ~n50837 & ~n50838 ;
  assign n50840 = ~n50834 & n50839 ;
  assign n50841 = n50809 & n50830 ;
  assign n50842 = ~n50815 & n50841 ;
  assign n50823 = n50816 & ~n50822 ;
  assign n50843 = decrypt_pad & ~\u0_uk_K_r14_reg[1]/NET0131  ;
  assign n50844 = ~decrypt_pad & ~\u0_uk_K_r14_reg[49]/NET0131  ;
  assign n50845 = ~n50843 & ~n50844 ;
  assign n50846 = \u0_R14_reg[31]/P0001  & ~n50845 ;
  assign n50847 = ~\u0_R14_reg[31]/P0001  & n50845 ;
  assign n50848 = ~n50846 & ~n50847 ;
  assign n50849 = ~n50823 & n50848 ;
  assign n50850 = ~n50842 & n50849 ;
  assign n50851 = n50840 & n50850 ;
  assign n50852 = ~n50815 & n50822 ;
  assign n50853 = n50836 & n50852 ;
  assign n50854 = ~n50848 & ~n50853 ;
  assign n50855 = n50815 & n50822 ;
  assign n50856 = ~n50815 & n50829 ;
  assign n50857 = ~n50809 & n50856 ;
  assign n50858 = ~n50855 & ~n50857 ;
  assign n50859 = n50854 & n50858 ;
  assign n50860 = ~n50851 & ~n50859 ;
  assign n50861 = decrypt_pad & ~\u0_uk_K_r14_reg[7]/NET0131  ;
  assign n50862 = ~decrypt_pad & ~\u0_uk_K_r14_reg[0]/NET0131  ;
  assign n50863 = ~n50861 & ~n50862 ;
  assign n50864 = \u0_R14_reg[32]/NET0131  & ~n50863 ;
  assign n50865 = ~\u0_R14_reg[32]/NET0131  & n50863 ;
  assign n50866 = ~n50864 & ~n50865 ;
  assign n50872 = ~n50853 & ~n50866 ;
  assign n50867 = n50809 & ~n50848 ;
  assign n50868 = ~n50829 & n50867 ;
  assign n50869 = n50822 & n50829 ;
  assign n50870 = n50809 & n50815 ;
  assign n50871 = n50869 & n50870 ;
  assign n50873 = ~n50868 & ~n50871 ;
  assign n50874 = n50872 & n50873 ;
  assign n50875 = ~n50860 & n50874 ;
  assign n50876 = ~n50809 & ~n50822 ;
  assign n50877 = ~n50829 & n50876 ;
  assign n50878 = ~n50841 & ~n50877 ;
  assign n50879 = n50854 & n50878 ;
  assign n50880 = ~n50836 & ~n50852 ;
  assign n50881 = ~n50853 & ~n50880 ;
  assign n50882 = n50848 & ~n50881 ;
  assign n50883 = n50840 & n50882 ;
  assign n50884 = ~n50879 & ~n50883 ;
  assign n50885 = ~n50809 & n50869 ;
  assign n50886 = n50815 & n50885 ;
  assign n50887 = n50866 & ~n50886 ;
  assign n50888 = ~n50884 & n50887 ;
  assign n50889 = ~n50875 & ~n50888 ;
  assign n50890 = ~\u0_L14_reg[5]/P0001  & ~n50889 ;
  assign n50891 = \u0_L14_reg[5]/P0001  & n50889 ;
  assign n50892 = ~n50890 & ~n50891 ;
  assign n50893 = decrypt_pad & ~\u0_uk_K_r14_reg[13]/NET0131  ;
  assign n50894 = ~decrypt_pad & ~\u0_uk_K_r14_reg[6]/NET0131  ;
  assign n50895 = ~n50893 & ~n50894 ;
  assign n50896 = \u0_R14_reg[4]/NET0131  & ~n50895 ;
  assign n50897 = ~\u0_R14_reg[4]/NET0131  & n50895 ;
  assign n50898 = ~n50896 & ~n50897 ;
  assign n50899 = decrypt_pad & ~\u0_uk_K_r14_reg[3]/NET0131  ;
  assign n50900 = ~decrypt_pad & ~\u0_uk_K_r14_reg[53]/NET0131  ;
  assign n50901 = ~n50899 & ~n50900 ;
  assign n50902 = \u0_R14_reg[3]/NET0131  & ~n50901 ;
  assign n50903 = ~\u0_R14_reg[3]/NET0131  & n50901 ;
  assign n50904 = ~n50902 & ~n50903 ;
  assign n50912 = decrypt_pad & ~\u0_uk_K_r14_reg[47]/NET0131  ;
  assign n50913 = ~decrypt_pad & ~\u0_uk_K_r14_reg[40]/NET0131  ;
  assign n50914 = ~n50912 & ~n50913 ;
  assign n50915 = \u0_R14_reg[32]/NET0131  & ~n50914 ;
  assign n50916 = ~\u0_R14_reg[32]/NET0131  & n50914 ;
  assign n50917 = ~n50915 & ~n50916 ;
  assign n50905 = decrypt_pad & ~\u0_uk_K_r14_reg[11]/NET0131  ;
  assign n50906 = ~decrypt_pad & ~\u0_uk_K_r14_reg[4]/NET0131  ;
  assign n50907 = ~n50905 & ~n50906 ;
  assign n50908 = \u0_R14_reg[1]/NET0131  & ~n50907 ;
  assign n50909 = ~\u0_R14_reg[1]/NET0131  & n50907 ;
  assign n50910 = ~n50908 & ~n50909 ;
  assign n50919 = decrypt_pad & ~\u0_uk_K_r14_reg[41]/NET0131  ;
  assign n50920 = ~decrypt_pad & ~\u0_uk_K_r14_reg[34]/NET0131  ;
  assign n50921 = ~n50919 & ~n50920 ;
  assign n50922 = \u0_R14_reg[5]/NET0131  & ~n50921 ;
  assign n50923 = ~\u0_R14_reg[5]/NET0131  & n50921 ;
  assign n50924 = ~n50922 & ~n50923 ;
  assign n50925 = n50910 & ~n50924 ;
  assign n50927 = decrypt_pad & ~\u0_uk_K_r14_reg[26]/NET0131  ;
  assign n50928 = ~decrypt_pad & ~\u0_uk_K_r14_reg[19]/NET0131  ;
  assign n50929 = ~n50927 & ~n50928 ;
  assign n50930 = \u0_R14_reg[2]/NET0131  & ~n50929 ;
  assign n50931 = ~\u0_R14_reg[2]/NET0131  & n50929 ;
  assign n50932 = ~n50930 & ~n50931 ;
  assign n50973 = n50925 & n50932 ;
  assign n50974 = n50917 & n50973 ;
  assign n50937 = n50910 & n50924 ;
  assign n50975 = ~n50917 & n50937 ;
  assign n50976 = ~n50974 & ~n50975 ;
  assign n50977 = n50904 & ~n50976 ;
  assign n50950 = n50904 & ~n50910 ;
  assign n50933 = ~n50917 & n50932 ;
  assign n50971 = ~n50924 & n50933 ;
  assign n50972 = n50950 & n50971 ;
  assign n50951 = n50917 & ~n50932 ;
  assign n50957 = ~n50910 & n50924 ;
  assign n50978 = n50951 & n50957 ;
  assign n50979 = ~n50972 & ~n50978 ;
  assign n50980 = ~n50977 & n50979 ;
  assign n50981 = n50898 & ~n50980 ;
  assign n50938 = n50917 & n50924 ;
  assign n50939 = ~n50904 & n50938 ;
  assign n50940 = ~n50937 & ~n50939 ;
  assign n50941 = n50932 & ~n50940 ;
  assign n50926 = ~n50917 & n50925 ;
  assign n50934 = n50924 & n50933 ;
  assign n50935 = ~n50926 & ~n50934 ;
  assign n50936 = n50904 & ~n50935 ;
  assign n50911 = ~n50904 & n50910 ;
  assign n50918 = n50911 & n50917 ;
  assign n50942 = ~n50910 & ~n50932 ;
  assign n50943 = ~n50924 & n50942 ;
  assign n50944 = ~n50918 & ~n50943 ;
  assign n50945 = ~n50936 & n50944 ;
  assign n50946 = ~n50941 & n50945 ;
  assign n50947 = ~n50898 & ~n50946 ;
  assign n50955 = n50932 & n50937 ;
  assign n50956 = n50917 & n50955 ;
  assign n50953 = n50925 & ~n50932 ;
  assign n50954 = n50917 & n50953 ;
  assign n50958 = ~n50917 & ~n50932 ;
  assign n50959 = n50957 & n50958 ;
  assign n50960 = ~n50954 & ~n50959 ;
  assign n50961 = ~n50956 & n50960 ;
  assign n50962 = ~n50904 & ~n50961 ;
  assign n50963 = ~n50925 & ~n50957 ;
  assign n50964 = ~n50917 & ~n50963 ;
  assign n50965 = n50917 & ~n50924 ;
  assign n50966 = ~n50910 & n50932 ;
  assign n50967 = n50965 & n50966 ;
  assign n50968 = ~n50964 & ~n50967 ;
  assign n50969 = n50898 & ~n50904 ;
  assign n50970 = ~n50968 & n50969 ;
  assign n50948 = n50904 & ~n50932 ;
  assign n50949 = n50926 & n50948 ;
  assign n50952 = n50950 & n50951 ;
  assign n50982 = ~n50949 & ~n50952 ;
  assign n50983 = ~n50970 & n50982 ;
  assign n50984 = ~n50962 & n50983 ;
  assign n50985 = ~n50947 & n50984 ;
  assign n50986 = ~n50981 & n50985 ;
  assign n50987 = \u0_L14_reg[23]/P0001  & ~n50986 ;
  assign n50988 = ~\u0_L14_reg[23]/P0001  & n50986 ;
  assign n50989 = ~n50987 & ~n50988 ;
  assign n50990 = ~n50815 & n50836 ;
  assign n50991 = ~n50822 & n50990 ;
  assign n50992 = ~n50829 & n50852 ;
  assign n50993 = n50809 & n50822 ;
  assign n50994 = ~n50823 & ~n50993 ;
  assign n50995 = ~n50992 & n50994 ;
  assign n50996 = n50848 & ~n50995 ;
  assign n50997 = ~n50991 & ~n50996 ;
  assign n50998 = ~n50866 & ~n50997 ;
  assign n51001 = ~n50836 & ~n50857 ;
  assign n51002 = n50822 & ~n51001 ;
  assign n51005 = n50830 & n50870 ;
  assign n50999 = n50829 & ~n50848 ;
  assign n51000 = n50835 & n50999 ;
  assign n51003 = ~n50815 & n50848 ;
  assign n51004 = n50876 & n51003 ;
  assign n51006 = ~n51000 & ~n51004 ;
  assign n51007 = ~n51005 & n51006 ;
  assign n51008 = ~n51002 & n51007 ;
  assign n51009 = n50866 & ~n51008 ;
  assign n51010 = n50816 & n50831 ;
  assign n51011 = ~n50841 & ~n51010 ;
  assign n51012 = ~n50834 & n51011 ;
  assign n51013 = ~n50848 & ~n51012 ;
  assign n51014 = ~n50822 & ~n50866 ;
  assign n51015 = n50867 & n51014 ;
  assign n51016 = n50816 & n50848 ;
  assign n51017 = n50832 & n51016 ;
  assign n51018 = ~n51015 & ~n51017 ;
  assign n51019 = ~n51013 & n51018 ;
  assign n51020 = ~n51009 & n51019 ;
  assign n51021 = ~n50998 & n51020 ;
  assign n51022 = ~\u0_L14_reg[15]/P0001  & ~n51021 ;
  assign n51023 = \u0_L14_reg[15]/P0001  & n51021 ;
  assign n51024 = ~n51022 & ~n51023 ;
  assign n51031 = ~n50809 & n50855 ;
  assign n51030 = n50809 & n50852 ;
  assign n51032 = ~n50877 & ~n51030 ;
  assign n51033 = ~n51031 & n51032 ;
  assign n51034 = ~n50848 & ~n51033 ;
  assign n51025 = ~n50809 & n50992 ;
  assign n51026 = n50822 & n50870 ;
  assign n51027 = ~n51025 & ~n51026 ;
  assign n51028 = n50848 & ~n51027 ;
  assign n51029 = ~n50829 & n50835 ;
  assign n51035 = ~n50842 & ~n51029 ;
  assign n51036 = ~n50886 & n51035 ;
  assign n51037 = ~n51028 & n51036 ;
  assign n51038 = ~n51034 & n51037 ;
  assign n51039 = n50866 & ~n51038 ;
  assign n51049 = n50848 & ~n50885 ;
  assign n51048 = n50815 & ~n50831 ;
  assign n51050 = ~n50992 & ~n51048 ;
  assign n51051 = n51049 & n51050 ;
  assign n51046 = ~n50809 & ~n50848 ;
  assign n51047 = n50852 & n51046 ;
  assign n51045 = n50870 & n50999 ;
  assign n51052 = ~n50838 & ~n51045 ;
  assign n51053 = ~n51047 & n51052 ;
  assign n51054 = ~n51051 & n51053 ;
  assign n51055 = ~n50866 & ~n51054 ;
  assign n51040 = n50830 & n51003 ;
  assign n51041 = n50822 & n50857 ;
  assign n51042 = ~n50837 & ~n50853 ;
  assign n51043 = ~n51041 & n51042 ;
  assign n51044 = ~n50848 & ~n51043 ;
  assign n51056 = ~n51040 & ~n51044 ;
  assign n51057 = ~n51055 & n51056 ;
  assign n51058 = ~n51039 & n51057 ;
  assign n51059 = \u0_L14_reg[27]/P0001  & n51058 ;
  assign n51060 = ~\u0_L14_reg[27]/P0001  & ~n51058 ;
  assign n51061 = ~n51059 & ~n51060 ;
  assign n51062 = decrypt_pad & ~\u0_uk_K_r14_reg[23]/NET0131  ;
  assign n51063 = ~decrypt_pad & ~\u0_uk_K_r14_reg[16]/NET0131  ;
  assign n51064 = ~n51062 & ~n51063 ;
  assign n51065 = \u0_R14_reg[20]/NET0131  & ~n51064 ;
  assign n51066 = ~\u0_R14_reg[20]/NET0131  & n51064 ;
  assign n51067 = ~n51065 & ~n51066 ;
  assign n51099 = decrypt_pad & ~\u0_uk_K_r14_reg[8]/NET0131  ;
  assign n51100 = ~decrypt_pad & ~\u0_uk_K_r14_reg[1]/NET0131  ;
  assign n51101 = ~n51099 & ~n51100 ;
  assign n51102 = \u0_R14_reg[19]/NET0131  & ~n51101 ;
  assign n51103 = ~\u0_R14_reg[19]/NET0131  & n51101 ;
  assign n51104 = ~n51102 & ~n51103 ;
  assign n51081 = decrypt_pad & ~\u0_uk_K_r14_reg[31]/NET0131  ;
  assign n51082 = ~decrypt_pad & ~\u0_uk_K_r14_reg[51]/NET0131  ;
  assign n51083 = ~n51081 & ~n51082 ;
  assign n51084 = \u0_R14_reg[17]/NET0131  & ~n51083 ;
  assign n51085 = ~\u0_R14_reg[17]/NET0131  & n51083 ;
  assign n51086 = ~n51084 & ~n51085 ;
  assign n51068 = decrypt_pad & ~\u0_uk_K_r14_reg[52]/NET0131  ;
  assign n51069 = ~decrypt_pad & ~\u0_uk_K_r14_reg[45]/NET0131  ;
  assign n51070 = ~n51068 & ~n51069 ;
  assign n51071 = \u0_R14_reg[21]/NET0131  & ~n51070 ;
  assign n51072 = ~\u0_R14_reg[21]/NET0131  & n51070 ;
  assign n51073 = ~n51071 & ~n51072 ;
  assign n51074 = decrypt_pad & ~\u0_uk_K_r14_reg[36]/NET0131  ;
  assign n51075 = ~decrypt_pad & ~\u0_uk_K_r14_reg[29]/NET0131  ;
  assign n51076 = ~n51074 & ~n51075 ;
  assign n51077 = \u0_R14_reg[16]/NET0131  & ~n51076 ;
  assign n51078 = ~\u0_R14_reg[16]/NET0131  & n51076 ;
  assign n51079 = ~n51077 & ~n51078 ;
  assign n51106 = n51073 & n51079 ;
  assign n51107 = ~n51086 & n51106 ;
  assign n51108 = ~n51073 & ~n51079 ;
  assign n51087 = decrypt_pad & ~\u0_uk_K_r14_reg[21]/NET0131  ;
  assign n51088 = ~decrypt_pad & ~\u0_uk_K_r14_reg[14]/NET0131  ;
  assign n51089 = ~n51087 & ~n51088 ;
  assign n51090 = \u0_R14_reg[18]/NET0131  & ~n51089 ;
  assign n51091 = ~\u0_R14_reg[18]/NET0131  & n51089 ;
  assign n51092 = ~n51090 & ~n51091 ;
  assign n51109 = n51073 & n51092 ;
  assign n51110 = ~n51108 & ~n51109 ;
  assign n51111 = ~n51107 & n51110 ;
  assign n51112 = ~n51104 & ~n51111 ;
  assign n51080 = ~n51073 & n51079 ;
  assign n51093 = ~n51086 & n51092 ;
  assign n51094 = ~n51080 & n51093 ;
  assign n51095 = n51080 & n51086 ;
  assign n51096 = n51073 & ~n51079 ;
  assign n51097 = ~n51092 & n51096 ;
  assign n51098 = ~n51095 & ~n51097 ;
  assign n51105 = ~n51098 & n51104 ;
  assign n51113 = ~n51094 & ~n51105 ;
  assign n51114 = ~n51112 & n51113 ;
  assign n51115 = ~n51067 & ~n51114 ;
  assign n51116 = ~n51086 & ~n51092 ;
  assign n51117 = n51080 & n51116 ;
  assign n51118 = n51104 & ~n51117 ;
  assign n51119 = n51093 & n51096 ;
  assign n51120 = n51118 & ~n51119 ;
  assign n51124 = ~n51086 & n51108 ;
  assign n51125 = ~n51092 & n51124 ;
  assign n51123 = n51092 & n51107 ;
  assign n51121 = n51086 & ~n51092 ;
  assign n51122 = n51080 & n51121 ;
  assign n51126 = ~n51104 & ~n51122 ;
  assign n51127 = ~n51123 & n51126 ;
  assign n51128 = ~n51125 & n51127 ;
  assign n51129 = ~n51120 & ~n51128 ;
  assign n51133 = n51086 & n51108 ;
  assign n51134 = n51079 & ~n51092 ;
  assign n51135 = n51073 & n51134 ;
  assign n51136 = ~n51133 & ~n51135 ;
  assign n51137 = n51104 & ~n51136 ;
  assign n51138 = n51106 & n51121 ;
  assign n51130 = n51080 & n51093 ;
  assign n51131 = n51086 & ~n51104 ;
  assign n51132 = n51096 & n51131 ;
  assign n51139 = ~n51130 & ~n51132 ;
  assign n51140 = ~n51138 & n51139 ;
  assign n51141 = ~n51137 & n51140 ;
  assign n51142 = n51067 & ~n51141 ;
  assign n51143 = ~n51129 & ~n51142 ;
  assign n51144 = ~n51115 & n51143 ;
  assign n51145 = \u0_L14_reg[3]/P0001  & n51144 ;
  assign n51146 = ~\u0_L14_reg[3]/P0001  & ~n51144 ;
  assign n51147 = ~n51145 & ~n51146 ;
  assign n51148 = ~n50932 & n50938 ;
  assign n51149 = ~n50934 & ~n51148 ;
  assign n51150 = n50911 & ~n51149 ;
  assign n51153 = ~n50917 & n50924 ;
  assign n51154 = ~n50910 & ~n50965 ;
  assign n51155 = ~n51153 & n51154 ;
  assign n51156 = ~n51148 & ~n51155 ;
  assign n51157 = ~n50942 & ~n51156 ;
  assign n51158 = n50925 & ~n50951 ;
  assign n51159 = ~n50957 & ~n51158 ;
  assign n51160 = n50904 & ~n51159 ;
  assign n51151 = ~n50938 & n50963 ;
  assign n51152 = ~n50904 & n51151 ;
  assign n51161 = ~n50898 & ~n51152 ;
  assign n51162 = ~n51160 & n51161 ;
  assign n51163 = ~n51157 & n51162 ;
  assign n51165 = n50917 & n50963 ;
  assign n51166 = ~n50964 & ~n51165 ;
  assign n51167 = n50932 & ~n51166 ;
  assign n51164 = n50948 & n51151 ;
  assign n51168 = n50898 & ~n50954 ;
  assign n51169 = ~n51164 & n51168 ;
  assign n51170 = ~n51167 & n51169 ;
  assign n51171 = ~n51163 & ~n51170 ;
  assign n51172 = ~n51150 & ~n51171 ;
  assign n51173 = \u0_L14_reg[9]/P0001  & n51172 ;
  assign n51174 = ~\u0_L14_reg[9]/P0001  & ~n51172 ;
  assign n51175 = ~n51173 & ~n51174 ;
  assign n51203 = decrypt_pad & ~\u0_uk_K_r14_reg[39]/P0001  ;
  assign n51204 = ~decrypt_pad & ~\u0_uk_K_r14_reg[32]/NET0131  ;
  assign n51205 = ~n51203 & ~n51204 ;
  assign n51206 = \u0_R14_reg[8]/NET0131  & ~n51205 ;
  assign n51207 = ~\u0_R14_reg[8]/NET0131  & n51205 ;
  assign n51208 = ~n51206 & ~n51207 ;
  assign n51196 = decrypt_pad & ~\u0_uk_K_r14_reg[48]/NET0131  ;
  assign n51197 = ~decrypt_pad & ~\u0_uk_K_r14_reg[41]/NET0131  ;
  assign n51198 = ~n51196 & ~n51197 ;
  assign n51199 = \u0_R14_reg[7]/NET0131  & ~n51198 ;
  assign n51200 = ~\u0_R14_reg[7]/NET0131  & n51198 ;
  assign n51201 = ~n51199 & ~n51200 ;
  assign n51189 = decrypt_pad & ~\u0_uk_K_r14_reg[6]/NET0131  ;
  assign n51190 = ~decrypt_pad & ~\u0_uk_K_r14_reg[24]/NET0131  ;
  assign n51191 = ~n51189 & ~n51190 ;
  assign n51192 = \u0_R14_reg[5]/NET0131  & ~n51191 ;
  assign n51193 = ~\u0_R14_reg[5]/NET0131  & n51191 ;
  assign n51194 = ~n51192 & ~n51193 ;
  assign n51176 = decrypt_pad & ~\u0_uk_K_r14_reg[27]/NET0131  ;
  assign n51177 = ~decrypt_pad & ~\u0_uk_K_r14_reg[20]/NET0131  ;
  assign n51178 = ~n51176 & ~n51177 ;
  assign n51179 = \u0_R14_reg[4]/NET0131  & ~n51178 ;
  assign n51180 = ~\u0_R14_reg[4]/NET0131  & n51178 ;
  assign n51181 = ~n51179 & ~n51180 ;
  assign n51182 = decrypt_pad & ~\u0_uk_K_r14_reg[19]/NET0131  ;
  assign n51183 = ~decrypt_pad & ~\u0_uk_K_r14_reg[12]/NET0131  ;
  assign n51184 = ~n51182 & ~n51183 ;
  assign n51185 = \u0_R14_reg[9]/NET0131  & ~n51184 ;
  assign n51186 = ~\u0_R14_reg[9]/NET0131  & n51184 ;
  assign n51187 = ~n51185 & ~n51186 ;
  assign n51238 = n51181 & ~n51187 ;
  assign n51239 = ~n51194 & n51238 ;
  assign n51210 = decrypt_pad & ~\u0_uk_K_r14_reg[54]/NET0131  ;
  assign n51211 = ~decrypt_pad & ~\u0_uk_K_r14_reg[47]/NET0131  ;
  assign n51212 = ~n51210 & ~n51211 ;
  assign n51213 = \u0_R14_reg[6]/NET0131  & ~n51212 ;
  assign n51214 = ~\u0_R14_reg[6]/NET0131  & n51212 ;
  assign n51215 = ~n51213 & ~n51214 ;
  assign n51240 = n51181 & ~n51215 ;
  assign n51241 = n51187 & n51240 ;
  assign n51242 = ~n51239 & ~n51241 ;
  assign n51243 = ~n51201 & ~n51242 ;
  assign n51234 = ~n51187 & n51194 ;
  assign n51188 = ~n51181 & n51187 ;
  assign n51235 = n51188 & ~n51194 ;
  assign n51236 = ~n51234 & ~n51235 ;
  assign n51237 = n51201 & ~n51236 ;
  assign n51244 = ~n51181 & n51215 ;
  assign n51245 = ~n51194 & n51244 ;
  assign n51246 = ~n51187 & n51245 ;
  assign n51247 = ~n51237 & ~n51246 ;
  assign n51248 = ~n51243 & n51247 ;
  assign n51249 = n51208 & ~n51248 ;
  assign n51218 = ~n51194 & ~n51215 ;
  assign n51219 = ~n51201 & n51215 ;
  assign n51220 = n51194 & n51219 ;
  assign n51221 = ~n51218 & ~n51220 ;
  assign n51222 = ~n51181 & ~n51221 ;
  assign n51209 = n51181 & n51187 ;
  assign n51227 = n51194 & n51209 ;
  assign n51228 = n51201 & n51227 ;
  assign n51216 = n51209 & n51215 ;
  assign n51217 = ~n51194 & n51216 ;
  assign n51223 = n51181 & n51194 ;
  assign n51224 = ~n51187 & n51215 ;
  assign n51225 = n51223 & n51224 ;
  assign n51226 = ~n51187 & n51218 ;
  assign n51229 = ~n51225 & ~n51226 ;
  assign n51230 = ~n51217 & n51229 ;
  assign n51231 = ~n51228 & n51230 ;
  assign n51232 = ~n51222 & n51231 ;
  assign n51233 = ~n51208 & ~n51232 ;
  assign n51195 = n51188 & n51194 ;
  assign n51202 = n51195 & ~n51201 ;
  assign n51250 = ~n51181 & n51234 ;
  assign n51251 = ~n51215 & n51250 ;
  assign n51252 = ~n51216 & ~n51251 ;
  assign n51253 = n51201 & ~n51252 ;
  assign n51254 = ~n51202 & ~n51253 ;
  assign n51255 = ~n51233 & n51254 ;
  assign n51256 = ~n51249 & n51255 ;
  assign n51257 = ~\u0_L14_reg[18]/P0001  & ~n51256 ;
  assign n51258 = \u0_L14_reg[18]/P0001  & n51256 ;
  assign n51259 = ~n51257 & ~n51258 ;
  assign n51287 = decrypt_pad & ~\u0_uk_K_r14_reg[17]/NET0131  ;
  assign n51288 = ~decrypt_pad & ~\u0_uk_K_r14_reg[10]/P0001  ;
  assign n51289 = ~n51287 & ~n51288 ;
  assign n51290 = \u0_R14_reg[12]/NET0131  & ~n51289 ;
  assign n51291 = ~\u0_R14_reg[12]/NET0131  & n51289 ;
  assign n51292 = ~n51290 & ~n51291 ;
  assign n51266 = decrypt_pad & ~\u0_uk_K_r14_reg[25]/NET0131  ;
  assign n51267 = ~decrypt_pad & ~\u0_uk_K_r14_reg[18]/NET0131  ;
  assign n51268 = ~n51266 & ~n51267 ;
  assign n51269 = \u0_R14_reg[9]/NET0131  & ~n51268 ;
  assign n51270 = ~\u0_R14_reg[9]/NET0131  & n51268 ;
  assign n51271 = ~n51269 & ~n51270 ;
  assign n51279 = decrypt_pad & ~\u0_uk_K_r14_reg[33]/NET0131  ;
  assign n51280 = ~decrypt_pad & ~\u0_uk_K_r14_reg[26]/NET0131  ;
  assign n51281 = ~n51279 & ~n51280 ;
  assign n51282 = \u0_R14_reg[10]/NET0131  & ~n51281 ;
  assign n51283 = ~\u0_R14_reg[10]/NET0131  & n51281 ;
  assign n51284 = ~n51282 & ~n51283 ;
  assign n51260 = decrypt_pad & ~\u0_uk_K_r14_reg[5]/NET0131  ;
  assign n51261 = ~decrypt_pad & ~\u0_uk_K_r14_reg[55]/NET0131  ;
  assign n51262 = ~n51260 & ~n51261 ;
  assign n51263 = \u0_R14_reg[13]/NET0131  & ~n51262 ;
  assign n51264 = ~\u0_R14_reg[13]/NET0131  & n51262 ;
  assign n51265 = ~n51263 & ~n51264 ;
  assign n51293 = decrypt_pad & ~\u0_uk_K_r14_reg[53]/NET0131  ;
  assign n51294 = ~decrypt_pad & ~\u0_uk_K_r14_reg[46]/NET0131  ;
  assign n51295 = ~n51293 & ~n51294 ;
  assign n51296 = \u0_R14_reg[8]/NET0131  & ~n51295 ;
  assign n51297 = ~\u0_R14_reg[8]/NET0131  & n51295 ;
  assign n51298 = ~n51296 & ~n51297 ;
  assign n51299 = ~n51265 & n51298 ;
  assign n51300 = ~n51284 & n51299 ;
  assign n51301 = ~n51271 & n51300 ;
  assign n51304 = ~n51265 & ~n51298 ;
  assign n51305 = n51284 & n51304 ;
  assign n51273 = decrypt_pad & ~\u0_uk_K_r14_reg[34]/NET0131  ;
  assign n51274 = ~decrypt_pad & ~\u0_uk_K_r14_reg[27]/NET0131  ;
  assign n51275 = ~n51273 & ~n51274 ;
  assign n51276 = \u0_R14_reg[11]/P0001  & ~n51275 ;
  assign n51277 = ~\u0_R14_reg[11]/P0001  & n51275 ;
  assign n51278 = ~n51276 & ~n51277 ;
  assign n51302 = n51265 & ~n51298 ;
  assign n51303 = ~n51284 & n51302 ;
  assign n51306 = n51278 & ~n51303 ;
  assign n51307 = ~n51305 & n51306 ;
  assign n51308 = ~n51301 & n51307 ;
  assign n51310 = n51271 & n51304 ;
  assign n51309 = n51284 & n51298 ;
  assign n51311 = ~n51278 & ~n51309 ;
  assign n51312 = ~n51310 & n51311 ;
  assign n51313 = ~n51308 & ~n51312 ;
  assign n51314 = n51292 & ~n51313 ;
  assign n51272 = ~n51265 & n51271 ;
  assign n51317 = ~n51272 & n51309 ;
  assign n51318 = n51271 & ~n51284 ;
  assign n51319 = ~n51265 & n51318 ;
  assign n51320 = ~n51317 & ~n51319 ;
  assign n51321 = n51278 & ~n51320 ;
  assign n51327 = ~n51272 & ~n51278 ;
  assign n51326 = ~n51271 & ~n51298 ;
  assign n51328 = ~n51309 & ~n51326 ;
  assign n51329 = n51327 & n51328 ;
  assign n51322 = ~n51271 & ~n51284 ;
  assign n51323 = n51265 & n51298 ;
  assign n51324 = ~n51304 & ~n51323 ;
  assign n51325 = n51322 & ~n51324 ;
  assign n51315 = ~n51271 & n51284 ;
  assign n51316 = n51302 & n51315 ;
  assign n51330 = ~n51292 & ~n51316 ;
  assign n51331 = ~n51325 & n51330 ;
  assign n51332 = ~n51329 & n51331 ;
  assign n51333 = ~n51321 & n51332 ;
  assign n51334 = ~n51314 & ~n51333 ;
  assign n51338 = n51265 & n51278 ;
  assign n51339 = ~n51271 & n51309 ;
  assign n51340 = n51338 & n51339 ;
  assign n51285 = ~n51278 & n51284 ;
  assign n51286 = n51272 & n51285 ;
  assign n51335 = n51284 & n51292 ;
  assign n51336 = n51271 & ~n51323 ;
  assign n51337 = n51335 & n51336 ;
  assign n51341 = ~n51286 & ~n51337 ;
  assign n51342 = ~n51340 & n51341 ;
  assign n51343 = ~n51334 & n51342 ;
  assign n51344 = \u0_L14_reg[30]/P0001  & ~n51343 ;
  assign n51345 = ~\u0_L14_reg[30]/P0001  & n51343 ;
  assign n51346 = ~n51344 & ~n51345 ;
  assign n51375 = ~n51299 & ~n51322 ;
  assign n51376 = ~n51278 & ~n51375 ;
  assign n51374 = n51278 & ~n51322 ;
  assign n51377 = ~n51302 & ~n51374 ;
  assign n51378 = ~n51376 & n51377 ;
  assign n51367 = ~n51271 & ~n51278 ;
  assign n51368 = n51303 & n51367 ;
  assign n51369 = ~n51301 & ~n51368 ;
  assign n51370 = ~n51271 & n51298 ;
  assign n51371 = n51278 & n51284 ;
  assign n51372 = ~n51304 & n51371 ;
  assign n51373 = ~n51370 & n51372 ;
  assign n51379 = n51369 & ~n51373 ;
  assign n51380 = ~n51378 & n51379 ;
  assign n51381 = n51292 & ~n51380 ;
  assign n51347 = n51304 & ~n51322 ;
  assign n51348 = ~n51303 & ~n51339 ;
  assign n51349 = ~n51347 & n51348 ;
  assign n51350 = n51278 & ~n51349 ;
  assign n51351 = ~n51265 & n51339 ;
  assign n51352 = ~n51350 & ~n51351 ;
  assign n51353 = ~n51292 & ~n51352 ;
  assign n51361 = n51284 & n51302 ;
  assign n51362 = n51272 & n51298 ;
  assign n51363 = ~n51361 & ~n51362 ;
  assign n51364 = ~n51325 & n51363 ;
  assign n51365 = ~n51278 & ~n51292 ;
  assign n51366 = ~n51364 & n51365 ;
  assign n51355 = n51271 & ~n51298 ;
  assign n51356 = n51278 & n51355 ;
  assign n51357 = ~n51284 & n51356 ;
  assign n51358 = n51265 & n51357 ;
  assign n51354 = n51278 & n51301 ;
  assign n51359 = n51271 & n51285 ;
  assign n51360 = n51323 & n51359 ;
  assign n51382 = ~n51354 & ~n51360 ;
  assign n51383 = ~n51358 & n51382 ;
  assign n51384 = ~n51366 & n51383 ;
  assign n51385 = ~n51353 & n51384 ;
  assign n51386 = ~n51381 & n51385 ;
  assign n51387 = \u0_L14_reg[24]/P0001  & n51386 ;
  assign n51388 = ~\u0_L14_reg[24]/P0001  & ~n51386 ;
  assign n51389 = ~n51387 & ~n51388 ;
  assign n51390 = ~n51355 & ~n51370 ;
  assign n51393 = n51265 & n51390 ;
  assign n51408 = ~n51356 & ~n51370 ;
  assign n51409 = ~n51265 & ~n51408 ;
  assign n51410 = ~n51393 & ~n51409 ;
  assign n51411 = ~n51284 & ~n51410 ;
  assign n51407 = n51271 & n51361 ;
  assign n51412 = ~n51300 & ~n51305 ;
  assign n51413 = ~n51278 & ~n51412 ;
  assign n51414 = ~n51407 & ~n51413 ;
  assign n51415 = ~n51411 & n51414 ;
  assign n51416 = n51292 & ~n51415 ;
  assign n51394 = ~n51284 & n51304 ;
  assign n51395 = ~n51393 & ~n51394 ;
  assign n51396 = ~n51278 & ~n51395 ;
  assign n51397 = ~n51271 & n51394 ;
  assign n51391 = n51338 & ~n51390 ;
  assign n51392 = n51278 & n51362 ;
  assign n51398 = ~n51391 & ~n51392 ;
  assign n51399 = ~n51397 & n51398 ;
  assign n51400 = ~n51396 & n51399 ;
  assign n51401 = ~n51292 & ~n51400 ;
  assign n51402 = n51284 & n51362 ;
  assign n51403 = ~n51271 & n51305 ;
  assign n51404 = ~n51402 & ~n51403 ;
  assign n51405 = n51278 & ~n51404 ;
  assign n51406 = n51309 & n51367 ;
  assign n51417 = ~n51405 & ~n51406 ;
  assign n51418 = ~n51401 & n51417 ;
  assign n51419 = ~n51416 & n51418 ;
  assign n51420 = \u0_L14_reg[16]/P0001  & n51419 ;
  assign n51421 = ~\u0_L14_reg[16]/P0001  & ~n51419 ;
  assign n51422 = ~n51420 & ~n51421 ;
  assign n51453 = decrypt_pad & ~\u0_uk_K_r13_reg[7]/NET0131  ;
  assign n51454 = ~decrypt_pad & ~\u0_uk_K_r13_reg[45]/NET0131  ;
  assign n51455 = ~n51453 & ~n51454 ;
  assign n51456 = \u0_R13_reg[27]/P0001  & ~n51455 ;
  assign n51457 = ~\u0_R13_reg[27]/P0001  & n51455 ;
  assign n51458 = ~n51456 & ~n51457 ;
  assign n51423 = decrypt_pad & ~\u0_uk_K_r13_reg[45]/NET0131  ;
  assign n51424 = ~decrypt_pad & ~\u0_uk_K_r13_reg[51]/NET0131  ;
  assign n51425 = ~n51423 & ~n51424 ;
  assign n51426 = \u0_R13_reg[29]/NET0131  & ~n51425 ;
  assign n51427 = ~\u0_R13_reg[29]/NET0131  & n51425 ;
  assign n51428 = ~n51426 & ~n51427 ;
  assign n51429 = decrypt_pad & ~\u0_uk_K_r13_reg[44]/NET0131  ;
  assign n51430 = ~decrypt_pad & ~\u0_uk_K_r13_reg[23]/NET0131  ;
  assign n51431 = ~n51429 & ~n51430 ;
  assign n51432 = \u0_R13_reg[25]/NET0131  & ~n51431 ;
  assign n51433 = ~\u0_R13_reg[25]/NET0131  & n51431 ;
  assign n51434 = ~n51432 & ~n51433 ;
  assign n51436 = decrypt_pad & ~\u0_uk_K_r13_reg[29]/NET0131  ;
  assign n51437 = ~decrypt_pad & ~\u0_uk_K_r13_reg[8]/NET0131  ;
  assign n51438 = ~n51436 & ~n51437 ;
  assign n51439 = \u0_R13_reg[26]/NET0131  & ~n51438 ;
  assign n51440 = ~\u0_R13_reg[26]/NET0131  & n51438 ;
  assign n51441 = ~n51439 & ~n51440 ;
  assign n51500 = ~n51434 & ~n51441 ;
  assign n51443 = decrypt_pad & ~\u0_uk_K_r13_reg[9]/NET0131  ;
  assign n51444 = ~decrypt_pad & ~\u0_uk_K_r13_reg[43]/NET0131  ;
  assign n51445 = ~n51443 & ~n51444 ;
  assign n51446 = \u0_R13_reg[24]/NET0131  & ~n51445 ;
  assign n51447 = ~\u0_R13_reg[24]/NET0131  & n51445 ;
  assign n51448 = ~n51446 & ~n51447 ;
  assign n51450 = ~n51434 & n51448 ;
  assign n51471 = n51434 & ~n51448 ;
  assign n51472 = ~n51450 & ~n51471 ;
  assign n51480 = ~n51441 & ~n51448 ;
  assign n51501 = ~n51472 & ~n51480 ;
  assign n51502 = ~n51500 & ~n51501 ;
  assign n51503 = ~n51428 & ~n51502 ;
  assign n51460 = ~n51434 & ~n51448 ;
  assign n51461 = n51428 & n51441 ;
  assign n51504 = n51460 & n51461 ;
  assign n51505 = ~n51503 & ~n51504 ;
  assign n51506 = n51458 & ~n51505 ;
  assign n51435 = n51428 & n51434 ;
  assign n51442 = n51435 & ~n51441 ;
  assign n51449 = n51442 & n51448 ;
  assign n51451 = n51441 & n51450 ;
  assign n51452 = ~n51449 & ~n51451 ;
  assign n51459 = ~n51452 & n51458 ;
  assign n51473 = n51441 & n51448 ;
  assign n51474 = n51428 & ~n51458 ;
  assign n51475 = ~n51473 & n51474 ;
  assign n51476 = ~n51472 & n51475 ;
  assign n51462 = ~n51428 & ~n51441 ;
  assign n51463 = ~n51461 & ~n51462 ;
  assign n51464 = n51460 & ~n51463 ;
  assign n51465 = decrypt_pad & ~\u0_uk_K_r13_reg[49]/NET0131  ;
  assign n51466 = ~decrypt_pad & ~\u0_uk_K_r13_reg[28]/NET0131  ;
  assign n51467 = ~n51465 & ~n51466 ;
  assign n51468 = \u0_R13_reg[28]/NET0131  & ~n51467 ;
  assign n51469 = ~\u0_R13_reg[28]/NET0131  & n51467 ;
  assign n51470 = ~n51468 & ~n51469 ;
  assign n51477 = ~n51464 & n51470 ;
  assign n51478 = ~n51476 & n51477 ;
  assign n51479 = ~n51459 & n51478 ;
  assign n51487 = ~n51428 & ~n51434 ;
  assign n51488 = ~n51448 & n51487 ;
  assign n51489 = n51441 & n51488 ;
  assign n51490 = ~n51428 & n51448 ;
  assign n51491 = n51434 & n51490 ;
  assign n51492 = n51428 & n51473 ;
  assign n51493 = ~n51491 & ~n51492 ;
  assign n51494 = ~n51489 & n51493 ;
  assign n51495 = ~n51458 & ~n51494 ;
  assign n51484 = n51448 & n51474 ;
  assign n51483 = ~n51450 & ~n51474 ;
  assign n51485 = ~n51441 & ~n51483 ;
  assign n51486 = ~n51484 & n51485 ;
  assign n51481 = ~n51473 & ~n51480 ;
  assign n51482 = n51435 & ~n51481 ;
  assign n51496 = ~n51470 & ~n51482 ;
  assign n51497 = ~n51486 & n51496 ;
  assign n51498 = ~n51495 & n51497 ;
  assign n51499 = ~n51479 & ~n51498 ;
  assign n51507 = n51434 & ~n51458 ;
  assign n51508 = ~n51481 & n51507 ;
  assign n51509 = ~n51499 & ~n51508 ;
  assign n51510 = ~n51506 & n51509 ;
  assign n51511 = \u0_L13_reg[22]/NET0131  & n51510 ;
  assign n51512 = ~\u0_L13_reg[22]/NET0131  & ~n51510 ;
  assign n51513 = ~n51511 & ~n51512 ;
  assign n51514 = decrypt_pad & ~\u0_uk_K_r13_reg[20]/NET0131  ;
  assign n51515 = ~decrypt_pad & ~\u0_uk_K_r13_reg[24]/NET0131  ;
  assign n51516 = ~n51514 & ~n51515 ;
  assign n51517 = \u0_R13_reg[4]/NET0131  & ~n51516 ;
  assign n51518 = ~\u0_R13_reg[4]/NET0131  & n51516 ;
  assign n51519 = ~n51517 & ~n51518 ;
  assign n51533 = decrypt_pad & ~\u0_uk_K_r13_reg[48]/NET0131  ;
  assign n51534 = ~decrypt_pad & ~\u0_uk_K_r13_reg[27]/NET0131  ;
  assign n51535 = ~n51533 & ~n51534 ;
  assign n51536 = \u0_R13_reg[5]/NET0131  & ~n51535 ;
  assign n51537 = ~\u0_R13_reg[5]/NET0131  & n51535 ;
  assign n51538 = ~n51536 & ~n51537 ;
  assign n51539 = decrypt_pad & ~\u0_uk_K_r13_reg[54]/NET0131  ;
  assign n51540 = ~decrypt_pad & ~\u0_uk_K_r13_reg[33]/NET0131  ;
  assign n51541 = ~n51539 & ~n51540 ;
  assign n51542 = \u0_R13_reg[32]/NET0131  & ~n51541 ;
  assign n51543 = ~\u0_R13_reg[32]/NET0131  & n51541 ;
  assign n51544 = ~n51542 & ~n51543 ;
  assign n51545 = ~n51538 & ~n51544 ;
  assign n51548 = decrypt_pad & ~\u0_uk_K_r13_reg[18]/NET0131  ;
  assign n51549 = ~decrypt_pad & ~\u0_uk_K_r13_reg[54]/NET0131  ;
  assign n51550 = ~n51548 & ~n51549 ;
  assign n51551 = \u0_R13_reg[1]/NET0131  & ~n51550 ;
  assign n51552 = ~\u0_R13_reg[1]/NET0131  & n51550 ;
  assign n51553 = ~n51551 & ~n51552 ;
  assign n51520 = decrypt_pad & ~\u0_uk_K_r13_reg[10]/NET0131  ;
  assign n51521 = ~decrypt_pad & ~\u0_uk_K_r13_reg[46]/NET0131  ;
  assign n51522 = ~n51520 & ~n51521 ;
  assign n51523 = \u0_R13_reg[3]/NET0131  & ~n51522 ;
  assign n51524 = ~\u0_R13_reg[3]/NET0131  & n51522 ;
  assign n51525 = ~n51523 & ~n51524 ;
  assign n51526 = decrypt_pad & ~\u0_uk_K_r13_reg[33]/NET0131  ;
  assign n51527 = ~decrypt_pad & ~\u0_uk_K_r13_reg[12]/NET0131  ;
  assign n51528 = ~n51526 & ~n51527 ;
  assign n51529 = \u0_R13_reg[2]/NET0131  & ~n51528 ;
  assign n51530 = ~\u0_R13_reg[2]/NET0131  & n51528 ;
  assign n51531 = ~n51529 & ~n51530 ;
  assign n51573 = n51525 & ~n51531 ;
  assign n51574 = n51553 & ~n51573 ;
  assign n51575 = ~n51544 & ~n51574 ;
  assign n51576 = ~n51531 & ~n51553 ;
  assign n51577 = ~n51538 & n51576 ;
  assign n51578 = ~n51575 & ~n51577 ;
  assign n51579 = ~n51545 & ~n51578 ;
  assign n51559 = n51538 & ~n51553 ;
  assign n51580 = n51531 & n51545 ;
  assign n51581 = ~n51559 & ~n51580 ;
  assign n51582 = n51525 & ~n51581 ;
  assign n51556 = n51544 & ~n51553 ;
  assign n51583 = ~n51525 & n51544 ;
  assign n51584 = n51531 & ~n51553 ;
  assign n51585 = ~n51583 & ~n51584 ;
  assign n51586 = ~n51556 & ~n51585 ;
  assign n51587 = ~n51582 & ~n51586 ;
  assign n51588 = ~n51579 & n51587 ;
  assign n51589 = n51519 & ~n51588 ;
  assign n51557 = ~n51538 & n51556 ;
  assign n51558 = n51531 & n51557 ;
  assign n51560 = ~n51531 & ~n51544 ;
  assign n51561 = ~n51559 & n51560 ;
  assign n51562 = ~n51558 & ~n51561 ;
  assign n51563 = ~n51525 & ~n51562 ;
  assign n51532 = n51525 & n51531 ;
  assign n51546 = n51538 & n51544 ;
  assign n51547 = ~n51545 & ~n51546 ;
  assign n51554 = n51547 & n51553 ;
  assign n51555 = n51532 & n51554 ;
  assign n51564 = ~n51525 & n51553 ;
  assign n51565 = n51546 & ~n51564 ;
  assign n51566 = ~n51538 & n51553 ;
  assign n51567 = ~n51544 & n51566 ;
  assign n51568 = ~n51565 & ~n51567 ;
  assign n51569 = ~n51531 & ~n51568 ;
  assign n51570 = ~n51555 & ~n51569 ;
  assign n51571 = ~n51563 & n51570 ;
  assign n51572 = ~n51519 & ~n51571 ;
  assign n51590 = n51525 & ~n51553 ;
  assign n51591 = ~n51531 & n51544 ;
  assign n51592 = ~n51580 & ~n51591 ;
  assign n51593 = n51590 & ~n51592 ;
  assign n51594 = n51546 & n51553 ;
  assign n51595 = n51531 & n51594 ;
  assign n51596 = ~n51531 & n51566 ;
  assign n51597 = n51538 & ~n51544 ;
  assign n51598 = n51584 & n51597 ;
  assign n51599 = ~n51596 & ~n51598 ;
  assign n51600 = ~n51595 & n51599 ;
  assign n51601 = ~n51525 & ~n51600 ;
  assign n51602 = ~n51593 & ~n51601 ;
  assign n51603 = ~n51572 & n51602 ;
  assign n51604 = ~n51589 & n51603 ;
  assign n51605 = ~\u0_L13_reg[31]/NET0131  & ~n51604 ;
  assign n51606 = \u0_L13_reg[31]/NET0131  & n51604 ;
  assign n51607 = ~n51605 & ~n51606 ;
  assign n51608 = decrypt_pad & ~\u0_uk_K_r13_reg[14]/NET0131  ;
  assign n51609 = ~decrypt_pad & ~\u0_uk_K_r13_reg[52]/P0001  ;
  assign n51610 = ~n51608 & ~n51609 ;
  assign n51611 = \u0_R13_reg[32]/NET0131  & ~n51610 ;
  assign n51612 = ~\u0_R13_reg[32]/NET0131  & n51610 ;
  assign n51613 = ~n51611 & ~n51612 ;
  assign n51647 = decrypt_pad & ~\u0_uk_K_r13_reg[8]/NET0131  ;
  assign n51648 = ~decrypt_pad & ~\u0_uk_K_r13_reg[42]/NET0131  ;
  assign n51649 = ~n51647 & ~n51648 ;
  assign n51650 = \u0_R13_reg[31]/NET0131  & ~n51649 ;
  assign n51651 = ~\u0_R13_reg[31]/NET0131  & n51649 ;
  assign n51652 = ~n51650 & ~n51651 ;
  assign n51626 = decrypt_pad & ~\u0_uk_K_r13_reg[50]/NET0131  ;
  assign n51627 = ~decrypt_pad & ~\u0_uk_K_r13_reg[29]/NET0131  ;
  assign n51628 = ~n51626 & ~n51627 ;
  assign n51629 = \u0_R13_reg[29]/NET0131  & ~n51628 ;
  assign n51630 = ~\u0_R13_reg[29]/NET0131  & n51628 ;
  assign n51631 = ~n51629 & ~n51630 ;
  assign n51633 = decrypt_pad & ~\u0_uk_K_r13_reg[35]/NET0131  ;
  assign n51634 = ~decrypt_pad & ~\u0_uk_K_r13_reg[14]/NET0131  ;
  assign n51635 = ~n51633 & ~n51634 ;
  assign n51636 = \u0_R13_reg[1]/NET0131  & ~n51635 ;
  assign n51637 = ~\u0_R13_reg[1]/NET0131  & n51635 ;
  assign n51638 = ~n51636 & ~n51637 ;
  assign n51614 = decrypt_pad & ~\u0_uk_K_r13_reg[51]/NET0131  ;
  assign n51615 = ~decrypt_pad & ~\u0_uk_K_r13_reg[30]/NET0131  ;
  assign n51616 = ~n51614 & ~n51615 ;
  assign n51617 = \u0_R13_reg[30]/NET0131  & ~n51616 ;
  assign n51618 = ~\u0_R13_reg[30]/NET0131  & n51616 ;
  assign n51619 = ~n51617 & ~n51618 ;
  assign n51620 = decrypt_pad & ~\u0_uk_K_r13_reg[23]/NET0131  ;
  assign n51621 = ~decrypt_pad & ~\u0_uk_K_r13_reg[2]/NET0131  ;
  assign n51622 = ~n51620 & ~n51621 ;
  assign n51623 = \u0_R13_reg[28]/NET0131  & ~n51622 ;
  assign n51624 = ~\u0_R13_reg[28]/NET0131  & n51622 ;
  assign n51625 = ~n51623 & ~n51624 ;
  assign n51654 = ~n51619 & n51625 ;
  assign n51656 = ~n51638 & n51654 ;
  assign n51657 = n51631 & n51656 ;
  assign n51668 = n51631 & ~n51638 ;
  assign n51669 = ~n51654 & ~n51668 ;
  assign n51670 = ~n51657 & ~n51669 ;
  assign n51671 = n51652 & ~n51670 ;
  assign n51672 = ~n51619 & ~n51631 ;
  assign n51673 = ~n51625 & n51672 ;
  assign n51674 = n51625 & ~n51631 ;
  assign n51675 = n51619 & n51674 ;
  assign n51676 = ~n51652 & ~n51675 ;
  assign n51677 = ~n51673 & n51676 ;
  assign n51678 = ~n51671 & ~n51677 ;
  assign n51659 = n51619 & ~n51625 ;
  assign n51679 = n51631 & n51659 ;
  assign n51680 = n51638 & n51679 ;
  assign n51681 = ~n51678 & ~n51680 ;
  assign n51682 = n51613 & ~n51681 ;
  assign n51641 = ~n51631 & ~n51638 ;
  assign n51642 = n51619 & n51641 ;
  assign n51643 = n51625 & n51642 ;
  assign n51644 = ~n51625 & n51638 ;
  assign n51645 = ~n51631 & n51644 ;
  assign n51646 = ~n51643 & ~n51645 ;
  assign n51653 = ~n51646 & n51652 ;
  assign n51632 = n51625 & n51631 ;
  assign n51639 = n51632 & n51638 ;
  assign n51640 = n51619 & n51639 ;
  assign n51655 = ~n51652 & n51654 ;
  assign n51663 = ~n51640 & ~n51655 ;
  assign n51660 = ~n51638 & ~n51659 ;
  assign n51658 = ~n51631 & n51638 ;
  assign n51661 = ~n51652 & ~n51658 ;
  assign n51662 = ~n51660 & n51661 ;
  assign n51664 = ~n51657 & ~n51662 ;
  assign n51665 = n51663 & n51664 ;
  assign n51666 = ~n51653 & n51665 ;
  assign n51667 = ~n51613 & ~n51666 ;
  assign n51683 = n51655 & n51668 ;
  assign n51684 = ~n51638 & n51679 ;
  assign n51685 = ~n51638 & n51673 ;
  assign n51686 = ~n51684 & ~n51685 ;
  assign n51687 = n51654 & n51658 ;
  assign n51688 = n51619 & n51645 ;
  assign n51689 = ~n51687 & ~n51688 ;
  assign n51690 = n51686 & n51689 ;
  assign n51691 = n51652 & ~n51690 ;
  assign n51692 = ~n51683 & ~n51691 ;
  assign n51693 = ~n51667 & n51692 ;
  assign n51694 = ~n51682 & n51693 ;
  assign n51695 = \u0_L13_reg[5]/NET0131  & ~n51694 ;
  assign n51696 = ~\u0_L13_reg[5]/NET0131  & n51694 ;
  assign n51697 = ~n51695 & ~n51696 ;
  assign n51704 = decrypt_pad & ~\u0_uk_K_r13_reg[27]/NET0131  ;
  assign n51705 = ~decrypt_pad & ~\u0_uk_K_r13_reg[6]/NET0131  ;
  assign n51706 = ~n51704 & ~n51705 ;
  assign n51707 = \u0_R13_reg[17]/NET0131  & ~n51706 ;
  assign n51708 = ~\u0_R13_reg[17]/NET0131  & n51706 ;
  assign n51709 = ~n51707 & ~n51708 ;
  assign n51710 = decrypt_pad & ~\u0_uk_K_r13_reg[5]/NET0131  ;
  assign n51711 = ~decrypt_pad & ~\u0_uk_K_r13_reg[41]/NET0131  ;
  assign n51712 = ~n51710 & ~n51711 ;
  assign n51713 = \u0_R13_reg[13]/NET0131  & ~n51712 ;
  assign n51714 = ~\u0_R13_reg[13]/NET0131  & n51712 ;
  assign n51715 = ~n51713 & ~n51714 ;
  assign n51698 = decrypt_pad & ~\u0_uk_K_r13_reg[11]/NET0131  ;
  assign n51699 = ~decrypt_pad & ~\u0_uk_K_r13_reg[47]/NET0131  ;
  assign n51700 = ~n51698 & ~n51699 ;
  assign n51701 = \u0_R13_reg[12]/NET0131  & ~n51700 ;
  assign n51702 = ~\u0_R13_reg[12]/NET0131  & n51700 ;
  assign n51703 = ~n51701 & ~n51702 ;
  assign n51718 = decrypt_pad & ~\u0_uk_K_r13_reg[6]/NET0131  ;
  assign n51719 = ~decrypt_pad & ~\u0_uk_K_r13_reg[10]/NET0131  ;
  assign n51720 = ~n51718 & ~n51719 ;
  assign n51721 = \u0_R13_reg[14]/NET0131  & ~n51720 ;
  assign n51722 = ~\u0_R13_reg[14]/NET0131  & n51720 ;
  assign n51723 = ~n51721 & ~n51722 ;
  assign n51749 = n51703 & ~n51723 ;
  assign n51750 = ~n51715 & n51749 ;
  assign n51751 = n51709 & n51750 ;
  assign n51733 = decrypt_pad & ~\u0_uk_K_r13_reg[39]/NET0131  ;
  assign n51734 = ~decrypt_pad & ~\u0_uk_K_r13_reg[18]/NET0131  ;
  assign n51735 = ~n51733 & ~n51734 ;
  assign n51736 = \u0_R13_reg[15]/NET0131  & ~n51735 ;
  assign n51737 = ~\u0_R13_reg[15]/NET0131  & n51735 ;
  assign n51738 = ~n51736 & ~n51737 ;
  assign n51746 = n51715 & n51738 ;
  assign n51747 = n51723 & n51746 ;
  assign n51748 = ~n51703 & n51747 ;
  assign n51752 = decrypt_pad & ~\u0_uk_K_r13_reg[47]/NET0131  ;
  assign n51753 = ~decrypt_pad & ~\u0_uk_K_r13_reg[26]/NET0131  ;
  assign n51754 = ~n51752 & ~n51753 ;
  assign n51755 = \u0_R13_reg[16]/NET0131  & ~n51754 ;
  assign n51756 = ~\u0_R13_reg[16]/NET0131  & n51754 ;
  assign n51757 = ~n51755 & ~n51756 ;
  assign n51758 = ~n51748 & ~n51757 ;
  assign n51759 = ~n51751 & n51758 ;
  assign n51729 = n51703 & ~n51709 ;
  assign n51742 = ~n51703 & n51709 ;
  assign n51743 = ~n51729 & ~n51742 ;
  assign n51725 = ~n51703 & ~n51715 ;
  assign n51740 = n51703 & n51715 ;
  assign n51741 = ~n51725 & ~n51740 ;
  assign n51744 = n51738 & ~n51741 ;
  assign n51745 = n51743 & n51744 ;
  assign n51716 = ~n51703 & ~n51709 ;
  assign n51717 = n51715 & n51716 ;
  assign n51724 = n51717 & n51723 ;
  assign n51726 = ~n51709 & ~n51723 ;
  assign n51727 = n51725 & n51726 ;
  assign n51728 = ~n51724 & ~n51727 ;
  assign n51730 = n51723 & n51729 ;
  assign n51731 = n51709 & ~n51715 ;
  assign n51732 = ~n51730 & ~n51731 ;
  assign n51739 = ~n51732 & ~n51738 ;
  assign n51760 = n51728 & ~n51739 ;
  assign n51761 = ~n51745 & n51760 ;
  assign n51762 = n51759 & n51761 ;
  assign n51768 = ~n51709 & n51725 ;
  assign n51769 = n51723 & ~n51768 ;
  assign n51767 = ~n51723 & ~n51741 ;
  assign n51770 = ~n51738 & ~n51767 ;
  assign n51771 = ~n51769 & n51770 ;
  assign n51763 = n51729 & n51746 ;
  assign n51764 = n51715 & n51742 ;
  assign n51765 = ~n51723 & n51764 ;
  assign n51766 = ~n51763 & ~n51765 ;
  assign n51774 = n51738 & n51742 ;
  assign n51775 = ~n51715 & n51774 ;
  assign n51772 = n51709 & n51723 ;
  assign n51773 = n51740 & n51772 ;
  assign n51776 = n51757 & ~n51773 ;
  assign n51777 = ~n51775 & n51776 ;
  assign n51778 = n51766 & n51777 ;
  assign n51779 = ~n51771 & n51778 ;
  assign n51780 = ~n51762 & ~n51779 ;
  assign n51785 = ~n51738 & n51765 ;
  assign n51781 = ~n51715 & n51738 ;
  assign n51782 = ~n51703 & n51726 ;
  assign n51783 = ~n51730 & ~n51782 ;
  assign n51784 = n51781 & ~n51783 ;
  assign n51786 = ~n51723 & n51763 ;
  assign n51787 = ~n51784 & ~n51786 ;
  assign n51788 = ~n51785 & n51787 ;
  assign n51789 = ~n51780 & n51788 ;
  assign n51790 = ~\u0_L13_reg[20]/NET0131  & ~n51789 ;
  assign n51791 = \u0_L13_reg[20]/NET0131  & n51789 ;
  assign n51792 = ~n51790 & ~n51791 ;
  assign n51850 = decrypt_pad & ~\u0_uk_K_r13_reg[42]/NET0131  ;
  assign n51851 = ~decrypt_pad & ~\u0_uk_K_r13_reg[21]/NET0131  ;
  assign n51852 = ~n51850 & ~n51851 ;
  assign n51853 = \u0_R13_reg[24]/NET0131  & ~n51852 ;
  assign n51854 = ~\u0_R13_reg[24]/NET0131  & n51852 ;
  assign n51855 = ~n51853 & ~n51854 ;
  assign n51819 = decrypt_pad & ~\u0_uk_K_r13_reg[31]/NET0131  ;
  assign n51820 = ~decrypt_pad & ~\u0_uk_K_r13_reg[37]/NET0131  ;
  assign n51821 = ~n51819 & ~n51820 ;
  assign n51822 = \u0_R13_reg[22]/P0001  & ~n51821 ;
  assign n51823 = ~\u0_R13_reg[22]/P0001  & n51821 ;
  assign n51824 = ~n51822 & ~n51823 ;
  assign n51793 = decrypt_pad & ~\u0_uk_K_r13_reg[36]/NET0131  ;
  assign n51794 = ~decrypt_pad & ~\u0_uk_K_r13_reg[15]/NET0131  ;
  assign n51795 = ~n51793 & ~n51794 ;
  assign n51796 = \u0_R13_reg[21]/NET0131  & ~n51795 ;
  assign n51797 = ~\u0_R13_reg[21]/NET0131  & n51795 ;
  assign n51798 = ~n51796 & ~n51797 ;
  assign n51806 = decrypt_pad & ~\u0_uk_K_r13_reg[21]/NET0131  ;
  assign n51807 = ~decrypt_pad & ~\u0_uk_K_r13_reg[0]/NET0131  ;
  assign n51808 = ~n51806 & ~n51807 ;
  assign n51809 = \u0_R13_reg[20]/NET0131  & ~n51808 ;
  assign n51810 = ~\u0_R13_reg[20]/NET0131  & n51808 ;
  assign n51811 = ~n51809 & ~n51810 ;
  assign n51835 = n51798 & ~n51811 ;
  assign n51799 = decrypt_pad & ~\u0_uk_K_r13_reg[37]/NET0131  ;
  assign n51800 = ~decrypt_pad & ~\u0_uk_K_r13_reg[16]/NET0131  ;
  assign n51801 = ~n51799 & ~n51800 ;
  assign n51802 = \u0_R13_reg[25]/NET0131  & ~n51801 ;
  assign n51803 = ~\u0_R13_reg[25]/NET0131  & n51801 ;
  assign n51804 = ~n51802 & ~n51803 ;
  assign n51863 = n51804 & n51811 ;
  assign n51877 = ~n51835 & ~n51863 ;
  assign n51878 = n51824 & ~n51877 ;
  assign n51813 = decrypt_pad & ~\u0_uk_K_r13_reg[16]/NET0131  ;
  assign n51814 = ~decrypt_pad & ~\u0_uk_K_r13_reg[50]/NET0131  ;
  assign n51815 = ~n51813 & ~n51814 ;
  assign n51816 = \u0_R13_reg[23]/NET0131  & ~n51815 ;
  assign n51817 = ~\u0_R13_reg[23]/NET0131  & n51815 ;
  assign n51818 = ~n51816 & ~n51817 ;
  assign n51874 = n51798 & n51804 ;
  assign n51875 = ~n51811 & n51874 ;
  assign n51876 = ~n51824 & ~n51875 ;
  assign n51879 = ~n51818 & ~n51876 ;
  assign n51880 = ~n51878 & n51879 ;
  assign n51840 = ~n51798 & n51811 ;
  assign n51867 = ~n51804 & n51840 ;
  assign n51868 = ~n51824 & n51867 ;
  assign n51836 = n51824 & n51835 ;
  assign n51866 = n51798 & n51863 ;
  assign n51869 = ~n51836 & ~n51866 ;
  assign n51870 = ~n51868 & n51869 ;
  assign n51871 = n51818 & ~n51870 ;
  assign n51844 = ~n51818 & ~n51824 ;
  assign n51872 = n51844 & n51863 ;
  assign n51873 = ~n51798 & n51872 ;
  assign n51881 = ~n51871 & ~n51873 ;
  assign n51882 = ~n51880 & n51881 ;
  assign n51883 = n51855 & ~n51882 ;
  assign n51805 = n51798 & ~n51804 ;
  assign n51812 = ~n51805 & n51811 ;
  assign n51825 = n51818 & ~n51824 ;
  assign n51826 = n51805 & ~n51824 ;
  assign n51827 = n51811 & n51826 ;
  assign n51828 = ~n51825 & ~n51827 ;
  assign n51829 = ~n51812 & ~n51828 ;
  assign n51830 = n51811 & ~n51824 ;
  assign n51837 = n51798 & n51830 ;
  assign n51838 = ~n51836 & ~n51837 ;
  assign n51839 = ~n51818 & ~n51838 ;
  assign n51831 = n51818 & ~n51830 ;
  assign n51832 = ~n51804 & ~n51811 ;
  assign n51833 = ~n51798 & ~n51832 ;
  assign n51834 = n51831 & n51833 ;
  assign n51841 = n51804 & n51824 ;
  assign n51842 = n51840 & n51841 ;
  assign n51843 = ~n51804 & n51811 ;
  assign n51845 = n51843 & n51844 ;
  assign n51846 = ~n51842 & ~n51845 ;
  assign n51847 = ~n51834 & n51846 ;
  assign n51848 = ~n51839 & n51847 ;
  assign n51849 = ~n51829 & n51848 ;
  assign n51856 = ~n51849 & ~n51855 ;
  assign n51859 = n51804 & ~n51811 ;
  assign n51860 = ~n51798 & n51859 ;
  assign n51861 = n51818 & ~n51860 ;
  assign n51862 = ~n51828 & ~n51861 ;
  assign n51857 = ~n51798 & n51832 ;
  assign n51858 = n51844 & n51857 ;
  assign n51864 = ~n51826 & ~n51863 ;
  assign n51865 = n51831 & ~n51864 ;
  assign n51884 = ~n51858 & ~n51865 ;
  assign n51885 = ~n51862 & n51884 ;
  assign n51886 = ~n51856 & n51885 ;
  assign n51887 = ~n51883 & n51886 ;
  assign n51888 = ~\u0_L13_reg[11]/NET0131  & n51887 ;
  assign n51889 = \u0_L13_reg[11]/NET0131  & ~n51887 ;
  assign n51890 = ~n51888 & ~n51889 ;
  assign n51904 = ~n51544 & ~n51576 ;
  assign n51905 = n51546 & n51576 ;
  assign n51906 = ~n51904 & ~n51905 ;
  assign n51907 = n51525 & ~n51906 ;
  assign n51910 = ~n51525 & ~n51591 ;
  assign n51911 = ~n51904 & n51910 ;
  assign n51903 = n51544 & n51596 ;
  assign n51908 = n51531 & n51538 ;
  assign n51909 = n51553 & n51908 ;
  assign n51912 = ~n51903 & ~n51909 ;
  assign n51913 = ~n51911 & n51912 ;
  assign n51914 = ~n51907 & n51913 ;
  assign n51915 = n51519 & ~n51914 ;
  assign n51893 = ~n51547 & ~n51553 ;
  assign n51894 = ~n51531 & n51545 ;
  assign n51895 = ~n51893 & ~n51894 ;
  assign n51896 = ~n51525 & ~n51895 ;
  assign n51897 = ~n51557 & ~n51594 ;
  assign n51898 = n51525 & ~n51897 ;
  assign n51891 = n51531 & n51566 ;
  assign n51892 = n51544 & n51891 ;
  assign n51899 = ~n51598 & ~n51892 ;
  assign n51900 = ~n51898 & n51899 ;
  assign n51901 = ~n51896 & n51900 ;
  assign n51902 = ~n51519 & ~n51901 ;
  assign n51916 = ~n51531 & n51597 ;
  assign n51917 = ~n51580 & ~n51916 ;
  assign n51918 = n51525 & n51553 ;
  assign n51919 = ~n51917 & n51918 ;
  assign n51920 = ~n51902 & ~n51919 ;
  assign n51921 = ~n51915 & n51920 ;
  assign n51922 = ~\u0_L13_reg[17]/NET0131  & ~n51921 ;
  assign n51923 = \u0_L13_reg[17]/NET0131  & n51921 ;
  assign n51924 = ~n51922 & ~n51923 ;
  assign n51941 = n51715 & ~n51723 ;
  assign n51942 = n51729 & ~n51941 ;
  assign n51943 = ~n51765 & ~n51942 ;
  assign n51944 = ~n51738 & ~n51943 ;
  assign n51938 = ~n51717 & ~n51751 ;
  assign n51939 = n51738 & ~n51938 ;
  assign n51940 = ~n51741 & n51772 ;
  assign n51945 = ~n51939 & ~n51940 ;
  assign n51946 = ~n51944 & n51945 ;
  assign n51947 = n51757 & ~n51946 ;
  assign n51929 = n51709 & ~n51723 ;
  assign n51930 = n51703 & ~n51929 ;
  assign n51933 = n51781 & n51930 ;
  assign n51934 = n51728 & ~n51933 ;
  assign n51925 = ~n51740 & ~n51774 ;
  assign n51926 = ~n51723 & ~n51925 ;
  assign n51927 = ~n51709 & ~n51715 ;
  assign n51928 = ~n51703 & ~n51927 ;
  assign n51931 = ~n51738 & ~n51928 ;
  assign n51932 = ~n51930 & n51931 ;
  assign n51935 = ~n51926 & ~n51932 ;
  assign n51936 = n51934 & n51935 ;
  assign n51937 = ~n51757 & ~n51936 ;
  assign n51948 = ~n51727 & ~n51940 ;
  assign n51949 = ~n51738 & ~n51948 ;
  assign n51950 = ~n51748 & ~n51786 ;
  assign n51951 = ~n51949 & n51950 ;
  assign n51952 = ~n51937 & n51951 ;
  assign n51953 = ~n51947 & n51952 ;
  assign n51954 = ~\u0_L13_reg[10]/NET0131  & ~n51953 ;
  assign n51955 = \u0_L13_reg[10]/NET0131  & n51953 ;
  assign n51956 = ~n51954 & ~n51955 ;
  assign n51958 = ~n51619 & n51668 ;
  assign n51959 = ~n51632 & ~n51645 ;
  assign n51960 = ~n51958 & n51959 ;
  assign n51961 = n51652 & ~n51960 ;
  assign n51957 = n51641 & n51654 ;
  assign n51962 = ~n51613 & ~n51957 ;
  assign n51963 = ~n51961 & n51962 ;
  assign n51968 = n51619 & ~n51652 ;
  assign n51969 = n51658 & n51968 ;
  assign n51964 = ~n51619 & n51632 ;
  assign n51970 = n51613 & ~n51964 ;
  assign n51971 = ~n51969 & n51970 ;
  assign n51966 = ~n51625 & n51641 ;
  assign n51967 = n51652 & n51966 ;
  assign n51965 = n51638 & n51675 ;
  assign n51972 = ~n51684 & ~n51965 ;
  assign n51973 = ~n51967 & n51972 ;
  assign n51974 = n51971 & n51973 ;
  assign n51975 = ~n51963 & ~n51974 ;
  assign n51976 = ~n51619 & n51631 ;
  assign n51977 = n51644 & n51976 ;
  assign n51978 = n51676 & ~n51977 ;
  assign n51979 = n51686 & n51978 ;
  assign n51980 = n51638 & n51673 ;
  assign n51981 = n51652 & ~n51680 ;
  assign n51982 = ~n51980 & n51981 ;
  assign n51983 = ~n51979 & ~n51982 ;
  assign n51984 = ~n51613 & ~n51652 ;
  assign n51985 = n51674 & n51984 ;
  assign n51986 = ~n51983 & ~n51985 ;
  assign n51987 = ~n51975 & n51986 ;
  assign n51988 = \u0_L13_reg[15]/P0001  & n51987 ;
  assign n51989 = ~\u0_L13_reg[15]/P0001  & ~n51987 ;
  assign n51990 = ~n51988 & ~n51989 ;
  assign n52015 = n51619 & n51632 ;
  assign n52013 = n51638 & n51672 ;
  assign n52014 = n51631 & n51644 ;
  assign n52016 = ~n52013 & ~n52014 ;
  assign n52017 = ~n52015 & n52016 ;
  assign n52018 = n51652 & ~n52017 ;
  assign n52009 = ~n51656 & ~n51965 ;
  assign n52010 = ~n51652 & ~n52009 ;
  assign n51994 = n51625 & n51668 ;
  assign n52011 = ~n51966 & ~n51994 ;
  assign n52012 = n51619 & ~n52011 ;
  assign n52019 = ~n51980 & ~n52012 ;
  assign n52020 = ~n52010 & n52019 ;
  assign n52021 = ~n52018 & n52020 ;
  assign n52022 = n51613 & ~n52021 ;
  assign n51992 = ~n51625 & ~n51652 ;
  assign n51993 = n51668 & n51992 ;
  assign n52000 = ~n51679 & ~n51993 ;
  assign n52001 = ~n51643 & n52000 ;
  assign n51991 = n51638 & n51655 ;
  assign n52002 = ~n51685 & ~n51991 ;
  assign n52003 = n52001 & n52002 ;
  assign n51995 = ~n51675 & ~n51994 ;
  assign n51996 = n51652 & ~n51995 ;
  assign n51997 = ~n51625 & n51968 ;
  assign n51998 = ~n51964 & ~n51997 ;
  assign n51999 = n51638 & ~n51998 ;
  assign n52004 = ~n51996 & ~n51999 ;
  assign n52005 = n52003 & n52004 ;
  assign n52006 = ~n51613 & ~n52005 ;
  assign n52007 = n51652 & n51673 ;
  assign n52008 = n51631 & n51991 ;
  assign n52023 = ~n52007 & ~n52008 ;
  assign n52024 = ~n52006 & n52023 ;
  assign n52025 = ~n52022 & n52024 ;
  assign n52026 = ~\u0_L13_reg[21]/NET0131  & ~n52025 ;
  assign n52027 = \u0_L13_reg[21]/NET0131  & n52025 ;
  assign n52028 = ~n52026 & ~n52027 ;
  assign n52029 = n51448 & ~n51458 ;
  assign n52030 = ~n51488 & ~n52029 ;
  assign n52031 = n51441 & ~n52030 ;
  assign n52036 = ~n51463 & ~n51472 ;
  assign n52034 = ~n51435 & ~n51487 ;
  assign n52035 = ~n51458 & ~n52034 ;
  assign n52032 = n51428 & n51458 ;
  assign n52033 = n51460 & n52032 ;
  assign n52037 = ~n51470 & ~n52033 ;
  assign n52038 = ~n52035 & n52037 ;
  assign n52039 = ~n52036 & n52038 ;
  assign n52040 = ~n52031 & n52039 ;
  assign n52042 = ~n51434 & ~n51462 ;
  assign n52043 = n51458 & ~n52042 ;
  assign n52044 = n51472 & ~n52043 ;
  assign n52045 = ~n52036 & ~n52044 ;
  assign n52041 = ~n51458 & n51504 ;
  assign n52046 = n51470 & ~n52041 ;
  assign n52047 = ~n52045 & n52046 ;
  assign n52048 = ~n52040 & ~n52047 ;
  assign n52049 = \u0_L13_reg[12]/NET0131  & n52048 ;
  assign n52050 = ~\u0_L13_reg[12]/NET0131  & ~n52048 ;
  assign n52051 = ~n52049 & ~n52050 ;
  assign n52052 = decrypt_pad & ~\u0_uk_K_r13_reg[30]/NET0131  ;
  assign n52053 = ~decrypt_pad & ~\u0_uk_K_r13_reg[9]/NET0131  ;
  assign n52054 = ~n52052 & ~n52053 ;
  assign n52055 = \u0_R13_reg[20]/NET0131  & ~n52054 ;
  assign n52056 = ~\u0_R13_reg[20]/NET0131  & n52054 ;
  assign n52057 = ~n52055 & ~n52056 ;
  assign n52087 = decrypt_pad & ~\u0_uk_K_r13_reg[15]/NET0131  ;
  assign n52088 = ~decrypt_pad & ~\u0_uk_K_r13_reg[49]/NET0131  ;
  assign n52089 = ~n52087 & ~n52088 ;
  assign n52090 = \u0_R13_reg[19]/NET0131  & ~n52089 ;
  assign n52091 = ~\u0_R13_reg[19]/NET0131  & n52089 ;
  assign n52092 = ~n52090 & ~n52091 ;
  assign n52071 = decrypt_pad & ~\u0_uk_K_r13_reg[0]/NET0131  ;
  assign n52072 = ~decrypt_pad & ~\u0_uk_K_r13_reg[38]/NET0131  ;
  assign n52073 = ~n52071 & ~n52072 ;
  assign n52074 = \u0_R13_reg[21]/NET0131  & ~n52073 ;
  assign n52075 = ~\u0_R13_reg[21]/NET0131  & n52073 ;
  assign n52076 = ~n52074 & ~n52075 ;
  assign n52064 = decrypt_pad & ~\u0_uk_K_r13_reg[43]/NET0131  ;
  assign n52065 = ~decrypt_pad & ~\u0_uk_K_r13_reg[22]/NET0131  ;
  assign n52066 = ~n52064 & ~n52065 ;
  assign n52067 = \u0_R13_reg[16]/NET0131  & ~n52066 ;
  assign n52068 = ~\u0_R13_reg[16]/NET0131  & n52066 ;
  assign n52069 = ~n52067 & ~n52068 ;
  assign n52079 = decrypt_pad & ~\u0_uk_K_r13_reg[28]/NET0131  ;
  assign n52080 = ~decrypt_pad & ~\u0_uk_K_r13_reg[7]/NET0131  ;
  assign n52081 = ~n52079 & ~n52080 ;
  assign n52082 = \u0_R13_reg[18]/NET0131  & ~n52081 ;
  assign n52083 = ~\u0_R13_reg[18]/NET0131  & n52081 ;
  assign n52084 = ~n52082 & ~n52083 ;
  assign n52094 = n52069 & n52084 ;
  assign n52095 = ~n52076 & ~n52094 ;
  assign n52058 = decrypt_pad & ~\u0_uk_K_r13_reg[38]/NET0131  ;
  assign n52059 = ~decrypt_pad & ~\u0_uk_K_r13_reg[44]/NET0131  ;
  assign n52060 = ~n52058 & ~n52059 ;
  assign n52061 = \u0_R13_reg[17]/NET0131  & ~n52060 ;
  assign n52062 = ~\u0_R13_reg[17]/NET0131  & n52060 ;
  assign n52063 = ~n52061 & ~n52062 ;
  assign n52101 = n52063 & ~n52084 ;
  assign n52102 = n52095 & ~n52101 ;
  assign n52099 = n52063 & n52069 ;
  assign n52100 = n52076 & n52099 ;
  assign n52103 = ~n52063 & ~n52069 ;
  assign n52104 = ~n52100 & ~n52103 ;
  assign n52105 = ~n52102 & n52104 ;
  assign n52106 = n52092 & ~n52105 ;
  assign n52070 = ~n52063 & n52069 ;
  assign n52077 = n52070 & n52076 ;
  assign n52078 = n52063 & ~n52069 ;
  assign n52085 = n52078 & ~n52084 ;
  assign n52086 = ~n52077 & ~n52085 ;
  assign n52093 = ~n52086 & ~n52092 ;
  assign n52096 = n52076 & n52084 ;
  assign n52097 = n52063 & ~n52096 ;
  assign n52098 = ~n52095 & n52097 ;
  assign n52107 = ~n52093 & ~n52098 ;
  assign n52108 = ~n52106 & n52107 ;
  assign n52109 = n52057 & ~n52108 ;
  assign n52125 = ~n52076 & n52103 ;
  assign n52126 = ~n52076 & n52099 ;
  assign n52127 = ~n52125 & ~n52126 ;
  assign n52128 = n52084 & ~n52127 ;
  assign n52129 = n52076 & n52103 ;
  assign n52130 = ~n52084 & n52129 ;
  assign n52131 = ~n52128 & ~n52130 ;
  assign n52132 = n52092 & ~n52131 ;
  assign n52113 = ~n52076 & n52092 ;
  assign n52114 = n52070 & ~n52076 ;
  assign n52115 = n52078 & n52084 ;
  assign n52116 = ~n52114 & ~n52115 ;
  assign n52117 = ~n52113 & ~n52116 ;
  assign n52119 = n52063 & ~n52076 ;
  assign n52120 = n52092 & ~n52119 ;
  assign n52118 = ~n52092 & ~n52103 ;
  assign n52121 = ~n52084 & ~n52118 ;
  assign n52122 = ~n52120 & n52121 ;
  assign n52123 = ~n52117 & ~n52122 ;
  assign n52124 = ~n52057 & ~n52123 ;
  assign n52110 = ~n52063 & n52084 ;
  assign n52111 = n52069 & ~n52092 ;
  assign n52112 = n52110 & n52111 ;
  assign n52133 = n52076 & ~n52084 ;
  assign n52134 = n52099 & n52133 ;
  assign n52135 = ~n52112 & ~n52134 ;
  assign n52136 = ~n52124 & n52135 ;
  assign n52137 = ~n52132 & n52136 ;
  assign n52138 = ~n52109 & n52137 ;
  assign n52139 = ~\u0_L13_reg[25]/NET0131  & ~n52138 ;
  assign n52140 = \u0_L13_reg[25]/NET0131  & n52138 ;
  assign n52141 = ~n52139 & ~n52140 ;
  assign n52146 = n51723 & n51725 ;
  assign n52147 = ~n51927 & ~n52146 ;
  assign n52148 = ~n51757 & ~n52147 ;
  assign n52142 = ~n51709 & ~n51741 ;
  assign n52143 = n51709 & ~n51740 ;
  assign n52144 = ~n51723 & ~n52143 ;
  assign n52145 = ~n52142 & n52144 ;
  assign n52149 = ~n51738 & ~n52145 ;
  assign n52150 = ~n52148 & n52149 ;
  assign n52151 = n51738 & ~n51751 ;
  assign n52152 = ~n51765 & n52151 ;
  assign n52153 = ~n52150 & ~n52152 ;
  assign n52154 = n51715 & ~n51783 ;
  assign n52157 = n51738 & n51768 ;
  assign n52163 = n51757 & ~n52157 ;
  assign n52164 = ~n52154 & n52163 ;
  assign n52155 = ~n51764 & ~n51774 ;
  assign n52156 = n51723 & ~n52155 ;
  assign n52158 = n51703 & n51709 ;
  assign n52159 = ~n51715 & n51929 ;
  assign n52160 = ~n52158 & ~n52159 ;
  assign n52161 = ~n51738 & ~n51749 ;
  assign n52162 = ~n52160 & n52161 ;
  assign n52165 = ~n52156 & ~n52162 ;
  assign n52166 = n52164 & n52165 ;
  assign n52167 = ~n51742 & n51747 ;
  assign n52168 = ~n51750 & ~n51757 ;
  assign n52169 = ~n52167 & n52168 ;
  assign n52170 = n51766 & n52169 ;
  assign n52171 = ~n52166 & ~n52170 ;
  assign n52172 = ~n52153 & ~n52171 ;
  assign n52173 = \u0_L13_reg[26]/NET0131  & n52172 ;
  assign n52174 = ~\u0_L13_reg[26]/NET0131  & ~n52172 ;
  assign n52175 = ~n52173 & ~n52174 ;
  assign n52176 = decrypt_pad & ~\u0_uk_K_r13_reg[46]/NET0131  ;
  assign n52177 = ~decrypt_pad & ~\u0_uk_K_r13_reg[25]/P0001  ;
  assign n52178 = ~n52176 & ~n52177 ;
  assign n52179 = \u0_R13_reg[8]/NET0131  & ~n52178 ;
  assign n52180 = ~\u0_R13_reg[8]/NET0131  & n52178 ;
  assign n52181 = ~n52179 & ~n52180 ;
  assign n52218 = decrypt_pad & ~\u0_uk_K_r13_reg[55]/NET0131  ;
  assign n52219 = ~decrypt_pad & ~\u0_uk_K_r13_reg[34]/NET0131  ;
  assign n52220 = ~n52218 & ~n52219 ;
  assign n52221 = \u0_R13_reg[7]/NET0131  & ~n52220 ;
  assign n52222 = ~\u0_R13_reg[7]/NET0131  & n52220 ;
  assign n52223 = ~n52221 & ~n52222 ;
  assign n52207 = decrypt_pad & ~\u0_uk_K_r13_reg[4]/NET0131  ;
  assign n52208 = ~decrypt_pad & ~\u0_uk_K_r13_reg[40]/NET0131  ;
  assign n52209 = ~n52207 & ~n52208 ;
  assign n52210 = \u0_R13_reg[6]/NET0131  & ~n52209 ;
  assign n52211 = ~\u0_R13_reg[6]/NET0131  & n52209 ;
  assign n52212 = ~n52210 & ~n52211 ;
  assign n52188 = decrypt_pad & ~\u0_uk_K_r13_reg[13]/NET0131  ;
  assign n52189 = ~decrypt_pad & ~\u0_uk_K_r13_reg[17]/NET0131  ;
  assign n52190 = ~n52188 & ~n52189 ;
  assign n52191 = \u0_R13_reg[5]/NET0131  & ~n52190 ;
  assign n52192 = ~\u0_R13_reg[5]/NET0131  & n52190 ;
  assign n52193 = ~n52191 & ~n52192 ;
  assign n52182 = decrypt_pad & ~\u0_uk_K_r13_reg[34]/NET0131  ;
  assign n52183 = ~decrypt_pad & ~\u0_uk_K_r13_reg[13]/NET0131  ;
  assign n52184 = ~n52182 & ~n52183 ;
  assign n52185 = \u0_R13_reg[4]/NET0131  & ~n52184 ;
  assign n52186 = ~\u0_R13_reg[4]/NET0131  & n52184 ;
  assign n52187 = ~n52185 & ~n52186 ;
  assign n52195 = decrypt_pad & ~\u0_uk_K_r13_reg[26]/NET0131  ;
  assign n52196 = ~decrypt_pad & ~\u0_uk_K_r13_reg[5]/NET0131  ;
  assign n52197 = ~n52195 & ~n52196 ;
  assign n52198 = \u0_R13_reg[9]/NET0131  & ~n52197 ;
  assign n52199 = ~\u0_R13_reg[9]/NET0131  & n52197 ;
  assign n52200 = ~n52198 & ~n52199 ;
  assign n52225 = ~n52187 & ~n52200 ;
  assign n52245 = n52193 & n52225 ;
  assign n52246 = n52212 & n52245 ;
  assign n52239 = n52187 & n52200 ;
  assign n52244 = n52193 & n52239 ;
  assign n52247 = ~n52193 & ~n52200 ;
  assign n52248 = n52187 & n52247 ;
  assign n52249 = ~n52244 & ~n52248 ;
  assign n52250 = ~n52246 & n52249 ;
  assign n52251 = n52223 & ~n52250 ;
  assign n52240 = ~n52193 & n52239 ;
  assign n52241 = ~n52223 & ~n52240 ;
  assign n52242 = n52187 & ~n52212 ;
  assign n52243 = ~n52241 & n52242 ;
  assign n52226 = ~n52212 & n52225 ;
  assign n52203 = ~n52187 & n52200 ;
  assign n52227 = n52193 & n52203 ;
  assign n52228 = ~n52226 & ~n52227 ;
  assign n52238 = ~n52223 & ~n52228 ;
  assign n52234 = ~n52193 & n52212 ;
  assign n52252 = n52203 & n52234 ;
  assign n52253 = ~n52238 & ~n52252 ;
  assign n52254 = ~n52243 & n52253 ;
  assign n52255 = ~n52251 & n52254 ;
  assign n52256 = n52181 & ~n52255 ;
  assign n52214 = ~n52193 & n52203 ;
  assign n52194 = n52187 & n52193 ;
  assign n52202 = n52187 & ~n52200 ;
  assign n52215 = n52202 & ~n52212 ;
  assign n52216 = ~n52194 & ~n52215 ;
  assign n52217 = ~n52214 & n52216 ;
  assign n52224 = ~n52217 & ~n52223 ;
  assign n52201 = n52194 & ~n52200 ;
  assign n52204 = ~n52193 & ~n52202 ;
  assign n52205 = ~n52203 & n52204 ;
  assign n52206 = ~n52201 & ~n52205 ;
  assign n52213 = ~n52206 & n52212 ;
  assign n52229 = n52223 & ~n52228 ;
  assign n52230 = ~n52213 & ~n52229 ;
  assign n52231 = ~n52224 & n52230 ;
  assign n52232 = ~n52181 & ~n52231 ;
  assign n52233 = n52201 & n52212 ;
  assign n52235 = ~n52187 & n52234 ;
  assign n52236 = ~n52233 & ~n52235 ;
  assign n52237 = ~n52223 & ~n52236 ;
  assign n52257 = ~n52232 & ~n52237 ;
  assign n52258 = ~n52256 & n52257 ;
  assign n52259 = ~\u0_L13_reg[28]/NET0131  & ~n52258 ;
  assign n52260 = \u0_L13_reg[28]/NET0131  & n52258 ;
  assign n52261 = ~n52259 & ~n52260 ;
  assign n52286 = n51824 & ~n51843 ;
  assign n52287 = ~n51859 & n52286 ;
  assign n52288 = ~n51857 & ~n52287 ;
  assign n52289 = ~n51818 & ~n52288 ;
  assign n52268 = n51798 & n51843 ;
  assign n52269 = n51824 & n52268 ;
  assign n52279 = ~n51804 & n51824 ;
  assign n52283 = n51835 & ~n52279 ;
  assign n52284 = ~n52269 & ~n52283 ;
  assign n52285 = n51818 & ~n52284 ;
  assign n52278 = ~n51824 & n51859 ;
  assign n52280 = ~n51811 & n52279 ;
  assign n52281 = ~n52278 & ~n52280 ;
  assign n52282 = ~n51798 & ~n52281 ;
  assign n52290 = n51846 & ~n52282 ;
  assign n52291 = ~n52285 & n52290 ;
  assign n52292 = ~n52289 & n52291 ;
  assign n52293 = n51855 & ~n52292 ;
  assign n52262 = ~n51866 & ~n51867 ;
  assign n52263 = ~n51798 & ~n51824 ;
  assign n52264 = ~n51836 & ~n52263 ;
  assign n52265 = ~n51804 & ~n52264 ;
  assign n52266 = n52262 & ~n52265 ;
  assign n52267 = n51818 & ~n52266 ;
  assign n52270 = ~n51824 & ~n51877 ;
  assign n52271 = ~n52269 & ~n52270 ;
  assign n52272 = ~n51818 & ~n52271 ;
  assign n52273 = n51824 & n51860 ;
  assign n52274 = ~n52272 & ~n52273 ;
  assign n52275 = ~n52267 & n52274 ;
  assign n52276 = ~n51855 & ~n52275 ;
  assign n52277 = n51825 & n51874 ;
  assign n52294 = ~n51868 & ~n52277 ;
  assign n52295 = ~n52276 & n52294 ;
  assign n52296 = ~n52293 & n52295 ;
  assign n52297 = \u0_L13_reg[29]/NET0131  & ~n52296 ;
  assign n52298 = ~\u0_L13_reg[29]/NET0131  & n52296 ;
  assign n52299 = ~n52297 & ~n52298 ;
  assign n52303 = ~n52194 & ~n52202 ;
  assign n52304 = n52212 & ~n52303 ;
  assign n52305 = ~n52214 & ~n52304 ;
  assign n52306 = ~n52223 & ~n52305 ;
  assign n52313 = n52193 & ~n52200 ;
  assign n52314 = ~n52214 & ~n52313 ;
  assign n52315 = ~n52212 & ~n52314 ;
  assign n52300 = n52212 & n52239 ;
  assign n52301 = ~n52193 & n52300 ;
  assign n52302 = n52223 & n52301 ;
  assign n52307 = ~n52193 & ~n52223 ;
  assign n52308 = n52200 & ~n52212 ;
  assign n52309 = n52307 & n52308 ;
  assign n52310 = n52203 & n52212 ;
  assign n52311 = n52193 & n52310 ;
  assign n52312 = ~n52309 & ~n52311 ;
  assign n52316 = ~n52302 & n52312 ;
  assign n52317 = ~n52315 & n52316 ;
  assign n52318 = ~n52306 & n52317 ;
  assign n52319 = ~n52181 & ~n52318 ;
  assign n52320 = n52193 & ~n52212 ;
  assign n52321 = ~n52234 & ~n52320 ;
  assign n52322 = n52239 & ~n52321 ;
  assign n52323 = ~n52215 & ~n52225 ;
  assign n52324 = ~n52320 & ~n52323 ;
  assign n52325 = ~n52322 & ~n52324 ;
  assign n52326 = n52181 & ~n52325 ;
  assign n52327 = n52203 & n52321 ;
  assign n52328 = ~n52223 & ~n52327 ;
  assign n52329 = ~n52326 & n52328 ;
  assign n52331 = n52216 & ~n52320 ;
  assign n52332 = n52181 & ~n52331 ;
  assign n52330 = ~n52200 & n52235 ;
  assign n52333 = n52194 & ~n52212 ;
  assign n52334 = n52223 & ~n52333 ;
  assign n52335 = ~n52330 & n52334 ;
  assign n52336 = ~n52332 & n52335 ;
  assign n52337 = ~n52329 & ~n52336 ;
  assign n52338 = ~n52319 & ~n52337 ;
  assign n52339 = \u0_L13_reg[2]/NET0131  & n52338 ;
  assign n52340 = ~\u0_L13_reg[2]/NET0131  & ~n52338 ;
  assign n52341 = ~n52339 & ~n52340 ;
  assign n52364 = ~n52084 & n52114 ;
  assign n52363 = n52084 & n52119 ;
  assign n52365 = ~n52129 & ~n52134 ;
  assign n52366 = ~n52363 & n52365 ;
  assign n52367 = ~n52364 & n52366 ;
  assign n52368 = ~n52092 & ~n52367 ;
  assign n52360 = ~n52086 & ~n52133 ;
  assign n52346 = n52076 & n52094 ;
  assign n52347 = ~n52085 & ~n52346 ;
  assign n52361 = ~n52125 & n52347 ;
  assign n52362 = n52092 & ~n52361 ;
  assign n52369 = ~n52360 & ~n52362 ;
  assign n52370 = ~n52368 & n52369 ;
  assign n52371 = ~n52057 & ~n52370 ;
  assign n52350 = n52076 & n52078 ;
  assign n52351 = ~n52125 & ~n52350 ;
  assign n52352 = ~n52092 & ~n52351 ;
  assign n52353 = ~n52077 & ~n52126 ;
  assign n52354 = ~n52352 & n52353 ;
  assign n52355 = ~n52084 & ~n52354 ;
  assign n52345 = ~n52076 & ~n52099 ;
  assign n52348 = n52092 & ~n52345 ;
  assign n52349 = n52347 & n52348 ;
  assign n52342 = n52084 & ~n52092 ;
  assign n52343 = n52100 & n52342 ;
  assign n52344 = n52084 & n52114 ;
  assign n52356 = ~n52343 & ~n52344 ;
  assign n52357 = ~n52349 & n52356 ;
  assign n52358 = ~n52355 & n52357 ;
  assign n52359 = n52057 & ~n52358 ;
  assign n52372 = ~n52099 & ~n52110 ;
  assign n52373 = n52095 & ~n52372 ;
  assign n52374 = n52092 & ~n52373 ;
  assign n52375 = n52084 & n52129 ;
  assign n52376 = ~n52069 & n52363 ;
  assign n52377 = ~n52375 & ~n52376 ;
  assign n52378 = ~n52092 & n52377 ;
  assign n52379 = ~n52374 & ~n52378 ;
  assign n52380 = ~n52359 & ~n52379 ;
  assign n52381 = ~n52371 & n52380 ;
  assign n52382 = ~\u0_L13_reg[14]/NET0131  & ~n52381 ;
  assign n52383 = \u0_L13_reg[14]/NET0131  & n52381 ;
  assign n52384 = ~n52382 & ~n52383 ;
  assign n52389 = ~n51826 & ~n51844 ;
  assign n52390 = ~n51811 & ~n52389 ;
  assign n52386 = ~n51804 & n51844 ;
  assign n52387 = ~n51841 & ~n52386 ;
  assign n52388 = n51798 & ~n52387 ;
  assign n52385 = n51825 & n51863 ;
  assign n52391 = n51855 & ~n52385 ;
  assign n52392 = ~n52388 & n52391 ;
  assign n52393 = ~n52390 & n52392 ;
  assign n52394 = n51818 & ~n52268 ;
  assign n52395 = ~n51842 & ~n52278 ;
  assign n52396 = n52394 & n52395 ;
  assign n52397 = n51798 & n51832 ;
  assign n52398 = ~n51818 & ~n52397 ;
  assign n52399 = ~n52273 & n52398 ;
  assign n52400 = ~n52396 & ~n52399 ;
  assign n52401 = ~n51855 & ~n51872 ;
  assign n52402 = ~n51868 & n52401 ;
  assign n52403 = ~n52400 & n52402 ;
  assign n52404 = ~n52393 & ~n52403 ;
  assign n52407 = ~n51818 & n52262 ;
  assign n52405 = ~n51857 & ~n51875 ;
  assign n52406 = n52394 & n52405 ;
  assign n52408 = n51824 & ~n52406 ;
  assign n52409 = ~n52407 & n52408 ;
  assign n52410 = n51832 & n51844 ;
  assign n52411 = ~n52409 & ~n52410 ;
  assign n52412 = ~n52404 & n52411 ;
  assign n52413 = ~\u0_L13_reg[4]/NET0131  & ~n52412 ;
  assign n52414 = \u0_L13_reg[4]/NET0131  & n52412 ;
  assign n52415 = ~n52413 & ~n52414 ;
  assign n52420 = n51715 & ~n51782 ;
  assign n52421 = n51738 & ~n51783 ;
  assign n52422 = ~n52420 & n52421 ;
  assign n52417 = ~n51726 & ~n51731 ;
  assign n52418 = n51703 & ~n51738 ;
  assign n52419 = ~n52417 & n52418 ;
  assign n52416 = ~n51743 & n51941 ;
  assign n52423 = ~n51773 & ~n52416 ;
  assign n52424 = ~n52419 & n52423 ;
  assign n52425 = ~n52422 & n52424 ;
  assign n52426 = ~n51757 & ~n52425 ;
  assign n52437 = n51715 & n51730 ;
  assign n52435 = ~n51709 & ~n51749 ;
  assign n52436 = n51781 & ~n52435 ;
  assign n52438 = ~n52146 & ~n52436 ;
  assign n52439 = ~n52437 & n52438 ;
  assign n52440 = n51757 & ~n52439 ;
  assign n52427 = ~n51724 & ~n51940 ;
  assign n52428 = n51738 & ~n52427 ;
  assign n52429 = n51723 & n52142 ;
  assign n52430 = ~n51729 & n51941 ;
  assign n52431 = ~n51764 & ~n52430 ;
  assign n52432 = n51757 & ~n52431 ;
  assign n52433 = ~n52429 & ~n52432 ;
  assign n52434 = ~n51738 & ~n52433 ;
  assign n52441 = ~n52428 & ~n52434 ;
  assign n52442 = ~n52440 & n52441 ;
  assign n52443 = ~n52426 & n52442 ;
  assign n52444 = ~\u0_L13_reg[1]/NET0131  & ~n52443 ;
  assign n52445 = \u0_L13_reg[1]/NET0131  & n52443 ;
  assign n52446 = ~n52444 & ~n52445 ;
  assign n52447 = n52194 & n52308 ;
  assign n52448 = ~n52233 & ~n52447 ;
  assign n52449 = ~n52212 & n52247 ;
  assign n52450 = n52187 & n52449 ;
  assign n52451 = ~n52245 & ~n52252 ;
  assign n52452 = ~n52450 & n52451 ;
  assign n52453 = ~n52181 & ~n52452 ;
  assign n52454 = n52448 & ~n52453 ;
  assign n52455 = ~n52223 & ~n52454 ;
  assign n52456 = ~n52200 & n52333 ;
  assign n52457 = ~n52205 & ~n52456 ;
  assign n52458 = n52223 & ~n52457 ;
  assign n52461 = n52212 & n52223 ;
  assign n52462 = n52187 & ~n52313 ;
  assign n52463 = n52461 & n52462 ;
  assign n52459 = ~n52187 & ~n52307 ;
  assign n52460 = n52308 & n52459 ;
  assign n52464 = ~n52181 & ~n52460 ;
  assign n52465 = ~n52463 & n52464 ;
  assign n52466 = ~n52458 & n52465 ;
  assign n52467 = n52212 & n52247 ;
  assign n52468 = n52241 & ~n52467 ;
  assign n52469 = n52223 & ~n52310 ;
  assign n52470 = ~n52449 & n52469 ;
  assign n52471 = ~n52468 & ~n52470 ;
  assign n52472 = n52193 & n52226 ;
  assign n52473 = n52181 & ~n52472 ;
  assign n52474 = n52312 & n52473 ;
  assign n52475 = n52448 & n52474 ;
  assign n52476 = ~n52471 & n52475 ;
  assign n52477 = ~n52466 & ~n52476 ;
  assign n52478 = ~n52455 & ~n52477 ;
  assign n52479 = ~\u0_L13_reg[13]/NET0131  & n52478 ;
  assign n52480 = \u0_L13_reg[13]/NET0131  & ~n52478 ;
  assign n52481 = ~n52479 & ~n52480 ;
  assign n52484 = ~n51805 & ~n51811 ;
  assign n52485 = n51818 & ~n51837 ;
  assign n52486 = ~n52484 & n52485 ;
  assign n52482 = ~n51818 & ~n52405 ;
  assign n52483 = n51824 & n51866 ;
  assign n52487 = ~n51855 & ~n52483 ;
  assign n52488 = ~n52482 & n52487 ;
  assign n52489 = ~n52486 & n52488 ;
  assign n52490 = ~n51837 & ~n51860 ;
  assign n52491 = n51818 & ~n52490 ;
  assign n52494 = ~n51826 & n51855 ;
  assign n52492 = n51835 & n51841 ;
  assign n52493 = ~n51818 & n51840 ;
  assign n52495 = ~n52492 & ~n52493 ;
  assign n52496 = n52494 & n52495 ;
  assign n52497 = ~n52282 & n52496 ;
  assign n52498 = ~n52491 & n52497 ;
  assign n52499 = ~n52489 & ~n52498 ;
  assign n52500 = ~n51862 & ~n51873 ;
  assign n52501 = ~n52499 & n52500 ;
  assign n52502 = ~\u0_L13_reg[19]/NET0131  & ~n52501 ;
  assign n52503 = \u0_L13_reg[19]/NET0131  & n52501 ;
  assign n52504 = ~n52502 & ~n52503 ;
  assign n52505 = ~n51559 & ~n51567 ;
  assign n52506 = ~n51544 & ~n52505 ;
  assign n52507 = ~n51558 & ~n52506 ;
  assign n52508 = ~n51525 & ~n52507 ;
  assign n52510 = n51525 & ~n51591 ;
  assign n52511 = n51554 & n52510 ;
  assign n52509 = n51580 & n51590 ;
  assign n52512 = ~n51905 & ~n52509 ;
  assign n52513 = ~n52511 & n52512 ;
  assign n52514 = ~n52508 & n52513 ;
  assign n52515 = n51519 & ~n52514 ;
  assign n52522 = n51532 & n51597 ;
  assign n52526 = ~n51577 & ~n51909 ;
  assign n52527 = ~n52522 & n52526 ;
  assign n52523 = n51525 & n51567 ;
  assign n52524 = ~n51553 & ~n51908 ;
  assign n52525 = n51583 & ~n52524 ;
  assign n52528 = ~n52523 & ~n52525 ;
  assign n52529 = n52527 & n52528 ;
  assign n52530 = ~n51519 & ~n52529 ;
  assign n52516 = ~n51556 & ~n51567 ;
  assign n52517 = n51573 & ~n52516 ;
  assign n52518 = n51559 & n51560 ;
  assign n52519 = ~n51595 & ~n52518 ;
  assign n52520 = ~n51903 & n52519 ;
  assign n52521 = ~n51525 & ~n52520 ;
  assign n52531 = ~n52517 & ~n52521 ;
  assign n52532 = ~n52530 & n52531 ;
  assign n52533 = ~n52515 & n52532 ;
  assign n52534 = \u0_L13_reg[23]/NET0131  & ~n52533 ;
  assign n52535 = ~\u0_L13_reg[23]/NET0131  & n52533 ;
  assign n52536 = ~n52534 & ~n52535 ;
  assign n52553 = ~n51625 & n51958 ;
  assign n52554 = ~n51639 & ~n52553 ;
  assign n52555 = n51652 & ~n52554 ;
  assign n52550 = ~n51673 & ~n51994 ;
  assign n52551 = ~n52014 & n52550 ;
  assign n52552 = ~n51652 & ~n52551 ;
  assign n52556 = ~n51643 & ~n52013 ;
  assign n52557 = ~n51680 & n52556 ;
  assign n52558 = ~n52552 & n52557 ;
  assign n52559 = ~n52555 & n52558 ;
  assign n52560 = n51613 & ~n52559 ;
  assign n52538 = n51652 & ~n51679 ;
  assign n52537 = n51638 & ~n51976 ;
  assign n52539 = ~n51958 & ~n52537 ;
  assign n52540 = n52538 & n52539 ;
  assign n52541 = n51625 & n51638 ;
  assign n52542 = n51968 & n52541 ;
  assign n52543 = ~n51993 & ~n52542 ;
  assign n52544 = ~n51688 & n52543 ;
  assign n52545 = ~n52540 & n52544 ;
  assign n52546 = ~n51613 & ~n52545 ;
  assign n52547 = ~n51684 & ~n51687 ;
  assign n52548 = ~n51652 & ~n52547 ;
  assign n52549 = n51642 & n51652 ;
  assign n52561 = ~n51683 & ~n52549 ;
  assign n52562 = ~n52548 & n52561 ;
  assign n52563 = ~n52546 & n52562 ;
  assign n52564 = ~n52560 & n52563 ;
  assign n52565 = \u0_L13_reg[27]/NET0131  & n52564 ;
  assign n52566 = ~\u0_L13_reg[27]/NET0131  & ~n52564 ;
  assign n52567 = ~n52565 & ~n52566 ;
  assign n52576 = n51441 & n51490 ;
  assign n52577 = ~n51442 & ~n51488 ;
  assign n52578 = ~n52576 & n52577 ;
  assign n52579 = n51458 & ~n52578 ;
  assign n52569 = n51428 & ~n51448 ;
  assign n52570 = ~n51490 & ~n52569 ;
  assign n52572 = ~n51472 & ~n51500 ;
  assign n52573 = n52570 & ~n52572 ;
  assign n52571 = ~n51500 & ~n52570 ;
  assign n52574 = ~n51458 & ~n52571 ;
  assign n52575 = ~n52573 & n52574 ;
  assign n52568 = n51441 & n51491 ;
  assign n52580 = n51470 & ~n52568 ;
  assign n52581 = ~n52575 & n52580 ;
  assign n52582 = ~n52579 & n52581 ;
  assign n52585 = n51428 & n51450 ;
  assign n52586 = n51448 & n51462 ;
  assign n52587 = ~n52585 & ~n52586 ;
  assign n52588 = n51458 & ~n52587 ;
  assign n52583 = n51434 & n51441 ;
  assign n52584 = n52570 & n52583 ;
  assign n52592 = ~n51470 & ~n52584 ;
  assign n52593 = ~n52588 & n52592 ;
  assign n52589 = n52035 & ~n52586 ;
  assign n52590 = ~n51463 & n51472 ;
  assign n52591 = n51481 & n52590 ;
  assign n52594 = ~n52589 & ~n52591 ;
  assign n52595 = n52593 & n52594 ;
  assign n52596 = ~n52582 & ~n52595 ;
  assign n52597 = n51458 & n51504 ;
  assign n52598 = n51441 & n51471 ;
  assign n52599 = ~n51449 & ~n52598 ;
  assign n52600 = ~n51458 & ~n52599 ;
  assign n52601 = ~n52597 & ~n52600 ;
  assign n52602 = ~n52596 & n52601 ;
  assign n52603 = \u0_L13_reg[32]/NET0131  & n52602 ;
  assign n52604 = ~\u0_L13_reg[32]/NET0131  & ~n52602 ;
  assign n52605 = ~n52603 & ~n52604 ;
  assign n52612 = decrypt_pad & ~\u0_uk_K_r13_reg[3]/NET0131  ;
  assign n52613 = ~decrypt_pad & ~\u0_uk_K_r13_reg[39]/NET0131  ;
  assign n52614 = ~n52612 & ~n52613 ;
  assign n52615 = \u0_R13_reg[8]/NET0131  & ~n52614 ;
  assign n52616 = ~\u0_R13_reg[8]/NET0131  & n52614 ;
  assign n52617 = ~n52615 & ~n52616 ;
  assign n52619 = decrypt_pad & ~\u0_uk_K_r13_reg[32]/NET0131  ;
  assign n52620 = ~decrypt_pad & ~\u0_uk_K_r13_reg[11]/NET0131  ;
  assign n52621 = ~n52619 & ~n52620 ;
  assign n52622 = \u0_R13_reg[9]/NET0131  & ~n52621 ;
  assign n52623 = ~\u0_R13_reg[9]/NET0131  & n52621 ;
  assign n52624 = ~n52622 & ~n52623 ;
  assign n52625 = decrypt_pad & ~\u0_uk_K_r13_reg[40]/NET0131  ;
  assign n52626 = ~decrypt_pad & ~\u0_uk_K_r13_reg[19]/NET0131  ;
  assign n52627 = ~n52625 & ~n52626 ;
  assign n52628 = \u0_R13_reg[10]/NET0131  & ~n52627 ;
  assign n52629 = ~\u0_R13_reg[10]/NET0131  & n52627 ;
  assign n52630 = ~n52628 & ~n52629 ;
  assign n52642 = n52624 & ~n52630 ;
  assign n52643 = ~n52617 & ~n52642 ;
  assign n52633 = decrypt_pad & ~\u0_uk_K_r13_reg[41]/NET0131  ;
  assign n52634 = ~decrypt_pad & ~\u0_uk_K_r13_reg[20]/NET0131  ;
  assign n52635 = ~n52633 & ~n52634 ;
  assign n52636 = \u0_R13_reg[11]/NET0131  & ~n52635 ;
  assign n52637 = ~\u0_R13_reg[11]/NET0131  & n52635 ;
  assign n52638 = ~n52636 & ~n52637 ;
  assign n52606 = decrypt_pad & ~\u0_uk_K_r13_reg[12]/NET0131  ;
  assign n52607 = ~decrypt_pad & ~\u0_uk_K_r13_reg[48]/NET0131  ;
  assign n52608 = ~n52606 & ~n52607 ;
  assign n52609 = \u0_R13_reg[13]/NET0131  & ~n52608 ;
  assign n52610 = ~\u0_R13_reg[13]/NET0131  & n52608 ;
  assign n52611 = ~n52609 & ~n52610 ;
  assign n52639 = n52611 & ~n52624 ;
  assign n52640 = ~n52611 & n52624 ;
  assign n52641 = ~n52639 & ~n52640 ;
  assign n52644 = ~n52638 & n52641 ;
  assign n52645 = ~n52643 & n52644 ;
  assign n52618 = ~n52611 & ~n52617 ;
  assign n52631 = n52624 & n52630 ;
  assign n52632 = n52618 & n52631 ;
  assign n52646 = decrypt_pad & ~\u0_uk_K_r13_reg[24]/NET0131  ;
  assign n52647 = ~decrypt_pad & ~\u0_uk_K_r13_reg[3]/NET0131  ;
  assign n52648 = ~n52646 & ~n52647 ;
  assign n52649 = \u0_R13_reg[12]/NET0131  & ~n52648 ;
  assign n52650 = ~\u0_R13_reg[12]/NET0131  & n52648 ;
  assign n52651 = ~n52649 & ~n52650 ;
  assign n52652 = ~n52632 & n52651 ;
  assign n52653 = ~n52645 & n52652 ;
  assign n52657 = n52611 & n52617 ;
  assign n52658 = ~n52618 & ~n52657 ;
  assign n52656 = ~n52624 & ~n52630 ;
  assign n52665 = n52611 & n52638 ;
  assign n52666 = n52656 & ~n52665 ;
  assign n52667 = n52658 & n52666 ;
  assign n52668 = n52617 & n52630 ;
  assign n52669 = n52640 & n52668 ;
  assign n52654 = ~n52617 & n52638 ;
  assign n52655 = n52642 & n52654 ;
  assign n52670 = ~n52651 & ~n52655 ;
  assign n52671 = ~n52669 & n52670 ;
  assign n52672 = ~n52667 & n52671 ;
  assign n52659 = ~n52656 & ~n52658 ;
  assign n52660 = ~n52631 & n52659 ;
  assign n52661 = n52611 & ~n52617 ;
  assign n52662 = n52630 & n52661 ;
  assign n52663 = n52624 & n52662 ;
  assign n52664 = ~n52638 & n52663 ;
  assign n52673 = ~n52660 & ~n52664 ;
  assign n52674 = n52672 & n52673 ;
  assign n52675 = ~n52653 & ~n52674 ;
  assign n52677 = ~n52618 & ~n52641 ;
  assign n52678 = ~n52662 & ~n52677 ;
  assign n52679 = n52651 & ~n52678 ;
  assign n52676 = n52630 & n52639 ;
  assign n52680 = n52618 & ~n52630 ;
  assign n52681 = ~n52624 & n52680 ;
  assign n52682 = ~n52676 & ~n52681 ;
  assign n52683 = ~n52679 & n52682 ;
  assign n52684 = n52638 & ~n52683 ;
  assign n52685 = ~n52675 & ~n52684 ;
  assign n52686 = ~\u0_L13_reg[6]/NET0131  & ~n52685 ;
  assign n52687 = \u0_L13_reg[6]/NET0131  & n52685 ;
  assign n52688 = ~n52686 & ~n52687 ;
  assign n52689 = n51458 & ~n51470 ;
  assign n52690 = n51441 & ~n51450 ;
  assign n52691 = n52570 & ~n52690 ;
  assign n52692 = ~n52570 & n52583 ;
  assign n52693 = ~n52691 & ~n52692 ;
  assign n52694 = n52689 & ~n52693 ;
  assign n52695 = ~n51487 & ~n52583 ;
  assign n52696 = n52570 & n52695 ;
  assign n52697 = ~n51458 & n51470 ;
  assign n52698 = ~n52689 & ~n52697 ;
  assign n52699 = ~n52692 & n52698 ;
  assign n52700 = ~n52696 & n52699 ;
  assign n52701 = ~n52694 & ~n52700 ;
  assign n52702 = ~n51489 & ~n52701 ;
  assign n52705 = ~n52576 & n52697 ;
  assign n52706 = ~n52598 & n52705 ;
  assign n52703 = ~n51434 & ~n51481 ;
  assign n52704 = n51434 & ~n52570 ;
  assign n52707 = ~n52703 & ~n52704 ;
  assign n52708 = n52706 & n52707 ;
  assign n52709 = ~n52702 & ~n52708 ;
  assign n52710 = ~\u0_L13_reg[7]/NET0131  & n52709 ;
  assign n52711 = \u0_L13_reg[7]/NET0131  & ~n52709 ;
  assign n52712 = ~n52710 & ~n52711 ;
  assign n52729 = ~n52069 & n52133 ;
  assign n52730 = ~n52077 & ~n52350 ;
  assign n52731 = ~n52729 & n52730 ;
  assign n52732 = ~n52092 & ~n52731 ;
  assign n52727 = ~n52100 & ~n52364 ;
  assign n52728 = n52092 & ~n52727 ;
  assign n52733 = ~n52085 & ~n52128 ;
  assign n52734 = ~n52728 & n52733 ;
  assign n52735 = ~n52732 & n52734 ;
  assign n52736 = ~n52057 & ~n52735 ;
  assign n52715 = ~n52077 & ~n52125 ;
  assign n52714 = ~n52077 & n52084 ;
  assign n52716 = n52092 & ~n52714 ;
  assign n52717 = ~n52715 & n52716 ;
  assign n52713 = ~n52084 & n52111 ;
  assign n52718 = n52377 & ~n52713 ;
  assign n52719 = ~n52717 & n52718 ;
  assign n52720 = n52057 & ~n52719 ;
  assign n52721 = ~n52092 & ~n52344 ;
  assign n52722 = n52092 & ~n52375 ;
  assign n52723 = n52076 & n52085 ;
  assign n52724 = ~n52363 & ~n52723 ;
  assign n52725 = n52722 & n52724 ;
  assign n52726 = ~n52721 & ~n52725 ;
  assign n52737 = ~n52720 & ~n52726 ;
  assign n52738 = ~n52736 & n52737 ;
  assign n52739 = ~\u0_L13_reg[8]/NET0131  & ~n52738 ;
  assign n52740 = \u0_L13_reg[8]/NET0131  & n52738 ;
  assign n52741 = ~n52739 & ~n52740 ;
  assign n52743 = n52618 & n52630 ;
  assign n52744 = ~n52630 & n52661 ;
  assign n52745 = ~n52743 & ~n52744 ;
  assign n52746 = ~n52624 & n52668 ;
  assign n52747 = n52618 & n52624 ;
  assign n52748 = ~n52746 & ~n52747 ;
  assign n52749 = n52745 & n52748 ;
  assign n52750 = ~n52651 & ~n52749 ;
  assign n52742 = n52642 & n52661 ;
  assign n52751 = ~n52611 & n52617 ;
  assign n52752 = n52656 & n52751 ;
  assign n52753 = n52638 & ~n52752 ;
  assign n52754 = ~n52742 & n52753 ;
  assign n52755 = ~n52750 & n52754 ;
  assign n52758 = ~n52630 & ~n52640 ;
  assign n52759 = n52658 & n52758 ;
  assign n52760 = ~n52651 & ~n52659 ;
  assign n52761 = ~n52759 & n52760 ;
  assign n52756 = n52624 & n52657 ;
  assign n52757 = n52630 & n52756 ;
  assign n52762 = ~n52638 & ~n52757 ;
  assign n52763 = ~n52761 & n52762 ;
  assign n52764 = ~n52755 & ~n52763 ;
  assign n52769 = ~n52656 & ~n52751 ;
  assign n52770 = ~n52638 & ~n52769 ;
  assign n52768 = n52638 & ~n52656 ;
  assign n52771 = ~n52661 & ~n52768 ;
  assign n52772 = ~n52770 & n52771 ;
  assign n52765 = n52624 & n52668 ;
  assign n52766 = ~n52662 & ~n52765 ;
  assign n52767 = n52638 & ~n52766 ;
  assign n52773 = ~n52667 & ~n52767 ;
  assign n52774 = ~n52772 & n52773 ;
  assign n52775 = n52651 & ~n52774 ;
  assign n52776 = ~n52764 & ~n52775 ;
  assign n52777 = ~\u0_L13_reg[24]/NET0131  & ~n52776 ;
  assign n52778 = \u0_L13_reg[24]/NET0131  & n52776 ;
  assign n52779 = ~n52777 & ~n52778 ;
  assign n52780 = ~n52624 & ~n52657 ;
  assign n52781 = ~n52756 & ~n52780 ;
  assign n52782 = ~n52618 & ~n52781 ;
  assign n52783 = n52638 & n52747 ;
  assign n52784 = ~n52782 & ~n52783 ;
  assign n52785 = ~n52630 & ~n52784 ;
  assign n52786 = ~n52630 & n52751 ;
  assign n52787 = ~n52743 & ~n52786 ;
  assign n52788 = ~n52638 & ~n52787 ;
  assign n52789 = n52651 & ~n52663 ;
  assign n52790 = ~n52788 & n52789 ;
  assign n52791 = ~n52785 & n52790 ;
  assign n52792 = ~n52617 & ~n52624 ;
  assign n52793 = n52611 & n52792 ;
  assign n52794 = ~n52680 & ~n52756 ;
  assign n52795 = ~n52793 & n52794 ;
  assign n52796 = ~n52638 & ~n52795 ;
  assign n52797 = n52638 & ~n52747 ;
  assign n52798 = n52781 & n52797 ;
  assign n52799 = ~n52651 & ~n52681 ;
  assign n52800 = ~n52798 & n52799 ;
  assign n52801 = ~n52796 & n52800 ;
  assign n52802 = ~n52791 & ~n52801 ;
  assign n52803 = ~n52638 & n52746 ;
  assign n52804 = ~n52624 & n52743 ;
  assign n52805 = ~n52669 & ~n52804 ;
  assign n52806 = n52638 & ~n52805 ;
  assign n52807 = ~n52803 & ~n52806 ;
  assign n52808 = ~n52802 & n52807 ;
  assign n52809 = ~\u0_L13_reg[16]/NET0131  & ~n52808 ;
  assign n52810 = \u0_L13_reg[16]/NET0131  & n52808 ;
  assign n52811 = ~n52809 & ~n52810 ;
  assign n52813 = ~n52630 & ~n52658 ;
  assign n52814 = ~n52662 & ~n52813 ;
  assign n52815 = ~n52624 & ~n52814 ;
  assign n52816 = ~n52640 & n52668 ;
  assign n52817 = ~n52611 & n52642 ;
  assign n52818 = ~n52816 & ~n52817 ;
  assign n52819 = n52638 & ~n52818 ;
  assign n52820 = ~n52638 & ~n52668 ;
  assign n52821 = ~n52640 & ~n52792 ;
  assign n52822 = n52820 & n52821 ;
  assign n52823 = ~n52819 & ~n52822 ;
  assign n52824 = ~n52815 & n52823 ;
  assign n52825 = ~n52651 & ~n52824 ;
  assign n52830 = n52745 & n52753 ;
  assign n52831 = ~n52747 & n52820 ;
  assign n52832 = n52651 & ~n52831 ;
  assign n52833 = ~n52830 & n52832 ;
  assign n52812 = n52665 & n52746 ;
  assign n52826 = ~n52611 & ~n52638 ;
  assign n52827 = ~n52651 & ~n52826 ;
  assign n52828 = n52631 & ~n52657 ;
  assign n52829 = ~n52827 & n52828 ;
  assign n52834 = ~n52812 & ~n52829 ;
  assign n52835 = ~n52833 & n52834 ;
  assign n52836 = ~n52825 & n52835 ;
  assign n52837 = \u0_L13_reg[30]/NET0131  & ~n52836 ;
  assign n52838 = ~\u0_L13_reg[30]/NET0131  & n52836 ;
  assign n52839 = ~n52837 & ~n52838 ;
  assign n52841 = ~n51891 & n52505 ;
  assign n52842 = n51525 & ~n52841 ;
  assign n52843 = ~n51546 & ~n51559 ;
  assign n52844 = ~n51566 & n52843 ;
  assign n52845 = ~n51525 & n52844 ;
  assign n52840 = n51531 & n51893 ;
  assign n52846 = ~n51531 & n51594 ;
  assign n52847 = ~n52840 & ~n52846 ;
  assign n52848 = ~n52845 & n52847 ;
  assign n52849 = ~n52842 & n52848 ;
  assign n52850 = ~n51519 & ~n52849 ;
  assign n52851 = ~n51544 & n51909 ;
  assign n52852 = ~n52846 & ~n52851 ;
  assign n52853 = ~n51525 & ~n52852 ;
  assign n52855 = n51531 & ~n51554 ;
  assign n52856 = ~n51893 & n52855 ;
  assign n52854 = n51573 & n52844 ;
  assign n52857 = ~n51903 & ~n52854 ;
  assign n52858 = ~n52856 & n52857 ;
  assign n52859 = n51519 & ~n52858 ;
  assign n52860 = ~n52853 & ~n52859 ;
  assign n52861 = ~n52850 & n52860 ;
  assign n52862 = ~\u0_L13_reg[9]/NET0131  & ~n52861 ;
  assign n52863 = \u0_L13_reg[9]/NET0131  & n52861 ;
  assign n52864 = ~n52862 & ~n52863 ;
  assign n52880 = ~n52069 & n52119 ;
  assign n52881 = n52069 & n52133 ;
  assign n52882 = ~n52880 & ~n52881 ;
  assign n52883 = n52092 & ~n52882 ;
  assign n52879 = ~n52092 & n52350 ;
  assign n52884 = ~n52134 & ~n52344 ;
  assign n52885 = ~n52879 & n52884 ;
  assign n52886 = ~n52883 & n52885 ;
  assign n52887 = n52057 & ~n52886 ;
  assign n52865 = ~n52364 & n52722 ;
  assign n52866 = ~n52084 & n52127 ;
  assign n52867 = ~n52714 & ~n52866 ;
  assign n52868 = ~n52092 & ~n52867 ;
  assign n52869 = ~n52865 & ~n52868 ;
  assign n52870 = ~n52126 & ~n52729 ;
  assign n52871 = n52092 & ~n52870 ;
  assign n52873 = n52076 & ~n52101 ;
  assign n52874 = n52069 & ~n52873 ;
  assign n52872 = n52092 & ~n52110 ;
  assign n52875 = ~n52729 & ~n52872 ;
  assign n52876 = ~n52874 & n52875 ;
  assign n52877 = ~n52871 & ~n52876 ;
  assign n52878 = ~n52057 & ~n52877 ;
  assign n52888 = ~n52869 & ~n52878 ;
  assign n52889 = ~n52887 & n52888 ;
  assign n52890 = ~\u0_L13_reg[3]/NET0131  & ~n52889 ;
  assign n52891 = \u0_L13_reg[3]/NET0131  & n52889 ;
  assign n52892 = ~n52890 & ~n52891 ;
  assign n52896 = n52223 & ~n52314 ;
  assign n52893 = n52200 & n52212 ;
  assign n52894 = ~n52223 & ~n52893 ;
  assign n52895 = n52462 & n52894 ;
  assign n52897 = n52181 & ~n52330 ;
  assign n52898 = ~n52895 & n52897 ;
  assign n52899 = ~n52896 & n52898 ;
  assign n52903 = ~n52181 & ~n52449 ;
  assign n52904 = ~n52233 & n52903 ;
  assign n52901 = ~n52187 & ~n52461 ;
  assign n52902 = n52321 & n52901 ;
  assign n52900 = n52223 & n52244 ;
  assign n52905 = ~n52301 & ~n52900 ;
  assign n52906 = ~n52902 & n52905 ;
  assign n52907 = n52904 & n52906 ;
  assign n52908 = ~n52899 & ~n52907 ;
  assign n52909 = ~n52300 & ~n52472 ;
  assign n52910 = n52223 & ~n52909 ;
  assign n52911 = ~n52223 & n52227 ;
  assign n52912 = ~n52910 & ~n52911 ;
  assign n52913 = ~n52908 & n52912 ;
  assign n52914 = \u0_L13_reg[18]/NET0131  & n52913 ;
  assign n52915 = ~\u0_L13_reg[18]/NET0131  & ~n52913 ;
  assign n52916 = ~n52914 & ~n52915 ;
  assign n52930 = decrypt_pad & ~\u0_uk_K_r12_reg[24]/NET0131  ;
  assign n52931 = ~decrypt_pad & ~\u0_uk_K_r12_reg[32]/NET0131  ;
  assign n52932 = ~n52930 & ~n52931 ;
  assign n52933 = \u0_R12_reg[3]/NET0131  & ~n52932 ;
  assign n52934 = ~\u0_R12_reg[3]/NET0131  & n52932 ;
  assign n52935 = ~n52933 & ~n52934 ;
  assign n52917 = decrypt_pad & ~\u0_uk_K_r12_reg[11]/NET0131  ;
  assign n52918 = ~decrypt_pad & ~\u0_uk_K_r12_reg[19]/NET0131  ;
  assign n52919 = ~n52917 & ~n52918 ;
  assign n52920 = \u0_R12_reg[32]/NET0131  & ~n52919 ;
  assign n52921 = ~\u0_R12_reg[32]/NET0131  & n52919 ;
  assign n52922 = ~n52920 & ~n52921 ;
  assign n52937 = decrypt_pad & ~\u0_uk_K_r12_reg[5]/NET0131  ;
  assign n52938 = ~decrypt_pad & ~\u0_uk_K_r12_reg[13]/NET0131  ;
  assign n52939 = ~n52937 & ~n52938 ;
  assign n52940 = \u0_R12_reg[5]/NET0131  & ~n52939 ;
  assign n52941 = ~\u0_R12_reg[5]/NET0131  & n52939 ;
  assign n52942 = ~n52940 & ~n52941 ;
  assign n52923 = decrypt_pad & ~\u0_uk_K_r12_reg[47]/NET0131  ;
  assign n52924 = ~decrypt_pad & ~\u0_uk_K_r12_reg[55]/NET0131  ;
  assign n52925 = ~n52923 & ~n52924 ;
  assign n52926 = \u0_R12_reg[2]/NET0131  & ~n52925 ;
  assign n52927 = ~\u0_R12_reg[2]/NET0131  & n52925 ;
  assign n52928 = ~n52926 & ~n52927 ;
  assign n52947 = decrypt_pad & ~\u0_uk_K_r12_reg[32]/NET0131  ;
  assign n52948 = ~decrypt_pad & ~\u0_uk_K_r12_reg[40]/NET0131  ;
  assign n52949 = ~n52947 & ~n52948 ;
  assign n52950 = \u0_R12_reg[1]/NET0131  & ~n52949 ;
  assign n52951 = ~\u0_R12_reg[1]/NET0131  & n52949 ;
  assign n52952 = ~n52950 & ~n52951 ;
  assign n52956 = n52928 & n52952 ;
  assign n52961 = ~n52942 & n52956 ;
  assign n52962 = n52922 & n52961 ;
  assign n52954 = n52922 & ~n52928 ;
  assign n52963 = n52942 & n52954 ;
  assign n52964 = ~n52962 & ~n52963 ;
  assign n52965 = n52935 & ~n52964 ;
  assign n52929 = ~n52922 & n52928 ;
  assign n52936 = n52929 & n52935 ;
  assign n52943 = n52936 & n52942 ;
  assign n52944 = ~n52922 & ~n52942 ;
  assign n52945 = ~n52928 & n52944 ;
  assign n52946 = ~n52943 & ~n52945 ;
  assign n52953 = ~n52946 & n52952 ;
  assign n52955 = ~n52929 & ~n52954 ;
  assign n52957 = n52942 & ~n52952 ;
  assign n52958 = ~n52935 & ~n52956 ;
  assign n52959 = ~n52957 & n52958 ;
  assign n52960 = n52955 & n52959 ;
  assign n52966 = n52954 & n52957 ;
  assign n52967 = ~n52960 & ~n52966 ;
  assign n52968 = ~n52953 & n52967 ;
  assign n52969 = ~n52965 & n52968 ;
  assign n52970 = decrypt_pad & ~\u0_uk_K_r12_reg[34]/NET0131  ;
  assign n52971 = ~decrypt_pad & ~\u0_uk_K_r12_reg[10]/P0001  ;
  assign n52972 = ~n52970 & ~n52971 ;
  assign n52973 = \u0_R12_reg[4]/NET0131  & ~n52972 ;
  assign n52974 = ~\u0_R12_reg[4]/NET0131  & n52972 ;
  assign n52975 = ~n52973 & ~n52974 ;
  assign n52976 = ~n52969 & ~n52975 ;
  assign n52990 = ~n52935 & n52952 ;
  assign n52977 = ~n52942 & ~n52952 ;
  assign n52991 = ~n52928 & n52977 ;
  assign n52992 = ~n52990 & ~n52991 ;
  assign n52993 = n52922 & ~n52992 ;
  assign n52987 = n52928 & n52944 ;
  assign n52988 = ~n52957 & ~n52987 ;
  assign n52989 = n52935 & ~n52988 ;
  assign n52994 = ~n52928 & n52935 ;
  assign n52995 = n52952 & ~n52994 ;
  assign n52982 = ~n52928 & ~n52942 ;
  assign n52996 = ~n52922 & ~n52982 ;
  assign n52997 = ~n52995 & n52996 ;
  assign n52998 = ~n52989 & ~n52997 ;
  assign n52999 = ~n52993 & n52998 ;
  assign n53000 = n52975 & ~n52999 ;
  assign n52983 = n52952 & n52982 ;
  assign n52979 = n52922 & n52942 ;
  assign n52980 = n52956 & n52979 ;
  assign n52981 = n52929 & n52957 ;
  assign n52984 = ~n52980 & ~n52981 ;
  assign n52985 = ~n52983 & n52984 ;
  assign n52986 = ~n52935 & ~n52985 ;
  assign n52978 = n52936 & n52977 ;
  assign n53001 = ~n52928 & ~n52952 ;
  assign n53002 = n52922 & n52935 ;
  assign n53003 = n53001 & n53002 ;
  assign n53004 = ~n52978 & ~n53003 ;
  assign n53005 = ~n52986 & n53004 ;
  assign n53006 = ~n53000 & n53005 ;
  assign n53007 = ~n52976 & n53006 ;
  assign n53008 = ~\u0_L12_reg[31]/NET0131  & ~n53007 ;
  assign n53009 = \u0_L12_reg[31]/NET0131  & n53007 ;
  assign n53010 = ~n53008 & ~n53009 ;
  assign n53011 = decrypt_pad & ~\u0_uk_K_r12_reg[1]/NET0131  ;
  assign n53012 = ~decrypt_pad & ~\u0_uk_K_r12_reg[7]/P0001  ;
  assign n53013 = ~n53011 & ~n53012 ;
  assign n53014 = \u0_R12_reg[24]/NET0131  & ~n53013 ;
  assign n53015 = ~\u0_R12_reg[24]/NET0131  & n53013 ;
  assign n53016 = ~n53014 & ~n53015 ;
  assign n53017 = decrypt_pad & ~\u0_uk_K_r12_reg[30]/NET0131  ;
  assign n53018 = ~decrypt_pad & ~\u0_uk_K_r12_reg[36]/NET0131  ;
  assign n53019 = ~n53017 & ~n53018 ;
  assign n53020 = \u0_R12_reg[23]/NET0131  & ~n53019 ;
  assign n53021 = ~\u0_R12_reg[23]/NET0131  & n53019 ;
  assign n53022 = ~n53020 & ~n53021 ;
  assign n53023 = decrypt_pad & ~\u0_uk_K_r12_reg[50]/NET0131  ;
  assign n53024 = ~decrypt_pad & ~\u0_uk_K_r12_reg[1]/NET0131  ;
  assign n53025 = ~n53023 & ~n53024 ;
  assign n53026 = \u0_R12_reg[21]/NET0131  & ~n53025 ;
  assign n53027 = ~\u0_R12_reg[21]/NET0131  & n53025 ;
  assign n53028 = ~n53026 & ~n53027 ;
  assign n53029 = decrypt_pad & ~\u0_uk_K_r12_reg[45]/NET0131  ;
  assign n53030 = ~decrypt_pad & ~\u0_uk_K_r12_reg[23]/NET0131  ;
  assign n53031 = ~n53029 & ~n53030 ;
  assign n53032 = \u0_R12_reg[22]/NET0131  & ~n53031 ;
  assign n53033 = ~\u0_R12_reg[22]/NET0131  & n53031 ;
  assign n53034 = ~n53032 & ~n53033 ;
  assign n53035 = ~n53028 & ~n53034 ;
  assign n53036 = decrypt_pad & ~\u0_uk_K_r12_reg[35]/NET0131  ;
  assign n53037 = ~decrypt_pad & ~\u0_uk_K_r12_reg[45]/NET0131  ;
  assign n53038 = ~n53036 & ~n53037 ;
  assign n53039 = \u0_R12_reg[20]/NET0131  & ~n53038 ;
  assign n53040 = ~\u0_R12_reg[20]/NET0131  & n53038 ;
  assign n53041 = ~n53039 & ~n53040 ;
  assign n53042 = decrypt_pad & ~\u0_uk_K_r12_reg[51]/NET0131  ;
  assign n53043 = ~decrypt_pad & ~\u0_uk_K_r12_reg[2]/NET0131  ;
  assign n53044 = ~n53042 & ~n53043 ;
  assign n53045 = \u0_R12_reg[25]/NET0131  & ~n53044 ;
  assign n53046 = ~\u0_R12_reg[25]/NET0131  & n53044 ;
  assign n53047 = ~n53045 & ~n53046 ;
  assign n53048 = n53041 & n53047 ;
  assign n53049 = n53035 & n53048 ;
  assign n53050 = n53028 & ~n53041 ;
  assign n53051 = n53034 & n53050 ;
  assign n53052 = ~n53035 & ~n53051 ;
  assign n53053 = ~n53034 & ~n53047 ;
  assign n53054 = ~n53048 & ~n53053 ;
  assign n53055 = n53052 & n53054 ;
  assign n53056 = ~n53049 & ~n53055 ;
  assign n53057 = ~n53022 & ~n53056 ;
  assign n53058 = ~n53028 & ~n53053 ;
  assign n53059 = n53022 & ~n53058 ;
  assign n53060 = ~n53034 & ~n53041 ;
  assign n53061 = n53028 & ~n53047 ;
  assign n53062 = n53041 & n53061 ;
  assign n53063 = ~n53060 & ~n53062 ;
  assign n53064 = n53059 & n53063 ;
  assign n53065 = ~n53057 & ~n53064 ;
  assign n53066 = n53016 & ~n53065 ;
  assign n53067 = ~n53022 & ~n53048 ;
  assign n53068 = ~n53028 & n53047 ;
  assign n53069 = ~n53028 & n53041 ;
  assign n53070 = ~n53068 & ~n53069 ;
  assign n53071 = ~n53067 & ~n53070 ;
  assign n53072 = ~n53022 & n53050 ;
  assign n53073 = ~n53071 & ~n53072 ;
  assign n53074 = n53034 & ~n53073 ;
  assign n53077 = n53041 & ~n53061 ;
  assign n53078 = n53022 & n53077 ;
  assign n53075 = n53041 & ~n53068 ;
  assign n53076 = ~n53022 & ~n53075 ;
  assign n53079 = ~n53034 & ~n53076 ;
  assign n53080 = ~n53078 & n53079 ;
  assign n53081 = ~n53074 & ~n53080 ;
  assign n53082 = ~n53016 & ~n53081 ;
  assign n53087 = ~n53041 & n53068 ;
  assign n53088 = n53022 & n53087 ;
  assign n53089 = ~n53022 & n53062 ;
  assign n53090 = ~n53088 & ~n53089 ;
  assign n53091 = ~n53034 & ~n53090 ;
  assign n53084 = ~n53041 & ~n53047 ;
  assign n53083 = ~n53022 & ~n53034 ;
  assign n53085 = ~n53028 & n53083 ;
  assign n53086 = n53084 & n53085 ;
  assign n53092 = n53034 & n53048 ;
  assign n53093 = n53050 & n53053 ;
  assign n53094 = ~n53092 & ~n53093 ;
  assign n53095 = n53022 & ~n53094 ;
  assign n53096 = ~n53086 & ~n53095 ;
  assign n53097 = ~n53091 & n53096 ;
  assign n53098 = ~n53082 & n53097 ;
  assign n53099 = ~n53066 & n53098 ;
  assign n53100 = \u0_L12_reg[11]/NET0131  & ~n53099 ;
  assign n53101 = ~\u0_L12_reg[11]/NET0131  & n53099 ;
  assign n53102 = ~n53100 & ~n53101 ;
  assign n53130 = decrypt_pad & ~\u0_uk_K_r12_reg[21]/NET0131  ;
  assign n53131 = ~decrypt_pad & ~\u0_uk_K_r12_reg[31]/NET0131  ;
  assign n53132 = ~n53130 & ~n53131 ;
  assign n53133 = \u0_R12_reg[27]/NET0131  & ~n53132 ;
  assign n53134 = ~\u0_R12_reg[27]/NET0131  & n53132 ;
  assign n53135 = ~n53133 & ~n53134 ;
  assign n53123 = decrypt_pad & ~\u0_uk_K_r12_reg[31]/NET0131  ;
  assign n53124 = ~decrypt_pad & ~\u0_uk_K_r12_reg[9]/NET0131  ;
  assign n53125 = ~n53123 & ~n53124 ;
  assign n53126 = \u0_R12_reg[25]/NET0131  & ~n53125 ;
  assign n53127 = ~\u0_R12_reg[25]/NET0131  & n53125 ;
  assign n53128 = ~n53126 & ~n53127 ;
  assign n53103 = decrypt_pad & ~\u0_uk_K_r12_reg[23]/NET0131  ;
  assign n53104 = ~decrypt_pad & ~\u0_uk_K_r12_reg[29]/NET0131  ;
  assign n53105 = ~n53103 & ~n53104 ;
  assign n53106 = \u0_R12_reg[24]/NET0131  & ~n53105 ;
  assign n53107 = ~\u0_R12_reg[24]/NET0131  & n53105 ;
  assign n53108 = ~n53106 & ~n53107 ;
  assign n53116 = decrypt_pad & ~\u0_uk_K_r12_reg[0]/NET0131  ;
  assign n53117 = ~decrypt_pad & ~\u0_uk_K_r12_reg[37]/NET0131  ;
  assign n53118 = ~n53116 & ~n53117 ;
  assign n53119 = \u0_R12_reg[29]/NET0131  & ~n53118 ;
  assign n53120 = ~\u0_R12_reg[29]/NET0131  & n53118 ;
  assign n53121 = ~n53119 & ~n53120 ;
  assign n53139 = n53108 & ~n53121 ;
  assign n53140 = n53128 & n53139 ;
  assign n53109 = decrypt_pad & ~\u0_uk_K_r12_reg[43]/NET0131  ;
  assign n53110 = ~decrypt_pad & ~\u0_uk_K_r12_reg[49]/NET0131  ;
  assign n53111 = ~n53109 & ~n53110 ;
  assign n53112 = \u0_R12_reg[26]/NET0131  & ~n53111 ;
  assign n53113 = ~\u0_R12_reg[26]/NET0131  & n53111 ;
  assign n53114 = ~n53112 & ~n53113 ;
  assign n53115 = n53108 & n53114 ;
  assign n53122 = n53115 & n53121 ;
  assign n53136 = ~n53121 & ~n53128 ;
  assign n53137 = ~n53108 & n53114 ;
  assign n53138 = n53136 & n53137 ;
  assign n53141 = ~n53122 & ~n53138 ;
  assign n53142 = ~n53140 & n53141 ;
  assign n53143 = ~n53135 & ~n53142 ;
  assign n53144 = ~n53108 & n53121 ;
  assign n53145 = ~n53128 & n53135 ;
  assign n53146 = n53144 & ~n53145 ;
  assign n53147 = n53108 & ~n53128 ;
  assign n53148 = n53121 & ~n53135 ;
  assign n53149 = n53147 & ~n53148 ;
  assign n53150 = ~n53146 & ~n53149 ;
  assign n53151 = ~n53114 & ~n53150 ;
  assign n53129 = n53122 & n53128 ;
  assign n53152 = decrypt_pad & ~\u0_uk_K_r12_reg[8]/NET0131  ;
  assign n53153 = ~decrypt_pad & ~\u0_uk_K_r12_reg[14]/NET0131  ;
  assign n53154 = ~n53152 & ~n53153 ;
  assign n53155 = \u0_R12_reg[28]/NET0131  & ~n53154 ;
  assign n53156 = ~\u0_R12_reg[28]/NET0131  & n53154 ;
  assign n53157 = ~n53155 & ~n53156 ;
  assign n53158 = ~n53129 & ~n53157 ;
  assign n53159 = ~n53151 & n53158 ;
  assign n53160 = ~n53143 & n53159 ;
  assign n53163 = n53114 & ~n53128 ;
  assign n53165 = n53121 & n53128 ;
  assign n53166 = ~n53114 & n53165 ;
  assign n53167 = ~n53163 & ~n53166 ;
  assign n53168 = n53108 & ~n53167 ;
  assign n53169 = n53135 & ~n53168 ;
  assign n53170 = n53121 & n53147 ;
  assign n53171 = ~n53114 & n53170 ;
  assign n53172 = ~n53108 & n53165 ;
  assign n53173 = ~n53135 & ~n53172 ;
  assign n53174 = ~n53171 & n53173 ;
  assign n53175 = ~n53169 & ~n53174 ;
  assign n53161 = ~n53108 & n53136 ;
  assign n53162 = ~n53114 & n53161 ;
  assign n53164 = n53144 & n53163 ;
  assign n53176 = n53157 & ~n53164 ;
  assign n53177 = ~n53162 & n53176 ;
  assign n53178 = ~n53175 & n53177 ;
  assign n53179 = ~n53160 & ~n53178 ;
  assign n53180 = ~n53114 & n53128 ;
  assign n53181 = ~n53108 & n53180 ;
  assign n53182 = n53108 & n53128 ;
  assign n53183 = n53114 & n53182 ;
  assign n53184 = ~n53135 & ~n53183 ;
  assign n53185 = ~n53181 & n53184 ;
  assign n53186 = n53128 & n53137 ;
  assign n53187 = ~n53121 & n53186 ;
  assign n53188 = ~n53164 & ~n53187 ;
  assign n53189 = n53136 & ~n53137 ;
  assign n53190 = n53135 & ~n53189 ;
  assign n53191 = n53188 & n53190 ;
  assign n53192 = ~n53185 & ~n53191 ;
  assign n53193 = ~n53179 & ~n53192 ;
  assign n53194 = \u0_L12_reg[22]/NET0131  & n53193 ;
  assign n53195 = ~\u0_L12_reg[22]/NET0131  & ~n53193 ;
  assign n53196 = ~n53194 & ~n53195 ;
  assign n53216 = ~n52944 & ~n52979 ;
  assign n53217 = ~n52952 & ~n53216 ;
  assign n53218 = ~n52945 & ~n53217 ;
  assign n53219 = ~n52935 & ~n53218 ;
  assign n53197 = ~n52942 & n52952 ;
  assign n53220 = ~n52957 & ~n53197 ;
  assign n53221 = n52922 & n53220 ;
  assign n53222 = n52935 & n53221 ;
  assign n53223 = ~n52962 & ~n52981 ;
  assign n53224 = ~n53222 & n53223 ;
  assign n53225 = ~n53219 & n53224 ;
  assign n53226 = ~n52975 & ~n53225 ;
  assign n53200 = ~n52922 & ~n53001 ;
  assign n53201 = ~n52966 & ~n53200 ;
  assign n53202 = n52935 & ~n53201 ;
  assign n53203 = ~n52935 & ~n52954 ;
  assign n53204 = ~n53200 & n53203 ;
  assign n53198 = n52954 & n53197 ;
  assign n53199 = n52942 & n52956 ;
  assign n53205 = ~n53198 & ~n53199 ;
  assign n53206 = ~n53204 & n53205 ;
  assign n53207 = ~n53202 & n53206 ;
  assign n53208 = n52975 & ~n53207 ;
  assign n53212 = ~n52922 & n53197 ;
  assign n53213 = n52928 & ~n53212 ;
  assign n53209 = ~n52922 & n52942 ;
  assign n53210 = n52952 & n53209 ;
  assign n53211 = ~n52928 & ~n53210 ;
  assign n53214 = n52935 & ~n53211 ;
  assign n53215 = ~n53213 & n53214 ;
  assign n53227 = ~n53208 & ~n53215 ;
  assign n53228 = ~n53226 & n53227 ;
  assign n53229 = ~\u0_L12_reg[17]/NET0131  & ~n53228 ;
  assign n53230 = \u0_L12_reg[17]/NET0131  & n53228 ;
  assign n53231 = ~n53229 & ~n53230 ;
  assign n53238 = decrypt_pad & ~\u0_uk_K_r12_reg[19]/NET0131  ;
  assign n53239 = ~decrypt_pad & ~\u0_uk_K_r12_reg[27]/NET0131  ;
  assign n53240 = ~n53238 & ~n53239 ;
  assign n53241 = \u0_R12_reg[13]/NET0131  & ~n53240 ;
  assign n53242 = ~\u0_R12_reg[13]/NET0131  & n53240 ;
  assign n53243 = ~n53241 & ~n53242 ;
  assign n53258 = decrypt_pad & ~\u0_uk_K_r12_reg[41]/NET0131  ;
  assign n53259 = ~decrypt_pad & ~\u0_uk_K_r12_reg[17]/NET0131  ;
  assign n53260 = ~n53258 & ~n53259 ;
  assign n53261 = \u0_R12_reg[17]/NET0131  & ~n53260 ;
  assign n53262 = ~\u0_R12_reg[17]/NET0131  & n53260 ;
  assign n53263 = ~n53261 & ~n53262 ;
  assign n53232 = decrypt_pad & ~\u0_uk_K_r12_reg[20]/NET0131  ;
  assign n53233 = ~decrypt_pad & ~\u0_uk_K_r12_reg[53]/NET0131  ;
  assign n53234 = ~n53232 & ~n53233 ;
  assign n53235 = \u0_R12_reg[14]/NET0131  & ~n53234 ;
  assign n53236 = ~\u0_R12_reg[14]/NET0131  & n53234 ;
  assign n53237 = ~n53235 & ~n53236 ;
  assign n53251 = decrypt_pad & ~\u0_uk_K_r12_reg[25]/NET0131  ;
  assign n53252 = ~decrypt_pad & ~\u0_uk_K_r12_reg[33]/NET0131  ;
  assign n53253 = ~n53251 & ~n53252 ;
  assign n53254 = \u0_R12_reg[12]/NET0131  & ~n53253 ;
  assign n53255 = ~\u0_R12_reg[12]/NET0131  & n53253 ;
  assign n53256 = ~n53254 & ~n53255 ;
  assign n53278 = n53237 & n53256 ;
  assign n53279 = n53263 & n53278 ;
  assign n53280 = n53243 & n53279 ;
  assign n53292 = decrypt_pad & ~\u0_uk_K_r12_reg[4]/NET0131  ;
  assign n53293 = ~decrypt_pad & ~\u0_uk_K_r12_reg[12]/NET0131  ;
  assign n53294 = ~n53292 & ~n53293 ;
  assign n53295 = \u0_R12_reg[16]/NET0131  & ~n53294 ;
  assign n53296 = ~\u0_R12_reg[16]/NET0131  & n53294 ;
  assign n53297 = ~n53295 & ~n53296 ;
  assign n53298 = ~n53280 & n53297 ;
  assign n53244 = decrypt_pad & ~\u0_uk_K_r12_reg[53]/NET0131  ;
  assign n53245 = ~decrypt_pad & ~\u0_uk_K_r12_reg[4]/NET0131  ;
  assign n53246 = ~n53244 & ~n53245 ;
  assign n53247 = \u0_R12_reg[15]/NET0131  & ~n53246 ;
  assign n53248 = ~\u0_R12_reg[15]/NET0131  & n53246 ;
  assign n53249 = ~n53247 & ~n53248 ;
  assign n53267 = ~n53237 & ~n53249 ;
  assign n53266 = n53243 & ~n53256 ;
  assign n53273 = ~n53243 & n53256 ;
  assign n53281 = ~n53266 & ~n53273 ;
  assign n53282 = n53267 & ~n53281 ;
  assign n53283 = ~n53256 & n53263 ;
  assign n53290 = n53249 & n53283 ;
  assign n53291 = ~n53243 & n53290 ;
  assign n53299 = ~n53282 & ~n53291 ;
  assign n53300 = n53298 & n53299 ;
  assign n53250 = n53243 & n53249 ;
  assign n53257 = n53250 & n53256 ;
  assign n53264 = n53257 & ~n53263 ;
  assign n53284 = n53243 & n53283 ;
  assign n53285 = ~n53237 & n53284 ;
  assign n53286 = ~n53264 & ~n53285 ;
  assign n53270 = ~n53243 & ~n53263 ;
  assign n53287 = ~n53256 & n53270 ;
  assign n53288 = ~n53249 & n53287 ;
  assign n53289 = n53237 & n53288 ;
  assign n53301 = n53286 & ~n53289 ;
  assign n53302 = n53300 & n53301 ;
  assign n53314 = n53237 & n53250 ;
  assign n53315 = ~n53256 & n53314 ;
  assign n53313 = n53249 & n53287 ;
  assign n53316 = ~n53297 & ~n53313 ;
  assign n53317 = ~n53315 & n53316 ;
  assign n53309 = ~n53243 & n53263 ;
  assign n53310 = ~n53263 & n53278 ;
  assign n53311 = ~n53309 & ~n53310 ;
  assign n53312 = ~n53249 & ~n53311 ;
  assign n53303 = ~n53237 & n53273 ;
  assign n53304 = ~n53257 & ~n53303 ;
  assign n53305 = n53263 & ~n53304 ;
  assign n53271 = ~n53237 & ~n53256 ;
  assign n53272 = n53270 & n53271 ;
  assign n53306 = ~n53263 & n53266 ;
  assign n53307 = n53237 & n53306 ;
  assign n53308 = ~n53272 & ~n53307 ;
  assign n53318 = ~n53305 & n53308 ;
  assign n53319 = ~n53312 & n53318 ;
  assign n53320 = n53317 & n53319 ;
  assign n53321 = ~n53302 & ~n53320 ;
  assign n53274 = ~n53263 & n53273 ;
  assign n53275 = n53237 & n53274 ;
  assign n53276 = ~n53272 & ~n53275 ;
  assign n53277 = n53249 & ~n53276 ;
  assign n53265 = ~n53237 & n53264 ;
  assign n53268 = n53263 & n53267 ;
  assign n53269 = n53266 & n53268 ;
  assign n53322 = ~n53265 & ~n53269 ;
  assign n53323 = ~n53277 & n53322 ;
  assign n53324 = ~n53321 & n53323 ;
  assign n53325 = ~\u0_L12_reg[20]/NET0131  & ~n53324 ;
  assign n53326 = \u0_L12_reg[20]/NET0131  & n53324 ;
  assign n53327 = ~n53325 & ~n53326 ;
  assign n53329 = ~n53047 & ~n53052 ;
  assign n53330 = ~n53061 & n53075 ;
  assign n53331 = ~n53329 & ~n53330 ;
  assign n53332 = n53022 & ~n53331 ;
  assign n53328 = n53034 & n53087 ;
  assign n53333 = n53034 & n53062 ;
  assign n53334 = ~n53034 & n53048 ;
  assign n53335 = n53028 & n53060 ;
  assign n53336 = ~n53334 & ~n53335 ;
  assign n53337 = ~n53333 & n53336 ;
  assign n53338 = ~n53022 & ~n53337 ;
  assign n53339 = ~n53328 & ~n53338 ;
  assign n53340 = ~n53332 & n53339 ;
  assign n53341 = ~n53016 & ~n53340 ;
  assign n53345 = n53034 & ~n53047 ;
  assign n53346 = n53050 & ~n53345 ;
  assign n53347 = ~n53333 & ~n53346 ;
  assign n53348 = n53022 & ~n53347 ;
  assign n53349 = n53034 & ~n53048 ;
  assign n53350 = ~n53084 & n53349 ;
  assign n53351 = ~n53059 & n53336 ;
  assign n53352 = ~n53350 & n53351 ;
  assign n53353 = ~n53348 & ~n53352 ;
  assign n53354 = n53016 & ~n53353 ;
  assign n53342 = n53028 & n53047 ;
  assign n53343 = n53022 & ~n53034 ;
  assign n53344 = n53342 & n53343 ;
  assign n53355 = n53053 & n53069 ;
  assign n53356 = ~n53344 & ~n53355 ;
  assign n53357 = ~n53354 & n53356 ;
  assign n53358 = ~n53341 & n53357 ;
  assign n53359 = \u0_L12_reg[29]/NET0131  & ~n53358 ;
  assign n53360 = ~\u0_L12_reg[29]/NET0131  & n53358 ;
  assign n53361 = ~n53359 & ~n53360 ;
  assign n53362 = decrypt_pad & ~\u0_uk_K_r12_reg[28]/NET0131  ;
  assign n53363 = ~decrypt_pad & ~\u0_uk_K_r12_reg[38]/NET0131  ;
  assign n53364 = ~n53362 & ~n53363 ;
  assign n53365 = \u0_R12_reg[32]/NET0131  & ~n53364 ;
  assign n53366 = ~\u0_R12_reg[32]/NET0131  & n53364 ;
  assign n53367 = ~n53365 & ~n53366 ;
  assign n53401 = decrypt_pad & ~\u0_uk_K_r12_reg[22]/NET0131  ;
  assign n53402 = ~decrypt_pad & ~\u0_uk_K_r12_reg[28]/NET0131  ;
  assign n53403 = ~n53401 & ~n53402 ;
  assign n53404 = \u0_R12_reg[31]/P0001  & ~n53403 ;
  assign n53405 = ~\u0_R12_reg[31]/P0001  & n53403 ;
  assign n53406 = ~n53404 & ~n53405 ;
  assign n53380 = decrypt_pad & ~\u0_uk_K_r12_reg[9]/NET0131  ;
  assign n53381 = ~decrypt_pad & ~\u0_uk_K_r12_reg[15]/NET0131  ;
  assign n53382 = ~n53380 & ~n53381 ;
  assign n53383 = \u0_R12_reg[29]/NET0131  & ~n53382 ;
  assign n53384 = ~\u0_R12_reg[29]/NET0131  & n53382 ;
  assign n53385 = ~n53383 & ~n53384 ;
  assign n53387 = decrypt_pad & ~\u0_uk_K_r12_reg[49]/NET0131  ;
  assign n53388 = ~decrypt_pad & ~\u0_uk_K_r12_reg[0]/NET0131  ;
  assign n53389 = ~n53387 & ~n53388 ;
  assign n53390 = \u0_R12_reg[1]/NET0131  & ~n53389 ;
  assign n53391 = ~\u0_R12_reg[1]/NET0131  & n53389 ;
  assign n53392 = ~n53390 & ~n53391 ;
  assign n53368 = decrypt_pad & ~\u0_uk_K_r12_reg[38]/NET0131  ;
  assign n53369 = ~decrypt_pad & ~\u0_uk_K_r12_reg[16]/NET0131  ;
  assign n53370 = ~n53368 & ~n53369 ;
  assign n53371 = \u0_R12_reg[30]/NET0131  & ~n53370 ;
  assign n53372 = ~\u0_R12_reg[30]/NET0131  & n53370 ;
  assign n53373 = ~n53371 & ~n53372 ;
  assign n53374 = decrypt_pad & ~\u0_uk_K_r12_reg[37]/NET0131  ;
  assign n53375 = ~decrypt_pad & ~\u0_uk_K_r12_reg[43]/NET0131  ;
  assign n53376 = ~n53374 & ~n53375 ;
  assign n53377 = \u0_R12_reg[28]/NET0131  & ~n53376 ;
  assign n53378 = ~\u0_R12_reg[28]/NET0131  & n53376 ;
  assign n53379 = ~n53377 & ~n53378 ;
  assign n53408 = ~n53373 & n53379 ;
  assign n53410 = ~n53392 & n53408 ;
  assign n53411 = n53385 & n53410 ;
  assign n53422 = n53385 & ~n53392 ;
  assign n53423 = ~n53408 & ~n53422 ;
  assign n53424 = ~n53411 & ~n53423 ;
  assign n53425 = n53406 & ~n53424 ;
  assign n53426 = ~n53373 & ~n53385 ;
  assign n53427 = ~n53379 & n53426 ;
  assign n53428 = n53379 & ~n53385 ;
  assign n53429 = n53373 & n53428 ;
  assign n53430 = ~n53406 & ~n53429 ;
  assign n53431 = ~n53427 & n53430 ;
  assign n53432 = ~n53425 & ~n53431 ;
  assign n53413 = n53373 & ~n53379 ;
  assign n53433 = n53385 & n53413 ;
  assign n53434 = n53392 & n53433 ;
  assign n53435 = ~n53432 & ~n53434 ;
  assign n53436 = n53367 & ~n53435 ;
  assign n53395 = ~n53385 & ~n53392 ;
  assign n53396 = n53373 & n53395 ;
  assign n53397 = n53379 & n53396 ;
  assign n53398 = ~n53379 & n53392 ;
  assign n53399 = ~n53385 & n53398 ;
  assign n53400 = ~n53397 & ~n53399 ;
  assign n53407 = ~n53400 & n53406 ;
  assign n53386 = n53379 & n53385 ;
  assign n53393 = n53386 & n53392 ;
  assign n53394 = n53373 & n53393 ;
  assign n53409 = ~n53406 & n53408 ;
  assign n53417 = ~n53394 & ~n53409 ;
  assign n53414 = ~n53392 & ~n53413 ;
  assign n53412 = ~n53385 & n53392 ;
  assign n53415 = ~n53406 & ~n53412 ;
  assign n53416 = ~n53414 & n53415 ;
  assign n53418 = ~n53411 & ~n53416 ;
  assign n53419 = n53417 & n53418 ;
  assign n53420 = ~n53407 & n53419 ;
  assign n53421 = ~n53367 & ~n53420 ;
  assign n53437 = n53409 & n53422 ;
  assign n53438 = ~n53392 & n53433 ;
  assign n53439 = ~n53392 & n53427 ;
  assign n53440 = ~n53438 & ~n53439 ;
  assign n53441 = n53408 & n53412 ;
  assign n53442 = n53373 & n53399 ;
  assign n53443 = ~n53441 & ~n53442 ;
  assign n53444 = n53440 & n53443 ;
  assign n53445 = n53406 & ~n53444 ;
  assign n53446 = ~n53437 & ~n53445 ;
  assign n53447 = ~n53421 & n53446 ;
  assign n53448 = ~n53436 & n53447 ;
  assign n53449 = \u0_L12_reg[5]/NET0131  & ~n53448 ;
  assign n53450 = ~\u0_L12_reg[5]/NET0131  & n53448 ;
  assign n53451 = ~n53449 & ~n53450 ;
  assign n53452 = decrypt_pad & ~\u0_uk_K_r12_reg[3]/NET0131  ;
  assign n53453 = ~decrypt_pad & ~\u0_uk_K_r12_reg[11]/NET0131  ;
  assign n53454 = ~n53452 & ~n53453 ;
  assign n53455 = \u0_R12_reg[8]/NET0131  & ~n53454 ;
  assign n53456 = ~\u0_R12_reg[8]/NET0131  & n53454 ;
  assign n53457 = ~n53455 & ~n53456 ;
  assign n53458 = decrypt_pad & ~\u0_uk_K_r12_reg[12]/NET0131  ;
  assign n53459 = ~decrypt_pad & ~\u0_uk_K_r12_reg[20]/NET0131  ;
  assign n53460 = ~n53458 & ~n53459 ;
  assign n53461 = \u0_R12_reg[7]/NET0131  & ~n53460 ;
  assign n53462 = ~\u0_R12_reg[7]/NET0131  & n53460 ;
  assign n53463 = ~n53461 & ~n53462 ;
  assign n53477 = decrypt_pad & ~\u0_uk_K_r12_reg[27]/NET0131  ;
  assign n53478 = ~decrypt_pad & ~\u0_uk_K_r12_reg[3]/NET0131  ;
  assign n53479 = ~n53477 & ~n53478 ;
  assign n53480 = \u0_R12_reg[5]/NET0131  & ~n53479 ;
  assign n53481 = ~\u0_R12_reg[5]/NET0131  & n53479 ;
  assign n53482 = ~n53480 & ~n53481 ;
  assign n53464 = decrypt_pad & ~\u0_uk_K_r12_reg[48]/NET0131  ;
  assign n53465 = ~decrypt_pad & ~\u0_uk_K_r12_reg[24]/NET0131  ;
  assign n53466 = ~n53464 & ~n53465 ;
  assign n53467 = \u0_R12_reg[4]/NET0131  & ~n53466 ;
  assign n53468 = ~\u0_R12_reg[4]/NET0131  & n53466 ;
  assign n53469 = ~n53467 & ~n53468 ;
  assign n53470 = decrypt_pad & ~\u0_uk_K_r12_reg[40]/NET0131  ;
  assign n53471 = ~decrypt_pad & ~\u0_uk_K_r12_reg[48]/NET0131  ;
  assign n53472 = ~n53470 & ~n53471 ;
  assign n53473 = \u0_R12_reg[9]/NET0131  & ~n53472 ;
  assign n53474 = ~\u0_R12_reg[9]/NET0131  & n53472 ;
  assign n53475 = ~n53473 & ~n53474 ;
  assign n53492 = ~n53469 & n53475 ;
  assign n53493 = ~n53482 & n53492 ;
  assign n53484 = decrypt_pad & ~\u0_uk_K_r12_reg[18]/NET0131  ;
  assign n53485 = ~decrypt_pad & ~\u0_uk_K_r12_reg[26]/NET0131  ;
  assign n53486 = ~n53484 & ~n53485 ;
  assign n53487 = \u0_R12_reg[6]/NET0131  & ~n53486 ;
  assign n53488 = ~\u0_R12_reg[6]/NET0131  & n53486 ;
  assign n53489 = ~n53487 & ~n53488 ;
  assign n53494 = n53469 & n53482 ;
  assign n53495 = n53469 & ~n53475 ;
  assign n53496 = ~n53494 & ~n53495 ;
  assign n53497 = n53489 & ~n53496 ;
  assign n53498 = ~n53493 & ~n53497 ;
  assign n53499 = ~n53463 & ~n53498 ;
  assign n53500 = ~n53475 & n53482 ;
  assign n53501 = ~n53493 & ~n53500 ;
  assign n53502 = ~n53489 & ~n53501 ;
  assign n53476 = n53469 & n53475 ;
  assign n53483 = n53476 & ~n53482 ;
  assign n53490 = n53483 & n53489 ;
  assign n53491 = n53463 & n53490 ;
  assign n53503 = ~n53463 & ~n53482 ;
  assign n53504 = n53475 & ~n53489 ;
  assign n53505 = n53503 & n53504 ;
  assign n53506 = n53482 & n53489 ;
  assign n53507 = n53492 & n53506 ;
  assign n53508 = ~n53505 & ~n53507 ;
  assign n53509 = ~n53491 & n53508 ;
  assign n53510 = ~n53502 & n53509 ;
  assign n53511 = ~n53499 & n53510 ;
  assign n53512 = ~n53457 & ~n53511 ;
  assign n53529 = ~n53469 & ~n53475 ;
  assign n53530 = ~n53490 & ~n53529 ;
  assign n53531 = n53457 & ~n53530 ;
  assign n53513 = ~n53482 & n53489 ;
  assign n53532 = n53492 & ~n53513 ;
  assign n53533 = ~n53531 & ~n53532 ;
  assign n53528 = n53482 & ~n53489 ;
  assign n53534 = ~n53463 & ~n53528 ;
  assign n53535 = ~n53533 & n53534 ;
  assign n53514 = ~n53475 & n53513 ;
  assign n53515 = ~n53469 & n53514 ;
  assign n53516 = ~n53489 & n53494 ;
  assign n53517 = ~n53515 & ~n53516 ;
  assign n53518 = n53463 & ~n53517 ;
  assign n53519 = ~n53482 & n53495 ;
  assign n53520 = n53476 & n53482 ;
  assign n53521 = ~n53519 & ~n53520 ;
  assign n53522 = ~n53489 & ~n53521 ;
  assign n53523 = ~n53469 & n53489 ;
  assign n53524 = n53463 & n53482 ;
  assign n53525 = ~n53523 & n53524 ;
  assign n53526 = ~n53522 & ~n53525 ;
  assign n53527 = n53457 & ~n53526 ;
  assign n53536 = ~n53518 & ~n53527 ;
  assign n53537 = ~n53535 & n53536 ;
  assign n53538 = ~n53512 & n53537 ;
  assign n53539 = \u0_L12_reg[2]/NET0131  & n53538 ;
  assign n53540 = ~\u0_L12_reg[2]/NET0131  & ~n53538 ;
  assign n53541 = ~n53539 & ~n53540 ;
  assign n53555 = ~n53028 & n53092 ;
  assign n53556 = ~n53060 & ~n53061 ;
  assign n53557 = ~n53084 & ~n53556 ;
  assign n53558 = ~n53555 & ~n53557 ;
  assign n53559 = ~n53016 & ~n53558 ;
  assign n53542 = ~n53047 & n53050 ;
  assign n53560 = n53070 & n53349 ;
  assign n53561 = ~n53542 & n53560 ;
  assign n53562 = ~n53559 & ~n53561 ;
  assign n53563 = n53022 & ~n53562 ;
  assign n53543 = ~n53334 & ~n53542 ;
  assign n53544 = ~n53328 & n53543 ;
  assign n53545 = ~n53022 & ~n53544 ;
  assign n53546 = ~n53355 & ~n53545 ;
  assign n53547 = ~n53016 & ~n53546 ;
  assign n53550 = ~n53077 & n53083 ;
  assign n53548 = n53022 & n53334 ;
  assign n53549 = n53034 & n53342 ;
  assign n53551 = ~n53093 & ~n53549 ;
  assign n53552 = ~n53548 & n53551 ;
  assign n53553 = ~n53550 & n53552 ;
  assign n53554 = n53016 & ~n53553 ;
  assign n53565 = ~n53053 & ~n53330 ;
  assign n53564 = ~n53034 & n53041 ;
  assign n53566 = ~n53022 & ~n53564 ;
  assign n53567 = ~n53565 & n53566 ;
  assign n53568 = ~n53554 & ~n53567 ;
  assign n53569 = ~n53547 & n53568 ;
  assign n53570 = ~n53563 & n53569 ;
  assign n53571 = ~\u0_L12_reg[4]/NET0131  & ~n53570 ;
  assign n53572 = \u0_L12_reg[4]/NET0131  & n53570 ;
  assign n53573 = ~n53571 & ~n53572 ;
  assign n53578 = ~n53114 & n53139 ;
  assign n53579 = ~n53122 & ~n53578 ;
  assign n53580 = ~n53128 & ~n53579 ;
  assign n53574 = n53135 & ~n53137 ;
  assign n53575 = ~n53136 & ~n53165 ;
  assign n53576 = ~n53115 & n53575 ;
  assign n53577 = ~n53574 & ~n53576 ;
  assign n53581 = ~n53121 & n53181 ;
  assign n53582 = n53144 & n53145 ;
  assign n53583 = ~n53157 & ~n53582 ;
  assign n53584 = ~n53581 & n53583 ;
  assign n53585 = ~n53577 & n53584 ;
  assign n53586 = ~n53580 & n53585 ;
  assign n53593 = ~n53162 & ~n53182 ;
  assign n53594 = n53135 & ~n53593 ;
  assign n53587 = ~n53170 & ~n53172 ;
  assign n53588 = ~n53114 & ~n53587 ;
  assign n53589 = ~n53139 & ~n53144 ;
  assign n53590 = ~n53108 & n53135 ;
  assign n53591 = n53163 & ~n53590 ;
  assign n53592 = ~n53589 & n53591 ;
  assign n53595 = n53157 & ~n53187 ;
  assign n53596 = ~n53592 & n53595 ;
  assign n53597 = ~n53588 & n53596 ;
  assign n53598 = ~n53594 & n53597 ;
  assign n53599 = ~n53586 & ~n53598 ;
  assign n53600 = \u0_L12_reg[12]/NET0131  & n53599 ;
  assign n53601 = ~\u0_L12_reg[12]/NET0131  & ~n53599 ;
  assign n53602 = ~n53600 & ~n53601 ;
  assign n53610 = n53256 & ~n53263 ;
  assign n53611 = ~n53237 & n53243 ;
  assign n53612 = n53610 & ~n53611 ;
  assign n53613 = ~n53285 & ~n53612 ;
  assign n53614 = ~n53249 & ~n53613 ;
  assign n53603 = n53237 & ~n53243 ;
  assign n53604 = ~n53256 & n53603 ;
  assign n53605 = n53263 & n53604 ;
  assign n53606 = ~n53280 & ~n53605 ;
  assign n53607 = n53263 & n53303 ;
  assign n53608 = ~n53306 & ~n53607 ;
  assign n53609 = n53249 & ~n53608 ;
  assign n53615 = n53606 & ~n53609 ;
  assign n53616 = ~n53614 & n53615 ;
  assign n53617 = n53297 & ~n53616 ;
  assign n53621 = ~n53237 & n53290 ;
  assign n53618 = ~n53270 & ~n53603 ;
  assign n53619 = n53249 & n53256 ;
  assign n53620 = ~n53618 & n53619 ;
  assign n53624 = ~n53288 & ~n53620 ;
  assign n53625 = ~n53621 & n53624 ;
  assign n53622 = ~n53268 & ~n53611 ;
  assign n53623 = n53256 & ~n53622 ;
  assign n53626 = n53308 & ~n53623 ;
  assign n53627 = n53625 & n53626 ;
  assign n53628 = ~n53297 & ~n53627 ;
  assign n53629 = ~n53272 & n53606 ;
  assign n53630 = ~n53249 & ~n53629 ;
  assign n53631 = ~n53265 & ~n53315 ;
  assign n53632 = ~n53630 & n53631 ;
  assign n53633 = ~n53628 & n53632 ;
  assign n53634 = ~n53617 & n53633 ;
  assign n53635 = ~\u0_L12_reg[10]/NET0131  & ~n53634 ;
  assign n53636 = \u0_L12_reg[10]/NET0131  & n53634 ;
  assign n53637 = ~n53635 & ~n53636 ;
  assign n53642 = ~n53463 & ~n53483 ;
  assign n53643 = ~n53514 & n53642 ;
  assign n53646 = n53475 & n53523 ;
  assign n53644 = ~n53482 & ~n53489 ;
  assign n53645 = ~n53475 & n53644 ;
  assign n53647 = n53463 & ~n53645 ;
  assign n53648 = ~n53646 & n53647 ;
  assign n53649 = ~n53643 & ~n53648 ;
  assign n53640 = n53482 & n53529 ;
  assign n53641 = ~n53489 & n53640 ;
  assign n53650 = n53457 & n53508 ;
  assign n53651 = ~n53641 & n53650 ;
  assign n53652 = ~n53649 & n53651 ;
  assign n53656 = ~n53469 & ~n53503 ;
  assign n53657 = n53504 & n53656 ;
  assign n53653 = n53463 & n53469 ;
  assign n53654 = n53489 & ~n53500 ;
  assign n53655 = n53653 & n53654 ;
  assign n53658 = ~n53457 & ~n53655 ;
  assign n53659 = ~n53657 & n53658 ;
  assign n53662 = ~n53463 & ~n53640 ;
  assign n53660 = n53492 & n53513 ;
  assign n53661 = n53495 & n53644 ;
  assign n53663 = ~n53660 & ~n53661 ;
  assign n53664 = n53662 & n53663 ;
  assign n53665 = n53659 & n53664 ;
  assign n53666 = ~n53652 & ~n53665 ;
  assign n53638 = n53495 & n53506 ;
  assign n53639 = n53475 & n53516 ;
  assign n53667 = ~n53638 & ~n53639 ;
  assign n53668 = ~n53666 & n53667 ;
  assign n53671 = ~n53476 & ~n53529 ;
  assign n53672 = ~n53482 & ~n53671 ;
  assign n53669 = ~n53489 & n53495 ;
  assign n53670 = n53482 & n53669 ;
  assign n53673 = n53463 & ~n53670 ;
  assign n53674 = ~n53672 & n53673 ;
  assign n53675 = n53659 & n53674 ;
  assign n53676 = ~n53668 & ~n53675 ;
  assign n53677 = ~\u0_L12_reg[13]/NET0131  & ~n53676 ;
  assign n53678 = \u0_L12_reg[13]/NET0131  & n53676 ;
  assign n53679 = ~n53677 & ~n53678 ;
  assign n53680 = decrypt_pad & ~\u0_uk_K_r12_reg[44]/P0001  ;
  assign n53681 = ~decrypt_pad & ~\u0_uk_K_r12_reg[50]/NET0131  ;
  assign n53682 = ~n53680 & ~n53681 ;
  assign n53683 = \u0_R12_reg[20]/NET0131  & ~n53682 ;
  assign n53684 = ~\u0_R12_reg[20]/NET0131  & n53682 ;
  assign n53685 = ~n53683 & ~n53684 ;
  assign n53705 = decrypt_pad & ~\u0_uk_K_r12_reg[42]/NET0131  ;
  assign n53706 = ~decrypt_pad & ~\u0_uk_K_r12_reg[52]/NET0131  ;
  assign n53707 = ~n53705 & ~n53706 ;
  assign n53708 = \u0_R12_reg[18]/NET0131  & ~n53707 ;
  assign n53709 = ~\u0_R12_reg[18]/NET0131  & n53707 ;
  assign n53710 = ~n53708 & ~n53709 ;
  assign n53712 = decrypt_pad & ~\u0_uk_K_r12_reg[52]/NET0131  ;
  assign n53713 = ~decrypt_pad & ~\u0_uk_K_r12_reg[30]/NET0131  ;
  assign n53714 = ~n53712 & ~n53713 ;
  assign n53715 = \u0_R12_reg[17]/NET0131  & ~n53714 ;
  assign n53716 = ~\u0_R12_reg[17]/NET0131  & n53714 ;
  assign n53717 = ~n53715 & ~n53716 ;
  assign n53718 = ~n53710 & n53717 ;
  assign n53692 = decrypt_pad & ~\u0_uk_K_r12_reg[2]/NET0131  ;
  assign n53693 = ~decrypt_pad & ~\u0_uk_K_r12_reg[8]/NET0131  ;
  assign n53694 = ~n53692 & ~n53693 ;
  assign n53695 = \u0_R12_reg[16]/NET0131  & ~n53694 ;
  assign n53696 = ~\u0_R12_reg[16]/NET0131  & n53694 ;
  assign n53697 = ~n53695 & ~n53696 ;
  assign n53745 = n53697 & ~n53717 ;
  assign n53746 = ~n53718 & ~n53745 ;
  assign n53698 = decrypt_pad & ~\u0_uk_K_r12_reg[14]/NET0131  ;
  assign n53699 = ~decrypt_pad & ~\u0_uk_K_r12_reg[51]/NET0131  ;
  assign n53700 = ~n53698 & ~n53699 ;
  assign n53701 = \u0_R12_reg[21]/NET0131  & ~n53700 ;
  assign n53702 = ~\u0_R12_reg[21]/NET0131  & n53700 ;
  assign n53703 = ~n53701 & ~n53702 ;
  assign n53726 = n53697 & ~n53703 ;
  assign n53747 = n53703 & ~n53710 ;
  assign n53748 = ~n53726 & ~n53747 ;
  assign n53749 = ~n53746 & n53748 ;
  assign n53704 = n53697 & n53703 ;
  assign n53750 = n53704 & n53717 ;
  assign n53751 = ~n53710 & n53750 ;
  assign n53686 = decrypt_pad & ~\u0_uk_K_r12_reg[29]/NET0131  ;
  assign n53687 = ~decrypt_pad & ~\u0_uk_K_r12_reg[35]/NET0131  ;
  assign n53688 = ~n53686 & ~n53687 ;
  assign n53689 = \u0_R12_reg[19]/NET0131  & ~n53688 ;
  assign n53690 = ~\u0_R12_reg[19]/NET0131  & n53688 ;
  assign n53691 = ~n53689 & ~n53690 ;
  assign n53752 = ~n53710 & ~n53717 ;
  assign n53753 = n53726 & n53752 ;
  assign n53756 = ~n53691 & ~n53753 ;
  assign n53721 = ~n53703 & n53717 ;
  assign n53754 = n53710 & n53721 ;
  assign n53731 = ~n53697 & ~n53717 ;
  assign n53755 = n53703 & n53731 ;
  assign n53757 = ~n53754 & ~n53755 ;
  assign n53758 = n53756 & n53757 ;
  assign n53759 = ~n53751 & n53758 ;
  assign n53732 = ~n53703 & n53731 ;
  assign n53762 = n53691 & ~n53732 ;
  assign n53760 = n53704 & n53710 ;
  assign n53761 = ~n53697 & n53718 ;
  assign n53763 = ~n53760 & ~n53761 ;
  assign n53764 = n53762 & n53763 ;
  assign n53765 = ~n53759 & ~n53764 ;
  assign n53766 = ~n53749 & ~n53765 ;
  assign n53767 = ~n53685 & ~n53766 ;
  assign n53722 = n53697 & n53721 ;
  assign n53711 = n53704 & ~n53710 ;
  assign n53719 = ~n53697 & n53703 ;
  assign n53720 = ~n53718 & n53719 ;
  assign n53723 = ~n53711 & ~n53720 ;
  assign n53724 = ~n53722 & n53723 ;
  assign n53725 = n53691 & ~n53724 ;
  assign n53730 = ~n53691 & ~n53710 ;
  assign n53733 = n53717 & n53719 ;
  assign n53734 = ~n53732 & ~n53733 ;
  assign n53735 = n53730 & ~n53734 ;
  assign n53736 = ~n53691 & n53710 ;
  assign n53737 = n53717 & ~n53736 ;
  assign n53727 = n53710 & ~n53717 ;
  assign n53738 = n53704 & ~n53727 ;
  assign n53739 = ~n53737 & n53738 ;
  assign n53728 = n53726 & n53727 ;
  assign n53729 = n53718 & n53726 ;
  assign n53740 = ~n53728 & ~n53729 ;
  assign n53741 = ~n53739 & n53740 ;
  assign n53742 = ~n53735 & n53741 ;
  assign n53743 = ~n53725 & n53742 ;
  assign n53744 = n53685 & ~n53743 ;
  assign n53768 = ~n53697 & n53721 ;
  assign n53769 = ~n53755 & ~n53768 ;
  assign n53770 = n53710 & ~n53769 ;
  assign n53771 = ~n53691 & ~n53770 ;
  assign n53772 = n53710 & n53732 ;
  assign n53773 = n53691 & ~n53729 ;
  assign n53774 = ~n53772 & n53773 ;
  assign n53775 = ~n53771 & ~n53774 ;
  assign n53776 = ~n53744 & ~n53775 ;
  assign n53777 = ~n53767 & n53776 ;
  assign n53778 = ~\u0_L12_reg[14]/NET0131  & ~n53777 ;
  assign n53779 = \u0_L12_reg[14]/NET0131  & n53777 ;
  assign n53780 = ~n53778 & ~n53779 ;
  assign n53782 = ~n53373 & n53422 ;
  assign n53783 = ~n53386 & ~n53399 ;
  assign n53784 = ~n53782 & n53783 ;
  assign n53785 = n53406 & ~n53784 ;
  assign n53781 = n53395 & n53408 ;
  assign n53786 = ~n53367 & ~n53781 ;
  assign n53787 = ~n53785 & n53786 ;
  assign n53792 = n53373 & ~n53406 ;
  assign n53793 = n53412 & n53792 ;
  assign n53788 = ~n53373 & n53386 ;
  assign n53794 = n53367 & ~n53788 ;
  assign n53795 = ~n53793 & n53794 ;
  assign n53790 = ~n53379 & n53395 ;
  assign n53791 = n53406 & n53790 ;
  assign n53789 = n53392 & n53429 ;
  assign n53796 = ~n53438 & ~n53789 ;
  assign n53797 = ~n53791 & n53796 ;
  assign n53798 = n53795 & n53797 ;
  assign n53799 = ~n53787 & ~n53798 ;
  assign n53800 = ~n53373 & n53385 ;
  assign n53801 = n53398 & n53800 ;
  assign n53802 = n53430 & ~n53801 ;
  assign n53803 = n53440 & n53802 ;
  assign n53804 = n53392 & n53427 ;
  assign n53805 = n53406 & ~n53434 ;
  assign n53806 = ~n53804 & n53805 ;
  assign n53807 = ~n53803 & ~n53806 ;
  assign n53808 = ~n53367 & ~n53406 ;
  assign n53809 = n53428 & n53808 ;
  assign n53810 = ~n53807 & ~n53809 ;
  assign n53811 = ~n53799 & n53810 ;
  assign n53812 = \u0_L12_reg[15]/P0001  & n53811 ;
  assign n53813 = ~\u0_L12_reg[15]/P0001  & ~n53811 ;
  assign n53814 = ~n53812 & ~n53813 ;
  assign n53828 = ~n53237 & ~n53263 ;
  assign n53829 = ~n53309 & ~n53828 ;
  assign n53830 = n53256 & ~n53829 ;
  assign n53831 = ~n53249 & ~n53830 ;
  assign n53832 = ~n53256 & n53828 ;
  assign n53833 = n53249 & ~n53832 ;
  assign n53834 = ~n53275 & n53833 ;
  assign n53835 = ~n53831 & ~n53834 ;
  assign n53836 = ~n53283 & ~n53610 ;
  assign n53837 = n53611 & ~n53836 ;
  assign n53838 = ~n53280 & ~n53837 ;
  assign n53839 = ~n53835 & n53838 ;
  assign n53840 = ~n53297 & ~n53839 ;
  assign n53822 = ~n53610 & n53611 ;
  assign n53823 = ~n53284 & ~n53822 ;
  assign n53824 = ~n53249 & ~n53823 ;
  assign n53817 = n53243 & n53310 ;
  assign n53825 = ~n53604 & ~n53817 ;
  assign n53826 = ~n53824 & n53825 ;
  assign n53827 = n53297 & ~n53826 ;
  assign n53815 = ~n53307 & n53606 ;
  assign n53816 = n53249 & ~n53815 ;
  assign n53819 = ~n53303 & ~n53309 ;
  assign n53820 = n53249 & n53297 ;
  assign n53821 = ~n53819 & n53820 ;
  assign n53818 = ~n53249 & n53817 ;
  assign n53841 = ~n53289 & ~n53818 ;
  assign n53842 = ~n53821 & n53841 ;
  assign n53843 = ~n53816 & n53842 ;
  assign n53844 = ~n53827 & n53843 ;
  assign n53845 = ~n53840 & n53844 ;
  assign n53846 = ~\u0_L12_reg[1]/NET0131  & ~n53845 ;
  assign n53847 = \u0_L12_reg[1]/NET0131  & n53845 ;
  assign n53848 = ~n53846 & ~n53847 ;
  assign n53873 = n53373 & n53386 ;
  assign n53871 = n53392 & n53426 ;
  assign n53872 = n53385 & n53398 ;
  assign n53874 = ~n53871 & ~n53872 ;
  assign n53875 = ~n53873 & n53874 ;
  assign n53876 = n53406 & ~n53875 ;
  assign n53867 = ~n53410 & ~n53789 ;
  assign n53868 = ~n53406 & ~n53867 ;
  assign n53852 = n53379 & n53422 ;
  assign n53869 = ~n53790 & ~n53852 ;
  assign n53870 = n53373 & ~n53869 ;
  assign n53877 = ~n53804 & ~n53870 ;
  assign n53878 = ~n53868 & n53877 ;
  assign n53879 = ~n53876 & n53878 ;
  assign n53880 = n53367 & ~n53879 ;
  assign n53850 = ~n53379 & ~n53406 ;
  assign n53851 = n53422 & n53850 ;
  assign n53858 = ~n53433 & ~n53851 ;
  assign n53859 = ~n53397 & n53858 ;
  assign n53849 = n53392 & n53409 ;
  assign n53860 = ~n53439 & ~n53849 ;
  assign n53861 = n53859 & n53860 ;
  assign n53853 = ~n53429 & ~n53852 ;
  assign n53854 = n53406 & ~n53853 ;
  assign n53855 = ~n53379 & n53792 ;
  assign n53856 = ~n53788 & ~n53855 ;
  assign n53857 = n53392 & ~n53856 ;
  assign n53862 = ~n53854 & ~n53857 ;
  assign n53863 = n53861 & n53862 ;
  assign n53864 = ~n53367 & ~n53863 ;
  assign n53865 = n53406 & n53427 ;
  assign n53866 = n53385 & n53849 ;
  assign n53881 = ~n53865 & ~n53866 ;
  assign n53882 = ~n53864 & n53881 ;
  assign n53883 = ~n53880 & n53882 ;
  assign n53884 = ~\u0_L12_reg[21]/NET0131  & ~n53883 ;
  assign n53885 = \u0_L12_reg[21]/NET0131  & n53883 ;
  assign n53886 = ~n53884 & ~n53885 ;
  assign n53888 = ~n53697 & n53710 ;
  assign n53889 = ~n53752 & ~n53888 ;
  assign n53890 = ~n53703 & ~n53889 ;
  assign n53891 = ~n53731 & ~n53750 ;
  assign n53892 = ~n53890 & n53891 ;
  assign n53893 = n53691 & ~n53892 ;
  assign n53894 = n53703 & n53745 ;
  assign n53895 = ~n53761 & ~n53894 ;
  assign n53896 = ~n53691 & ~n53895 ;
  assign n53887 = n53717 & n53747 ;
  assign n53897 = n53710 & n53722 ;
  assign n53898 = ~n53887 & ~n53897 ;
  assign n53899 = ~n53896 & n53898 ;
  assign n53900 = ~n53893 & n53899 ;
  assign n53901 = n53685 & ~n53900 ;
  assign n53913 = ~n53772 & ~n53897 ;
  assign n53914 = ~n53697 & n53747 ;
  assign n53915 = ~n53717 & n53914 ;
  assign n53916 = n53913 & ~n53915 ;
  assign n53917 = n53691 & ~n53916 ;
  assign n53903 = n53717 & ~n53888 ;
  assign n53902 = ~n53717 & ~n53726 ;
  assign n53904 = n53691 & ~n53703 ;
  assign n53905 = ~n53902 & ~n53904 ;
  assign n53906 = ~n53903 & n53905 ;
  assign n53908 = n53691 & ~n53721 ;
  assign n53907 = ~n53691 & ~n53731 ;
  assign n53909 = ~n53710 & ~n53907 ;
  assign n53910 = ~n53908 & n53909 ;
  assign n53911 = ~n53906 & ~n53910 ;
  assign n53912 = ~n53685 & ~n53911 ;
  assign n53918 = n53736 & n53745 ;
  assign n53919 = ~n53751 & ~n53918 ;
  assign n53920 = ~n53912 & n53919 ;
  assign n53921 = ~n53917 & n53920 ;
  assign n53922 = ~n53901 & n53921 ;
  assign n53923 = ~\u0_L12_reg[25]/NET0131  & ~n53922 ;
  assign n53924 = \u0_L12_reg[25]/NET0131  & n53922 ;
  assign n53925 = ~n53923 & ~n53924 ;
  assign n53926 = n53266 & n53828 ;
  assign n53932 = n53297 & ~n53926 ;
  assign n53933 = ~n53313 & n53932 ;
  assign n53934 = ~n53817 & n53933 ;
  assign n53927 = n53271 & n53309 ;
  assign n53928 = ~n53279 & ~n53927 ;
  assign n53929 = ~n53249 & ~n53928 ;
  assign n53930 = ~n53284 & ~n53290 ;
  assign n53931 = n53237 & ~n53930 ;
  assign n53935 = ~n53929 & ~n53931 ;
  assign n53936 = n53934 & n53935 ;
  assign n53937 = ~n53283 & n53314 ;
  assign n53938 = ~n53297 & ~n53303 ;
  assign n53939 = ~n53937 & n53938 ;
  assign n53940 = n53286 & n53939 ;
  assign n53941 = ~n53936 & ~n53940 ;
  assign n53944 = n53243 & n53836 ;
  assign n53945 = ~n53274 & ~n53944 ;
  assign n53946 = ~n53237 & ~n53945 ;
  assign n53942 = ~n53270 & ~n53604 ;
  assign n53943 = ~n53297 & ~n53942 ;
  assign n53947 = ~n53249 & ~n53943 ;
  assign n53948 = ~n53946 & n53947 ;
  assign n53949 = n53249 & ~n53285 ;
  assign n53950 = ~n53607 & n53949 ;
  assign n53951 = ~n53948 & ~n53950 ;
  assign n53952 = ~n53941 & ~n53951 ;
  assign n53953 = ~\u0_L12_reg[26]/NET0131  & ~n53952 ;
  assign n53954 = \u0_L12_reg[26]/NET0131  & n53952 ;
  assign n53955 = ~n53953 & ~n53954 ;
  assign n53956 = ~n53745 & ~n53752 ;
  assign n53957 = n53691 & ~n53719 ;
  assign n53958 = ~n53726 & n53957 ;
  assign n53959 = ~n53956 & n53958 ;
  assign n53960 = n53697 & n53730 ;
  assign n53961 = n53685 & ~n53960 ;
  assign n53962 = ~n53770 & n53961 ;
  assign n53963 = ~n53959 & n53962 ;
  assign n53964 = n53691 & ~n53753 ;
  assign n53965 = ~n53750 & n53964 ;
  assign n53966 = n53719 & ~n53727 ;
  assign n53967 = ~n53691 & ~n53894 ;
  assign n53968 = ~n53966 & n53967 ;
  assign n53969 = ~n53965 & ~n53968 ;
  assign n53970 = ~n53685 & ~n53761 ;
  assign n53971 = n53913 & n53970 ;
  assign n53972 = ~n53969 & n53971 ;
  assign n53973 = ~n53963 & ~n53972 ;
  assign n53974 = ~n53691 & n53728 ;
  assign n53976 = n53718 & n53719 ;
  assign n53975 = n53719 & n53727 ;
  assign n53977 = ~n53754 & ~n53975 ;
  assign n53978 = ~n53976 & n53977 ;
  assign n53979 = n53691 & ~n53978 ;
  assign n53980 = ~n53974 & ~n53979 ;
  assign n53981 = ~n53973 & n53980 ;
  assign n53982 = ~\u0_L12_reg[8]/NET0131  & ~n53981 ;
  assign n53983 = \u0_L12_reg[8]/NET0131  & n53981 ;
  assign n53984 = ~n53982 & ~n53983 ;
  assign n54002 = ~n52922 & ~n53220 ;
  assign n54003 = n52922 & n52928 ;
  assign n54004 = n52977 & n54003 ;
  assign n54005 = ~n54002 & ~n54004 ;
  assign n54006 = n52975 & ~n54005 ;
  assign n54001 = n53001 & n53209 ;
  assign n54007 = ~n52980 & ~n53198 ;
  assign n54008 = ~n54001 & n54007 ;
  assign n54009 = ~n54006 & n54008 ;
  assign n54010 = ~n52935 & ~n54009 ;
  assign n53986 = ~n52962 & ~n53210 ;
  assign n53987 = n52935 & ~n53986 ;
  assign n53988 = ~n52966 & n52975 ;
  assign n53989 = ~n52978 & n53988 ;
  assign n53990 = ~n53987 & n53989 ;
  assign n53995 = ~n52975 & ~n52991 ;
  assign n53996 = ~n53199 & n53995 ;
  assign n53994 = n52935 & n53212 ;
  assign n53991 = ~n52935 & ~n52977 ;
  assign n53992 = n52922 & ~n53001 ;
  assign n53993 = n53991 & n53992 ;
  assign n53997 = ~n52943 & ~n53993 ;
  assign n53998 = ~n53994 & n53997 ;
  assign n53999 = n53996 & n53998 ;
  assign n54000 = ~n53990 & ~n53999 ;
  assign n53985 = n52994 & n53212 ;
  assign n54011 = ~n53003 & ~n53985 ;
  assign n54012 = ~n54000 & n54011 ;
  assign n54013 = ~n54010 & n54012 ;
  assign n54014 = \u0_L12_reg[23]/NET0131  & ~n54013 ;
  assign n54015 = ~\u0_L12_reg[23]/NET0131  & n54013 ;
  assign n54016 = ~n54014 & ~n54015 ;
  assign n54017 = ~n53022 & ~n53069 ;
  assign n54018 = n53028 & n53564 ;
  assign n54019 = n53022 & ~n54018 ;
  assign n54020 = ~n54017 & ~n54019 ;
  assign n54021 = ~n53041 & ~n53061 ;
  assign n54022 = ~n53068 & n54021 ;
  assign n54023 = n53034 & ~n53088 ;
  assign n54024 = ~n54022 & n54023 ;
  assign n54025 = ~n53034 & ~n53061 ;
  assign n54026 = ~n53087 & n54025 ;
  assign n54027 = ~n54024 & ~n54026 ;
  assign n54028 = ~n54020 & ~n54027 ;
  assign n54029 = n53016 & ~n54028 ;
  assign n54033 = n54019 & ~n54021 ;
  assign n54034 = n53041 & n53549 ;
  assign n54035 = ~n54033 & ~n54034 ;
  assign n54036 = ~n53016 & ~n54035 ;
  assign n54030 = ~n53016 & n54022 ;
  assign n54031 = ~n53049 & ~n54030 ;
  assign n54032 = ~n53022 & ~n54031 ;
  assign n54037 = ~n53091 & ~n54032 ;
  assign n54038 = ~n54036 & n54037 ;
  assign n54039 = ~n54029 & n54038 ;
  assign n54040 = ~\u0_L12_reg[19]/P0001  & ~n54039 ;
  assign n54041 = \u0_L12_reg[19]/P0001  & n54039 ;
  assign n54042 = ~n54040 & ~n54041 ;
  assign n54061 = n53489 & n53640 ;
  assign n54062 = n53521 & ~n54061 ;
  assign n54063 = n53463 & ~n54062 ;
  assign n54046 = ~n53489 & n53529 ;
  assign n54047 = n53482 & n53492 ;
  assign n54048 = ~n54046 & ~n54047 ;
  assign n54060 = ~n53463 & ~n54048 ;
  assign n54058 = ~n53483 & ~n53653 ;
  assign n54059 = ~n53489 & ~n54058 ;
  assign n54064 = ~n53660 & ~n54059 ;
  assign n54065 = ~n54060 & n54064 ;
  assign n54066 = ~n54063 & n54065 ;
  assign n54067 = n53457 & ~n54066 ;
  assign n54043 = ~n53482 & n53523 ;
  assign n54044 = ~n53638 & ~n54043 ;
  assign n54045 = ~n53463 & ~n54044 ;
  assign n54049 = n53463 & n54048 ;
  assign n54050 = ~n53463 & ~n53494 ;
  assign n54051 = ~n53493 & n54050 ;
  assign n54052 = ~n53669 & n54051 ;
  assign n54053 = ~n54049 & ~n54052 ;
  assign n54054 = n53513 & ~n53671 ;
  assign n54055 = ~n53638 & ~n54054 ;
  assign n54056 = ~n54053 & n54055 ;
  assign n54057 = ~n53457 & ~n54056 ;
  assign n54068 = ~n54045 & ~n54057 ;
  assign n54069 = ~n54067 & n54068 ;
  assign n54070 = ~\u0_L12_reg[28]/NET0131  & ~n54069 ;
  assign n54071 = \u0_L12_reg[28]/NET0131  & n54069 ;
  assign n54072 = ~n54070 & ~n54071 ;
  assign n54089 = ~n53379 & n53782 ;
  assign n54090 = ~n53393 & ~n54089 ;
  assign n54091 = n53406 & ~n54090 ;
  assign n54086 = ~n53427 & ~n53852 ;
  assign n54087 = ~n53872 & n54086 ;
  assign n54088 = ~n53406 & ~n54087 ;
  assign n54092 = ~n53397 & ~n53871 ;
  assign n54093 = ~n53434 & n54092 ;
  assign n54094 = ~n54088 & n54093 ;
  assign n54095 = ~n54091 & n54094 ;
  assign n54096 = n53367 & ~n54095 ;
  assign n54074 = n53406 & ~n53433 ;
  assign n54073 = n53392 & ~n53800 ;
  assign n54075 = ~n53782 & ~n54073 ;
  assign n54076 = n54074 & n54075 ;
  assign n54077 = n53379 & n53392 ;
  assign n54078 = n53792 & n54077 ;
  assign n54079 = ~n53851 & ~n54078 ;
  assign n54080 = ~n53442 & n54079 ;
  assign n54081 = ~n54076 & n54080 ;
  assign n54082 = ~n53367 & ~n54081 ;
  assign n54083 = ~n53438 & ~n53441 ;
  assign n54084 = ~n53406 & ~n54083 ;
  assign n54085 = n53396 & n53406 ;
  assign n54097 = ~n53437 & ~n54085 ;
  assign n54098 = ~n54084 & n54097 ;
  assign n54099 = ~n54082 & n54098 ;
  assign n54100 = ~n54096 & n54099 ;
  assign n54101 = \u0_L12_reg[27]/NET0131  & n54100 ;
  assign n54102 = ~\u0_L12_reg[27]/NET0131  & ~n54100 ;
  assign n54103 = ~n54101 & ~n54102 ;
  assign n54120 = ~n53114 & ~n53128 ;
  assign n54122 = n53575 & ~n54120 ;
  assign n54123 = n53589 & ~n54122 ;
  assign n54121 = ~n53589 & ~n54120 ;
  assign n54124 = n53157 & ~n54121 ;
  assign n54125 = ~n54123 & n54124 ;
  assign n54126 = n53108 & n53166 ;
  assign n54127 = ~n53186 & ~n54126 ;
  assign n54128 = ~n54125 & n54127 ;
  assign n54129 = ~n53135 & ~n54128 ;
  assign n54104 = ~n53575 & ~n53578 ;
  assign n54105 = ~n53135 & ~n54104 ;
  assign n54106 = n53135 & ~n53170 ;
  assign n54107 = ~n53578 & n54106 ;
  assign n54108 = ~n54105 & ~n54107 ;
  assign n54109 = n53128 & ~n53579 ;
  assign n54110 = n53188 & ~n54109 ;
  assign n54111 = ~n54108 & n54110 ;
  assign n54112 = ~n53157 & ~n54111 ;
  assign n54113 = n53135 & n53164 ;
  assign n54114 = n53114 & n53139 ;
  assign n54115 = ~n53161 & ~n53166 ;
  assign n54116 = ~n54114 & n54115 ;
  assign n54117 = ~n53148 & n53157 ;
  assign n54118 = ~n53184 & n54117 ;
  assign n54119 = ~n54116 & n54118 ;
  assign n54130 = ~n54113 & ~n54119 ;
  assign n54131 = ~n54112 & n54130 ;
  assign n54132 = ~n54129 & n54131 ;
  assign n54133 = \u0_L12_reg[32]/NET0131  & n54132 ;
  assign n54134 = ~\u0_L12_reg[32]/NET0131  & ~n54132 ;
  assign n54135 = ~n54133 & ~n54134 ;
  assign n54137 = n53685 & ~n53728 ;
  assign n54138 = ~n53733 & ~n53751 ;
  assign n54139 = n54137 & n54138 ;
  assign n54140 = ~n53726 & n53727 ;
  assign n54141 = ~n53685 & ~n54140 ;
  assign n54142 = ~n53748 & ~n53894 ;
  assign n54143 = n54141 & n54142 ;
  assign n54144 = ~n54139 & ~n54143 ;
  assign n54136 = n53748 & ~n53956 ;
  assign n54145 = ~n53691 & ~n53729 ;
  assign n54146 = ~n54136 & n54145 ;
  assign n54147 = ~n54144 & n54146 ;
  assign n54148 = ~n53722 & ~n53914 ;
  assign n54149 = n54141 & n54148 ;
  assign n54150 = ~n53711 & ~n53768 ;
  assign n54151 = n54137 & n54150 ;
  assign n54152 = ~n54149 & ~n54151 ;
  assign n54153 = n53964 & ~n53975 ;
  assign n54154 = ~n54152 & n54153 ;
  assign n54155 = ~n54147 & ~n54154 ;
  assign n54156 = ~\u0_L12_reg[3]/NET0131  & n54155 ;
  assign n54157 = \u0_L12_reg[3]/NET0131  & ~n54155 ;
  assign n54158 = ~n54156 & ~n54157 ;
  assign n54159 = decrypt_pad & ~\u0_uk_K_r12_reg[13]/NET0131  ;
  assign n54160 = ~decrypt_pad & ~\u0_uk_K_r12_reg[46]/NET0131  ;
  assign n54161 = ~n54159 & ~n54160 ;
  assign n54162 = \u0_R12_reg[12]/NET0131  & ~n54161 ;
  assign n54163 = ~\u0_R12_reg[12]/NET0131  & n54161 ;
  assign n54164 = ~n54162 & ~n54163 ;
  assign n54165 = decrypt_pad & ~\u0_uk_K_r12_reg[46]/NET0131  ;
  assign n54166 = ~decrypt_pad & ~\u0_uk_K_r12_reg[54]/NET0131  ;
  assign n54167 = ~n54165 & ~n54166 ;
  assign n54168 = \u0_R12_reg[9]/NET0131  & ~n54167 ;
  assign n54169 = ~\u0_R12_reg[9]/NET0131  & n54167 ;
  assign n54170 = ~n54168 & ~n54169 ;
  assign n54171 = decrypt_pad & ~\u0_uk_K_r12_reg[54]/NET0131  ;
  assign n54172 = ~decrypt_pad & ~\u0_uk_K_r12_reg[5]/NET0131  ;
  assign n54173 = ~n54171 & ~n54172 ;
  assign n54174 = \u0_R12_reg[10]/NET0131  & ~n54173 ;
  assign n54175 = ~\u0_R12_reg[10]/NET0131  & n54173 ;
  assign n54176 = ~n54174 & ~n54175 ;
  assign n54177 = n54170 & n54176 ;
  assign n54178 = decrypt_pad & ~\u0_uk_K_r12_reg[17]/NET0131  ;
  assign n54179 = ~decrypt_pad & ~\u0_uk_K_r12_reg[25]/NET0131  ;
  assign n54180 = ~n54178 & ~n54179 ;
  assign n54181 = \u0_R12_reg[8]/NET0131  & ~n54180 ;
  assign n54182 = ~\u0_R12_reg[8]/NET0131  & n54180 ;
  assign n54183 = ~n54181 & ~n54182 ;
  assign n54184 = decrypt_pad & ~\u0_uk_K_r12_reg[55]/NET0131  ;
  assign n54185 = ~decrypt_pad & ~\u0_uk_K_r12_reg[6]/NET0131  ;
  assign n54186 = ~n54184 & ~n54185 ;
  assign n54187 = \u0_R12_reg[11]/NET0131  & ~n54186 ;
  assign n54188 = ~\u0_R12_reg[11]/NET0131  & n54186 ;
  assign n54189 = ~n54187 & ~n54188 ;
  assign n54190 = ~n54183 & n54189 ;
  assign n54191 = decrypt_pad & ~\u0_uk_K_r12_reg[26]/NET0131  ;
  assign n54192 = ~decrypt_pad & ~\u0_uk_K_r12_reg[34]/NET0131  ;
  assign n54193 = ~n54191 & ~n54192 ;
  assign n54194 = \u0_R12_reg[13]/NET0131  & ~n54193 ;
  assign n54195 = ~\u0_R12_reg[13]/NET0131  & n54193 ;
  assign n54196 = ~n54194 & ~n54195 ;
  assign n54197 = ~n54183 & n54196 ;
  assign n54198 = n54183 & ~n54196 ;
  assign n54199 = ~n54197 & ~n54198 ;
  assign n54200 = ~n54190 & ~n54199 ;
  assign n54201 = n54177 & n54200 ;
  assign n54202 = n54170 & ~n54176 ;
  assign n54203 = n54190 & n54202 ;
  assign n54208 = ~n54201 & ~n54203 ;
  assign n54204 = ~n54170 & ~n54176 ;
  assign n54205 = n54199 & ~n54204 ;
  assign n54206 = ~n54177 & n54205 ;
  assign n54207 = n54200 & n54204 ;
  assign n54209 = ~n54206 & ~n54207 ;
  assign n54210 = n54208 & n54209 ;
  assign n54211 = ~n54164 & ~n54210 ;
  assign n54215 = ~n54170 & n54196 ;
  assign n54227 = n54176 & n54197 ;
  assign n54228 = n54170 & n54198 ;
  assign n54229 = ~n54227 & ~n54228 ;
  assign n54230 = ~n54215 & n54229 ;
  assign n54231 = n54164 & n54189 ;
  assign n54232 = ~n54230 & n54231 ;
  assign n54216 = n54176 & n54215 ;
  assign n54212 = ~n54183 & ~n54196 ;
  assign n54217 = ~n54176 & n54212 ;
  assign n54218 = ~n54170 & n54217 ;
  assign n54219 = ~n54216 & ~n54218 ;
  assign n54220 = n54189 & ~n54219 ;
  assign n54213 = n54164 & n54177 ;
  assign n54214 = n54212 & n54213 ;
  assign n54222 = n54170 & ~n54196 ;
  assign n54223 = ~n54189 & ~n54222 ;
  assign n54221 = ~n54183 & ~n54202 ;
  assign n54224 = n54164 & ~n54215 ;
  assign n54225 = ~n54221 & n54224 ;
  assign n54226 = n54223 & n54225 ;
  assign n54233 = ~n54214 & ~n54226 ;
  assign n54234 = ~n54220 & n54233 ;
  assign n54235 = ~n54232 & n54234 ;
  assign n54236 = ~n54211 & n54235 ;
  assign n54237 = ~\u0_L12_reg[6]/NET0131  & ~n54236 ;
  assign n54238 = \u0_L12_reg[6]/NET0131  & n54236 ;
  assign n54239 = ~n54237 & ~n54238 ;
  assign n54242 = ~n53221 & ~n54002 ;
  assign n54243 = n52928 & ~n54242 ;
  assign n54240 = ~n52979 & n52994 ;
  assign n54241 = n53220 & n54240 ;
  assign n54244 = n52975 & ~n53198 ;
  assign n54245 = ~n54241 & n54244 ;
  assign n54246 = ~n54243 & n54245 ;
  assign n54249 = ~n53210 & n53991 ;
  assign n54250 = n52935 & ~n52957 ;
  assign n54251 = ~n52961 & n54250 ;
  assign n54252 = ~n53212 & n54251 ;
  assign n54253 = ~n54249 & ~n54252 ;
  assign n54247 = n52928 & n53217 ;
  assign n54248 = n52952 & n52963 ;
  assign n54254 = ~n52975 & ~n54248 ;
  assign n54255 = ~n54247 & n54254 ;
  assign n54256 = ~n54253 & n54255 ;
  assign n54257 = ~n54246 & ~n54256 ;
  assign n54258 = n52942 & n52990 ;
  assign n54259 = ~n52955 & n54258 ;
  assign n54260 = ~n54257 & ~n54259 ;
  assign n54261 = ~\u0_L12_reg[9]/NET0131  & ~n54260 ;
  assign n54262 = \u0_L12_reg[9]/NET0131  & n54260 ;
  assign n54263 = ~n54261 & ~n54262 ;
  assign n54265 = ~n53108 & ~n53163 ;
  assign n54266 = ~n53180 & n54265 ;
  assign n54264 = n53128 & ~n53589 ;
  assign n54267 = ~n54114 & ~n54264 ;
  assign n54268 = ~n54266 & n54267 ;
  assign n54269 = ~n53135 & ~n54268 ;
  assign n54272 = ~n53114 & n53589 ;
  assign n54273 = ~n53136 & n54272 ;
  assign n54274 = n53135 & n54273 ;
  assign n54270 = ~n53170 & ~n54264 ;
  assign n54271 = n53114 & ~n54270 ;
  assign n54275 = n53157 & ~n54271 ;
  assign n54276 = ~n54274 & n54275 ;
  assign n54277 = ~n54269 & n54276 ;
  assign n54278 = n53114 & n54264 ;
  assign n54279 = n54106 & ~n54272 ;
  assign n54280 = ~n54278 & n54279 ;
  assign n54281 = ~n53157 & ~n54280 ;
  assign n54282 = ~n54277 & ~n54281 ;
  assign n54283 = ~n53135 & n54271 ;
  assign n54284 = ~n53135 & n54273 ;
  assign n54285 = ~n53138 & ~n54284 ;
  assign n54286 = ~n53135 & n53157 ;
  assign n54287 = ~n54285 & ~n54286 ;
  assign n54288 = ~n54283 & ~n54287 ;
  assign n54289 = ~n54282 & n54288 ;
  assign n54290 = ~\u0_L12_reg[7]/NET0131  & ~n54289 ;
  assign n54291 = \u0_L12_reg[7]/NET0131  & n54289 ;
  assign n54292 = ~n54290 & ~n54291 ;
  assign n54294 = n54183 & n54196 ;
  assign n54295 = n54170 & n54294 ;
  assign n54296 = ~n54170 & ~n54294 ;
  assign n54297 = ~n54295 & ~n54296 ;
  assign n54298 = ~n54212 & ~n54297 ;
  assign n54299 = n54190 & n54222 ;
  assign n54300 = ~n54298 & ~n54299 ;
  assign n54301 = ~n54176 & ~n54300 ;
  assign n54302 = n54176 & n54212 ;
  assign n54303 = ~n54176 & n54198 ;
  assign n54304 = ~n54302 & ~n54303 ;
  assign n54305 = ~n54189 & ~n54304 ;
  assign n54293 = n54177 & n54197 ;
  assign n54306 = n54164 & ~n54293 ;
  assign n54307 = ~n54305 & n54306 ;
  assign n54308 = ~n54301 & n54307 ;
  assign n54311 = ~n54170 & ~n54183 ;
  assign n54312 = n54196 & n54311 ;
  assign n54313 = ~n54217 & ~n54295 ;
  assign n54314 = ~n54312 & n54313 ;
  assign n54315 = ~n54189 & ~n54314 ;
  assign n54309 = n54189 & ~n54212 ;
  assign n54310 = n54297 & n54309 ;
  assign n54316 = ~n54164 & ~n54218 ;
  assign n54317 = ~n54310 & n54316 ;
  assign n54318 = ~n54315 & n54317 ;
  assign n54319 = ~n54308 & ~n54318 ;
  assign n54320 = n54176 & n54183 ;
  assign n54321 = ~n54170 & n54320 ;
  assign n54322 = ~n54189 & n54321 ;
  assign n54323 = ~n54170 & n54302 ;
  assign n54324 = n54176 & n54228 ;
  assign n54325 = ~n54323 & ~n54324 ;
  assign n54326 = n54189 & ~n54325 ;
  assign n54327 = ~n54322 & ~n54326 ;
  assign n54328 = ~n54319 & n54327 ;
  assign n54329 = ~\u0_L12_reg[16]/NET0131  & ~n54328 ;
  assign n54330 = \u0_L12_reg[16]/NET0131  & n54328 ;
  assign n54331 = ~n54329 & ~n54330 ;
  assign n54342 = ~n54196 & n54321 ;
  assign n54343 = ~n54176 & n54197 ;
  assign n54344 = ~n54302 & ~n54343 ;
  assign n54345 = n54170 & n54212 ;
  assign n54346 = ~n54321 & ~n54345 ;
  assign n54347 = n54344 & n54346 ;
  assign n54348 = n54189 & ~n54347 ;
  assign n54349 = ~n54342 & ~n54348 ;
  assign n54350 = ~n54164 & ~n54349 ;
  assign n54332 = n54189 & ~n54197 ;
  assign n54333 = n54204 & n54332 ;
  assign n54338 = ~n54207 & ~n54333 ;
  assign n54334 = n54170 & n54320 ;
  assign n54335 = ~n54227 & ~n54334 ;
  assign n54336 = n54189 & ~n54335 ;
  assign n54337 = ~n54189 & n54205 ;
  assign n54339 = ~n54336 & ~n54337 ;
  assign n54340 = n54338 & n54339 ;
  assign n54341 = n54164 & ~n54340 ;
  assign n54357 = n54199 & n54204 ;
  assign n54358 = n54229 & ~n54357 ;
  assign n54359 = ~n54164 & ~n54189 ;
  assign n54360 = ~n54358 & n54359 ;
  assign n54351 = ~n54170 & n54303 ;
  assign n54352 = n54170 & n54343 ;
  assign n54353 = ~n54351 & ~n54352 ;
  assign n54354 = n54189 & ~n54353 ;
  assign n54355 = n54176 & ~n54189 ;
  assign n54356 = n54295 & n54355 ;
  assign n54361 = ~n54354 & ~n54356 ;
  assign n54362 = ~n54360 & n54361 ;
  assign n54363 = ~n54341 & n54362 ;
  assign n54364 = ~n54350 & n54363 ;
  assign n54365 = ~\u0_L12_reg[24]/NET0131  & ~n54364 ;
  assign n54366 = \u0_L12_reg[24]/NET0131  & n54364 ;
  assign n54367 = ~n54365 & ~n54366 ;
  assign n54369 = ~n54320 & ~n54345 ;
  assign n54370 = n54164 & ~n54369 ;
  assign n54371 = ~n54189 & ~n54370 ;
  assign n54372 = n54189 & n54344 ;
  assign n54373 = ~n54351 & n54372 ;
  assign n54374 = n54164 & ~n54373 ;
  assign n54375 = n54215 & n54320 ;
  assign n54376 = ~n54374 & ~n54375 ;
  assign n54377 = ~n54371 & ~n54376 ;
  assign n54378 = ~n54222 & n54320 ;
  assign n54379 = ~n54196 & n54202 ;
  assign n54380 = ~n54378 & ~n54379 ;
  assign n54381 = n54189 & ~n54380 ;
  assign n54384 = ~n54170 & n54227 ;
  assign n54382 = ~n54311 & ~n54320 ;
  assign n54383 = n54223 & n54382 ;
  assign n54385 = ~n54357 & ~n54383 ;
  assign n54386 = ~n54384 & n54385 ;
  assign n54387 = ~n54381 & n54386 ;
  assign n54388 = ~n54164 & ~n54387 ;
  assign n54368 = n54213 & ~n54294 ;
  assign n54389 = n54222 & n54355 ;
  assign n54390 = ~n54368 & ~n54389 ;
  assign n54391 = ~n54388 & n54390 ;
  assign n54392 = ~n54377 & n54391 ;
  assign n54393 = \u0_L12_reg[30]/NET0131  & ~n54392 ;
  assign n54394 = ~\u0_L12_reg[30]/NET0131  & n54392 ;
  assign n54395 = ~n54393 & ~n54394 ;
  assign n54397 = n53469 & n53504 ;
  assign n54398 = ~n53519 & ~n54397 ;
  assign n54399 = ~n53463 & ~n54398 ;
  assign n54396 = n53463 & ~n53501 ;
  assign n54400 = n53457 & ~n53515 ;
  assign n54401 = ~n54396 & n54400 ;
  assign n54402 = ~n54399 & n54401 ;
  assign n54404 = ~n53463 & n53506 ;
  assign n54405 = ~n53644 & ~n54404 ;
  assign n54406 = ~n53469 & ~n54405 ;
  assign n54407 = ~n53457 & ~n53638 ;
  assign n54408 = ~n53645 & n54407 ;
  assign n54403 = n53463 & n53520 ;
  assign n54409 = ~n53490 & ~n54403 ;
  assign n54410 = n54408 & n54409 ;
  assign n54411 = ~n54406 & n54410 ;
  assign n54412 = ~n54402 & ~n54411 ;
  assign n54413 = ~n53463 & n54047 ;
  assign n54414 = n53476 & n53489 ;
  assign n54415 = ~n53641 & ~n54414 ;
  assign n54416 = n53463 & ~n54415 ;
  assign n54417 = ~n54413 & ~n54416 ;
  assign n54418 = ~n54412 & n54417 ;
  assign n54419 = \u0_L12_reg[18]/NET0131  & n54418 ;
  assign n54420 = ~\u0_L12_reg[18]/NET0131  & ~n54418 ;
  assign n54421 = ~n54419 & ~n54420 ;
  assign n54422 = decrypt_pad & ~\u0_uk_K_r11_reg[22]/NET0131  ;
  assign n54423 = ~decrypt_pad & ~\u0_uk_K_r11_reg[0]/NET0131  ;
  assign n54424 = ~n54422 & ~n54423 ;
  assign n54425 = \u0_R11_reg[28]/NET0131  & ~n54424 ;
  assign n54426 = ~\u0_R11_reg[28]/NET0131  & n54424 ;
  assign n54427 = ~n54425 & ~n54426 ;
  assign n54428 = decrypt_pad & ~\u0_uk_K_r11_reg[2]/NET0131  ;
  assign n54429 = ~decrypt_pad & ~\u0_uk_K_r11_reg[35]/NET0131  ;
  assign n54430 = ~n54428 & ~n54429 ;
  assign n54431 = \u0_R11_reg[26]/NET0131  & ~n54430 ;
  assign n54432 = ~\u0_R11_reg[26]/NET0131  & n54430 ;
  assign n54433 = ~n54431 & ~n54432 ;
  assign n54447 = decrypt_pad & ~\u0_uk_K_r11_reg[14]/NET0131  ;
  assign n54448 = ~decrypt_pad & ~\u0_uk_K_r11_reg[23]/NET0131  ;
  assign n54449 = ~n54447 & ~n54448 ;
  assign n54450 = \u0_R11_reg[29]/NET0131  & ~n54449 ;
  assign n54451 = ~\u0_R11_reg[29]/NET0131  & n54449 ;
  assign n54452 = ~n54450 & ~n54451 ;
  assign n54474 = ~n54433 & ~n54452 ;
  assign n54458 = decrypt_pad & ~\u0_uk_K_r11_reg[35]/NET0131  ;
  assign n54459 = ~decrypt_pad & ~\u0_uk_K_r11_reg[44]/NET0131  ;
  assign n54460 = ~n54458 & ~n54459 ;
  assign n54461 = \u0_R11_reg[27]/NET0131  & ~n54460 ;
  assign n54462 = ~\u0_R11_reg[27]/NET0131  & n54460 ;
  assign n54463 = ~n54461 & ~n54462 ;
  assign n54441 = decrypt_pad & ~\u0_uk_K_r11_reg[45]/NET0131  ;
  assign n54442 = ~decrypt_pad & ~\u0_uk_K_r11_reg[50]/NET0131  ;
  assign n54443 = ~n54441 & ~n54442 ;
  assign n54444 = \u0_R11_reg[25]/NET0131  & ~n54443 ;
  assign n54445 = ~\u0_R11_reg[25]/NET0131  & n54443 ;
  assign n54446 = ~n54444 & ~n54445 ;
  assign n54472 = n54433 & n54446 ;
  assign n54490 = ~n54463 & ~n54472 ;
  assign n54491 = ~n54474 & n54490 ;
  assign n54434 = decrypt_pad & ~\u0_uk_K_r11_reg[37]/NET0131  ;
  assign n54435 = ~decrypt_pad & ~\u0_uk_K_r11_reg[15]/NET0131  ;
  assign n54436 = ~n54434 & ~n54435 ;
  assign n54437 = \u0_R11_reg[24]/NET0131  & ~n54436 ;
  assign n54438 = ~\u0_R11_reg[24]/NET0131  & n54436 ;
  assign n54439 = ~n54437 & ~n54438 ;
  assign n54471 = ~n54433 & ~n54446 ;
  assign n54489 = n54463 & ~n54471 ;
  assign n54492 = n54439 & ~n54489 ;
  assign n54493 = ~n54491 & n54492 ;
  assign n54455 = n54433 & ~n54446 ;
  assign n54486 = ~n54452 & n54455 ;
  assign n54487 = ~n54439 & n54486 ;
  assign n54488 = ~n54463 & n54487 ;
  assign n54440 = ~n54433 & ~n54439 ;
  assign n54482 = n54433 & n54439 ;
  assign n54483 = ~n54440 & ~n54482 ;
  assign n54494 = ~n54446 & n54463 ;
  assign n54495 = n54452 & ~n54494 ;
  assign n54496 = ~n54483 & n54495 ;
  assign n54497 = ~n54488 & ~n54496 ;
  assign n54498 = ~n54493 & n54497 ;
  assign n54499 = ~n54427 & ~n54498 ;
  assign n54464 = n54439 & n54452 ;
  assign n54465 = ~n54446 & n54464 ;
  assign n54466 = ~n54433 & n54465 ;
  assign n54467 = n54446 & n54452 ;
  assign n54468 = ~n54439 & n54467 ;
  assign n54469 = ~n54466 & ~n54468 ;
  assign n54470 = ~n54463 & ~n54469 ;
  assign n54473 = ~n54471 & ~n54472 ;
  assign n54475 = n54439 & n54463 ;
  assign n54476 = ~n54474 & n54475 ;
  assign n54477 = n54473 & n54476 ;
  assign n54453 = ~n54446 & ~n54452 ;
  assign n54454 = n54440 & n54453 ;
  assign n54456 = ~n54439 & n54452 ;
  assign n54457 = n54455 & n54456 ;
  assign n54478 = ~n54454 & ~n54457 ;
  assign n54479 = ~n54477 & n54478 ;
  assign n54480 = ~n54470 & n54479 ;
  assign n54481 = n54427 & ~n54480 ;
  assign n54500 = ~n54439 & ~n54452 ;
  assign n54501 = n54472 & n54500 ;
  assign n54502 = ~n54457 & ~n54501 ;
  assign n54503 = n54439 & n54453 ;
  assign n54504 = n54502 & ~n54503 ;
  assign n54505 = n54463 & ~n54504 ;
  assign n54484 = n54446 & ~n54463 ;
  assign n54485 = ~n54483 & n54484 ;
  assign n54506 = n54474 & n54494 ;
  assign n54507 = ~n54485 & ~n54506 ;
  assign n54508 = ~n54505 & n54507 ;
  assign n54509 = ~n54481 & n54508 ;
  assign n54510 = ~n54499 & n54509 ;
  assign n54511 = ~\u0_L11_reg[22]/NET0131  & ~n54510 ;
  assign n54512 = \u0_L11_reg[22]/NET0131  & n54510 ;
  assign n54513 = ~n54511 & ~n54512 ;
  assign n54514 = decrypt_pad & ~\u0_uk_K_r11_reg[13]/NET0131  ;
  assign n54515 = ~decrypt_pad & ~\u0_uk_K_r11_reg[18]/NET0131  ;
  assign n54516 = ~n54514 & ~n54515 ;
  assign n54517 = \u0_R11_reg[3]/NET0131  & ~n54516 ;
  assign n54518 = ~\u0_R11_reg[3]/NET0131  & n54516 ;
  assign n54519 = ~n54517 & ~n54518 ;
  assign n54526 = decrypt_pad & ~\u0_uk_K_r11_reg[19]/NET0131  ;
  assign n54527 = ~decrypt_pad & ~\u0_uk_K_r11_reg[24]/NET0131  ;
  assign n54528 = ~n54526 & ~n54527 ;
  assign n54529 = \u0_R11_reg[5]/NET0131  & ~n54528 ;
  assign n54530 = ~\u0_R11_reg[5]/NET0131  & n54528 ;
  assign n54531 = ~n54529 & ~n54530 ;
  assign n54533 = decrypt_pad & ~\u0_uk_K_r11_reg[46]/NET0131  ;
  assign n54534 = ~decrypt_pad & ~\u0_uk_K_r11_reg[26]/NET0131  ;
  assign n54535 = ~n54533 & ~n54534 ;
  assign n54536 = \u0_R11_reg[1]/NET0131  & ~n54535 ;
  assign n54537 = ~\u0_R11_reg[1]/NET0131  & n54535 ;
  assign n54538 = ~n54536 & ~n54537 ;
  assign n54540 = n54531 & ~n54538 ;
  assign n54520 = decrypt_pad & ~\u0_uk_K_r11_reg[4]/NET0131  ;
  assign n54521 = ~decrypt_pad & ~\u0_uk_K_r11_reg[41]/NET0131  ;
  assign n54522 = ~n54520 & ~n54521 ;
  assign n54523 = \u0_R11_reg[2]/NET0131  & ~n54522 ;
  assign n54524 = ~\u0_R11_reg[2]/NET0131  & n54522 ;
  assign n54525 = ~n54523 & ~n54524 ;
  assign n54541 = decrypt_pad & ~\u0_uk_K_r11_reg[25]/NET0131  ;
  assign n54542 = ~decrypt_pad & ~\u0_uk_K_r11_reg[5]/NET0131  ;
  assign n54543 = ~n54541 & ~n54542 ;
  assign n54544 = \u0_R11_reg[32]/NET0131  & ~n54543 ;
  assign n54545 = ~\u0_R11_reg[32]/NET0131  & n54543 ;
  assign n54546 = ~n54544 & ~n54545 ;
  assign n54547 = n54525 & ~n54546 ;
  assign n54574 = ~n54531 & n54547 ;
  assign n54575 = ~n54540 & ~n54574 ;
  assign n54576 = n54519 & ~n54575 ;
  assign n54583 = n54538 & ~n54546 ;
  assign n54584 = ~n54519 & n54538 ;
  assign n54585 = ~n54547 & ~n54584 ;
  assign n54586 = ~n54583 & ~n54585 ;
  assign n54580 = n54531 & ~n54546 ;
  assign n54572 = n54519 & ~n54525 ;
  assign n54581 = n54538 & ~n54572 ;
  assign n54582 = n54580 & ~n54581 ;
  assign n54555 = decrypt_pad & ~\u0_uk_K_r11_reg[48]/NET0131  ;
  assign n54556 = ~decrypt_pad & ~\u0_uk_K_r11_reg[53]/P0001  ;
  assign n54557 = ~n54555 & ~n54556 ;
  assign n54558 = \u0_R11_reg[4]/NET0131  & ~n54557 ;
  assign n54559 = ~\u0_R11_reg[4]/NET0131  & n54557 ;
  assign n54560 = ~n54558 & ~n54559 ;
  assign n54577 = ~n54525 & ~n54538 ;
  assign n54578 = ~n54531 & n54546 ;
  assign n54579 = n54577 & n54578 ;
  assign n54587 = n54560 & ~n54579 ;
  assign n54588 = ~n54582 & n54587 ;
  assign n54589 = ~n54586 & n54588 ;
  assign n54590 = ~n54576 & n54589 ;
  assign n54594 = n54531 & n54546 ;
  assign n54595 = ~n54584 & n54594 ;
  assign n54596 = ~n54531 & n54583 ;
  assign n54597 = ~n54595 & ~n54596 ;
  assign n54598 = ~n54525 & ~n54597 ;
  assign n54591 = ~n54578 & ~n54580 ;
  assign n54562 = n54525 & n54538 ;
  assign n54592 = n54519 & n54562 ;
  assign n54593 = ~n54591 & n54592 ;
  assign n54599 = ~n54560 & ~n54593 ;
  assign n54600 = ~n54598 & n54599 ;
  assign n54601 = ~n54590 & ~n54600 ;
  assign n54549 = ~n54538 & n54546 ;
  assign n54550 = ~n54531 & n54549 ;
  assign n54551 = n54525 & n54550 ;
  assign n54552 = ~n54525 & ~n54546 ;
  assign n54553 = ~n54540 & n54552 ;
  assign n54554 = ~n54551 & ~n54553 ;
  assign n54561 = ~n54554 & ~n54560 ;
  assign n54563 = n54531 & n54562 ;
  assign n54564 = n54546 & n54563 ;
  assign n54532 = ~n54525 & ~n54531 ;
  assign n54539 = n54532 & n54538 ;
  assign n54548 = n54540 & n54547 ;
  assign n54565 = ~n54539 & ~n54548 ;
  assign n54566 = ~n54564 & n54565 ;
  assign n54567 = ~n54561 & n54566 ;
  assign n54568 = ~n54519 & ~n54567 ;
  assign n54569 = ~n54531 & ~n54538 ;
  assign n54570 = n54519 & n54547 ;
  assign n54571 = n54569 & n54570 ;
  assign n54573 = n54549 & n54572 ;
  assign n54602 = ~n54571 & ~n54573 ;
  assign n54603 = ~n54568 & n54602 ;
  assign n54604 = ~n54601 & n54603 ;
  assign n54605 = ~\u0_L11_reg[31]/NET0131  & ~n54604 ;
  assign n54606 = \u0_L11_reg[31]/NET0131  & n54604 ;
  assign n54607 = ~n54605 & ~n54606 ;
  assign n54647 = decrypt_pad & ~\u0_uk_K_r11_reg[15]/NET0131  ;
  assign n54648 = ~decrypt_pad & ~\u0_uk_K_r11_reg[52]/NET0131  ;
  assign n54649 = ~n54647 & ~n54648 ;
  assign n54650 = \u0_R11_reg[24]/NET0131  & ~n54649 ;
  assign n54651 = ~\u0_R11_reg[24]/NET0131  & n54649 ;
  assign n54652 = ~n54650 & ~n54651 ;
  assign n54608 = decrypt_pad & ~\u0_uk_K_r11_reg[0]/NET0131  ;
  assign n54609 = ~decrypt_pad & ~\u0_uk_K_r11_reg[9]/NET0131  ;
  assign n54610 = ~n54608 & ~n54609 ;
  assign n54611 = \u0_R11_reg[22]/NET0131  & ~n54610 ;
  assign n54612 = ~\u0_R11_reg[22]/NET0131  & n54610 ;
  assign n54613 = ~n54611 & ~n54612 ;
  assign n54614 = decrypt_pad & ~\u0_uk_K_r11_reg[9]/NET0131  ;
  assign n54615 = ~decrypt_pad & ~\u0_uk_K_r11_reg[42]/NET0131  ;
  assign n54616 = ~n54614 & ~n54615 ;
  assign n54617 = \u0_R11_reg[21]/NET0131  & ~n54616 ;
  assign n54618 = ~\u0_R11_reg[21]/NET0131  & n54616 ;
  assign n54619 = ~n54617 & ~n54618 ;
  assign n54620 = decrypt_pad & ~\u0_uk_K_r11_reg[49]/NET0131  ;
  assign n54621 = ~decrypt_pad & ~\u0_uk_K_r11_reg[31]/NET0131  ;
  assign n54622 = ~n54620 & ~n54621 ;
  assign n54623 = \u0_R11_reg[20]/NET0131  & ~n54622 ;
  assign n54624 = ~\u0_R11_reg[20]/NET0131  & n54622 ;
  assign n54625 = ~n54623 & ~n54624 ;
  assign n54626 = n54619 & ~n54625 ;
  assign n54634 = decrypt_pad & ~\u0_uk_K_r11_reg[38]/NET0131  ;
  assign n54635 = ~decrypt_pad & ~\u0_uk_K_r11_reg[43]/NET0131  ;
  assign n54636 = ~n54634 & ~n54635 ;
  assign n54637 = \u0_R11_reg[25]/NET0131  & ~n54636 ;
  assign n54638 = ~\u0_R11_reg[25]/NET0131  & n54636 ;
  assign n54639 = ~n54637 & ~n54638 ;
  assign n54641 = n54625 & n54639 ;
  assign n54683 = ~n54626 & ~n54641 ;
  assign n54684 = n54613 & ~n54683 ;
  assign n54627 = decrypt_pad & ~\u0_uk_K_r11_reg[44]/NET0131  ;
  assign n54628 = ~decrypt_pad & ~\u0_uk_K_r11_reg[22]/NET0131  ;
  assign n54629 = ~n54627 & ~n54628 ;
  assign n54630 = \u0_R11_reg[23]/NET0131  & ~n54629 ;
  assign n54631 = ~\u0_R11_reg[23]/NET0131  & n54629 ;
  assign n54632 = ~n54630 & ~n54631 ;
  assign n54681 = n54626 & n54639 ;
  assign n54682 = ~n54613 & ~n54681 ;
  assign n54685 = ~n54632 & ~n54682 ;
  assign n54686 = ~n54684 & n54685 ;
  assign n54663 = ~n54613 & ~n54632 ;
  assign n54679 = n54641 & n54663 ;
  assign n54680 = ~n54619 & n54679 ;
  assign n54687 = ~n54613 & ~n54639 ;
  assign n54688 = ~n54619 & ~n54687 ;
  assign n54689 = n54632 & ~n54688 ;
  assign n54672 = n54619 & n54625 ;
  assign n54673 = ~n54639 & n54672 ;
  assign n54690 = ~n54613 & ~n54625 ;
  assign n54691 = ~n54673 & ~n54690 ;
  assign n54692 = n54689 & n54691 ;
  assign n54693 = ~n54680 & ~n54692 ;
  assign n54694 = ~n54686 & n54693 ;
  assign n54695 = n54652 & ~n54694 ;
  assign n54656 = n54619 & ~n54639 ;
  assign n54657 = n54625 & ~n54656 ;
  assign n54658 = n54632 & ~n54657 ;
  assign n54653 = ~n54619 & n54639 ;
  assign n54654 = n54625 & ~n54653 ;
  assign n54655 = ~n54632 & n54654 ;
  assign n54659 = ~n54613 & ~n54655 ;
  assign n54660 = ~n54658 & n54659 ;
  assign n54642 = ~n54632 & ~n54641 ;
  assign n54640 = ~n54625 & ~n54639 ;
  assign n54643 = ~n54619 & ~n54640 ;
  assign n54644 = ~n54642 & n54643 ;
  assign n54633 = n54626 & ~n54632 ;
  assign n54645 = n54613 & ~n54633 ;
  assign n54646 = ~n54644 & n54645 ;
  assign n54661 = ~n54646 & ~n54652 ;
  assign n54662 = ~n54660 & n54661 ;
  assign n54675 = ~n54625 & n54653 ;
  assign n54676 = n54632 & ~n54675 ;
  assign n54674 = ~n54632 & ~n54673 ;
  assign n54677 = ~n54613 & ~n54674 ;
  assign n54678 = ~n54676 & n54677 ;
  assign n54664 = ~n54619 & n54640 ;
  assign n54665 = n54663 & n54664 ;
  assign n54666 = n54613 & n54625 ;
  assign n54667 = n54626 & ~n54639 ;
  assign n54668 = ~n54666 & ~n54667 ;
  assign n54669 = n54613 & ~n54639 ;
  assign n54670 = n54632 & ~n54669 ;
  assign n54671 = ~n54668 & n54670 ;
  assign n54696 = ~n54665 & ~n54671 ;
  assign n54697 = ~n54678 & n54696 ;
  assign n54698 = ~n54662 & n54697 ;
  assign n54699 = ~n54695 & n54698 ;
  assign n54700 = \u0_L11_reg[11]/P0001  & ~n54699 ;
  assign n54701 = ~\u0_L11_reg[11]/P0001  & n54699 ;
  assign n54702 = ~n54700 & ~n54701 ;
  assign n54755 = decrypt_pad & ~\u0_uk_K_r11_reg[42]/NET0131  ;
  assign n54756 = ~decrypt_pad & ~\u0_uk_K_r11_reg[51]/NET0131  ;
  assign n54757 = ~n54755 & ~n54756 ;
  assign n54758 = \u0_R11_reg[32]/NET0131  & ~n54757 ;
  assign n54759 = ~\u0_R11_reg[32]/NET0131  & n54757 ;
  assign n54760 = ~n54758 & ~n54759 ;
  assign n54733 = decrypt_pad & ~\u0_uk_K_r11_reg[36]/NET0131  ;
  assign n54734 = ~decrypt_pad & ~\u0_uk_K_r11_reg[14]/NET0131  ;
  assign n54735 = ~n54733 & ~n54734 ;
  assign n54736 = \u0_R11_reg[31]/P0001  & ~n54735 ;
  assign n54737 = ~\u0_R11_reg[31]/P0001  & n54735 ;
  assign n54738 = ~n54736 & ~n54737 ;
  assign n54703 = decrypt_pad & ~\u0_uk_K_r11_reg[52]/NET0131  ;
  assign n54704 = ~decrypt_pad & ~\u0_uk_K_r11_reg[2]/NET0131  ;
  assign n54705 = ~n54703 & ~n54704 ;
  assign n54706 = \u0_R11_reg[30]/NET0131  & ~n54705 ;
  assign n54707 = ~\u0_R11_reg[30]/NET0131  & n54705 ;
  assign n54708 = ~n54706 & ~n54707 ;
  assign n54709 = decrypt_pad & ~\u0_uk_K_r11_reg[23]/NET0131  ;
  assign n54710 = ~decrypt_pad & ~\u0_uk_K_r11_reg[1]/NET0131  ;
  assign n54711 = ~n54709 & ~n54710 ;
  assign n54712 = \u0_R11_reg[29]/NET0131  & ~n54711 ;
  assign n54713 = ~\u0_R11_reg[29]/NET0131  & n54711 ;
  assign n54714 = ~n54712 & ~n54713 ;
  assign n54722 = decrypt_pad & ~\u0_uk_K_r11_reg[51]/NET0131  ;
  assign n54723 = ~decrypt_pad & ~\u0_uk_K_r11_reg[29]/NET0131  ;
  assign n54724 = ~n54722 & ~n54723 ;
  assign n54725 = \u0_R11_reg[28]/NET0131  & ~n54724 ;
  assign n54726 = ~\u0_R11_reg[28]/NET0131  & n54724 ;
  assign n54727 = ~n54725 & ~n54726 ;
  assign n54768 = ~n54714 & n54727 ;
  assign n54716 = decrypt_pad & ~\u0_uk_K_r11_reg[8]/NET0131  ;
  assign n54717 = ~decrypt_pad & ~\u0_uk_K_r11_reg[45]/NET0131  ;
  assign n54718 = ~n54716 & ~n54717 ;
  assign n54719 = \u0_R11_reg[1]/NET0131  & ~n54718 ;
  assign n54720 = ~\u0_R11_reg[1]/NET0131  & n54718 ;
  assign n54721 = ~n54719 & ~n54720 ;
  assign n54769 = n54721 & n54727 ;
  assign n54770 = ~n54768 & ~n54769 ;
  assign n54771 = ~n54708 & ~n54770 ;
  assign n54766 = ~n54721 & ~n54727 ;
  assign n54767 = n54714 & n54766 ;
  assign n54741 = n54708 & n54714 ;
  assign n54772 = ~n54721 & n54741 ;
  assign n54773 = ~n54767 & ~n54772 ;
  assign n54774 = ~n54771 & n54773 ;
  assign n54775 = n54738 & ~n54774 ;
  assign n54762 = ~n54708 & ~n54714 ;
  assign n54763 = ~n54727 & n54762 ;
  assign n54764 = ~n54738 & n54763 ;
  assign n54742 = n54721 & n54741 ;
  assign n54765 = ~n54727 & n54742 ;
  assign n54776 = ~n54764 & ~n54765 ;
  assign n54777 = ~n54775 & n54776 ;
  assign n54778 = n54760 & ~n54777 ;
  assign n54743 = ~n54708 & n54714 ;
  assign n54744 = ~n54721 & n54743 ;
  assign n54740 = ~n54708 & ~n54738 ;
  assign n54745 = ~n54740 & ~n54742 ;
  assign n54746 = ~n54744 & n54745 ;
  assign n54747 = n54727 & ~n54746 ;
  assign n54715 = n54708 & ~n54714 ;
  assign n54728 = ~n54721 & n54727 ;
  assign n54729 = n54715 & n54728 ;
  assign n54730 = n54721 & ~n54727 ;
  assign n54731 = ~n54714 & n54730 ;
  assign n54732 = ~n54729 & ~n54731 ;
  assign n54739 = ~n54732 & n54738 ;
  assign n54748 = ~n54728 & ~n54738 ;
  assign n54749 = ~n54714 & n54721 ;
  assign n54750 = ~n54708 & ~n54721 ;
  assign n54751 = ~n54749 & ~n54750 ;
  assign n54752 = n54748 & n54751 ;
  assign n54753 = ~n54739 & ~n54752 ;
  assign n54754 = ~n54747 & n54753 ;
  assign n54761 = ~n54754 & ~n54760 ;
  assign n54785 = ~n54727 & n54772 ;
  assign n54786 = n54762 & n54769 ;
  assign n54787 = ~n54785 & ~n54786 ;
  assign n54788 = n54708 & n54731 ;
  assign n54789 = ~n54714 & n54766 ;
  assign n54790 = ~n54708 & n54789 ;
  assign n54791 = ~n54788 & ~n54790 ;
  assign n54792 = n54787 & n54791 ;
  assign n54793 = n54738 & ~n54792 ;
  assign n54779 = n54708 & ~n54738 ;
  assign n54780 = n54760 & n54768 ;
  assign n54781 = n54779 & n54780 ;
  assign n54782 = n54714 & n54727 ;
  assign n54783 = ~n54721 & n54782 ;
  assign n54784 = n54740 & n54783 ;
  assign n54794 = ~n54781 & ~n54784 ;
  assign n54795 = ~n54793 & n54794 ;
  assign n54796 = ~n54761 & n54795 ;
  assign n54797 = ~n54778 & n54796 ;
  assign n54798 = \u0_L11_reg[5]/NET0131  & ~n54797 ;
  assign n54799 = ~\u0_L11_reg[5]/NET0131  & n54797 ;
  assign n54800 = ~n54798 & ~n54799 ;
  assign n54830 = decrypt_pad & ~\u0_uk_K_r11_reg[10]/NET0131  ;
  assign n54831 = ~decrypt_pad & ~\u0_uk_K_r11_reg[47]/NET0131  ;
  assign n54832 = ~n54830 & ~n54831 ;
  assign n54833 = \u0_R11_reg[15]/NET0131  & ~n54832 ;
  assign n54834 = ~\u0_R11_reg[15]/NET0131  & n54832 ;
  assign n54835 = ~n54833 & ~n54834 ;
  assign n54801 = decrypt_pad & ~\u0_uk_K_r11_reg[33]/NET0131  ;
  assign n54802 = ~decrypt_pad & ~\u0_uk_K_r11_reg[13]/NET0131  ;
  assign n54803 = ~n54801 & ~n54802 ;
  assign n54804 = \u0_R11_reg[13]/NET0131  & ~n54803 ;
  assign n54805 = ~\u0_R11_reg[13]/NET0131  & n54803 ;
  assign n54806 = ~n54804 & ~n54805 ;
  assign n54814 = decrypt_pad & ~\u0_uk_K_r11_reg[55]/NET0131  ;
  assign n54815 = ~decrypt_pad & ~\u0_uk_K_r11_reg[3]/NET0131  ;
  assign n54816 = ~n54814 & ~n54815 ;
  assign n54817 = \u0_R11_reg[17]/NET0131  & ~n54816 ;
  assign n54818 = ~\u0_R11_reg[17]/NET0131  & n54816 ;
  assign n54819 = ~n54817 & ~n54818 ;
  assign n54851 = ~n54806 & n54819 ;
  assign n54807 = decrypt_pad & ~\u0_uk_K_r11_reg[34]/NET0131  ;
  assign n54808 = ~decrypt_pad & ~\u0_uk_K_r11_reg[39]/NET0131  ;
  assign n54809 = ~n54807 & ~n54808 ;
  assign n54810 = \u0_R11_reg[14]/NET0131  & ~n54809 ;
  assign n54811 = ~\u0_R11_reg[14]/NET0131  & n54809 ;
  assign n54812 = ~n54810 & ~n54811 ;
  assign n54820 = decrypt_pad & ~\u0_uk_K_r11_reg[39]/NET0131  ;
  assign n54821 = ~decrypt_pad & ~\u0_uk_K_r11_reg[19]/NET0131  ;
  assign n54822 = ~n54820 & ~n54821 ;
  assign n54823 = \u0_R11_reg[12]/NET0131  & ~n54822 ;
  assign n54824 = ~\u0_R11_reg[12]/NET0131  & n54822 ;
  assign n54825 = ~n54823 & ~n54824 ;
  assign n54826 = ~n54819 & n54825 ;
  assign n54852 = n54812 & n54826 ;
  assign n54853 = ~n54851 & ~n54852 ;
  assign n54854 = ~n54835 & ~n54853 ;
  assign n54836 = ~n54819 & n54835 ;
  assign n54856 = ~n54806 & ~n54825 ;
  assign n54857 = n54836 & n54856 ;
  assign n54845 = decrypt_pad & ~\u0_uk_K_r11_reg[18]/NET0131  ;
  assign n54846 = ~decrypt_pad & ~\u0_uk_K_r11_reg[55]/NET0131  ;
  assign n54847 = ~n54845 & ~n54846 ;
  assign n54848 = \u0_R11_reg[16]/NET0131  & ~n54847 ;
  assign n54849 = ~\u0_R11_reg[16]/NET0131  & n54847 ;
  assign n54850 = ~n54848 & ~n54849 ;
  assign n54840 = ~n54812 & n54825 ;
  assign n54855 = n54840 & n54851 ;
  assign n54867 = ~n54850 & ~n54855 ;
  assign n54868 = ~n54857 & n54867 ;
  assign n54858 = n54806 & n54835 ;
  assign n54841 = n54812 & ~n54825 ;
  assign n54859 = n54819 & n54825 ;
  assign n54860 = ~n54841 & ~n54859 ;
  assign n54861 = n54858 & ~n54860 ;
  assign n54862 = n54806 & ~n54819 ;
  assign n54863 = n54841 & n54862 ;
  assign n54864 = ~n54812 & ~n54819 ;
  assign n54865 = n54856 & n54864 ;
  assign n54866 = ~n54863 & ~n54865 ;
  assign n54869 = ~n54861 & n54866 ;
  assign n54870 = n54868 & n54869 ;
  assign n54871 = ~n54854 & n54870 ;
  assign n54872 = ~n54835 & n54856 ;
  assign n54873 = ~n54819 & n54872 ;
  assign n54874 = n54812 & n54873 ;
  assign n54875 = n54806 & n54825 ;
  assign n54876 = n54812 & n54819 ;
  assign n54877 = ~n54836 & ~n54876 ;
  assign n54878 = n54875 & ~n54877 ;
  assign n54885 = n54850 & ~n54878 ;
  assign n54827 = n54819 & ~n54825 ;
  assign n54813 = n54806 & ~n54812 ;
  assign n54879 = ~n54806 & n54835 ;
  assign n54880 = ~n54813 & ~n54879 ;
  assign n54881 = n54827 & ~n54880 ;
  assign n54882 = ~n54856 & ~n54875 ;
  assign n54883 = ~n54812 & ~n54835 ;
  assign n54884 = n54882 & n54883 ;
  assign n54886 = ~n54881 & ~n54884 ;
  assign n54887 = n54885 & n54886 ;
  assign n54888 = ~n54874 & n54887 ;
  assign n54889 = ~n54871 & ~n54888 ;
  assign n54828 = ~n54826 & ~n54827 ;
  assign n54829 = n54813 & ~n54828 ;
  assign n54837 = n54819 & ~n54835 ;
  assign n54838 = ~n54836 & ~n54837 ;
  assign n54839 = n54829 & ~n54838 ;
  assign n54842 = ~n54840 & ~n54841 ;
  assign n54843 = n54836 & n54842 ;
  assign n54844 = ~n54806 & n54843 ;
  assign n54890 = ~n54839 & ~n54844 ;
  assign n54891 = ~n54889 & n54890 ;
  assign n54892 = ~\u0_L11_reg[20]/NET0131  & ~n54891 ;
  assign n54893 = \u0_L11_reg[20]/NET0131  & n54891 ;
  assign n54894 = ~n54892 & ~n54893 ;
  assign n54895 = n54806 & ~n54835 ;
  assign n54909 = n54812 & ~n54827 ;
  assign n54910 = ~n54826 & ~n54909 ;
  assign n54911 = n54895 & n54910 ;
  assign n54907 = n54812 & ~n54882 ;
  assign n54908 = ~n54859 & n54907 ;
  assign n54912 = ~n54819 & ~n54840 ;
  assign n54913 = n54879 & ~n54912 ;
  assign n54914 = ~n54908 & ~n54913 ;
  assign n54915 = ~n54911 & n54914 ;
  assign n54916 = n54850 & ~n54915 ;
  assign n54897 = n54806 & ~n54864 ;
  assign n54898 = n54843 & ~n54897 ;
  assign n54900 = ~n54851 & ~n54864 ;
  assign n54901 = n54825 & ~n54835 ;
  assign n54902 = ~n54900 & n54901 ;
  assign n54899 = n54875 & n54876 ;
  assign n54903 = ~n54829 & ~n54899 ;
  assign n54904 = ~n54902 & n54903 ;
  assign n54905 = ~n54898 & n54904 ;
  assign n54906 = ~n54850 & ~n54905 ;
  assign n54917 = n54819 & n54907 ;
  assign n54918 = ~n54863 & ~n54917 ;
  assign n54919 = n54835 & ~n54918 ;
  assign n54896 = n54852 & n54895 ;
  assign n54920 = ~n54874 & ~n54896 ;
  assign n54921 = ~n54919 & n54920 ;
  assign n54922 = ~n54906 & n54921 ;
  assign n54923 = ~n54916 & n54922 ;
  assign n54924 = ~\u0_L11_reg[1]/NET0131  & ~n54923 ;
  assign n54925 = \u0_L11_reg[1]/NET0131  & n54923 ;
  assign n54926 = ~n54924 & ~n54925 ;
  assign n54947 = ~n54813 & n54826 ;
  assign n54948 = n54813 & n54827 ;
  assign n54949 = ~n54947 & ~n54948 ;
  assign n54950 = ~n54835 & ~n54949 ;
  assign n54944 = n54835 & ~n54876 ;
  assign n54945 = n54828 & n54944 ;
  assign n54946 = n54882 & n54945 ;
  assign n54951 = ~n54917 & ~n54946 ;
  assign n54952 = ~n54950 & n54951 ;
  assign n54953 = n54850 & ~n54952 ;
  assign n54928 = ~n54812 & n54819 ;
  assign n54933 = ~n54825 & n54835 ;
  assign n54934 = n54928 & n54933 ;
  assign n54935 = n54866 & ~n54934 ;
  assign n54931 = ~n54806 & ~n54837 ;
  assign n54932 = n54840 & ~n54931 ;
  assign n54927 = n54825 & n54835 ;
  assign n54929 = ~n54806 & n54927 ;
  assign n54930 = ~n54928 & n54929 ;
  assign n54936 = ~n54873 & ~n54930 ;
  assign n54937 = ~n54932 & n54936 ;
  assign n54938 = n54935 & n54937 ;
  assign n54939 = ~n54850 & ~n54938 ;
  assign n54940 = ~n54865 & ~n54917 ;
  assign n54941 = ~n54835 & ~n54940 ;
  assign n54942 = n54858 & ~n54928 ;
  assign n54943 = ~n54842 & n54942 ;
  assign n54954 = ~n54941 & ~n54943 ;
  assign n54955 = ~n54939 & n54954 ;
  assign n54956 = ~n54953 & n54955 ;
  assign n54957 = ~\u0_L11_reg[10]/NET0131  & ~n54956 ;
  assign n54958 = \u0_L11_reg[10]/NET0131  & n54956 ;
  assign n54959 = ~n54957 & ~n54958 ;
  assign n54997 = decrypt_pad & ~\u0_uk_K_r11_reg[17]/NET0131  ;
  assign n54998 = ~decrypt_pad & ~\u0_uk_K_r11_reg[54]/NET0131  ;
  assign n54999 = ~n54997 & ~n54998 ;
  assign n55000 = \u0_R11_reg[8]/NET0131  & ~n54999 ;
  assign n55001 = ~\u0_R11_reg[8]/NET0131  & n54999 ;
  assign n55002 = ~n55000 & ~n55001 ;
  assign n54990 = decrypt_pad & ~\u0_uk_K_r11_reg[26]/NET0131  ;
  assign n54991 = ~decrypt_pad & ~\u0_uk_K_r11_reg[6]/NET0131  ;
  assign n54992 = ~n54990 & ~n54991 ;
  assign n54993 = \u0_R11_reg[7]/NET0131  & ~n54992 ;
  assign n54994 = ~\u0_R11_reg[7]/NET0131  & n54992 ;
  assign n54995 = ~n54993 & ~n54994 ;
  assign n54960 = decrypt_pad & ~\u0_uk_K_r11_reg[32]/NET0131  ;
  assign n54961 = ~decrypt_pad & ~\u0_uk_K_r11_reg[12]/NET0131  ;
  assign n54962 = ~n54960 & ~n54961 ;
  assign n54963 = \u0_R11_reg[6]/NET0131  & ~n54962 ;
  assign n54964 = ~\u0_R11_reg[6]/NET0131  & n54962 ;
  assign n54965 = ~n54963 & ~n54964 ;
  assign n54973 = decrypt_pad & ~\u0_uk_K_r11_reg[5]/NET0131  ;
  assign n54974 = ~decrypt_pad & ~\u0_uk_K_r11_reg[10]/NET0131  ;
  assign n54975 = ~n54973 & ~n54974 ;
  assign n54976 = \u0_R11_reg[4]/NET0131  & ~n54975 ;
  assign n54977 = ~\u0_R11_reg[4]/NET0131  & n54975 ;
  assign n54978 = ~n54976 & ~n54977 ;
  assign n54966 = decrypt_pad & ~\u0_uk_K_r11_reg[41]/NET0131  ;
  assign n54967 = ~decrypt_pad & ~\u0_uk_K_r11_reg[46]/NET0131  ;
  assign n54968 = ~n54966 & ~n54967 ;
  assign n54969 = \u0_R11_reg[5]/NET0131  & ~n54968 ;
  assign n54970 = ~\u0_R11_reg[5]/NET0131  & n54968 ;
  assign n54971 = ~n54969 & ~n54970 ;
  assign n54980 = decrypt_pad & ~\u0_uk_K_r11_reg[54]/NET0131  ;
  assign n54981 = ~decrypt_pad & ~\u0_uk_K_r11_reg[34]/NET0131  ;
  assign n54982 = ~n54980 & ~n54981 ;
  assign n54983 = \u0_R11_reg[9]/NET0131  & ~n54982 ;
  assign n54984 = ~\u0_R11_reg[9]/NET0131  & n54982 ;
  assign n54985 = ~n54983 & ~n54984 ;
  assign n54986 = n54971 & ~n54985 ;
  assign n55026 = ~n54978 & n54986 ;
  assign n55027 = n54965 & n55026 ;
  assign n55007 = ~n54971 & n54985 ;
  assign n55028 = ~n54986 & ~n55007 ;
  assign n55029 = n54978 & n55028 ;
  assign n55030 = ~n55027 & ~n55029 ;
  assign n55031 = n54995 & ~n55030 ;
  assign n55003 = ~n54978 & ~n54985 ;
  assign n55013 = ~n54965 & n55003 ;
  assign n55014 = ~n54978 & n54985 ;
  assign n55015 = n54971 & n55014 ;
  assign n55016 = ~n55013 & ~n55015 ;
  assign n55025 = ~n54995 & ~n55016 ;
  assign n55004 = n54978 & n54985 ;
  assign n55010 = ~n54971 & n55004 ;
  assign n55022 = n54978 & n54995 ;
  assign n55023 = ~n55010 & ~n55022 ;
  assign n55024 = ~n54965 & ~n55023 ;
  assign n55032 = n54965 & n55014 ;
  assign n55033 = ~n54971 & n55032 ;
  assign n55034 = ~n55024 & ~n55033 ;
  assign n55035 = ~n55025 & n55034 ;
  assign n55036 = ~n55031 & n55035 ;
  assign n55037 = n55002 & ~n55036 ;
  assign n54972 = n54965 & ~n54971 ;
  assign n54979 = n54972 & ~n54978 ;
  assign n54987 = n54965 & n54978 ;
  assign n54988 = n54986 & n54987 ;
  assign n54989 = ~n54979 & ~n54988 ;
  assign n54996 = ~n54989 & ~n54995 ;
  assign n55017 = n54995 & ~n55016 ;
  assign n55008 = ~n54972 & n54978 ;
  assign n55009 = ~n55007 & ~n55008 ;
  assign n55011 = ~n54995 & ~n55010 ;
  assign n55012 = ~n55009 & n55011 ;
  assign n55005 = ~n55003 & ~n55004 ;
  assign n55006 = n54972 & ~n55005 ;
  assign n55018 = ~n54988 & ~n55006 ;
  assign n55019 = ~n55012 & n55018 ;
  assign n55020 = ~n55017 & n55019 ;
  assign n55021 = ~n55002 & ~n55020 ;
  assign n55038 = ~n54996 & ~n55021 ;
  assign n55039 = ~n55037 & n55038 ;
  assign n55040 = ~\u0_L11_reg[28]/NET0131  & ~n55039 ;
  assign n55041 = \u0_L11_reg[28]/NET0131  & n55039 ;
  assign n55042 = ~n55040 & ~n55041 ;
  assign n55049 = ~n54748 & ~n54779 ;
  assign n55050 = n54708 & n54768 ;
  assign n55051 = n54721 & n55050 ;
  assign n55052 = ~n55049 & ~n55051 ;
  assign n55053 = n54727 & n54741 ;
  assign n55056 = n54738 & ~n55053 ;
  assign n55054 = ~n54708 & n54749 ;
  assign n55055 = n54714 & n54730 ;
  assign n55057 = ~n55054 & ~n55055 ;
  assign n55058 = n55056 & n55057 ;
  assign n55059 = ~n55052 & ~n55058 ;
  assign n55047 = ~n54783 & ~n54789 ;
  assign n55048 = n54708 & ~n55047 ;
  assign n55046 = n54721 & n54763 ;
  assign n55060 = n54760 & ~n55046 ;
  assign n55061 = ~n55048 & n55060 ;
  assign n55062 = ~n55059 & n55061 ;
  assign n55071 = ~n54729 & ~n54760 ;
  assign n55044 = n54740 & n54769 ;
  assign n55065 = ~n54727 & n54741 ;
  assign n55072 = ~n55044 & ~n55065 ;
  assign n55073 = n55071 & n55072 ;
  assign n55070 = ~n54738 & n54767 ;
  assign n55074 = ~n54790 & ~n55070 ;
  assign n55075 = n55073 & n55074 ;
  assign n55063 = ~n54783 & ~n55050 ;
  assign n55064 = n54738 & ~n55063 ;
  assign n55066 = ~n54727 & n54779 ;
  assign n55067 = n54727 & n54743 ;
  assign n55068 = ~n55066 & ~n55067 ;
  assign n55069 = n54721 & ~n55068 ;
  assign n55076 = ~n55064 & ~n55069 ;
  assign n55077 = n55075 & n55076 ;
  assign n55078 = ~n55062 & ~n55077 ;
  assign n55043 = n54738 & n54763 ;
  assign n55045 = n54714 & n55044 ;
  assign n55079 = ~n55043 & ~n55045 ;
  assign n55080 = ~n55078 & n55079 ;
  assign n55081 = ~\u0_L11_reg[21]/NET0131  & ~n55080 ;
  assign n55082 = \u0_L11_reg[21]/NET0131  & n55080 ;
  assign n55083 = ~n55081 & ~n55082 ;
  assign n55085 = n54439 & n54446 ;
  assign n55086 = ~n54454 & ~n55085 ;
  assign n55087 = n54463 & ~n55086 ;
  assign n55091 = n54427 & ~n54501 ;
  assign n55092 = ~n54466 & n55091 ;
  assign n55084 = n54457 & ~n54463 ;
  assign n55088 = ~n54467 & ~n54482 ;
  assign n55089 = ~n54464 & ~n54472 ;
  assign n55090 = ~n55088 & n55089 ;
  assign n55093 = ~n55084 & ~n55090 ;
  assign n55094 = n55092 & n55093 ;
  assign n55095 = ~n55087 & n55094 ;
  assign n55099 = n54446 & n54500 ;
  assign n55100 = ~n54503 & ~n55099 ;
  assign n55101 = ~n54433 & ~n55100 ;
  assign n55096 = n54433 & n54465 ;
  assign n55097 = ~n54472 & ~n54494 ;
  assign n55098 = n54456 & ~n55097 ;
  assign n55105 = ~n55096 & ~n55098 ;
  assign n55106 = ~n55101 & n55105 ;
  assign n55102 = ~n54453 & n55088 ;
  assign n55103 = ~n54463 & ~n55102 ;
  assign n55104 = ~n54427 & ~n54487 ;
  assign n55107 = ~n55103 & n55104 ;
  assign n55108 = n55106 & n55107 ;
  assign n55109 = ~n55095 & ~n55108 ;
  assign n55110 = \u0_L11_reg[12]/NET0131  & n55109 ;
  assign n55111 = ~\u0_L11_reg[12]/NET0131  & ~n55109 ;
  assign n55112 = ~n55110 & ~n55111 ;
  assign n55132 = ~n54538 & n54591 ;
  assign n55133 = n54532 & ~n54546 ;
  assign n55134 = ~n55132 & ~n55133 ;
  assign n55135 = ~n54519 & ~n55134 ;
  assign n55136 = n54538 & n54546 ;
  assign n55137 = n54531 & n55136 ;
  assign n55138 = ~n54550 & ~n55137 ;
  assign n55139 = n54519 & ~n55138 ;
  assign n55131 = n54562 & n54578 ;
  assign n55140 = ~n54548 & ~n55131 ;
  assign n55141 = ~n55139 & n55140 ;
  assign n55142 = ~n55135 & n55141 ;
  assign n55143 = ~n54560 & ~n55142 ;
  assign n55113 = n54538 & n54580 ;
  assign n55114 = ~n54525 & n55113 ;
  assign n55115 = ~n54531 & n54562 ;
  assign n55116 = ~n54546 & n55115 ;
  assign n55117 = ~n55114 & ~n55116 ;
  assign n55118 = n54519 & ~n55117 ;
  assign n55120 = ~n54546 & ~n54577 ;
  assign n55121 = n54577 & n54594 ;
  assign n55122 = ~n55120 & ~n55121 ;
  assign n55123 = n54519 & ~n55122 ;
  assign n55124 = ~n54525 & n54546 ;
  assign n55125 = ~n54519 & ~n55124 ;
  assign n55126 = ~n55120 & n55125 ;
  assign n55119 = n54539 & n54546 ;
  assign n55127 = ~n54563 & ~n55119 ;
  assign n55128 = ~n55126 & n55127 ;
  assign n55129 = ~n55123 & n55128 ;
  assign n55130 = n54560 & ~n55129 ;
  assign n55144 = ~n55118 & ~n55130 ;
  assign n55145 = ~n55143 & n55144 ;
  assign n55146 = ~\u0_L11_reg[17]/NET0131  & ~n55145 ;
  assign n55147 = \u0_L11_reg[17]/NET0131  & n55145 ;
  assign n55148 = ~n55146 & ~n55147 ;
  assign n55149 = decrypt_pad & ~\u0_uk_K_r11_reg[31]/NET0131  ;
  assign n55150 = ~decrypt_pad & ~\u0_uk_K_r11_reg[36]/NET0131  ;
  assign n55151 = ~n55149 & ~n55150 ;
  assign n55152 = \u0_R11_reg[20]/NET0131  & ~n55151 ;
  assign n55153 = ~\u0_R11_reg[20]/NET0131  & n55151 ;
  assign n55154 = ~n55152 & ~n55153 ;
  assign n55184 = decrypt_pad & ~\u0_uk_K_r11_reg[43]/NET0131  ;
  assign n55185 = ~decrypt_pad & ~\u0_uk_K_r11_reg[21]/NET0131  ;
  assign n55186 = ~n55184 & ~n55185 ;
  assign n55187 = \u0_R11_reg[19]/NET0131  & ~n55186 ;
  assign n55188 = ~\u0_R11_reg[19]/NET0131  & n55186 ;
  assign n55189 = ~n55187 & ~n55188 ;
  assign n55168 = decrypt_pad & ~\u0_uk_K_r11_reg[28]/NET0131  ;
  assign n55169 = ~decrypt_pad & ~\u0_uk_K_r11_reg[37]/NET0131  ;
  assign n55170 = ~n55168 & ~n55169 ;
  assign n55171 = \u0_R11_reg[21]/NET0131  & ~n55170 ;
  assign n55172 = ~\u0_R11_reg[21]/NET0131  & n55170 ;
  assign n55173 = ~n55171 & ~n55172 ;
  assign n55161 = decrypt_pad & ~\u0_uk_K_r11_reg[16]/NET0131  ;
  assign n55162 = ~decrypt_pad & ~\u0_uk_K_r11_reg[49]/NET0131  ;
  assign n55163 = ~n55161 & ~n55162 ;
  assign n55164 = \u0_R11_reg[16]/NET0131  & ~n55163 ;
  assign n55165 = ~\u0_R11_reg[16]/NET0131  & n55163 ;
  assign n55166 = ~n55164 & ~n55165 ;
  assign n55176 = decrypt_pad & ~\u0_uk_K_r11_reg[1]/NET0131  ;
  assign n55177 = ~decrypt_pad & ~\u0_uk_K_r11_reg[38]/NET0131  ;
  assign n55178 = ~n55176 & ~n55177 ;
  assign n55179 = \u0_R11_reg[18]/NET0131  & ~n55178 ;
  assign n55180 = ~\u0_R11_reg[18]/NET0131  & n55178 ;
  assign n55181 = ~n55179 & ~n55180 ;
  assign n55191 = n55166 & n55181 ;
  assign n55192 = ~n55173 & ~n55191 ;
  assign n55155 = decrypt_pad & ~\u0_uk_K_r11_reg[7]/NET0131  ;
  assign n55156 = ~decrypt_pad & ~\u0_uk_K_r11_reg[16]/NET0131  ;
  assign n55157 = ~n55155 & ~n55156 ;
  assign n55158 = \u0_R11_reg[17]/NET0131  & ~n55157 ;
  assign n55159 = ~\u0_R11_reg[17]/NET0131  & n55157 ;
  assign n55160 = ~n55158 & ~n55159 ;
  assign n55198 = n55160 & ~n55181 ;
  assign n55199 = n55192 & ~n55198 ;
  assign n55196 = n55160 & n55166 ;
  assign n55197 = n55173 & n55196 ;
  assign n55200 = ~n55160 & ~n55166 ;
  assign n55201 = ~n55197 & ~n55200 ;
  assign n55202 = ~n55199 & n55201 ;
  assign n55203 = n55189 & ~n55202 ;
  assign n55167 = ~n55160 & n55166 ;
  assign n55174 = n55167 & n55173 ;
  assign n55175 = n55160 & ~n55166 ;
  assign n55182 = n55175 & ~n55181 ;
  assign n55183 = ~n55174 & ~n55182 ;
  assign n55190 = ~n55183 & ~n55189 ;
  assign n55193 = n55173 & n55181 ;
  assign n55194 = n55160 & ~n55193 ;
  assign n55195 = ~n55192 & n55194 ;
  assign n55204 = ~n55190 & ~n55195 ;
  assign n55205 = ~n55203 & n55204 ;
  assign n55206 = n55154 & ~n55205 ;
  assign n55222 = ~n55173 & n55200 ;
  assign n55223 = ~n55173 & n55196 ;
  assign n55224 = ~n55222 & ~n55223 ;
  assign n55225 = n55181 & ~n55224 ;
  assign n55226 = n55173 & n55200 ;
  assign n55227 = ~n55181 & n55226 ;
  assign n55228 = ~n55225 & ~n55227 ;
  assign n55229 = n55189 & ~n55228 ;
  assign n55210 = ~n55173 & n55189 ;
  assign n55211 = n55167 & ~n55173 ;
  assign n55212 = n55175 & n55181 ;
  assign n55213 = ~n55211 & ~n55212 ;
  assign n55214 = ~n55210 & ~n55213 ;
  assign n55216 = n55160 & ~n55173 ;
  assign n55217 = n55189 & ~n55216 ;
  assign n55215 = ~n55189 & ~n55200 ;
  assign n55218 = ~n55181 & ~n55215 ;
  assign n55219 = ~n55217 & n55218 ;
  assign n55220 = ~n55214 & ~n55219 ;
  assign n55221 = ~n55154 & ~n55220 ;
  assign n55207 = ~n55160 & n55181 ;
  assign n55208 = n55166 & ~n55189 ;
  assign n55209 = n55207 & n55208 ;
  assign n55230 = n55173 & ~n55181 ;
  assign n55231 = n55196 & n55230 ;
  assign n55232 = ~n55209 & ~n55231 ;
  assign n55233 = ~n55221 & n55232 ;
  assign n55234 = ~n55229 & n55233 ;
  assign n55235 = ~n55206 & n55234 ;
  assign n55236 = ~\u0_L11_reg[25]/NET0131  & ~n55235 ;
  assign n55237 = \u0_L11_reg[25]/NET0131  & n55235 ;
  assign n55238 = ~n55236 & ~n55237 ;
  assign n55243 = n54654 & ~n54656 ;
  assign n55244 = n54619 & ~n54669 ;
  assign n55245 = ~n54672 & ~n54688 ;
  assign n55246 = ~n55244 & n55245 ;
  assign n55247 = ~n55243 & ~n55246 ;
  assign n55248 = n54632 & ~n55247 ;
  assign n55239 = ~n54613 & ~n54683 ;
  assign n55240 = n54669 & n54672 ;
  assign n55241 = ~n55239 & ~n55240 ;
  assign n55242 = ~n54632 & ~n55241 ;
  assign n55249 = n54613 & n54675 ;
  assign n55250 = ~n55242 & ~n55249 ;
  assign n55251 = ~n55248 & n55250 ;
  assign n55252 = ~n54652 & ~n55251 ;
  assign n55255 = n54626 & ~n54669 ;
  assign n55256 = ~n55240 & ~n55255 ;
  assign n55257 = n54632 & ~n55256 ;
  assign n55258 = n54613 & ~n54640 ;
  assign n55259 = ~n54641 & n55258 ;
  assign n55260 = ~n54689 & ~n55239 ;
  assign n55261 = ~n55259 & n55260 ;
  assign n55262 = ~n55257 & ~n55261 ;
  assign n55263 = n54652 & ~n55262 ;
  assign n55253 = ~n54619 & n54625 ;
  assign n55254 = n54687 & n55253 ;
  assign n55264 = n54619 & n54639 ;
  assign n55265 = ~n54613 & n54632 ;
  assign n55266 = n55264 & n55265 ;
  assign n55267 = ~n55254 & ~n55266 ;
  assign n55268 = ~n55263 & n55267 ;
  assign n55269 = ~n55252 & n55268 ;
  assign n55270 = \u0_L11_reg[29]/NET0131  & ~n55269 ;
  assign n55271 = ~\u0_L11_reg[29]/NET0131  & n55269 ;
  assign n55272 = ~n55270 & ~n55271 ;
  assign n55277 = ~n54965 & n55029 ;
  assign n55273 = n54971 & n54978 ;
  assign n55274 = ~n54965 & n54971 ;
  assign n55275 = ~n55273 & ~n55274 ;
  assign n55276 = n54995 & ~n55275 ;
  assign n55278 = n55002 & ~n55276 ;
  assign n55279 = ~n55277 & n55278 ;
  assign n55280 = ~n54971 & ~n54995 ;
  assign n55281 = ~n54965 & n54985 ;
  assign n55282 = n55280 & n55281 ;
  assign n55283 = n54965 & n55015 ;
  assign n55284 = ~n55282 & ~n55283 ;
  assign n55289 = n54985 & n54995 ;
  assign n55290 = ~n54971 & n54987 ;
  assign n55291 = n55289 & n55290 ;
  assign n55292 = ~n55002 & ~n55291 ;
  assign n55293 = n55284 & n55292 ;
  assign n55285 = ~n54987 & ~n55007 ;
  assign n55286 = n55011 & ~n55285 ;
  assign n55287 = ~n55004 & ~n55028 ;
  assign n55288 = ~n54965 & n55287 ;
  assign n55294 = ~n55286 & ~n55288 ;
  assign n55295 = n55293 & n55294 ;
  assign n55296 = ~n55279 & ~n55295 ;
  assign n55297 = ~n54972 & n55014 ;
  assign n55298 = n55002 & ~n55005 ;
  assign n55299 = ~n55008 & n55298 ;
  assign n55300 = ~n55297 & ~n55299 ;
  assign n55301 = ~n55274 & ~n55300 ;
  assign n55302 = ~n54995 & ~n55301 ;
  assign n55303 = n54979 & ~n54985 ;
  assign n55304 = n54978 & n55274 ;
  assign n55305 = n54995 & ~n55304 ;
  assign n55306 = ~n55303 & n55305 ;
  assign n55307 = ~n55302 & ~n55306 ;
  assign n55308 = ~n55296 & ~n55307 ;
  assign n55309 = \u0_L11_reg[2]/NET0131  & n55308 ;
  assign n55310 = ~\u0_L11_reg[2]/NET0131  & ~n55308 ;
  assign n55311 = ~n55309 & ~n55310 ;
  assign n55334 = ~n55181 & n55211 ;
  assign n55333 = n55181 & n55216 ;
  assign n55335 = ~n55226 & ~n55231 ;
  assign n55336 = ~n55333 & n55335 ;
  assign n55337 = ~n55334 & n55336 ;
  assign n55338 = ~n55189 & ~n55337 ;
  assign n55330 = ~n55183 & ~n55230 ;
  assign n55316 = n55173 & n55191 ;
  assign n55317 = ~n55182 & ~n55316 ;
  assign n55331 = ~n55222 & n55317 ;
  assign n55332 = n55189 & ~n55331 ;
  assign n55339 = ~n55330 & ~n55332 ;
  assign n55340 = ~n55338 & n55339 ;
  assign n55341 = ~n55154 & ~n55340 ;
  assign n55320 = n55173 & n55175 ;
  assign n55321 = ~n55222 & ~n55320 ;
  assign n55322 = ~n55189 & ~n55321 ;
  assign n55323 = ~n55174 & ~n55223 ;
  assign n55324 = ~n55322 & n55323 ;
  assign n55325 = ~n55181 & ~n55324 ;
  assign n55315 = ~n55173 & ~n55196 ;
  assign n55318 = n55189 & ~n55315 ;
  assign n55319 = n55317 & n55318 ;
  assign n55312 = n55181 & ~n55189 ;
  assign n55313 = n55197 & n55312 ;
  assign n55314 = n55181 & n55211 ;
  assign n55326 = ~n55313 & ~n55314 ;
  assign n55327 = ~n55319 & n55326 ;
  assign n55328 = ~n55325 & n55327 ;
  assign n55329 = n55154 & ~n55328 ;
  assign n55342 = ~n55196 & ~n55207 ;
  assign n55343 = n55192 & ~n55342 ;
  assign n55344 = n55189 & ~n55343 ;
  assign n55345 = n55181 & n55226 ;
  assign n55346 = ~n55166 & n55333 ;
  assign n55347 = ~n55345 & ~n55346 ;
  assign n55348 = ~n55189 & n55347 ;
  assign n55349 = ~n55344 & ~n55348 ;
  assign n55350 = ~n55329 & ~n55349 ;
  assign n55351 = ~n55341 & n55350 ;
  assign n55352 = ~\u0_L11_reg[14]/NET0131  & ~n55351 ;
  assign n55353 = \u0_L11_reg[14]/NET0131  & n55351 ;
  assign n55354 = ~n55352 & ~n55353 ;
  assign n55362 = ~n54666 & ~n54690 ;
  assign n55363 = n54639 & ~n54672 ;
  assign n55364 = ~n55362 & n55363 ;
  assign n55365 = n54632 & ~n54673 ;
  assign n55366 = ~n55364 & n55365 ;
  assign n55367 = ~n54632 & ~n54667 ;
  assign n55368 = ~n55249 & n55367 ;
  assign n55369 = ~n55366 & ~n55368 ;
  assign n55370 = ~n54679 & ~n55254 ;
  assign n55371 = ~n55369 & n55370 ;
  assign n55372 = ~n54652 & ~n55371 ;
  assign n55356 = ~n54613 & ~n54640 ;
  assign n55357 = n55244 & ~n55356 ;
  assign n55355 = ~n54657 & n54663 ;
  assign n55358 = n54641 & n55265 ;
  assign n55359 = ~n55355 & ~n55358 ;
  assign n55360 = ~n55357 & n55359 ;
  assign n55361 = n54652 & ~n55360 ;
  assign n55373 = n54613 & ~n55243 ;
  assign n55374 = ~n54632 & ~n55356 ;
  assign n55375 = ~n55373 & n55374 ;
  assign n55376 = ~n54625 & ~n54653 ;
  assign n55377 = ~n54656 & n55376 ;
  assign n55378 = ~n54673 & ~n55377 ;
  assign n55379 = n54613 & n54632 ;
  assign n55380 = ~n55378 & n55379 ;
  assign n55381 = ~n55375 & ~n55380 ;
  assign n55382 = ~n55361 & n55381 ;
  assign n55383 = ~n55372 & n55382 ;
  assign n55384 = ~\u0_L11_reg[4]/NET0131  & ~n55383 ;
  assign n55385 = \u0_L11_reg[4]/NET0131  & n55383 ;
  assign n55386 = ~n55384 & ~n55385 ;
  assign n55387 = ~n54744 & ~n54782 ;
  assign n55388 = ~n54731 & n55387 ;
  assign n55389 = n54738 & ~n55388 ;
  assign n55390 = n54750 & n54768 ;
  assign n55391 = ~n55389 & ~n55390 ;
  assign n55392 = ~n54760 & ~n55391 ;
  assign n55402 = n54749 & n54779 ;
  assign n55404 = ~n55067 & ~n55402 ;
  assign n55405 = ~n54785 & n55404 ;
  assign n55403 = n54738 & n54789 ;
  assign n55406 = ~n55051 & ~n55403 ;
  assign n55407 = n55405 & n55406 ;
  assign n55408 = n54760 & ~n55407 ;
  assign n55393 = n54730 & n54743 ;
  assign n55394 = ~n55050 & ~n55393 ;
  assign n55395 = ~n54785 & n55394 ;
  assign n55396 = ~n54790 & n55395 ;
  assign n55397 = ~n54738 & ~n55396 ;
  assign n55398 = ~n54765 & ~n55046 ;
  assign n55399 = n54738 & ~n55398 ;
  assign n55400 = ~n54738 & ~n54760 ;
  assign n55401 = n54768 & n55400 ;
  assign n55409 = ~n55399 & ~n55401 ;
  assign n55410 = ~n55397 & n55409 ;
  assign n55411 = ~n55408 & n55410 ;
  assign n55412 = ~n55392 & n55411 ;
  assign n55413 = \u0_L11_reg[15]/P0001  & n55412 ;
  assign n55414 = ~\u0_L11_reg[15]/P0001  & ~n55412 ;
  assign n55415 = ~n55413 & ~n55414 ;
  assign n55416 = ~n54763 & ~n54783 ;
  assign n55417 = ~n55055 & n55416 ;
  assign n55418 = ~n54738 & ~n55417 ;
  assign n55419 = ~n54728 & n54738 ;
  assign n55420 = ~n55387 & n55419 ;
  assign n55421 = ~n54729 & ~n55054 ;
  assign n55422 = ~n54765 & n55421 ;
  assign n55423 = ~n55420 & n55422 ;
  assign n55424 = ~n55418 & n55423 ;
  assign n55425 = n54760 & ~n55424 ;
  assign n55427 = n54738 & ~n54744 ;
  assign n55426 = n54721 & ~n54743 ;
  assign n55428 = ~n55065 & ~n55426 ;
  assign n55429 = n55427 & n55428 ;
  assign n55430 = ~n54788 & ~n55429 ;
  assign n55431 = ~n54760 & ~n55430 ;
  assign n55437 = ~n54738 & ~n54787 ;
  assign n55432 = n54769 & n54779 ;
  assign n55433 = ~n55070 & ~n55432 ;
  assign n55434 = ~n54760 & ~n55433 ;
  assign n55435 = ~n54721 & n54738 ;
  assign n55436 = n54715 & n55435 ;
  assign n55438 = ~n54784 & ~n55436 ;
  assign n55439 = ~n55434 & n55438 ;
  assign n55440 = ~n55437 & n55439 ;
  assign n55441 = ~n55431 & n55440 ;
  assign n55442 = ~n55425 & n55441 ;
  assign n55443 = ~\u0_L11_reg[27]/NET0131  & ~n55442 ;
  assign n55444 = \u0_L11_reg[27]/NET0131  & n55442 ;
  assign n55445 = ~n55443 & ~n55444 ;
  assign n55462 = ~n55166 & n55230 ;
  assign n55463 = ~n55174 & ~n55320 ;
  assign n55464 = ~n55462 & n55463 ;
  assign n55465 = ~n55189 & ~n55464 ;
  assign n55460 = ~n55197 & ~n55334 ;
  assign n55461 = n55189 & ~n55460 ;
  assign n55466 = ~n55182 & ~n55225 ;
  assign n55467 = ~n55461 & n55466 ;
  assign n55468 = ~n55465 & n55467 ;
  assign n55469 = ~n55154 & ~n55468 ;
  assign n55448 = ~n55174 & ~n55222 ;
  assign n55447 = ~n55174 & n55181 ;
  assign n55449 = n55189 & ~n55447 ;
  assign n55450 = ~n55448 & n55449 ;
  assign n55446 = ~n55181 & n55208 ;
  assign n55451 = n55347 & ~n55446 ;
  assign n55452 = ~n55450 & n55451 ;
  assign n55453 = n55154 & ~n55452 ;
  assign n55454 = ~n55189 & ~n55314 ;
  assign n55455 = n55189 & ~n55345 ;
  assign n55456 = n55173 & n55182 ;
  assign n55457 = ~n55333 & ~n55456 ;
  assign n55458 = n55455 & n55457 ;
  assign n55459 = ~n55454 & ~n55458 ;
  assign n55470 = ~n55453 & ~n55459 ;
  assign n55471 = ~n55469 & n55470 ;
  assign n55472 = ~\u0_L11_reg[8]/NET0131  & ~n55471 ;
  assign n55473 = \u0_L11_reg[8]/NET0131  & n55471 ;
  assign n55474 = ~n55472 & ~n55473 ;
  assign n55476 = n54632 & n54672 ;
  assign n55477 = ~n54656 & ~n55476 ;
  assign n55478 = ~n54613 & ~n55477 ;
  assign n55475 = n54613 & n55377 ;
  assign n55479 = n54613 & ~n54632 ;
  assign n55480 = n54675 & ~n55479 ;
  assign n55481 = ~n54632 & n55253 ;
  assign n55482 = ~n55480 & ~n55481 ;
  assign n55483 = ~n55475 & n55482 ;
  assign n55484 = ~n55478 & n55483 ;
  assign n55485 = n54652 & ~n55484 ;
  assign n55488 = n54666 & n55264 ;
  assign n55489 = ~n54632 & ~n55488 ;
  assign n55490 = ~n55377 & n55489 ;
  assign n55486 = n54632 & ~n55253 ;
  assign n55487 = n54668 & n55486 ;
  assign n55491 = ~n54652 & ~n55487 ;
  assign n55492 = ~n55490 & n55491 ;
  assign n55493 = ~n54678 & ~n54680 ;
  assign n55494 = ~n55492 & n55493 ;
  assign n55495 = ~n55485 & n55494 ;
  assign n55496 = ~\u0_L11_reg[19]/NET0131  & ~n55495 ;
  assign n55497 = \u0_L11_reg[19]/NET0131  & n55495 ;
  assign n55498 = ~n55496 & ~n55497 ;
  assign n55499 = ~n54540 & ~n54596 ;
  assign n55500 = ~n54546 & ~n55499 ;
  assign n55501 = ~n54551 & ~n55500 ;
  assign n55502 = ~n54519 & ~n55501 ;
  assign n55503 = ~n55113 & ~n55131 ;
  assign n55504 = n54519 & ~n55503 ;
  assign n55505 = ~n54571 & ~n55121 ;
  assign n55506 = ~n55504 & n55505 ;
  assign n55507 = ~n55502 & n55506 ;
  assign n55508 = n54560 & ~n55507 ;
  assign n55522 = n54577 & n54580 ;
  assign n55523 = ~n54564 & ~n55522 ;
  assign n55524 = ~n55119 & n55523 ;
  assign n55525 = ~n54519 & ~n55524 ;
  assign n55509 = n54525 & n54594 ;
  assign n55510 = ~n55136 & ~n55509 ;
  assign n55511 = ~n54519 & ~n55510 ;
  assign n55512 = n54519 & n54583 ;
  assign n55513 = ~n54531 & ~n54577 ;
  assign n55514 = ~n55512 & n55513 ;
  assign n55515 = n54531 & ~n54562 ;
  assign n55516 = ~n54570 & n55515 ;
  assign n55517 = ~n55514 & ~n55516 ;
  assign n55518 = ~n55511 & ~n55517 ;
  assign n55519 = ~n54560 & ~n55518 ;
  assign n55520 = ~n54549 & ~n54596 ;
  assign n55521 = n54572 & ~n55520 ;
  assign n55526 = ~n55519 & ~n55521 ;
  assign n55527 = ~n55525 & n55526 ;
  assign n55528 = ~n55508 & n55527 ;
  assign n55529 = \u0_L11_reg[23]/NET0131  & ~n55528 ;
  assign n55530 = ~\u0_L11_reg[23]/NET0131  & n55528 ;
  assign n55531 = ~n55529 & ~n55530 ;
  assign n55532 = n54985 & n55304 ;
  assign n55533 = ~n54988 & ~n55532 ;
  assign n55534 = ~n54971 & ~n54985 ;
  assign n55535 = ~n54965 & n55534 ;
  assign n55536 = n54978 & n55535 ;
  assign n55537 = ~n55026 & ~n55033 ;
  assign n55538 = ~n55536 & n55537 ;
  assign n55539 = ~n55002 & ~n55538 ;
  assign n55540 = n55533 & ~n55539 ;
  assign n55541 = ~n54995 & ~n55540 ;
  assign n55542 = n54965 & n55534 ;
  assign n55543 = n55011 & ~n55542 ;
  assign n55544 = n54995 & ~n55032 ;
  assign n55545 = ~n55535 & n55544 ;
  assign n55546 = ~n55543 & ~n55545 ;
  assign n55547 = n54971 & n55013 ;
  assign n55548 = n55002 & ~n55547 ;
  assign n55549 = n55284 & n55548 ;
  assign n55550 = n55533 & n55549 ;
  assign n55551 = ~n55546 & n55550 ;
  assign n55555 = n55005 & ~n55304 ;
  assign n55554 = n54971 & ~n55005 ;
  assign n55556 = n54995 & ~n55554 ;
  assign n55557 = ~n55555 & n55556 ;
  assign n55558 = ~n54978 & ~n55280 ;
  assign n55559 = n55281 & n55558 ;
  assign n55552 = n54965 & ~n54986 ;
  assign n55553 = n55022 & n55552 ;
  assign n55560 = ~n55002 & ~n55553 ;
  assign n55561 = ~n55559 & n55560 ;
  assign n55562 = ~n55557 & n55561 ;
  assign n55563 = ~n55551 & ~n55562 ;
  assign n55564 = ~n55541 & ~n55563 ;
  assign n55565 = ~\u0_L11_reg[13]/NET0131  & n55564 ;
  assign n55566 = \u0_L11_reg[13]/NET0131  & ~n55564 ;
  assign n55567 = ~n55565 & ~n55566 ;
  assign n55602 = decrypt_pad & ~\u0_uk_K_r11_reg[12]/NET0131  ;
  assign n55603 = ~decrypt_pad & ~\u0_uk_K_r11_reg[17]/NET0131  ;
  assign n55604 = ~n55602 & ~n55603 ;
  assign n55605 = \u0_R11_reg[11]/P0001  & ~n55604 ;
  assign n55606 = ~\u0_R11_reg[11]/P0001  & n55604 ;
  assign n55607 = ~n55605 & ~n55606 ;
  assign n55568 = decrypt_pad & ~\u0_uk_K_r11_reg[27]/P0001  ;
  assign n55569 = ~decrypt_pad & ~\u0_uk_K_r11_reg[32]/NET0131  ;
  assign n55570 = ~n55568 & ~n55569 ;
  assign n55571 = \u0_R11_reg[12]/NET0131  & ~n55570 ;
  assign n55572 = ~\u0_R11_reg[12]/NET0131  & n55570 ;
  assign n55573 = ~n55571 & ~n55572 ;
  assign n55581 = decrypt_pad & ~\u0_uk_K_r11_reg[40]/NET0131  ;
  assign n55582 = ~decrypt_pad & ~\u0_uk_K_r11_reg[20]/NET0131  ;
  assign n55583 = ~n55581 & ~n55582 ;
  assign n55584 = \u0_R11_reg[13]/NET0131  & ~n55583 ;
  assign n55585 = ~\u0_R11_reg[13]/NET0131  & n55583 ;
  assign n55586 = ~n55584 & ~n55585 ;
  assign n55594 = decrypt_pad & ~\u0_uk_K_r11_reg[3]/NET0131  ;
  assign n55595 = ~decrypt_pad & ~\u0_uk_K_r11_reg[40]/NET0131  ;
  assign n55596 = ~n55594 & ~n55595 ;
  assign n55597 = \u0_R11_reg[9]/NET0131  & ~n55596 ;
  assign n55598 = ~\u0_R11_reg[9]/NET0131  & n55596 ;
  assign n55599 = ~n55597 & ~n55598 ;
  assign n55610 = n55586 & ~n55599 ;
  assign n55574 = decrypt_pad & ~\u0_uk_K_r11_reg[11]/NET0131  ;
  assign n55575 = ~decrypt_pad & ~\u0_uk_K_r11_reg[48]/NET0131  ;
  assign n55576 = ~n55574 & ~n55575 ;
  assign n55577 = \u0_R11_reg[10]/NET0131  & ~n55576 ;
  assign n55578 = ~\u0_R11_reg[10]/NET0131  & n55576 ;
  assign n55579 = ~n55577 & ~n55578 ;
  assign n55587 = decrypt_pad & ~\u0_uk_K_r11_reg[6]/NET0131  ;
  assign n55588 = ~decrypt_pad & ~\u0_uk_K_r11_reg[11]/NET0131  ;
  assign n55589 = ~n55587 & ~n55588 ;
  assign n55590 = \u0_R11_reg[8]/NET0131  & ~n55589 ;
  assign n55591 = ~\u0_R11_reg[8]/NET0131  & n55589 ;
  assign n55592 = ~n55590 & ~n55591 ;
  assign n55611 = n55586 & ~n55592 ;
  assign n55612 = n55579 & n55611 ;
  assign n55613 = ~n55586 & n55592 ;
  assign n55614 = n55599 & n55613 ;
  assign n55615 = ~n55612 & ~n55614 ;
  assign n55616 = ~n55610 & n55615 ;
  assign n55617 = n55573 & ~n55616 ;
  assign n55593 = ~n55586 & ~n55592 ;
  assign n55608 = ~n55579 & ~n55599 ;
  assign n55609 = n55593 & n55608 ;
  assign n55618 = n55579 & ~n55599 ;
  assign n55619 = n55586 & n55618 ;
  assign n55620 = ~n55609 & ~n55619 ;
  assign n55621 = ~n55617 & n55620 ;
  assign n55622 = n55607 & ~n55621 ;
  assign n55625 = ~n55579 & n55599 ;
  assign n55626 = ~n55618 & ~n55625 ;
  assign n55623 = n55586 & n55592 ;
  assign n55624 = ~n55593 & ~n55623 ;
  assign n55627 = ~n55592 & n55607 ;
  assign n55631 = n55624 & ~n55627 ;
  assign n55632 = n55626 & ~n55631 ;
  assign n55628 = n55599 & n55627 ;
  assign n55629 = n55624 & ~n55626 ;
  assign n55630 = ~n55628 & n55629 ;
  assign n55633 = ~n55573 & ~n55630 ;
  assign n55634 = ~n55632 & n55633 ;
  assign n55580 = n55573 & n55579 ;
  assign n55600 = n55593 & n55599 ;
  assign n55601 = n55580 & n55600 ;
  assign n55636 = n55592 & ~n55610 ;
  assign n55637 = ~n55625 & ~n55636 ;
  assign n55635 = ~n55586 & n55599 ;
  assign n55638 = n55573 & ~n55607 ;
  assign n55639 = ~n55635 & n55638 ;
  assign n55640 = ~n55637 & n55639 ;
  assign n55641 = ~n55601 & ~n55640 ;
  assign n55642 = ~n55634 & n55641 ;
  assign n55643 = ~n55622 & n55642 ;
  assign n55644 = ~\u0_L11_reg[6]/NET0131  & ~n55643 ;
  assign n55645 = \u0_L11_reg[6]/NET0131  & n55643 ;
  assign n55646 = ~n55644 & ~n55645 ;
  assign n55647 = n54433 & ~n54452 ;
  assign n55648 = n54439 & n55647 ;
  assign n55651 = n54463 & ~n55648 ;
  assign n55649 = ~n54433 & n54467 ;
  assign n55650 = ~n54446 & n54500 ;
  assign n55652 = ~n55649 & ~n55650 ;
  assign n55653 = n55651 & n55652 ;
  assign n55654 = ~n54464 & ~n54500 ;
  assign n55655 = n54471 & n55654 ;
  assign n55656 = ~n54463 & ~n55099 ;
  assign n55657 = ~n55096 & n55656 ;
  assign n55658 = ~n55655 & n55657 ;
  assign n55659 = ~n55653 & ~n55658 ;
  assign n55660 = n55085 & n55647 ;
  assign n55661 = ~n55659 & ~n55660 ;
  assign n55662 = n54427 & ~n55661 ;
  assign n55667 = ~n54467 & ~n54486 ;
  assign n55668 = ~n55650 & n55667 ;
  assign n55669 = ~n54463 & ~n55668 ;
  assign n55663 = ~n54446 & ~n54463 ;
  assign n55664 = n54439 & ~n55647 ;
  assign n55665 = ~n55663 & n55664 ;
  assign n55666 = ~n55649 & n55665 ;
  assign n55670 = n54502 & ~n55666 ;
  assign n55671 = ~n55669 & n55670 ;
  assign n55672 = ~n54427 & ~n55671 ;
  assign n55673 = n54457 & n54463 ;
  assign n55674 = ~n54474 & n54484 ;
  assign n55675 = n54483 & n55674 ;
  assign n55676 = ~n55673 & ~n55675 ;
  assign n55677 = ~n55672 & n55676 ;
  assign n55678 = ~n55662 & n55677 ;
  assign n55679 = \u0_L11_reg[32]/NET0131  & n55678 ;
  assign n55680 = ~\u0_L11_reg[32]/NET0131  & ~n55678 ;
  assign n55681 = ~n55679 & ~n55680 ;
  assign n55684 = ~n54439 & ~n54473 ;
  assign n55682 = ~n54446 & ~n54482 ;
  assign n55683 = n55654 & ~n55682 ;
  assign n55685 = n54427 & ~n54463 ;
  assign n55686 = ~n55683 & n55685 ;
  assign n55687 = ~n55684 & n55686 ;
  assign n55688 = ~n54433 & ~n55654 ;
  assign n55689 = ~n54453 & n55688 ;
  assign n55690 = n54472 & n55654 ;
  assign n55691 = ~n54427 & n54463 ;
  assign n55692 = ~n55685 & ~n55691 ;
  assign n55693 = ~n54487 & n55692 ;
  assign n55694 = ~n55690 & n55693 ;
  assign n55695 = ~n55689 & n55694 ;
  assign n55696 = ~n55687 & ~n55695 ;
  assign n55697 = ~n55096 & ~n55696 ;
  assign n55698 = ~n54465 & ~n55688 ;
  assign n55699 = ~n55690 & n55698 ;
  assign n55700 = n54463 & n55104 ;
  assign n55701 = ~n55699 & n55700 ;
  assign n55702 = ~n55697 & ~n55701 ;
  assign n55703 = ~\u0_L11_reg[7]/NET0131  & n55702 ;
  assign n55704 = \u0_L11_reg[7]/NET0131  & ~n55702 ;
  assign n55705 = ~n55703 & ~n55704 ;
  assign n55720 = n55607 & ~n55611 ;
  assign n55721 = ~n55631 & ~n55720 ;
  assign n55722 = n55608 & ~n55721 ;
  assign n55723 = ~n55607 & ~n55608 ;
  assign n55724 = ~n55624 & n55723 ;
  assign n55725 = ~n55722 & ~n55724 ;
  assign n55726 = n55573 & ~n55725 ;
  assign n55709 = n55579 & n55593 ;
  assign n55710 = ~n55579 & n55611 ;
  assign n55711 = ~n55709 & ~n55710 ;
  assign n55712 = n55592 & n55618 ;
  assign n55713 = ~n55600 & ~n55712 ;
  assign n55714 = n55711 & n55713 ;
  assign n55715 = n55607 & ~n55714 ;
  assign n55716 = ~n55599 & n55613 ;
  assign n55717 = n55579 & n55716 ;
  assign n55718 = ~n55715 & ~n55717 ;
  assign n55719 = ~n55573 & ~n55718 ;
  assign n55727 = n55599 & n55611 ;
  assign n55728 = ~n55716 & ~n55727 ;
  assign n55729 = ~n55579 & ~n55728 ;
  assign n55730 = n55579 & n55592 ;
  assign n55731 = n55599 & n55730 ;
  assign n55732 = ~n55612 & ~n55731 ;
  assign n55733 = n55573 & ~n55732 ;
  assign n55734 = ~n55729 & ~n55733 ;
  assign n55735 = n55607 & ~n55734 ;
  assign n55706 = n55599 & n55623 ;
  assign n55707 = n55579 & ~n55607 ;
  assign n55708 = n55706 & n55707 ;
  assign n55736 = n55608 & ~n55624 ;
  assign n55737 = n55615 & ~n55736 ;
  assign n55738 = ~n55573 & ~n55607 ;
  assign n55739 = ~n55737 & n55738 ;
  assign n55740 = ~n55708 & ~n55739 ;
  assign n55741 = ~n55735 & n55740 ;
  assign n55742 = ~n55719 & n55741 ;
  assign n55743 = ~n55726 & n55742 ;
  assign n55744 = ~\u0_L11_reg[24]/NET0131  & ~n55743 ;
  assign n55745 = \u0_L11_reg[24]/NET0131  & n55743 ;
  assign n55746 = ~n55744 & ~n55745 ;
  assign n55750 = n55608 & n55613 ;
  assign n55751 = n55711 & ~n55750 ;
  assign n55752 = n55607 & ~n55751 ;
  assign n55748 = ~n55600 & ~n55730 ;
  assign n55749 = ~n55607 & ~n55748 ;
  assign n55753 = n55573 & ~n55749 ;
  assign n55754 = ~n55752 & n55753 ;
  assign n55757 = ~n55635 & n55730 ;
  assign n55756 = ~n55586 & n55625 ;
  assign n55758 = n55607 & ~n55756 ;
  assign n55759 = ~n55757 & n55758 ;
  assign n55760 = ~n55579 & n55592 ;
  assign n55761 = ~n55635 & n55760 ;
  assign n55762 = ~n55607 & ~n55727 ;
  assign n55763 = ~n55761 & n55762 ;
  assign n55764 = ~n55759 & ~n55763 ;
  assign n55755 = ~n55599 & n55612 ;
  assign n55765 = ~n55573 & ~n55736 ;
  assign n55766 = ~n55755 & n55765 ;
  assign n55767 = ~n55764 & n55766 ;
  assign n55768 = ~n55754 & ~n55767 ;
  assign n55771 = n55607 & n55618 ;
  assign n55772 = n55623 & n55771 ;
  assign n55747 = n55635 & n55707 ;
  assign n55769 = n55580 & n55599 ;
  assign n55770 = ~n55623 & n55769 ;
  assign n55773 = ~n55747 & ~n55770 ;
  assign n55774 = ~n55772 & n55773 ;
  assign n55775 = ~n55768 & n55774 ;
  assign n55776 = \u0_L11_reg[30]/NET0131  & ~n55775 ;
  assign n55777 = ~\u0_L11_reg[30]/NET0131  & n55775 ;
  assign n55778 = ~n55776 & ~n55777 ;
  assign n55794 = ~n55166 & n55216 ;
  assign n55795 = n55166 & n55230 ;
  assign n55796 = ~n55794 & ~n55795 ;
  assign n55797 = n55189 & ~n55796 ;
  assign n55793 = ~n55189 & n55320 ;
  assign n55798 = ~n55231 & ~n55314 ;
  assign n55799 = ~n55793 & n55798 ;
  assign n55800 = ~n55797 & n55799 ;
  assign n55801 = n55154 & ~n55800 ;
  assign n55779 = ~n55334 & n55455 ;
  assign n55780 = ~n55181 & n55224 ;
  assign n55781 = ~n55447 & ~n55780 ;
  assign n55782 = ~n55189 & ~n55781 ;
  assign n55783 = ~n55779 & ~n55782 ;
  assign n55784 = ~n55223 & ~n55462 ;
  assign n55785 = n55189 & ~n55784 ;
  assign n55787 = n55173 & ~n55198 ;
  assign n55788 = n55166 & ~n55787 ;
  assign n55786 = n55189 & ~n55207 ;
  assign n55789 = ~n55462 & ~n55786 ;
  assign n55790 = ~n55788 & n55789 ;
  assign n55791 = ~n55785 & ~n55790 ;
  assign n55792 = ~n55154 & ~n55791 ;
  assign n55802 = ~n55783 & ~n55792 ;
  assign n55803 = ~n55801 & n55802 ;
  assign n55804 = ~\u0_L11_reg[3]/NET0131  & ~n55803 ;
  assign n55805 = \u0_L11_reg[3]/NET0131  & n55803 ;
  assign n55806 = ~n55804 & ~n55805 ;
  assign n55821 = n55138 & ~n55500 ;
  assign n55822 = n54525 & ~n55821 ;
  assign n55811 = ~n54569 & ~n55113 ;
  assign n55820 = n54572 & ~n55811 ;
  assign n55823 = ~n55119 & ~n55820 ;
  assign n55824 = ~n55822 & n55823 ;
  assign n55825 = n54560 & ~n55824 ;
  assign n55807 = ~n54525 & n55137 ;
  assign n55808 = ~n54546 & n54563 ;
  assign n55809 = ~n55807 & ~n55808 ;
  assign n55810 = ~n54519 & ~n55809 ;
  assign n55813 = ~n55115 & n55499 ;
  assign n55814 = n54519 & ~n55813 ;
  assign n55815 = n54525 & n55132 ;
  assign n55812 = ~n54519 & ~n55811 ;
  assign n55816 = ~n55807 & ~n55812 ;
  assign n55817 = ~n55815 & n55816 ;
  assign n55818 = ~n55814 & n55817 ;
  assign n55819 = ~n54560 & ~n55818 ;
  assign n55826 = ~n55810 & ~n55819 ;
  assign n55827 = ~n55825 & n55826 ;
  assign n55828 = ~\u0_L11_reg[9]/NET0131  & ~n55827 ;
  assign n55829 = \u0_L11_reg[9]/NET0131  & n55827 ;
  assign n55830 = ~n55828 & ~n55829 ;
  assign n55837 = ~n55599 & ~n55623 ;
  assign n55838 = ~n55593 & ~n55706 ;
  assign n55839 = ~n55837 & n55838 ;
  assign n55840 = n55607 & n55839 ;
  assign n55833 = ~n55599 & n55611 ;
  assign n55832 = ~n55579 & n55593 ;
  assign n55834 = ~n55706 & ~n55832 ;
  assign n55835 = ~n55833 & n55834 ;
  assign n55836 = ~n55607 & ~n55835 ;
  assign n55841 = ~n55609 & ~n55836 ;
  assign n55842 = ~n55840 & n55841 ;
  assign n55843 = ~n55573 & ~n55842 ;
  assign n55848 = n55599 & n55607 ;
  assign n55849 = n55593 & ~n55848 ;
  assign n55850 = ~n55579 & ~n55849 ;
  assign n55851 = ~n55839 & n55850 ;
  assign n55844 = ~n55579 & n55613 ;
  assign n55845 = ~n55709 & ~n55844 ;
  assign n55846 = ~n55607 & ~n55845 ;
  assign n55847 = n55579 & n55727 ;
  assign n55852 = ~n55846 & ~n55847 ;
  assign n55853 = ~n55851 & n55852 ;
  assign n55854 = n55573 & ~n55853 ;
  assign n55831 = ~n55607 & n55712 ;
  assign n55855 = n55593 & n55618 ;
  assign n55856 = ~n55586 & n55731 ;
  assign n55857 = ~n55855 & ~n55856 ;
  assign n55858 = n55607 & ~n55857 ;
  assign n55859 = ~n55831 & ~n55858 ;
  assign n55860 = ~n55854 & n55859 ;
  assign n55861 = ~n55843 & n55860 ;
  assign n55862 = ~\u0_L11_reg[16]/NET0131  & ~n55861 ;
  assign n55863 = \u0_L11_reg[16]/NET0131  & n55861 ;
  assign n55864 = ~n55862 & ~n55863 ;
  assign n55881 = n55002 & n55287 ;
  assign n55882 = n54965 & n55004 ;
  assign n55883 = ~n55547 & ~n55882 ;
  assign n55884 = ~n55881 & n55883 ;
  assign n55885 = n54995 & ~n55884 ;
  assign n55869 = ~n54972 & ~n54978 ;
  assign n55868 = n54965 & n54995 ;
  assign n55870 = ~n55274 & ~n55868 ;
  assign n55871 = n55869 & n55870 ;
  assign n55867 = n54987 & ~n55028 ;
  assign n55866 = n55273 & n55289 ;
  assign n55872 = ~n55535 & ~n55866 ;
  assign n55873 = ~n55867 & n55872 ;
  assign n55874 = ~n55871 & n55873 ;
  assign n55875 = ~n55002 & ~n55874 ;
  assign n55865 = n55002 & n55303 ;
  assign n55876 = ~n55281 & ~n55534 ;
  assign n55877 = n54978 & n55002 ;
  assign n55878 = ~n55876 & n55877 ;
  assign n55879 = ~n55015 & ~n55878 ;
  assign n55880 = ~n54995 & ~n55879 ;
  assign n55886 = ~n55865 & ~n55880 ;
  assign n55887 = ~n55875 & n55886 ;
  assign n55888 = ~n55885 & n55887 ;
  assign n55889 = \u0_L11_reg[18]/NET0131  & n55888 ;
  assign n55890 = ~\u0_L11_reg[18]/NET0131  & ~n55888 ;
  assign n55891 = ~n55889 & ~n55890 ;
  assign n55892 = decrypt_pad & ~\u0_uk_K_r10_reg[5]/NET0131  ;
  assign n55893 = ~decrypt_pad & ~\u0_uk_K_r10_reg[39]/NET0131  ;
  assign n55894 = ~n55892 & ~n55893 ;
  assign n55895 = \u0_R10_reg[4]/NET0131  & ~n55894 ;
  assign n55896 = ~\u0_R10_reg[4]/NET0131  & n55894 ;
  assign n55897 = ~n55895 & ~n55896 ;
  assign n55911 = decrypt_pad & ~\u0_uk_K_r10_reg[39]/NET0131  ;
  assign n55912 = ~decrypt_pad & ~\u0_uk_K_r10_reg[48]/NET0131  ;
  assign n55913 = ~n55911 & ~n55912 ;
  assign n55914 = \u0_R10_reg[32]/NET0131  & ~n55913 ;
  assign n55915 = ~\u0_R10_reg[32]/NET0131  & n55913 ;
  assign n55916 = ~n55914 & ~n55915 ;
  assign n55917 = decrypt_pad & ~\u0_uk_K_r10_reg[33]/NET0131  ;
  assign n55918 = ~decrypt_pad & ~\u0_uk_K_r10_reg[10]/NET0131  ;
  assign n55919 = ~n55917 & ~n55918 ;
  assign n55920 = \u0_R10_reg[5]/NET0131  & ~n55919 ;
  assign n55921 = ~\u0_R10_reg[5]/NET0131  & n55919 ;
  assign n55922 = ~n55920 & ~n55921 ;
  assign n55924 = ~n55916 & ~n55922 ;
  assign n55898 = decrypt_pad & ~\u0_uk_K_r10_reg[27]/NET0131  ;
  assign n55899 = ~decrypt_pad & ~\u0_uk_K_r10_reg[4]/NET0131  ;
  assign n55900 = ~n55898 & ~n55899 ;
  assign n55901 = \u0_R10_reg[3]/NET0131  & ~n55900 ;
  assign n55902 = ~\u0_R10_reg[3]/NET0131  & n55900 ;
  assign n55903 = ~n55901 & ~n55902 ;
  assign n55904 = decrypt_pad & ~\u0_uk_K_r10_reg[18]/NET0131  ;
  assign n55905 = ~decrypt_pad & ~\u0_uk_K_r10_reg[27]/NET0131  ;
  assign n55906 = ~n55904 & ~n55905 ;
  assign n55907 = \u0_R10_reg[2]/NET0131  & ~n55906 ;
  assign n55908 = ~\u0_R10_reg[2]/NET0131  & n55906 ;
  assign n55909 = ~n55907 & ~n55908 ;
  assign n55934 = ~n55909 & ~n55916 ;
  assign n55955 = n55903 & n55934 ;
  assign n55925 = decrypt_pad & ~\u0_uk_K_r10_reg[3]/NET0131  ;
  assign n55926 = ~decrypt_pad & ~\u0_uk_K_r10_reg[12]/NET0131  ;
  assign n55927 = ~n55925 & ~n55926 ;
  assign n55928 = \u0_R10_reg[1]/NET0131  & ~n55927 ;
  assign n55929 = ~\u0_R10_reg[1]/NET0131  & n55927 ;
  assign n55930 = ~n55928 & ~n55929 ;
  assign n55937 = ~n55922 & ~n55930 ;
  assign n55953 = ~n55909 & n55937 ;
  assign n55954 = ~n55916 & ~n55930 ;
  assign n55956 = ~n55953 & ~n55954 ;
  assign n55957 = ~n55955 & n55956 ;
  assign n55958 = ~n55924 & ~n55957 ;
  assign n55935 = n55922 & ~n55930 ;
  assign n55959 = n55909 & n55924 ;
  assign n55960 = ~n55935 & ~n55959 ;
  assign n55961 = n55903 & ~n55960 ;
  assign n55951 = ~n55903 & n55916 ;
  assign n55952 = n55930 & n55951 ;
  assign n55962 = n55909 & n55954 ;
  assign n55963 = ~n55952 & ~n55962 ;
  assign n55964 = ~n55961 & n55963 ;
  assign n55965 = ~n55958 & n55964 ;
  assign n55966 = n55897 & ~n55965 ;
  assign n55923 = n55916 & n55922 ;
  assign n55942 = ~n55903 & n55930 ;
  assign n55943 = n55923 & ~n55942 ;
  assign n55944 = ~n55922 & n55930 ;
  assign n55945 = ~n55916 & n55944 ;
  assign n55946 = ~n55943 & ~n55945 ;
  assign n55947 = ~n55909 & ~n55946 ;
  assign n55910 = n55903 & n55909 ;
  assign n55931 = ~n55924 & n55930 ;
  assign n55932 = ~n55923 & n55931 ;
  assign n55933 = n55910 & n55932 ;
  assign n55936 = n55934 & ~n55935 ;
  assign n55938 = n55909 & n55916 ;
  assign n55939 = n55937 & n55938 ;
  assign n55940 = ~n55936 & ~n55939 ;
  assign n55941 = ~n55903 & ~n55940 ;
  assign n55948 = ~n55933 & ~n55941 ;
  assign n55949 = ~n55947 & n55948 ;
  assign n55950 = ~n55897 & ~n55949 ;
  assign n55970 = n55909 & n55922 ;
  assign n55971 = n55930 & n55970 ;
  assign n55972 = n55916 & n55971 ;
  assign n55973 = ~n55944 & ~n55970 ;
  assign n55974 = n55909 & ~n55954 ;
  assign n55975 = ~n55973 & ~n55974 ;
  assign n55976 = ~n55972 & ~n55975 ;
  assign n55977 = ~n55903 & ~n55976 ;
  assign n55967 = ~n55909 & ~n55930 ;
  assign n55968 = n55903 & n55916 ;
  assign n55969 = n55967 & n55968 ;
  assign n55978 = n55910 & ~n55930 ;
  assign n55979 = n55924 & n55978 ;
  assign n55980 = ~n55969 & ~n55979 ;
  assign n55981 = ~n55977 & n55980 ;
  assign n55982 = ~n55950 & n55981 ;
  assign n55983 = ~n55966 & n55982 ;
  assign n55984 = ~\u0_L10_reg[31]/NET0131  & ~n55983 ;
  assign n55985 = \u0_L10_reg[31]/NET0131  & n55983 ;
  assign n55986 = ~n55984 & ~n55985 ;
  assign n55993 = decrypt_pad & ~\u0_uk_K_r10_reg[16]/NET0131  ;
  assign n55994 = ~decrypt_pad & ~\u0_uk_K_r10_reg[21]/NET0131  ;
  assign n55995 = ~n55993 & ~n55994 ;
  assign n55996 = \u0_R10_reg[26]/NET0131  & ~n55995 ;
  assign n55997 = ~\u0_R10_reg[26]/NET0131  & n55995 ;
  assign n55998 = ~n55996 & ~n55997 ;
  assign n56001 = decrypt_pad & ~\u0_uk_K_r10_reg[0]/NET0131  ;
  assign n56002 = ~decrypt_pad & ~\u0_uk_K_r10_reg[36]/NET0131  ;
  assign n56003 = ~n56001 & ~n56002 ;
  assign n56004 = \u0_R10_reg[25]/NET0131  & ~n56003 ;
  assign n56005 = ~\u0_R10_reg[25]/NET0131  & n56003 ;
  assign n56006 = ~n56004 & ~n56005 ;
  assign n55987 = decrypt_pad & ~\u0_uk_K_r10_reg[51]/NET0131  ;
  assign n55988 = ~decrypt_pad & ~\u0_uk_K_r10_reg[1]/NET0131  ;
  assign n55989 = ~n55987 & ~n55988 ;
  assign n55990 = \u0_R10_reg[24]/NET0131  & ~n55989 ;
  assign n55991 = ~\u0_R10_reg[24]/NET0131  & n55989 ;
  assign n55992 = ~n55990 & ~n55991 ;
  assign n56009 = decrypt_pad & ~\u0_uk_K_r10_reg[28]/NET0131  ;
  assign n56010 = ~decrypt_pad & ~\u0_uk_K_r10_reg[9]/NET0131  ;
  assign n56011 = ~n56009 & ~n56010 ;
  assign n56012 = \u0_R10_reg[29]/NET0131  & ~n56011 ;
  assign n56013 = ~\u0_R10_reg[29]/NET0131  & n56011 ;
  assign n56014 = ~n56012 & ~n56013 ;
  assign n56015 = n55992 & n56014 ;
  assign n56016 = ~n56006 & n56015 ;
  assign n56017 = ~n55998 & n56016 ;
  assign n56018 = ~n55992 & n56014 ;
  assign n56019 = n56006 & n56018 ;
  assign n56020 = ~n56017 & ~n56019 ;
  assign n56021 = decrypt_pad & ~\u0_uk_K_r10_reg[36]/NET0131  ;
  assign n56022 = ~decrypt_pad & ~\u0_uk_K_r10_reg[45]/P0001  ;
  assign n56023 = ~n56021 & ~n56022 ;
  assign n56024 = \u0_R10_reg[28]/NET0131  & ~n56023 ;
  assign n56025 = ~\u0_R10_reg[28]/NET0131  & n56023 ;
  assign n56026 = ~n56024 & ~n56025 ;
  assign n56027 = ~n56020 & n56026 ;
  assign n56000 = n55992 & ~n55998 ;
  assign n55999 = ~n55992 & n55998 ;
  assign n56007 = ~n55999 & n56006 ;
  assign n56008 = ~n56000 & n56007 ;
  assign n56028 = decrypt_pad & ~\u0_uk_K_r10_reg[49]/NET0131  ;
  assign n56029 = ~decrypt_pad & ~\u0_uk_K_r10_reg[30]/NET0131  ;
  assign n56030 = ~n56028 & ~n56029 ;
  assign n56031 = \u0_R10_reg[27]/NET0131  & ~n56030 ;
  assign n56032 = ~\u0_R10_reg[27]/NET0131  & n56030 ;
  assign n56033 = ~n56031 & ~n56032 ;
  assign n56034 = ~n56008 & ~n56033 ;
  assign n56035 = ~n56027 & n56034 ;
  assign n56036 = n55998 & ~n56006 ;
  assign n56037 = n56018 & n56036 ;
  assign n56038 = n55999 & n56006 ;
  assign n56039 = ~n56014 & n56038 ;
  assign n56040 = ~n56037 & ~n56039 ;
  assign n56041 = ~n56006 & ~n56014 ;
  assign n56042 = ~n55999 & n56041 ;
  assign n56043 = n56033 & ~n56042 ;
  assign n56044 = n56040 & n56043 ;
  assign n56045 = ~n56035 & ~n56044 ;
  assign n56055 = n56018 & ~n56033 ;
  assign n56051 = n55992 & ~n56014 ;
  assign n56056 = n55992 & n56033 ;
  assign n56057 = ~n56051 & ~n56056 ;
  assign n56058 = ~n56006 & ~n56057 ;
  assign n56059 = ~n56055 & ~n56058 ;
  assign n56060 = ~n55998 & ~n56059 ;
  assign n56046 = n55998 & n56015 ;
  assign n56052 = ~n56033 & n56051 ;
  assign n56053 = ~n56046 & ~n56052 ;
  assign n56054 = n56006 & ~n56053 ;
  assign n56047 = ~n55992 & ~n56014 ;
  assign n56048 = n56036 & n56047 ;
  assign n56049 = ~n56046 & ~n56048 ;
  assign n56050 = ~n56033 & ~n56049 ;
  assign n56061 = n56006 & n56014 ;
  assign n56062 = ~n55998 & n56061 ;
  assign n56063 = ~n55992 & n56062 ;
  assign n56064 = ~n56026 & ~n56063 ;
  assign n56065 = ~n56050 & n56064 ;
  assign n56066 = ~n56054 & n56065 ;
  assign n56067 = ~n56060 & n56066 ;
  assign n56071 = ~n56036 & ~n56062 ;
  assign n56072 = n56056 & ~n56071 ;
  assign n56068 = ~n55998 & ~n56006 ;
  assign n56069 = ~n55992 & n56068 ;
  assign n56070 = ~n56014 & n56069 ;
  assign n56073 = n56026 & ~n56037 ;
  assign n56074 = ~n56070 & n56073 ;
  assign n56075 = ~n56072 & n56074 ;
  assign n56076 = ~n56067 & ~n56075 ;
  assign n56077 = ~n56045 & ~n56076 ;
  assign n56078 = ~\u0_L10_reg[22]/NET0131  & ~n56077 ;
  assign n56079 = \u0_L10_reg[22]/NET0131  & n56077 ;
  assign n56080 = ~n56078 & ~n56079 ;
  assign n56137 = decrypt_pad & ~\u0_uk_K_r10_reg[29]/NET0131  ;
  assign n56138 = ~decrypt_pad & ~\u0_uk_K_r10_reg[38]/NET0131  ;
  assign n56139 = ~n56137 & ~n56138 ;
  assign n56140 = \u0_R10_reg[24]/NET0131  & ~n56139 ;
  assign n56141 = ~\u0_R10_reg[24]/NET0131  & n56139 ;
  assign n56142 = ~n56140 & ~n56141 ;
  assign n56081 = decrypt_pad & ~\u0_uk_K_r10_reg[31]/NET0131  ;
  assign n56082 = ~decrypt_pad & ~\u0_uk_K_r10_reg[8]/NET0131  ;
  assign n56083 = ~n56081 & ~n56082 ;
  assign n56084 = \u0_R10_reg[23]/NET0131  & ~n56083 ;
  assign n56085 = ~\u0_R10_reg[23]/NET0131  & n56083 ;
  assign n56086 = ~n56084 & ~n56085 ;
  assign n56087 = decrypt_pad & ~\u0_uk_K_r10_reg[14]/NET0131  ;
  assign n56088 = ~decrypt_pad & ~\u0_uk_K_r10_reg[50]/NET0131  ;
  assign n56089 = ~n56087 & ~n56088 ;
  assign n56090 = \u0_R10_reg[22]/NET0131  & ~n56089 ;
  assign n56091 = ~\u0_R10_reg[22]/NET0131  & n56089 ;
  assign n56092 = ~n56090 & ~n56091 ;
  assign n56094 = decrypt_pad & ~\u0_uk_K_r10_reg[8]/NET0131  ;
  assign n56095 = ~decrypt_pad & ~\u0_uk_K_r10_reg[44]/NET0131  ;
  assign n56096 = ~n56094 & ~n56095 ;
  assign n56097 = \u0_R10_reg[20]/NET0131  & ~n56096 ;
  assign n56098 = ~\u0_R10_reg[20]/NET0131  & n56096 ;
  assign n56099 = ~n56097 & ~n56098 ;
  assign n56100 = decrypt_pad & ~\u0_uk_K_r10_reg[23]/NET0131  ;
  assign n56101 = ~decrypt_pad & ~\u0_uk_K_r10_reg[28]/NET0131  ;
  assign n56102 = ~n56100 & ~n56101 ;
  assign n56103 = \u0_R10_reg[21]/NET0131  & ~n56102 ;
  assign n56104 = ~\u0_R10_reg[21]/NET0131  & n56102 ;
  assign n56105 = ~n56103 & ~n56104 ;
  assign n56120 = ~n56099 & n56105 ;
  assign n56121 = n56092 & n56120 ;
  assign n56147 = ~n56092 & n56099 ;
  assign n56160 = n56105 & n56147 ;
  assign n56161 = ~n56121 & ~n56160 ;
  assign n56162 = ~n56086 & ~n56161 ;
  assign n56093 = ~n56086 & ~n56092 ;
  assign n56107 = decrypt_pad & ~\u0_uk_K_r10_reg[52]/NET0131  ;
  assign n56108 = ~decrypt_pad & ~\u0_uk_K_r10_reg[29]/NET0131  ;
  assign n56109 = ~n56107 & ~n56108 ;
  assign n56110 = \u0_R10_reg[25]/NET0131  & ~n56109 ;
  assign n56111 = ~\u0_R10_reg[25]/NET0131  & n56109 ;
  assign n56112 = ~n56110 & ~n56111 ;
  assign n56114 = n56099 & ~n56112 ;
  assign n56156 = n56093 & n56114 ;
  assign n56152 = n56092 & n56099 ;
  assign n56157 = n56112 & n56152 ;
  assign n56158 = ~n56105 & n56157 ;
  assign n56159 = ~n56156 & ~n56158 ;
  assign n56145 = n56105 & ~n56112 ;
  assign n56146 = n56099 & ~n56145 ;
  assign n56148 = n56086 & ~n56092 ;
  assign n56149 = ~n56147 & ~n56148 ;
  assign n56150 = ~n56146 & ~n56149 ;
  assign n56151 = ~n56099 & n56112 ;
  assign n56153 = ~n56151 & ~n56152 ;
  assign n56154 = n56086 & ~n56105 ;
  assign n56155 = ~n56153 & n56154 ;
  assign n56163 = ~n56150 & ~n56155 ;
  assign n56164 = n56159 & n56163 ;
  assign n56165 = ~n56162 & n56164 ;
  assign n56166 = ~n56142 & ~n56165 ;
  assign n56118 = n56099 & n56112 ;
  assign n56127 = ~n56118 & ~n56120 ;
  assign n56128 = n56092 & ~n56127 ;
  assign n56131 = n56099 & ~n56105 ;
  assign n56132 = n56112 & n56131 ;
  assign n56129 = n56105 & n56112 ;
  assign n56130 = ~n56099 & n56129 ;
  assign n56133 = ~n56092 & ~n56130 ;
  assign n56134 = ~n56132 & n56133 ;
  assign n56135 = ~n56128 & ~n56134 ;
  assign n56136 = ~n56086 & ~n56135 ;
  assign n56122 = ~n56105 & n56114 ;
  assign n56123 = ~n56092 & n56122 ;
  assign n56119 = n56105 & n56118 ;
  assign n56124 = n56086 & ~n56119 ;
  assign n56125 = ~n56121 & n56124 ;
  assign n56126 = ~n56123 & n56125 ;
  assign n56143 = ~n56126 & n56142 ;
  assign n56144 = ~n56136 & n56143 ;
  assign n56167 = ~n56099 & n56145 ;
  assign n56168 = ~n56092 & n56167 ;
  assign n56169 = ~n56157 & ~n56168 ;
  assign n56170 = n56086 & ~n56169 ;
  assign n56106 = ~n56099 & ~n56105 ;
  assign n56113 = n56106 & ~n56112 ;
  assign n56115 = n56105 & n56114 ;
  assign n56116 = ~n56113 & ~n56115 ;
  assign n56117 = n56093 & ~n56116 ;
  assign n56171 = ~n56105 & n56151 ;
  assign n56172 = n56148 & n56171 ;
  assign n56173 = ~n56117 & ~n56172 ;
  assign n56174 = ~n56170 & n56173 ;
  assign n56175 = ~n56144 & n56174 ;
  assign n56176 = ~n56166 & n56175 ;
  assign n56177 = ~\u0_L10_reg[11]/NET0131  & n56176 ;
  assign n56178 = \u0_L10_reg[11]/NET0131  & ~n56176 ;
  assign n56179 = ~n56177 & ~n56178 ;
  assign n56193 = ~n55923 & ~n55924 ;
  assign n56194 = ~n55930 & ~n56193 ;
  assign n56195 = ~n55909 & n55924 ;
  assign n56196 = ~n56194 & ~n56195 ;
  assign n56197 = ~n55903 & ~n56196 ;
  assign n56198 = ~n55935 & ~n55944 ;
  assign n56199 = n55968 & n56198 ;
  assign n56192 = n55954 & n55970 ;
  assign n56200 = n55938 & n55944 ;
  assign n56201 = ~n56192 & ~n56200 ;
  assign n56202 = ~n56199 & n56201 ;
  assign n56203 = ~n56197 & n56202 ;
  assign n56204 = ~n55897 & ~n56203 ;
  assign n56182 = ~n55916 & ~n55967 ;
  assign n56183 = n55923 & n55967 ;
  assign n56184 = ~n56182 & ~n56183 ;
  assign n56185 = n55903 & ~n56184 ;
  assign n56180 = ~n55909 & n55916 ;
  assign n56186 = ~n55903 & ~n56180 ;
  assign n56187 = ~n56182 & n56186 ;
  assign n56181 = n55944 & n56180 ;
  assign n56188 = ~n55971 & ~n56181 ;
  assign n56189 = ~n56187 & n56188 ;
  assign n56190 = ~n56185 & n56189 ;
  assign n56191 = n55897 & ~n56190 ;
  assign n56205 = n55922 & n55934 ;
  assign n56206 = ~n55959 & ~n56205 ;
  assign n56207 = n55903 & n55930 ;
  assign n56208 = ~n56206 & n56207 ;
  assign n56209 = ~n56191 & ~n56208 ;
  assign n56210 = ~n56204 & n56209 ;
  assign n56211 = ~\u0_L10_reg[17]/NET0131  & ~n56210 ;
  assign n56212 = \u0_L10_reg[17]/NET0131  & n56210 ;
  assign n56213 = ~n56211 & ~n56212 ;
  assign n56214 = decrypt_pad & ~\u0_uk_K_r10_reg[24]/NET0131  ;
  assign n56215 = ~decrypt_pad & ~\u0_uk_K_r10_reg[33]/NET0131  ;
  assign n56216 = ~n56214 & ~n56215 ;
  assign n56217 = \u0_R10_reg[15]/NET0131  & ~n56216 ;
  assign n56218 = ~\u0_R10_reg[15]/NET0131  & n56216 ;
  assign n56219 = ~n56217 & ~n56218 ;
  assign n56220 = decrypt_pad & ~\u0_uk_K_r10_reg[47]/NET0131  ;
  assign n56221 = ~decrypt_pad & ~\u0_uk_K_r10_reg[24]/NET0131  ;
  assign n56222 = ~n56220 & ~n56221 ;
  assign n56223 = \u0_R10_reg[13]/NET0131  & ~n56222 ;
  assign n56224 = ~\u0_R10_reg[13]/NET0131  & n56222 ;
  assign n56225 = ~n56223 & ~n56224 ;
  assign n56262 = n56219 & n56225 ;
  assign n56227 = decrypt_pad & ~\u0_uk_K_r10_reg[53]/NET0131  ;
  assign n56228 = ~decrypt_pad & ~\u0_uk_K_r10_reg[5]/NET0131  ;
  assign n56229 = ~n56227 & ~n56228 ;
  assign n56230 = \u0_R10_reg[12]/NET0131  & ~n56229 ;
  assign n56231 = ~\u0_R10_reg[12]/NET0131  & n56229 ;
  assign n56232 = ~n56230 & ~n56231 ;
  assign n56233 = decrypt_pad & ~\u0_uk_K_r10_reg[12]/NET0131  ;
  assign n56234 = ~decrypt_pad & ~\u0_uk_K_r10_reg[46]/NET0131  ;
  assign n56235 = ~n56233 & ~n56234 ;
  assign n56236 = \u0_R10_reg[17]/NET0131  & ~n56235 ;
  assign n56237 = ~\u0_R10_reg[17]/NET0131  & n56235 ;
  assign n56238 = ~n56236 & ~n56237 ;
  assign n56239 = n56232 & ~n56238 ;
  assign n56240 = decrypt_pad & ~\u0_uk_K_r10_reg[48]/NET0131  ;
  assign n56241 = ~decrypt_pad & ~\u0_uk_K_r10_reg[25]/NET0131  ;
  assign n56242 = ~n56240 & ~n56241 ;
  assign n56243 = \u0_R10_reg[14]/NET0131  & ~n56242 ;
  assign n56244 = ~\u0_R10_reg[14]/NET0131  & n56242 ;
  assign n56245 = ~n56243 & ~n56244 ;
  assign n56261 = ~n56232 & ~n56245 ;
  assign n56263 = ~n56239 & ~n56261 ;
  assign n56264 = n56262 & n56263 ;
  assign n56269 = decrypt_pad & ~\u0_uk_K_r10_reg[32]/NET0131  ;
  assign n56270 = ~decrypt_pad & ~\u0_uk_K_r10_reg[41]/P0001  ;
  assign n56271 = ~n56269 & ~n56270 ;
  assign n56272 = \u0_R10_reg[16]/NET0131  & ~n56271 ;
  assign n56273 = ~\u0_R10_reg[16]/NET0131  & n56271 ;
  assign n56274 = ~n56272 & ~n56273 ;
  assign n56275 = ~n56264 & ~n56274 ;
  assign n56254 = ~n56225 & ~n56238 ;
  assign n56255 = ~n56232 & n56254 ;
  assign n56265 = n56219 & n56255 ;
  assign n56266 = ~n56225 & n56232 ;
  assign n56267 = ~n56245 & n56266 ;
  assign n56268 = n56238 & n56267 ;
  assign n56276 = ~n56265 & ~n56268 ;
  assign n56277 = n56275 & n56276 ;
  assign n56251 = n56225 & ~n56232 ;
  assign n56252 = ~n56238 & n56251 ;
  assign n56253 = n56245 & n56252 ;
  assign n56256 = ~n56245 & n56255 ;
  assign n56257 = ~n56253 & ~n56256 ;
  assign n56246 = n56239 & n56245 ;
  assign n56258 = ~n56225 & n56238 ;
  assign n56259 = ~n56246 & ~n56258 ;
  assign n56260 = ~n56219 & ~n56259 ;
  assign n56278 = n56257 & ~n56260 ;
  assign n56279 = n56277 & n56278 ;
  assign n56291 = ~n56251 & ~n56266 ;
  assign n56292 = ~n56219 & ~n56245 ;
  assign n56293 = ~n56291 & n56292 ;
  assign n56284 = n56239 & n56262 ;
  assign n56226 = n56219 & ~n56225 ;
  assign n56282 = ~n56232 & n56238 ;
  assign n56283 = n56226 & n56282 ;
  assign n56294 = n56274 & ~n56283 ;
  assign n56295 = ~n56284 & n56294 ;
  assign n56296 = ~n56293 & n56295 ;
  assign n56280 = ~n56219 & n56255 ;
  assign n56281 = n56245 & n56280 ;
  assign n56285 = n56225 & ~n56245 ;
  assign n56286 = n56282 & n56285 ;
  assign n56287 = n56232 & n56238 ;
  assign n56288 = n56225 & n56287 ;
  assign n56289 = n56245 & n56288 ;
  assign n56290 = ~n56286 & ~n56289 ;
  assign n56297 = ~n56281 & n56290 ;
  assign n56298 = n56296 & n56297 ;
  assign n56299 = ~n56279 & ~n56298 ;
  assign n56247 = ~n56238 & ~n56245 ;
  assign n56248 = ~n56232 & n56247 ;
  assign n56249 = ~n56246 & ~n56248 ;
  assign n56250 = n56226 & ~n56249 ;
  assign n56300 = ~n56219 & n56286 ;
  assign n56301 = n56239 & n56285 ;
  assign n56302 = n56219 & n56301 ;
  assign n56303 = ~n56300 & ~n56302 ;
  assign n56304 = ~n56250 & n56303 ;
  assign n56305 = ~n56299 & n56304 ;
  assign n56306 = ~\u0_L10_reg[20]/NET0131  & ~n56305 ;
  assign n56307 = \u0_L10_reg[20]/NET0131  & n56305 ;
  assign n56308 = ~n56306 & ~n56307 ;
  assign n56331 = n56092 & ~n56151 ;
  assign n56332 = ~n56114 & n56331 ;
  assign n56333 = ~n56113 & ~n56332 ;
  assign n56334 = ~n56086 & ~n56333 ;
  assign n56316 = n56145 & n56152 ;
  assign n56324 = n56092 & ~n56112 ;
  assign n56328 = n56120 & ~n56324 ;
  assign n56329 = ~n56316 & ~n56328 ;
  assign n56330 = n56086 & ~n56329 ;
  assign n56325 = ~n56092 & n56112 ;
  assign n56326 = ~n56324 & ~n56325 ;
  assign n56327 = n56106 & ~n56326 ;
  assign n56335 = n56159 & ~n56327 ;
  assign n56336 = ~n56330 & n56335 ;
  assign n56337 = ~n56334 & n56336 ;
  assign n56338 = n56142 & ~n56337 ;
  assign n56309 = ~n56119 & ~n56122 ;
  assign n56310 = ~n56092 & ~n56105 ;
  assign n56311 = ~n56121 & ~n56310 ;
  assign n56312 = ~n56112 & ~n56311 ;
  assign n56313 = n56309 & ~n56312 ;
  assign n56314 = n56086 & ~n56313 ;
  assign n56315 = ~n56092 & ~n56127 ;
  assign n56317 = ~n56315 & ~n56316 ;
  assign n56318 = ~n56086 & ~n56317 ;
  assign n56319 = n56092 & n56171 ;
  assign n56320 = ~n56318 & ~n56319 ;
  assign n56321 = ~n56314 & n56320 ;
  assign n56322 = ~n56142 & ~n56321 ;
  assign n56323 = n56129 & n56148 ;
  assign n56339 = ~n56123 & ~n56323 ;
  assign n56340 = ~n56322 & n56339 ;
  assign n56341 = ~n56338 & n56340 ;
  assign n56342 = \u0_L10_reg[29]/NET0131  & ~n56341 ;
  assign n56343 = ~\u0_L10_reg[29]/NET0131  & n56341 ;
  assign n56344 = ~n56342 & ~n56343 ;
  assign n56345 = decrypt_pad & ~\u0_uk_K_r10_reg[7]/NET0131  ;
  assign n56346 = ~decrypt_pad & ~\u0_uk_K_r10_reg[43]/NET0131  ;
  assign n56347 = ~n56345 & ~n56346 ;
  assign n56348 = \u0_R10_reg[30]/NET0131  & ~n56347 ;
  assign n56349 = ~\u0_R10_reg[30]/NET0131  & n56347 ;
  assign n56350 = ~n56348 & ~n56349 ;
  assign n56351 = decrypt_pad & ~\u0_uk_K_r10_reg[37]/NET0131  ;
  assign n56352 = ~decrypt_pad & ~\u0_uk_K_r10_reg[42]/NET0131  ;
  assign n56353 = ~n56351 & ~n56352 ;
  assign n56354 = \u0_R10_reg[29]/NET0131  & ~n56353 ;
  assign n56355 = ~\u0_R10_reg[29]/NET0131  & n56353 ;
  assign n56356 = ~n56354 & ~n56355 ;
  assign n56357 = decrypt_pad & ~\u0_uk_K_r10_reg[22]/NET0131  ;
  assign n56358 = ~decrypt_pad & ~\u0_uk_K_r10_reg[31]/NET0131  ;
  assign n56359 = ~n56357 & ~n56358 ;
  assign n56360 = \u0_R10_reg[1]/NET0131  & ~n56359 ;
  assign n56361 = ~\u0_R10_reg[1]/NET0131  & n56359 ;
  assign n56362 = ~n56360 & ~n56361 ;
  assign n56363 = n56356 & n56362 ;
  assign n56364 = decrypt_pad & ~\u0_uk_K_r10_reg[38]/NET0131  ;
  assign n56365 = ~decrypt_pad & ~\u0_uk_K_r10_reg[15]/NET0131  ;
  assign n56366 = ~n56364 & ~n56365 ;
  assign n56367 = \u0_R10_reg[28]/NET0131  & ~n56366 ;
  assign n56368 = ~\u0_R10_reg[28]/NET0131  & n56366 ;
  assign n56369 = ~n56367 & ~n56368 ;
  assign n56370 = n56363 & ~n56369 ;
  assign n56371 = n56350 & n56370 ;
  assign n56372 = ~n56350 & n56369 ;
  assign n56373 = n56356 & ~n56362 ;
  assign n56374 = ~n56372 & ~n56373 ;
  assign n56375 = ~n56362 & n56372 ;
  assign n56376 = n56356 & n56375 ;
  assign n56377 = ~n56374 & ~n56376 ;
  assign n56378 = decrypt_pad & ~\u0_uk_K_r10_reg[50]/NET0131  ;
  assign n56379 = ~decrypt_pad & ~\u0_uk_K_r10_reg[0]/NET0131  ;
  assign n56380 = ~n56378 & ~n56379 ;
  assign n56381 = \u0_R10_reg[31]/P0001  & ~n56380 ;
  assign n56382 = ~\u0_R10_reg[31]/P0001  & n56380 ;
  assign n56383 = ~n56381 & ~n56382 ;
  assign n56384 = ~n56377 & n56383 ;
  assign n56385 = ~n56350 & ~n56356 ;
  assign n56386 = ~n56369 & n56385 ;
  assign n56387 = ~n56356 & n56369 ;
  assign n56388 = n56350 & n56387 ;
  assign n56389 = ~n56383 & ~n56388 ;
  assign n56390 = ~n56386 & n56389 ;
  assign n56391 = ~n56384 & ~n56390 ;
  assign n56392 = ~n56371 & ~n56391 ;
  assign n56393 = decrypt_pad & ~\u0_uk_K_r10_reg[1]/NET0131  ;
  assign n56394 = ~decrypt_pad & ~\u0_uk_K_r10_reg[37]/NET0131  ;
  assign n56395 = ~n56393 & ~n56394 ;
  assign n56396 = \u0_R10_reg[32]/NET0131  & ~n56395 ;
  assign n56397 = ~\u0_R10_reg[32]/NET0131  & n56395 ;
  assign n56398 = ~n56396 & ~n56397 ;
  assign n56399 = ~n56392 & n56398 ;
  assign n56415 = ~n56362 & n56388 ;
  assign n56407 = n56362 & ~n56369 ;
  assign n56408 = ~n56356 & n56407 ;
  assign n56416 = n56383 & ~n56408 ;
  assign n56417 = ~n56415 & n56416 ;
  assign n56402 = n56350 & ~n56362 ;
  assign n56403 = ~n56369 & n56402 ;
  assign n56418 = ~n56363 & ~n56383 ;
  assign n56419 = ~n56403 & n56418 ;
  assign n56420 = ~n56417 & ~n56419 ;
  assign n56421 = n56356 & n56369 ;
  assign n56422 = n56350 & n56421 ;
  assign n56423 = n56362 & n56422 ;
  assign n56400 = n56372 & ~n56383 ;
  assign n56424 = ~n56376 & ~n56400 ;
  assign n56425 = ~n56423 & n56424 ;
  assign n56426 = ~n56420 & n56425 ;
  assign n56427 = ~n56398 & ~n56426 ;
  assign n56401 = n56373 & n56400 ;
  assign n56404 = n56356 & n56403 ;
  assign n56405 = ~n56362 & n56386 ;
  assign n56406 = ~n56404 & ~n56405 ;
  assign n56409 = n56350 & n56408 ;
  assign n56410 = ~n56356 & n56362 ;
  assign n56411 = n56372 & n56410 ;
  assign n56412 = ~n56409 & ~n56411 ;
  assign n56413 = n56406 & n56412 ;
  assign n56414 = n56383 & ~n56413 ;
  assign n56428 = ~n56401 & ~n56414 ;
  assign n56429 = ~n56427 & n56428 ;
  assign n56430 = ~n56399 & n56429 ;
  assign n56431 = \u0_L10_reg[5]/NET0131  & ~n56430 ;
  assign n56432 = ~\u0_L10_reg[5]/NET0131  & n56430 ;
  assign n56433 = ~n56431 & ~n56432 ;
  assign n56436 = ~n56093 & ~n56168 ;
  assign n56437 = ~n56146 & ~n56436 ;
  assign n56435 = n56092 & n56129 ;
  assign n56434 = n56118 & n56148 ;
  assign n56438 = n56142 & ~n56434 ;
  assign n56439 = ~n56435 & n56438 ;
  assign n56440 = ~n56437 & n56439 ;
  assign n56441 = ~n56099 & n56325 ;
  assign n56442 = n56086 & ~n56115 ;
  assign n56443 = ~n56441 & n56442 ;
  assign n56444 = ~n56158 & n56443 ;
  assign n56445 = ~n56086 & ~n56167 ;
  assign n56446 = ~n56319 & n56445 ;
  assign n56447 = ~n56444 & ~n56446 ;
  assign n56448 = n56093 & n56118 ;
  assign n56449 = ~n56142 & ~n56448 ;
  assign n56450 = ~n56123 & n56449 ;
  assign n56451 = ~n56447 & n56450 ;
  assign n56452 = ~n56440 & ~n56451 ;
  assign n56453 = n56092 & n56309 ;
  assign n56454 = ~n56086 & ~n56147 ;
  assign n56455 = ~n56325 & n56454 ;
  assign n56456 = ~n56453 & n56455 ;
  assign n56457 = n56116 & ~n56130 ;
  assign n56458 = n56086 & n56092 ;
  assign n56459 = ~n56457 & n56458 ;
  assign n56460 = ~n56456 & ~n56459 ;
  assign n56461 = ~n56452 & n56460 ;
  assign n56462 = ~\u0_L10_reg[4]/NET0131  & ~n56461 ;
  assign n56463 = \u0_L10_reg[4]/NET0131  & n56461 ;
  assign n56464 = ~n56462 & ~n56463 ;
  assign n56465 = decrypt_pad & ~\u0_uk_K_r10_reg[6]/NET0131  ;
  assign n56466 = ~decrypt_pad & ~\u0_uk_K_r10_reg[40]/NET0131  ;
  assign n56467 = ~n56465 & ~n56466 ;
  assign n56468 = \u0_R10_reg[8]/NET0131  & ~n56467 ;
  assign n56469 = ~\u0_R10_reg[8]/NET0131  & n56467 ;
  assign n56470 = ~n56468 & ~n56469 ;
  assign n56471 = decrypt_pad & ~\u0_uk_K_r10_reg[46]/NET0131  ;
  assign n56472 = ~decrypt_pad & ~\u0_uk_K_r10_reg[55]/NET0131  ;
  assign n56473 = ~n56471 & ~n56472 ;
  assign n56474 = \u0_R10_reg[6]/NET0131  & ~n56473 ;
  assign n56475 = ~\u0_R10_reg[6]/NET0131  & n56473 ;
  assign n56476 = ~n56474 & ~n56475 ;
  assign n56477 = decrypt_pad & ~\u0_uk_K_r10_reg[11]/NET0131  ;
  assign n56478 = ~decrypt_pad & ~\u0_uk_K_r10_reg[20]/NET0131  ;
  assign n56479 = ~n56477 & ~n56478 ;
  assign n56480 = \u0_R10_reg[9]/NET0131  & ~n56479 ;
  assign n56481 = ~\u0_R10_reg[9]/NET0131  & n56479 ;
  assign n56482 = ~n56480 & ~n56481 ;
  assign n56483 = ~n56476 & n56482 ;
  assign n56484 = decrypt_pad & ~\u0_uk_K_r10_reg[55]/NET0131  ;
  assign n56485 = ~decrypt_pad & ~\u0_uk_K_r10_reg[32]/NET0131  ;
  assign n56486 = ~n56484 & ~n56485 ;
  assign n56487 = \u0_R10_reg[5]/NET0131  & ~n56486 ;
  assign n56488 = ~\u0_R10_reg[5]/NET0131  & n56486 ;
  assign n56489 = ~n56487 & ~n56488 ;
  assign n56490 = decrypt_pad & ~\u0_uk_K_r10_reg[40]/NET0131  ;
  assign n56491 = ~decrypt_pad & ~\u0_uk_K_r10_reg[17]/NET0131  ;
  assign n56492 = ~n56490 & ~n56491 ;
  assign n56493 = \u0_R10_reg[7]/NET0131  & ~n56492 ;
  assign n56494 = ~\u0_R10_reg[7]/NET0131  & n56492 ;
  assign n56495 = ~n56493 & ~n56494 ;
  assign n56496 = ~n56489 & ~n56495 ;
  assign n56497 = n56483 & n56496 ;
  assign n56498 = decrypt_pad & ~\u0_uk_K_r10_reg[19]/NET0131  ;
  assign n56499 = ~decrypt_pad & ~\u0_uk_K_r10_reg[53]/NET0131  ;
  assign n56500 = ~n56498 & ~n56499 ;
  assign n56501 = \u0_R10_reg[4]/NET0131  & ~n56500 ;
  assign n56502 = ~\u0_R10_reg[4]/NET0131  & n56500 ;
  assign n56503 = ~n56501 & ~n56502 ;
  assign n56504 = n56482 & ~n56503 ;
  assign n56505 = n56489 & n56504 ;
  assign n56506 = n56476 & n56505 ;
  assign n56507 = ~n56497 & ~n56506 ;
  assign n56509 = n56482 & ~n56489 ;
  assign n56514 = n56476 & n56503 ;
  assign n56515 = n56509 & n56514 ;
  assign n56516 = n56495 & n56515 ;
  assign n56521 = n56507 & ~n56516 ;
  assign n56508 = n56482 & n56503 ;
  assign n56510 = ~n56482 & n56489 ;
  assign n56511 = ~n56509 & ~n56510 ;
  assign n56512 = ~n56508 & ~n56511 ;
  assign n56513 = ~n56476 & n56512 ;
  assign n56517 = ~n56489 & n56508 ;
  assign n56518 = ~n56495 & ~n56517 ;
  assign n56519 = ~n56509 & ~n56514 ;
  assign n56520 = n56518 & ~n56519 ;
  assign n56522 = ~n56513 & ~n56520 ;
  assign n56523 = n56521 & n56522 ;
  assign n56524 = ~n56470 & ~n56523 ;
  assign n56526 = ~n56482 & ~n56503 ;
  assign n56543 = ~n56515 & ~n56526 ;
  assign n56544 = n56470 & ~n56543 ;
  assign n56525 = n56476 & ~n56489 ;
  assign n56545 = n56504 & ~n56525 ;
  assign n56546 = ~n56544 & ~n56545 ;
  assign n56542 = ~n56476 & n56489 ;
  assign n56547 = ~n56495 & ~n56542 ;
  assign n56548 = ~n56546 & n56547 ;
  assign n56527 = n56525 & n56526 ;
  assign n56528 = n56489 & n56503 ;
  assign n56529 = ~n56476 & n56528 ;
  assign n56530 = ~n56527 & ~n56529 ;
  assign n56531 = n56495 & ~n56530 ;
  assign n56532 = ~n56482 & ~n56489 ;
  assign n56533 = ~n56476 & n56532 ;
  assign n56534 = n56503 & n56533 ;
  assign n56535 = n56476 & ~n56503 ;
  assign n56536 = n56489 & n56495 ;
  assign n56537 = ~n56535 & n56536 ;
  assign n56538 = n56483 & n56528 ;
  assign n56539 = ~n56537 & ~n56538 ;
  assign n56540 = ~n56534 & n56539 ;
  assign n56541 = n56470 & ~n56540 ;
  assign n56549 = ~n56531 & ~n56541 ;
  assign n56550 = ~n56548 & n56549 ;
  assign n56551 = ~n56524 & n56550 ;
  assign n56552 = \u0_L10_reg[2]/NET0131  & n56551 ;
  assign n56553 = ~\u0_L10_reg[2]/NET0131  & ~n56551 ;
  assign n56554 = ~n56552 & ~n56553 ;
  assign n56555 = ~n56350 & n56373 ;
  assign n56556 = ~n56408 & ~n56421 ;
  assign n56557 = ~n56555 & n56556 ;
  assign n56558 = n56383 & ~n56557 ;
  assign n56559 = ~n56356 & n56375 ;
  assign n56560 = ~n56398 & ~n56559 ;
  assign n56561 = ~n56558 & n56560 ;
  assign n56562 = ~n56350 & n56356 ;
  assign n56563 = n56369 & n56562 ;
  assign n56570 = n56398 & ~n56563 ;
  assign n56564 = ~n56362 & ~n56369 ;
  assign n56565 = ~n56356 & n56383 ;
  assign n56566 = n56564 & n56565 ;
  assign n56567 = n56350 & ~n56383 ;
  assign n56568 = n56410 & n56567 ;
  assign n56571 = ~n56566 & ~n56568 ;
  assign n56572 = n56570 & n56571 ;
  assign n56569 = n56362 & n56388 ;
  assign n56573 = ~n56404 & ~n56569 ;
  assign n56574 = n56572 & n56573 ;
  assign n56575 = ~n56561 & ~n56574 ;
  assign n56576 = n56407 & n56562 ;
  assign n56577 = n56389 & ~n56576 ;
  assign n56578 = n56406 & n56577 ;
  assign n56579 = ~n56350 & n56408 ;
  assign n56580 = ~n56371 & n56383 ;
  assign n56581 = ~n56579 & n56580 ;
  assign n56582 = ~n56578 & ~n56581 ;
  assign n56583 = ~n56383 & ~n56398 ;
  assign n56584 = n56387 & n56583 ;
  assign n56585 = ~n56582 & ~n56584 ;
  assign n56586 = ~n56575 & n56585 ;
  assign n56587 = \u0_L10_reg[15]/P0001  & n56586 ;
  assign n56588 = ~\u0_L10_reg[15]/P0001  & ~n56586 ;
  assign n56589 = ~n56587 & ~n56588 ;
  assign n56596 = ~n56369 & ~n56383 ;
  assign n56597 = n56373 & n56596 ;
  assign n56603 = ~n56398 & ~n56597 ;
  assign n56604 = ~n56405 & n56603 ;
  assign n56601 = n56362 & n56372 ;
  assign n56602 = ~n56565 & n56601 ;
  assign n56605 = ~n56415 & ~n56602 ;
  assign n56606 = n56604 & n56605 ;
  assign n56592 = n56356 & ~n56369 ;
  assign n56593 = ~n56383 & n56407 ;
  assign n56594 = ~n56592 & ~n56593 ;
  assign n56595 = n56350 & ~n56594 ;
  assign n56598 = n56369 & n56373 ;
  assign n56599 = ~n56388 & ~n56598 ;
  assign n56600 = n56383 & ~n56599 ;
  assign n56607 = ~n56595 & ~n56600 ;
  assign n56608 = n56606 & n56607 ;
  assign n56609 = ~n56375 & ~n56383 ;
  assign n56610 = ~n56569 & n56609 ;
  assign n56612 = ~n56370 & n56383 ;
  assign n56611 = n56362 & n56385 ;
  assign n56613 = ~n56422 & ~n56611 ;
  assign n56614 = n56612 & n56613 ;
  assign n56615 = ~n56610 & ~n56614 ;
  assign n56616 = ~n56362 & ~n56592 ;
  assign n56617 = n56350 & ~n56387 ;
  assign n56618 = n56616 & n56617 ;
  assign n56619 = n56398 & ~n56579 ;
  assign n56620 = ~n56618 & n56619 ;
  assign n56621 = ~n56615 & n56620 ;
  assign n56622 = ~n56608 & ~n56621 ;
  assign n56590 = n56383 & n56386 ;
  assign n56591 = n56363 & n56400 ;
  assign n56623 = ~n56590 & ~n56591 ;
  assign n56624 = ~n56622 & n56623 ;
  assign n56625 = ~\u0_L10_reg[21]/NET0131  & ~n56624 ;
  assign n56626 = \u0_L10_reg[21]/NET0131  & n56624 ;
  assign n56627 = ~n56625 & ~n56626 ;
  assign n56683 = decrypt_pad & ~\u0_uk_K_r10_reg[45]/P0001  ;
  assign n56684 = ~decrypt_pad & ~\u0_uk_K_r10_reg[22]/NET0131  ;
  assign n56685 = ~n56683 & ~n56684 ;
  assign n56686 = \u0_R10_reg[20]/NET0131  & ~n56685 ;
  assign n56687 = ~\u0_R10_reg[20]/NET0131  & n56685 ;
  assign n56688 = ~n56686 & ~n56687 ;
  assign n56628 = decrypt_pad & ~\u0_uk_K_r10_reg[2]/NET0131  ;
  assign n56629 = ~decrypt_pad & ~\u0_uk_K_r10_reg[7]/NET0131  ;
  assign n56630 = ~n56628 & ~n56629 ;
  assign n56631 = \u0_R10_reg[19]/NET0131  & ~n56630 ;
  assign n56632 = ~\u0_R10_reg[19]/NET0131  & n56630 ;
  assign n56633 = ~n56631 & ~n56632 ;
  assign n56640 = decrypt_pad & ~\u0_uk_K_r10_reg[21]/NET0131  ;
  assign n56641 = ~decrypt_pad & ~\u0_uk_K_r10_reg[2]/NET0131  ;
  assign n56642 = ~n56640 & ~n56641 ;
  assign n56643 = \u0_R10_reg[17]/NET0131  & ~n56642 ;
  assign n56644 = ~\u0_R10_reg[17]/NET0131  & n56642 ;
  assign n56645 = ~n56643 & ~n56644 ;
  assign n56653 = decrypt_pad & ~\u0_uk_K_r10_reg[30]/NET0131  ;
  assign n56654 = ~decrypt_pad & ~\u0_uk_K_r10_reg[35]/NET0131  ;
  assign n56655 = ~n56653 & ~n56654 ;
  assign n56656 = \u0_R10_reg[16]/NET0131  & ~n56655 ;
  assign n56657 = ~\u0_R10_reg[16]/NET0131  & n56655 ;
  assign n56658 = ~n56656 & ~n56657 ;
  assign n56634 = decrypt_pad & ~\u0_uk_K_r10_reg[15]/NET0131  ;
  assign n56635 = ~decrypt_pad & ~\u0_uk_K_r10_reg[51]/NET0131  ;
  assign n56636 = ~n56634 & ~n56635 ;
  assign n56637 = \u0_R10_reg[18]/NET0131  & ~n56636 ;
  assign n56638 = ~\u0_R10_reg[18]/NET0131  & n56636 ;
  assign n56639 = ~n56637 & ~n56638 ;
  assign n56646 = decrypt_pad & ~\u0_uk_K_r10_reg[42]/NET0131  ;
  assign n56647 = ~decrypt_pad & ~\u0_uk_K_r10_reg[23]/NET0131  ;
  assign n56648 = ~n56646 & ~n56647 ;
  assign n56649 = \u0_R10_reg[21]/NET0131  & ~n56648 ;
  assign n56650 = ~\u0_R10_reg[21]/NET0131  & n56648 ;
  assign n56651 = ~n56649 & ~n56650 ;
  assign n56695 = ~n56639 & ~n56651 ;
  assign n56696 = n56658 & ~n56695 ;
  assign n56697 = ~n56645 & ~n56696 ;
  assign n56661 = ~n56651 & ~n56658 ;
  assign n56662 = n56639 & n56661 ;
  assign n56698 = n56651 & n56658 ;
  assign n56699 = n56645 & n56698 ;
  assign n56700 = ~n56662 & ~n56699 ;
  assign n56701 = ~n56697 & n56700 ;
  assign n56702 = n56633 & ~n56701 ;
  assign n56671 = n56645 & ~n56658 ;
  assign n56703 = ~n56639 & n56671 ;
  assign n56704 = ~n56645 & n56698 ;
  assign n56705 = ~n56703 & ~n56704 ;
  assign n56706 = ~n56633 & ~n56705 ;
  assign n56652 = n56645 & ~n56651 ;
  assign n56659 = n56652 & n56658 ;
  assign n56660 = n56639 & n56659 ;
  assign n56665 = ~n56639 & n56651 ;
  assign n56690 = n56645 & n56665 ;
  assign n56707 = ~n56660 & ~n56690 ;
  assign n56708 = ~n56706 & n56707 ;
  assign n56709 = ~n56702 & n56708 ;
  assign n56710 = n56688 & ~n56709 ;
  assign n56670 = n56633 & ~n56651 ;
  assign n56672 = n56639 & n56671 ;
  assign n56673 = ~n56651 & n56658 ;
  assign n56674 = ~n56645 & n56673 ;
  assign n56675 = ~n56672 & ~n56674 ;
  assign n56676 = ~n56670 & ~n56675 ;
  assign n56679 = n56633 & ~n56652 ;
  assign n56677 = ~n56645 & ~n56658 ;
  assign n56678 = ~n56633 & ~n56677 ;
  assign n56680 = ~n56639 & ~n56678 ;
  assign n56681 = ~n56679 & n56680 ;
  assign n56682 = ~n56676 & ~n56681 ;
  assign n56689 = ~n56682 & ~n56688 ;
  assign n56663 = ~n56645 & n56662 ;
  assign n56664 = ~n56660 & ~n56663 ;
  assign n56666 = ~n56658 & n56665 ;
  assign n56667 = ~n56645 & n56666 ;
  assign n56668 = n56664 & ~n56667 ;
  assign n56669 = n56633 & ~n56668 ;
  assign n56691 = ~n56633 & n56639 ;
  assign n56692 = ~n56645 & n56691 ;
  assign n56693 = ~n56690 & ~n56692 ;
  assign n56694 = n56658 & ~n56693 ;
  assign n56711 = ~n56669 & ~n56694 ;
  assign n56712 = ~n56689 & n56711 ;
  assign n56713 = ~n56710 & n56712 ;
  assign n56714 = ~\u0_L10_reg[25]/NET0131  & ~n56713 ;
  assign n56715 = \u0_L10_reg[25]/NET0131  & n56713 ;
  assign n56716 = ~n56714 & ~n56715 ;
  assign n56722 = ~n56160 & ~n56171 ;
  assign n56723 = n56086 & ~n56722 ;
  assign n56720 = n56105 & ~n56325 ;
  assign n56721 = ~n56331 & n56720 ;
  assign n56719 = ~n56086 & n56131 ;
  assign n56724 = n56142 & ~n56719 ;
  assign n56725 = ~n56327 & n56724 ;
  assign n56726 = ~n56721 & n56725 ;
  assign n56727 = ~n56723 & n56726 ;
  assign n56729 = ~n56086 & ~n56113 ;
  assign n56730 = ~n56130 & n56729 ;
  assign n56731 = n56086 & ~n56131 ;
  assign n56732 = ~n56152 & n56731 ;
  assign n56733 = ~n56167 & n56732 ;
  assign n56734 = ~n56730 & ~n56733 ;
  assign n56728 = n56099 & n56435 ;
  assign n56735 = ~n56142 & ~n56728 ;
  assign n56736 = ~n56734 & n56735 ;
  assign n56737 = ~n56727 & ~n56736 ;
  assign n56717 = ~n56115 & ~n56132 ;
  assign n56718 = n56093 & ~n56717 ;
  assign n56738 = ~n56172 & ~n56718 ;
  assign n56739 = ~n56737 & n56738 ;
  assign n56740 = ~\u0_L10_reg[19]/NET0131  & ~n56739 ;
  assign n56741 = \u0_L10_reg[19]/NET0131  & n56739 ;
  assign n56742 = ~n56740 & ~n56741 ;
  assign n56761 = ~n56247 & ~n56258 ;
  assign n56762 = n56232 & ~n56761 ;
  assign n56763 = ~n56219 & ~n56762 ;
  assign n56764 = ~n56225 & n56246 ;
  assign n56765 = n56219 & ~n56248 ;
  assign n56766 = ~n56764 & n56765 ;
  assign n56767 = ~n56763 & ~n56766 ;
  assign n56768 = n56290 & ~n56301 ;
  assign n56769 = ~n56767 & n56768 ;
  assign n56770 = ~n56274 & ~n56769 ;
  assign n56755 = n56245 & ~n56282 ;
  assign n56752 = ~n56219 & n56225 ;
  assign n56756 = ~n56239 & n56752 ;
  assign n56757 = ~n56755 & n56756 ;
  assign n56743 = ~n56232 & n56245 ;
  assign n56744 = ~n56225 & n56743 ;
  assign n56754 = n56225 & n56246 ;
  assign n56758 = ~n56744 & ~n56754 ;
  assign n56759 = ~n56757 & n56758 ;
  assign n56760 = n56274 & ~n56759 ;
  assign n56745 = n56238 & n56744 ;
  assign n56746 = ~n56289 & ~n56745 ;
  assign n56747 = ~n56253 & n56746 ;
  assign n56748 = n56219 & ~n56747 ;
  assign n56749 = ~n56258 & ~n56267 ;
  assign n56750 = n56219 & n56274 ;
  assign n56751 = ~n56749 & n56750 ;
  assign n56753 = n56246 & n56752 ;
  assign n56771 = ~n56281 & ~n56753 ;
  assign n56772 = ~n56751 & n56771 ;
  assign n56773 = ~n56748 & n56772 ;
  assign n56774 = ~n56760 & n56773 ;
  assign n56775 = ~n56770 & n56774 ;
  assign n56776 = ~\u0_L10_reg[1]/NET0131  & ~n56775 ;
  assign n56777 = \u0_L10_reg[1]/NET0131  & n56775 ;
  assign n56778 = ~n56776 & ~n56777 ;
  assign n56779 = n55934 & n55935 ;
  assign n56780 = ~n56181 & ~n56779 ;
  assign n56781 = ~n55903 & ~n56780 ;
  assign n56782 = n55903 & ~n55954 ;
  assign n56783 = ~n55931 & n56782 ;
  assign n56784 = ~n55972 & ~n56783 ;
  assign n56785 = ~n56781 & n56784 ;
  assign n56786 = ~n55910 & ~n56785 ;
  assign n56787 = n55932 & ~n56180 ;
  assign n56788 = n55903 & ~n56787 ;
  assign n56789 = ~n55916 & ~n56198 ;
  assign n56790 = ~n55903 & ~n55939 ;
  assign n56791 = ~n56789 & n56790 ;
  assign n56792 = ~n56788 & ~n56791 ;
  assign n56793 = n55897 & ~n56183 ;
  assign n56794 = ~n55979 & n56793 ;
  assign n56795 = ~n56792 & n56794 ;
  assign n56800 = ~n55897 & ~n55953 ;
  assign n56801 = ~n55971 & n56800 ;
  assign n56796 = ~n55937 & n55951 ;
  assign n56797 = ~n55967 & n56796 ;
  assign n56798 = n55903 & ~n55916 ;
  assign n56799 = ~n55973 & n56798 ;
  assign n56802 = ~n56797 & ~n56799 ;
  assign n56803 = n56801 & n56802 ;
  assign n56804 = ~n56795 & ~n56803 ;
  assign n56805 = ~n56786 & ~n56804 ;
  assign n56806 = \u0_L10_reg[23]/NET0131  & ~n56805 ;
  assign n56807 = ~\u0_L10_reg[23]/NET0131  & n56805 ;
  assign n56808 = ~n56806 & ~n56807 ;
  assign n56812 = ~n56476 & n56526 ;
  assign n56813 = ~n56505 & ~n56812 ;
  assign n56814 = n56495 & n56813 ;
  assign n56818 = ~n56489 & n56535 ;
  assign n56819 = ~n56495 & ~n56818 ;
  assign n56816 = ~n56482 & n56503 ;
  assign n56817 = ~n56476 & n56816 ;
  assign n56815 = ~n56489 & n56504 ;
  assign n56820 = ~n56528 & ~n56815 ;
  assign n56821 = ~n56817 & n56820 ;
  assign n56822 = n56819 & n56821 ;
  assign n56823 = ~n56814 & ~n56822 ;
  assign n56810 = ~n56508 & ~n56526 ;
  assign n56811 = n56525 & ~n56810 ;
  assign n56809 = n56510 & n56514 ;
  assign n56824 = ~n56470 & ~n56809 ;
  assign n56825 = ~n56811 & n56824 ;
  assign n56826 = ~n56823 & n56825 ;
  assign n56832 = n56503 & n56511 ;
  assign n56831 = n56510 & n56535 ;
  assign n56833 = n56495 & ~n56831 ;
  assign n56834 = ~n56832 & n56833 ;
  assign n56835 = ~n56809 & n56813 ;
  assign n56836 = n56819 & n56835 ;
  assign n56837 = ~n56834 & ~n56836 ;
  assign n56827 = n56495 & n56503 ;
  assign n56828 = ~n56517 & ~n56827 ;
  assign n56829 = ~n56476 & ~n56828 ;
  assign n56830 = n56504 & n56525 ;
  assign n56838 = n56470 & ~n56830 ;
  assign n56839 = ~n56829 & n56838 ;
  assign n56840 = ~n56837 & n56839 ;
  assign n56841 = ~n56826 & ~n56840 ;
  assign n56842 = ~\u0_L10_reg[28]/NET0131  & n56841 ;
  assign n56843 = \u0_L10_reg[28]/NET0131  & ~n56841 ;
  assign n56844 = ~n56842 & ~n56843 ;
  assign n56869 = n56651 & n56671 ;
  assign n56870 = ~n56666 & ~n56704 ;
  assign n56871 = ~n56869 & n56870 ;
  assign n56872 = ~n56633 & ~n56871 ;
  assign n56866 = ~n56639 & n56674 ;
  assign n56867 = ~n56699 & ~n56866 ;
  assign n56868 = n56633 & ~n56867 ;
  assign n56873 = n56664 & ~n56703 ;
  assign n56874 = ~n56868 & n56873 ;
  assign n56875 = ~n56872 & n56874 ;
  assign n56876 = ~n56688 & ~n56875 ;
  assign n56845 = n56639 & ~n56645 ;
  assign n56846 = n56673 & n56845 ;
  assign n56847 = ~n56633 & ~n56846 ;
  assign n56848 = n56639 & n56651 ;
  assign n56849 = n56677 & n56848 ;
  assign n56850 = n56633 & ~n56849 ;
  assign n56851 = n56639 & n56652 ;
  assign n56852 = n56665 & n56671 ;
  assign n56853 = ~n56851 & ~n56852 ;
  assign n56854 = n56850 & n56853 ;
  assign n56855 = ~n56847 & ~n56854 ;
  assign n56859 = ~n56849 & ~n56851 ;
  assign n56860 = ~n56658 & ~n56859 ;
  assign n56856 = n56677 & n56695 ;
  assign n56857 = ~n56704 & ~n56856 ;
  assign n56858 = n56633 & ~n56857 ;
  assign n56861 = ~n56633 & ~n56639 ;
  assign n56862 = n56658 & n56861 ;
  assign n56863 = ~n56858 & ~n56862 ;
  assign n56864 = ~n56860 & n56863 ;
  assign n56865 = n56688 & ~n56864 ;
  assign n56877 = ~n56855 & ~n56865 ;
  assign n56878 = ~n56876 & n56877 ;
  assign n56879 = ~\u0_L10_reg[8]/NET0131  & ~n56878 ;
  assign n56880 = \u0_L10_reg[8]/NET0131  & n56878 ;
  assign n56881 = ~n56879 & ~n56880 ;
  assign n56882 = n55992 & n56006 ;
  assign n56883 = ~n56070 & ~n56882 ;
  assign n56884 = n56033 & ~n56883 ;
  assign n56885 = ~n56051 & ~n56055 ;
  assign n56886 = n56036 & ~n56885 ;
  assign n56887 = ~n56017 & n56026 ;
  assign n56888 = ~n56039 & ~n56063 ;
  assign n56889 = n56887 & n56888 ;
  assign n56890 = ~n56886 & n56889 ;
  assign n56891 = ~n56884 & n56890 ;
  assign n56892 = ~n56041 & ~n56061 ;
  assign n56893 = ~n55992 & n56892 ;
  assign n56894 = ~n56056 & ~n56893 ;
  assign n56895 = n55998 & ~n56894 ;
  assign n56897 = ~n56033 & ~n56892 ;
  assign n56896 = n56006 & n56047 ;
  assign n56898 = ~n55998 & ~n56896 ;
  assign n56899 = ~n56897 & n56898 ;
  assign n56900 = ~n56895 & ~n56899 ;
  assign n56902 = n56018 & n56033 ;
  assign n56901 = ~n55998 & n56051 ;
  assign n56903 = ~n56046 & ~n56901 ;
  assign n56904 = ~n56902 & n56903 ;
  assign n56905 = ~n56006 & ~n56904 ;
  assign n56906 = ~n56026 & ~n56905 ;
  assign n56907 = ~n56900 & n56906 ;
  assign n56908 = ~n56891 & ~n56907 ;
  assign n56909 = \u0_L10_reg[12]/NET0131  & n56908 ;
  assign n56910 = ~\u0_L10_reg[12]/NET0131  & ~n56908 ;
  assign n56911 = ~n56909 & ~n56910 ;
  assign n56926 = ~n56252 & ~n56268 ;
  assign n56927 = n56219 & ~n56926 ;
  assign n56928 = n56239 & ~n56285 ;
  assign n56929 = ~n56286 & ~n56928 ;
  assign n56930 = ~n56219 & ~n56929 ;
  assign n56931 = n56746 & ~n56930 ;
  assign n56932 = ~n56927 & n56931 ;
  assign n56933 = n56274 & ~n56932 ;
  assign n56914 = ~n56245 & ~n56254 ;
  assign n56915 = ~n56226 & ~n56914 ;
  assign n56912 = n56219 & ~n56245 ;
  assign n56913 = n56258 & n56912 ;
  assign n56916 = n56232 & ~n56913 ;
  assign n56917 = ~n56915 & n56916 ;
  assign n56918 = n56282 & n56912 ;
  assign n56919 = ~n56280 & ~n56918 ;
  assign n56920 = n56257 & n56919 ;
  assign n56921 = ~n56917 & n56920 ;
  assign n56922 = ~n56274 & ~n56921 ;
  assign n56923 = ~n56256 & n56746 ;
  assign n56924 = ~n56219 & ~n56923 ;
  assign n56925 = n56262 & n56743 ;
  assign n56934 = ~n56302 & ~n56925 ;
  assign n56935 = ~n56924 & n56934 ;
  assign n56936 = ~n56922 & n56935 ;
  assign n56937 = ~n56933 & n56936 ;
  assign n56938 = ~\u0_L10_reg[10]/NET0131  & ~n56937 ;
  assign n56939 = \u0_L10_reg[10]/NET0131  & n56937 ;
  assign n56940 = ~n56938 & ~n56939 ;
  assign n56941 = ~n56538 & ~n56809 ;
  assign n56942 = ~n56503 & n56510 ;
  assign n56943 = ~n56830 & ~n56942 ;
  assign n56944 = ~n56534 & n56943 ;
  assign n56945 = ~n56470 & ~n56944 ;
  assign n56946 = n56941 & ~n56945 ;
  assign n56947 = ~n56495 & ~n56946 ;
  assign n56953 = ~n56489 & n56810 ;
  assign n56952 = n56489 & ~n56817 ;
  assign n56954 = n56495 & ~n56952 ;
  assign n56955 = ~n56953 & n56954 ;
  assign n56950 = ~n56476 & ~n56496 ;
  assign n56951 = n56504 & n56950 ;
  assign n56948 = n56476 & ~n56510 ;
  assign n56949 = n56827 & n56948 ;
  assign n56956 = ~n56470 & ~n56949 ;
  assign n56957 = ~n56951 & n56956 ;
  assign n56958 = ~n56955 & n56957 ;
  assign n56959 = ~n56482 & n56525 ;
  assign n56960 = n56518 & ~n56959 ;
  assign n56961 = n56476 & n56504 ;
  assign n56962 = n56495 & ~n56533 ;
  assign n56963 = ~n56961 & n56962 ;
  assign n56964 = ~n56960 & ~n56963 ;
  assign n56965 = ~n56476 & n56942 ;
  assign n56966 = n56470 & n56941 ;
  assign n56967 = ~n56965 & n56966 ;
  assign n56968 = n56507 & n56967 ;
  assign n56969 = ~n56964 & n56968 ;
  assign n56970 = ~n56958 & ~n56969 ;
  assign n56971 = ~n56947 & ~n56970 ;
  assign n56972 = ~\u0_L10_reg[13]/NET0131  & n56971 ;
  assign n56973 = \u0_L10_reg[13]/NET0131  & ~n56971 ;
  assign n56974 = ~n56972 & ~n56973 ;
  assign n56981 = n56651 & n56677 ;
  assign n56998 = ~n56659 & ~n56981 ;
  assign n56996 = ~n56658 & n56848 ;
  assign n56997 = ~n56639 & n56698 ;
  assign n56999 = ~n56996 & ~n56997 ;
  assign n57000 = n56998 & n56999 ;
  assign n57001 = n56633 & ~n57000 ;
  assign n56977 = ~n56645 & n56661 ;
  assign n56990 = ~n56869 & ~n56977 ;
  assign n56991 = n56861 & ~n56990 ;
  assign n56994 = ~n56645 & ~n56848 ;
  assign n56995 = n56696 & n56994 ;
  assign n56992 = n56691 & n56699 ;
  assign n56993 = ~n56639 & n56659 ;
  assign n57002 = ~n56992 & ~n56993 ;
  assign n57003 = ~n56995 & n57002 ;
  assign n57004 = ~n56991 & n57003 ;
  assign n57005 = ~n57001 & n57004 ;
  assign n57006 = n56688 & ~n57005 ;
  assign n56975 = ~n56665 & ~n56705 ;
  assign n56978 = n56633 & ~n56703 ;
  assign n56976 = n56639 & n56698 ;
  assign n56979 = ~n56976 & ~n56977 ;
  assign n56980 = n56978 & n56979 ;
  assign n56983 = ~n56633 & ~n56851 ;
  assign n56984 = ~n56981 & n56983 ;
  assign n56982 = n56658 & n56690 ;
  assign n56985 = ~n56866 & ~n56982 ;
  assign n56986 = n56984 & n56985 ;
  assign n56987 = ~n56980 & ~n56986 ;
  assign n56988 = ~n56975 & ~n56987 ;
  assign n56989 = ~n56688 & ~n56988 ;
  assign n57007 = ~n56633 & n56860 ;
  assign n57008 = ~n56663 & ~n56993 ;
  assign n57009 = n56633 & ~n57008 ;
  assign n57010 = ~n57007 & ~n57009 ;
  assign n57011 = ~n56989 & n57010 ;
  assign n57012 = ~n57006 & n57011 ;
  assign n57013 = ~\u0_L10_reg[14]/NET0131  & ~n57012 ;
  assign n57014 = \u0_L10_reg[14]/NET0131  & n57012 ;
  assign n57015 = ~n57013 & ~n57014 ;
  assign n57032 = n55909 & ~n55932 ;
  assign n57033 = ~n56194 & n57032 ;
  assign n57019 = ~n55923 & n56198 ;
  assign n57030 = n55903 & ~n55909 ;
  assign n57031 = n57019 & n57030 ;
  assign n57034 = ~n56181 & ~n57031 ;
  assign n57035 = ~n57033 & n57034 ;
  assign n57036 = n55897 & ~n57035 ;
  assign n57016 = n55930 & n56180 ;
  assign n57017 = n55903 & ~n56198 ;
  assign n57018 = ~n57016 & n57017 ;
  assign n57022 = n55922 & n57016 ;
  assign n57023 = ~n57018 & ~n57022 ;
  assign n57020 = ~n55903 & n57019 ;
  assign n57021 = n55909 & n56194 ;
  assign n57024 = ~n57020 & ~n57021 ;
  assign n57025 = n57023 & n57024 ;
  assign n57026 = ~n55897 & ~n57025 ;
  assign n57027 = ~n55916 & n55971 ;
  assign n57028 = ~n57022 & ~n57027 ;
  assign n57029 = ~n55903 & ~n57028 ;
  assign n57037 = ~n57026 & ~n57029 ;
  assign n57038 = ~n57036 & n57037 ;
  assign n57039 = ~\u0_L10_reg[9]/NET0131  & ~n57038 ;
  assign n57040 = \u0_L10_reg[9]/NET0131  & n57038 ;
  assign n57041 = ~n57039 & ~n57040 ;
  assign n57058 = ~n56370 & ~n56386 ;
  assign n57059 = ~n56598 & n57058 ;
  assign n57060 = ~n56383 & ~n57059 ;
  assign n57061 = ~n56371 & ~n56611 ;
  assign n57049 = n56362 & n56369 ;
  assign n57054 = ~n56564 & ~n57049 ;
  assign n57055 = n56356 & n56383 ;
  assign n57056 = ~n56402 & n57055 ;
  assign n57057 = ~n57054 & n57056 ;
  assign n57062 = ~n56415 & ~n57057 ;
  assign n57063 = n57061 & n57062 ;
  assign n57064 = ~n57060 & n57063 ;
  assign n57065 = n56398 & ~n57064 ;
  assign n57042 = ~n56562 & ~n56616 ;
  assign n57043 = n56383 & ~n56555 ;
  assign n57044 = ~n57042 & n57043 ;
  assign n57045 = ~n56409 & ~n57044 ;
  assign n57046 = ~n56398 & ~n57045 ;
  assign n57047 = ~n56404 & ~n56411 ;
  assign n57048 = ~n56383 & ~n57047 ;
  assign n57050 = n56567 & n57049 ;
  assign n57051 = ~n56597 & ~n57050 ;
  assign n57052 = ~n56398 & ~n57051 ;
  assign n57053 = n56402 & n56565 ;
  assign n57066 = ~n56401 & ~n57053 ;
  assign n57067 = ~n57052 & n57066 ;
  assign n57068 = ~n57048 & n57067 ;
  assign n57069 = ~n57046 & n57068 ;
  assign n57070 = ~n57065 & n57069 ;
  assign n57071 = ~\u0_L10_reg[27]/NET0131  & ~n57070 ;
  assign n57072 = \u0_L10_reg[27]/NET0131  & n57070 ;
  assign n57073 = ~n57071 & ~n57072 ;
  assign n57081 = ~n56015 & ~n56047 ;
  assign n57082 = ~n55998 & ~n57081 ;
  assign n57083 = ~n56016 & ~n56068 ;
  assign n57084 = ~n57082 & ~n57083 ;
  assign n57085 = ~n56896 & ~n57084 ;
  assign n57086 = ~n56033 & ~n57085 ;
  assign n57074 = n55998 & ~n56014 ;
  assign n57075 = ~n56006 & ~n56033 ;
  assign n57076 = n55992 & ~n57075 ;
  assign n57077 = n57074 & n57076 ;
  assign n57078 = ~n56006 & n56047 ;
  assign n57079 = ~n56062 & ~n57078 ;
  assign n57080 = n56033 & ~n57079 ;
  assign n57087 = ~n57077 & ~n57080 ;
  assign n57088 = ~n57086 & n57087 ;
  assign n57089 = n56026 & ~n57088 ;
  assign n57095 = ~n56062 & ~n57074 ;
  assign n57096 = n57076 & n57095 ;
  assign n57094 = n56897 & ~n56901 ;
  assign n57097 = n56040 & ~n57094 ;
  assign n57098 = ~n57096 & n57097 ;
  assign n57099 = ~n56026 & ~n57098 ;
  assign n57090 = n56033 & n56037 ;
  assign n57091 = n55992 & n56062 ;
  assign n57092 = ~n56038 & ~n57091 ;
  assign n57093 = ~n56033 & ~n57092 ;
  assign n57100 = ~n57090 & ~n57093 ;
  assign n57101 = ~n57099 & n57100 ;
  assign n57102 = ~n57089 & n57101 ;
  assign n57103 = \u0_L10_reg[32]/NET0131  & n57102 ;
  assign n57104 = ~\u0_L10_reg[32]/NET0131  & ~n57102 ;
  assign n57105 = ~n57103 & ~n57104 ;
  assign n57112 = decrypt_pad & ~\u0_uk_K_r10_reg[26]/NET0131  ;
  assign n57113 = ~decrypt_pad & ~\u0_uk_K_r10_reg[3]/NET0131  ;
  assign n57114 = ~n57112 & ~n57113 ;
  assign n57115 = \u0_R10_reg[11]/NET0131  & ~n57114 ;
  assign n57116 = ~\u0_R10_reg[11]/NET0131  & n57114 ;
  assign n57117 = ~n57115 & ~n57116 ;
  assign n57106 = decrypt_pad & ~\u0_uk_K_r10_reg[41]/P0001  ;
  assign n57107 = ~decrypt_pad & ~\u0_uk_K_r10_reg[18]/NET0131  ;
  assign n57108 = ~n57106 & ~n57107 ;
  assign n57109 = \u0_R10_reg[12]/NET0131  & ~n57108 ;
  assign n57110 = ~\u0_R10_reg[12]/NET0131  & n57108 ;
  assign n57111 = ~n57109 & ~n57110 ;
  assign n57118 = decrypt_pad & ~\u0_uk_K_r10_reg[54]/NET0131  ;
  assign n57119 = ~decrypt_pad & ~\u0_uk_K_r10_reg[6]/NET0131  ;
  assign n57120 = ~n57118 & ~n57119 ;
  assign n57121 = \u0_R10_reg[13]/NET0131  & ~n57120 ;
  assign n57122 = ~\u0_R10_reg[13]/NET0131  & n57120 ;
  assign n57123 = ~n57121 & ~n57122 ;
  assign n57131 = decrypt_pad & ~\u0_uk_K_r10_reg[17]/NET0131  ;
  assign n57132 = ~decrypt_pad & ~\u0_uk_K_r10_reg[26]/NET0131  ;
  assign n57133 = ~n57131 & ~n57132 ;
  assign n57134 = \u0_R10_reg[9]/NET0131  & ~n57133 ;
  assign n57135 = ~\u0_R10_reg[9]/NET0131  & n57133 ;
  assign n57136 = ~n57134 & ~n57135 ;
  assign n57176 = n57123 & ~n57136 ;
  assign n57124 = decrypt_pad & ~\u0_uk_K_r10_reg[20]/NET0131  ;
  assign n57125 = ~decrypt_pad & ~\u0_uk_K_r10_reg[54]/NET0131  ;
  assign n57126 = ~n57124 & ~n57125 ;
  assign n57127 = \u0_R10_reg[8]/NET0131  & ~n57126 ;
  assign n57128 = ~\u0_R10_reg[8]/NET0131  & n57126 ;
  assign n57129 = ~n57127 & ~n57128 ;
  assign n57156 = ~n57123 & n57136 ;
  assign n57157 = n57129 & n57156 ;
  assign n57130 = n57123 & ~n57129 ;
  assign n57138 = decrypt_pad & ~\u0_uk_K_r10_reg[25]/NET0131  ;
  assign n57139 = ~decrypt_pad & ~\u0_uk_K_r10_reg[34]/NET0131  ;
  assign n57140 = ~n57138 & ~n57139 ;
  assign n57141 = \u0_R10_reg[10]/NET0131  & ~n57140 ;
  assign n57142 = ~\u0_R10_reg[10]/NET0131  & n57140 ;
  assign n57143 = ~n57141 & ~n57142 ;
  assign n57178 = n57130 & n57143 ;
  assign n57179 = ~n57157 & ~n57178 ;
  assign n57180 = ~n57176 & n57179 ;
  assign n57181 = n57111 & ~n57180 ;
  assign n57177 = n57143 & n57176 ;
  assign n57148 = ~n57123 & ~n57129 ;
  assign n57182 = ~n57143 & n57148 ;
  assign n57183 = ~n57136 & n57182 ;
  assign n57184 = ~n57177 & ~n57183 ;
  assign n57185 = ~n57181 & n57184 ;
  assign n57186 = n57117 & ~n57185 ;
  assign n57149 = n57123 & n57129 ;
  assign n57150 = ~n57148 & ~n57149 ;
  assign n57147 = ~n57136 & ~n57143 ;
  assign n57153 = n57117 & ~n57129 ;
  assign n57159 = n57147 & ~n57153 ;
  assign n57160 = n57150 & n57159 ;
  assign n57154 = n57136 & ~n57143 ;
  assign n57155 = n57153 & n57154 ;
  assign n57158 = n57143 & n57157 ;
  assign n57161 = ~n57155 & ~n57158 ;
  assign n57162 = ~n57160 & n57161 ;
  assign n57137 = n57130 & n57136 ;
  assign n57144 = n57137 & n57143 ;
  assign n57145 = ~n57117 & n57144 ;
  assign n57146 = n57136 & n57143 ;
  assign n57151 = ~n57147 & ~n57150 ;
  assign n57152 = ~n57146 & n57151 ;
  assign n57163 = ~n57145 & ~n57152 ;
  assign n57164 = n57162 & n57163 ;
  assign n57165 = ~n57111 & ~n57164 ;
  assign n57166 = n57111 & n57146 ;
  assign n57167 = n57148 & n57166 ;
  assign n57168 = n57123 & n57154 ;
  assign n57169 = n57129 & ~n57136 ;
  assign n57170 = ~n57123 & n57169 ;
  assign n57171 = n57136 & n57149 ;
  assign n57172 = ~n57170 & ~n57171 ;
  assign n57173 = ~n57168 & n57172 ;
  assign n57174 = n57111 & ~n57117 ;
  assign n57175 = ~n57173 & n57174 ;
  assign n57187 = ~n57167 & ~n57175 ;
  assign n57188 = ~n57165 & n57187 ;
  assign n57189 = ~n57186 & n57188 ;
  assign n57190 = ~\u0_L10_reg[6]/NET0131  & ~n57189 ;
  assign n57191 = \u0_L10_reg[6]/NET0131  & n57189 ;
  assign n57192 = ~n57190 & ~n57191 ;
  assign n57193 = n56850 & ~n56866 ;
  assign n57194 = n56639 & n56704 ;
  assign n57195 = ~n56633 & ~n56856 ;
  assign n57196 = ~n56993 & n57195 ;
  assign n57197 = ~n57194 & n57196 ;
  assign n57198 = ~n57193 & ~n57197 ;
  assign n57199 = ~n56633 & ~n56661 ;
  assign n57200 = ~n56848 & n57199 ;
  assign n57201 = ~n56704 & n57200 ;
  assign n57202 = n56633 & ~n56659 ;
  assign n57203 = ~n56666 & n57202 ;
  assign n57204 = ~n57201 & ~n57203 ;
  assign n57205 = ~n56673 & n56845 ;
  assign n57206 = ~n56688 & ~n57205 ;
  assign n57207 = ~n57204 & n57206 ;
  assign n57208 = n56645 & n56661 ;
  assign n57209 = ~n56997 & ~n57208 ;
  assign n57210 = n56633 & ~n57209 ;
  assign n57211 = ~n56633 & n56869 ;
  assign n57212 = n56688 & ~n56846 ;
  assign n57213 = ~n56982 & n57212 ;
  assign n57214 = ~n57211 & n57213 ;
  assign n57215 = ~n57210 & n57214 ;
  assign n57216 = ~n57207 & ~n57215 ;
  assign n57217 = ~n57198 & ~n57216 ;
  assign n57218 = ~\u0_L10_reg[3]/NET0131  & ~n57217 ;
  assign n57219 = \u0_L10_reg[3]/NET0131  & n57217 ;
  assign n57220 = ~n57218 & ~n57219 ;
  assign n57221 = n56006 & n57081 ;
  assign n57222 = n55992 & n57074 ;
  assign n57223 = ~n56038 & ~n56069 ;
  assign n57224 = ~n57222 & n57223 ;
  assign n57225 = ~n57221 & n57224 ;
  assign n57226 = ~n56033 & ~n57225 ;
  assign n57229 = ~n56016 & ~n57221 ;
  assign n57230 = n55998 & ~n57229 ;
  assign n57227 = ~n56041 & n57082 ;
  assign n57228 = n56033 & n57227 ;
  assign n57231 = n56026 & ~n57228 ;
  assign n57232 = ~n57230 & n57231 ;
  assign n57233 = ~n57226 & n57232 ;
  assign n57234 = n55998 & n57221 ;
  assign n57235 = ~n56016 & n56033 ;
  assign n57236 = ~n57082 & n57235 ;
  assign n57237 = ~n57234 & n57236 ;
  assign n57238 = ~n56026 & ~n57237 ;
  assign n57239 = ~n57233 & ~n57238 ;
  assign n57240 = n56033 & ~n56048 ;
  assign n57241 = ~n56048 & ~n57227 ;
  assign n57242 = ~n56026 & ~n57241 ;
  assign n57243 = ~n56033 & ~n57230 ;
  assign n57244 = ~n57242 & n57243 ;
  assign n57245 = ~n57240 & ~n57244 ;
  assign n57246 = ~n57239 & ~n57245 ;
  assign n57247 = ~\u0_L10_reg[7]/NET0131  & ~n57246 ;
  assign n57248 = \u0_L10_reg[7]/NET0131  & n57246 ;
  assign n57249 = ~n57247 & ~n57248 ;
  assign n57262 = ~n56525 & ~n56536 ;
  assign n57264 = n56508 & ~n57262 ;
  assign n57258 = ~n56503 & ~n56542 ;
  assign n57263 = n57258 & n57262 ;
  assign n57265 = ~n56533 & ~n56809 ;
  assign n57266 = ~n57263 & n57265 ;
  assign n57267 = ~n57264 & n57266 ;
  assign n57268 = ~n56470 & ~n57267 ;
  assign n57255 = n56495 & n56512 ;
  assign n57256 = ~n56527 & ~n57255 ;
  assign n57257 = n56470 & ~n57256 ;
  assign n57250 = ~n56483 & ~n56532 ;
  assign n57251 = n56470 & n56503 ;
  assign n57252 = ~n57250 & n57251 ;
  assign n57253 = ~n56505 & ~n57252 ;
  assign n57254 = ~n56495 & ~n57253 ;
  assign n57259 = ~n56483 & n56495 ;
  assign n57260 = ~n56816 & n57259 ;
  assign n57261 = ~n57258 & n57260 ;
  assign n57269 = ~n57254 & ~n57261 ;
  assign n57270 = ~n57257 & n57269 ;
  assign n57271 = ~n57268 & n57270 ;
  assign n57272 = \u0_L10_reg[18]/NET0131  & n57271 ;
  assign n57273 = ~\u0_L10_reg[18]/NET0131  & ~n57271 ;
  assign n57274 = ~n57272 & ~n57273 ;
  assign n57275 = n57130 & ~n57136 ;
  assign n57292 = n57153 & n57156 ;
  assign n57293 = ~n57275 & ~n57292 ;
  assign n57294 = n57172 & n57293 ;
  assign n57295 = ~n57143 & ~n57294 ;
  assign n57286 = n57143 & n57148 ;
  assign n57296 = n57129 & ~n57143 ;
  assign n57297 = ~n57123 & n57296 ;
  assign n57298 = ~n57286 & ~n57297 ;
  assign n57299 = ~n57117 & ~n57298 ;
  assign n57300 = ~n57144 & ~n57299 ;
  assign n57301 = ~n57295 & n57300 ;
  assign n57302 = n57111 & ~n57301 ;
  assign n57276 = ~n57171 & ~n57182 ;
  assign n57277 = ~n57275 & n57276 ;
  assign n57278 = ~n57117 & ~n57277 ;
  assign n57279 = ~n57136 & ~n57149 ;
  assign n57280 = n57117 & ~n57148 ;
  assign n57281 = ~n57171 & n57280 ;
  assign n57282 = ~n57279 & n57281 ;
  assign n57283 = ~n57183 & ~n57282 ;
  assign n57284 = ~n57278 & n57283 ;
  assign n57285 = ~n57111 & ~n57284 ;
  assign n57287 = ~n57136 & n57286 ;
  assign n57288 = ~n57158 & ~n57287 ;
  assign n57289 = n57117 & ~n57288 ;
  assign n57290 = ~n57117 & n57143 ;
  assign n57291 = n57169 & n57290 ;
  assign n57303 = ~n57289 & ~n57291 ;
  assign n57304 = ~n57285 & n57303 ;
  assign n57305 = ~n57302 & n57304 ;
  assign n57306 = ~\u0_L10_reg[16]/NET0131  & ~n57305 ;
  assign n57307 = \u0_L10_reg[16]/NET0131  & n57305 ;
  assign n57308 = ~n57306 & ~n57307 ;
  assign n57325 = ~n57117 & n57151 ;
  assign n57319 = n57129 & n57146 ;
  assign n57320 = ~n57178 & ~n57319 ;
  assign n57321 = n57117 & ~n57320 ;
  assign n57322 = n57117 & ~n57143 ;
  assign n57323 = ~n57130 & ~n57136 ;
  assign n57324 = n57322 & n57323 ;
  assign n57326 = ~n57160 & ~n57324 ;
  assign n57327 = ~n57321 & n57326 ;
  assign n57328 = ~n57325 & n57327 ;
  assign n57329 = n57111 & ~n57328 ;
  assign n57309 = n57130 & ~n57143 ;
  assign n57310 = ~n57286 & ~n57309 ;
  assign n57311 = n57136 & n57148 ;
  assign n57312 = n57143 & n57169 ;
  assign n57313 = ~n57311 & ~n57312 ;
  assign n57314 = n57310 & n57313 ;
  assign n57315 = n57117 & ~n57314 ;
  assign n57316 = n57143 & n57170 ;
  assign n57317 = ~n57315 & ~n57316 ;
  assign n57318 = ~n57111 & ~n57317 ;
  assign n57333 = n57147 & ~n57150 ;
  assign n57334 = n57179 & ~n57333 ;
  assign n57335 = ~n57111 & ~n57117 ;
  assign n57336 = ~n57334 & n57335 ;
  assign n57330 = n57171 & n57290 ;
  assign n57331 = ~n57137 & ~n57170 ;
  assign n57332 = n57322 & ~n57331 ;
  assign n57337 = ~n57330 & ~n57332 ;
  assign n57338 = ~n57336 & n57337 ;
  assign n57339 = ~n57318 & n57338 ;
  assign n57340 = ~n57329 & n57339 ;
  assign n57341 = ~\u0_L10_reg[24]/NET0131  & ~n57340 ;
  assign n57342 = \u0_L10_reg[24]/NET0131  & n57340 ;
  assign n57343 = ~n57341 & ~n57342 ;
  assign n57349 = n57143 & n57275 ;
  assign n57353 = ~n57111 & ~n57333 ;
  assign n57354 = ~n57349 & n57353 ;
  assign n57344 = n57129 & n57143 ;
  assign n57345 = ~n57156 & n57344 ;
  assign n57346 = ~n57123 & n57154 ;
  assign n57347 = ~n57345 & ~n57346 ;
  assign n57348 = n57117 & ~n57347 ;
  assign n57350 = ~n57156 & n57296 ;
  assign n57351 = ~n57137 & ~n57350 ;
  assign n57352 = ~n57117 & ~n57351 ;
  assign n57355 = ~n57348 & ~n57352 ;
  assign n57356 = n57354 & n57355 ;
  assign n57359 = ~n57143 & n57170 ;
  assign n57360 = n57310 & ~n57359 ;
  assign n57361 = n57117 & ~n57360 ;
  assign n57357 = ~n57311 & ~n57344 ;
  assign n57358 = ~n57117 & ~n57357 ;
  assign n57362 = n57111 & ~n57358 ;
  assign n57363 = ~n57361 & n57362 ;
  assign n57364 = ~n57356 & ~n57363 ;
  assign n57367 = n57117 & n57176 ;
  assign n57368 = n57344 & n57367 ;
  assign n57365 = ~n57149 & n57166 ;
  assign n57366 = n57156 & n57290 ;
  assign n57369 = ~n57365 & ~n57366 ;
  assign n57370 = ~n57368 & n57369 ;
  assign n57371 = ~n57364 & n57370 ;
  assign n57372 = \u0_L10_reg[30]/NET0131  & ~n57371 ;
  assign n57373 = ~\u0_L10_reg[30]/NET0131  & n57371 ;
  assign n57374 = ~n57372 & ~n57373 ;
  assign n57375 = decrypt_pad & ~\u0_uk_K_r9_reg[8]/NET0131  ;
  assign n57376 = ~decrypt_pad & ~\u0_uk_K_r9_reg[16]/NET0131  ;
  assign n57377 = ~n57375 & ~n57376 ;
  assign n57378 = \u0_R9_reg[27]/NET0131  & ~n57377 ;
  assign n57379 = ~\u0_R9_reg[27]/NET0131  & n57377 ;
  assign n57380 = ~n57378 & ~n57379 ;
  assign n57381 = decrypt_pad & ~\u0_uk_K_r9_reg[30]/NET0131  ;
  assign n57382 = ~decrypt_pad & ~\u0_uk_K_r9_reg[7]/NET0131  ;
  assign n57383 = ~n57381 & ~n57382 ;
  assign n57384 = \u0_R9_reg[26]/NET0131  & ~n57383 ;
  assign n57385 = ~\u0_R9_reg[26]/NET0131  & n57383 ;
  assign n57386 = ~n57384 & ~n57385 ;
  assign n57394 = decrypt_pad & ~\u0_uk_K_r9_reg[38]/NET0131  ;
  assign n57395 = ~decrypt_pad & ~\u0_uk_K_r9_reg[42]/NET0131  ;
  assign n57396 = ~n57394 & ~n57395 ;
  assign n57397 = \u0_R9_reg[24]/NET0131  & ~n57396 ;
  assign n57398 = ~\u0_R9_reg[24]/NET0131  & n57396 ;
  assign n57399 = ~n57397 & ~n57398 ;
  assign n57387 = decrypt_pad & ~\u0_uk_K_r9_reg[14]/NET0131  ;
  assign n57388 = ~decrypt_pad & ~\u0_uk_K_r9_reg[22]/NET0131  ;
  assign n57389 = ~n57387 & ~n57388 ;
  assign n57390 = \u0_R9_reg[25]/NET0131  & ~n57389 ;
  assign n57391 = ~\u0_R9_reg[25]/NET0131  & n57389 ;
  assign n57392 = ~n57390 & ~n57391 ;
  assign n57400 = decrypt_pad & ~\u0_uk_K_r9_reg[42]/NET0131  ;
  assign n57401 = ~decrypt_pad & ~\u0_uk_K_r9_reg[50]/NET0131  ;
  assign n57402 = ~n57400 & ~n57401 ;
  assign n57403 = \u0_R9_reg[29]/NET0131  & ~n57402 ;
  assign n57404 = ~\u0_R9_reg[29]/NET0131  & n57402 ;
  assign n57405 = ~n57403 & ~n57404 ;
  assign n57412 = ~n57392 & ~n57405 ;
  assign n57413 = ~n57399 & n57412 ;
  assign n57414 = n57386 & n57413 ;
  assign n57393 = n57386 & ~n57392 ;
  assign n57406 = n57399 & ~n57405 ;
  assign n57407 = ~n57393 & n57406 ;
  assign n57408 = ~n57386 & ~n57399 ;
  assign n57409 = n57386 & n57399 ;
  assign n57410 = ~n57408 & ~n57409 ;
  assign n57411 = n57405 & ~n57410 ;
  assign n57415 = ~n57407 & ~n57411 ;
  assign n57416 = ~n57414 & n57415 ;
  assign n57417 = ~n57380 & ~n57416 ;
  assign n57418 = n57380 & n57399 ;
  assign n57419 = ~n57386 & ~n57392 ;
  assign n57420 = n57418 & n57419 ;
  assign n57421 = n57392 & n57411 ;
  assign n57422 = ~n57420 & ~n57421 ;
  assign n57423 = ~n57417 & n57422 ;
  assign n57424 = decrypt_pad & ~\u0_uk_K_r9_reg[50]/NET0131  ;
  assign n57425 = ~decrypt_pad & ~\u0_uk_K_r9_reg[31]/P0001  ;
  assign n57426 = ~n57424 & ~n57425 ;
  assign n57427 = \u0_R9_reg[28]/NET0131  & ~n57426 ;
  assign n57428 = ~\u0_R9_reg[28]/NET0131  & n57426 ;
  assign n57429 = ~n57427 & ~n57428 ;
  assign n57430 = ~n57423 & ~n57429 ;
  assign n57432 = n57392 & n57405 ;
  assign n57448 = ~n57399 & n57432 ;
  assign n57450 = n57386 & ~n57448 ;
  assign n57446 = ~n57392 & n57405 ;
  assign n57447 = n57399 & n57446 ;
  assign n57449 = ~n57447 & ~n57448 ;
  assign n57451 = ~n57380 & ~n57449 ;
  assign n57452 = ~n57450 & n57451 ;
  assign n57440 = ~n57386 & n57432 ;
  assign n57441 = ~n57393 & ~n57440 ;
  assign n57442 = n57418 & ~n57441 ;
  assign n57443 = ~n57386 & n57413 ;
  assign n57444 = ~n57399 & n57405 ;
  assign n57445 = n57393 & n57444 ;
  assign n57453 = ~n57443 & ~n57445 ;
  assign n57454 = ~n57442 & n57453 ;
  assign n57455 = ~n57452 & n57454 ;
  assign n57456 = n57429 & ~n57455 ;
  assign n57431 = n57386 & ~n57399 ;
  assign n57433 = ~n57412 & ~n57432 ;
  assign n57434 = n57431 & n57433 ;
  assign n57435 = n57412 & ~n57431 ;
  assign n57436 = ~n57434 & ~n57435 ;
  assign n57437 = n57380 & ~n57436 ;
  assign n57438 = ~n57380 & n57392 ;
  assign n57439 = ~n57410 & n57438 ;
  assign n57457 = ~n57437 & ~n57439 ;
  assign n57458 = ~n57456 & n57457 ;
  assign n57459 = ~n57430 & n57458 ;
  assign n57460 = ~\u0_L9_reg[22]/NET0131  & ~n57459 ;
  assign n57461 = \u0_L9_reg[22]/NET0131  & n57459 ;
  assign n57462 = ~n57460 & ~n57461 ;
  assign n57490 = decrypt_pad & ~\u0_uk_K_r9_reg[19]/NET0131  ;
  assign n57491 = ~decrypt_pad & ~\u0_uk_K_r9_reg[25]/NET0131  ;
  assign n57492 = ~n57490 & ~n57491 ;
  assign n57493 = \u0_R9_reg[4]/NET0131  & ~n57492 ;
  assign n57494 = ~\u0_R9_reg[4]/NET0131  & n57492 ;
  assign n57495 = ~n57493 & ~n57494 ;
  assign n57463 = decrypt_pad & ~\u0_uk_K_r9_reg[41]/NET0131  ;
  assign n57464 = ~decrypt_pad & ~\u0_uk_K_r9_reg[47]/NET0131  ;
  assign n57465 = ~n57463 & ~n57464 ;
  assign n57466 = \u0_R9_reg[3]/NET0131  & ~n57465 ;
  assign n57467 = ~\u0_R9_reg[3]/NET0131  & n57465 ;
  assign n57468 = ~n57466 & ~n57467 ;
  assign n57482 = decrypt_pad & ~\u0_uk_K_r9_reg[17]/NET0131  ;
  assign n57483 = ~decrypt_pad & ~\u0_uk_K_r9_reg[55]/NET0131  ;
  assign n57484 = ~n57482 & ~n57483 ;
  assign n57485 = \u0_R9_reg[1]/NET0131  & ~n57484 ;
  assign n57486 = ~\u0_R9_reg[1]/NET0131  & n57484 ;
  assign n57487 = ~n57485 & ~n57486 ;
  assign n57497 = decrypt_pad & ~\u0_uk_K_r9_reg[47]/NET0131  ;
  assign n57498 = ~decrypt_pad & ~\u0_uk_K_r9_reg[53]/NET0131  ;
  assign n57499 = ~n57497 & ~n57498 ;
  assign n57500 = \u0_R9_reg[5]/NET0131  & ~n57499 ;
  assign n57501 = ~\u0_R9_reg[5]/NET0131  & n57499 ;
  assign n57502 = ~n57500 & ~n57501 ;
  assign n57510 = ~n57487 & n57502 ;
  assign n57469 = decrypt_pad & ~\u0_uk_K_r9_reg[32]/NET0131  ;
  assign n57470 = ~decrypt_pad & ~\u0_uk_K_r9_reg[13]/NET0131  ;
  assign n57471 = ~n57469 & ~n57470 ;
  assign n57472 = \u0_R9_reg[2]/NET0131  & ~n57471 ;
  assign n57473 = ~\u0_R9_reg[2]/NET0131  & n57471 ;
  assign n57474 = ~n57472 & ~n57473 ;
  assign n57476 = decrypt_pad & ~\u0_uk_K_r9_reg[53]/NET0131  ;
  assign n57477 = ~decrypt_pad & ~\u0_uk_K_r9_reg[34]/NET0131  ;
  assign n57478 = ~n57476 & ~n57477 ;
  assign n57479 = \u0_R9_reg[32]/NET0131  & ~n57478 ;
  assign n57480 = ~\u0_R9_reg[32]/NET0131  & n57478 ;
  assign n57481 = ~n57479 & ~n57480 ;
  assign n57528 = n57474 & ~n57481 ;
  assign n57529 = ~n57502 & n57528 ;
  assign n57530 = ~n57510 & ~n57529 ;
  assign n57531 = n57468 & ~n57530 ;
  assign n57515 = ~n57468 & n57487 ;
  assign n57524 = ~n57487 & ~n57502 ;
  assign n57525 = ~n57474 & n57524 ;
  assign n57526 = ~n57515 & ~n57525 ;
  assign n57527 = n57481 & ~n57526 ;
  assign n57475 = n57468 & ~n57474 ;
  assign n57533 = ~n57475 & n57487 ;
  assign n57532 = ~n57474 & ~n57502 ;
  assign n57534 = ~n57481 & ~n57532 ;
  assign n57535 = ~n57533 & n57534 ;
  assign n57536 = ~n57527 & ~n57535 ;
  assign n57537 = ~n57531 & n57536 ;
  assign n57538 = n57495 & ~n57537 ;
  assign n57488 = n57481 & ~n57487 ;
  assign n57508 = n57488 & ~n57502 ;
  assign n57509 = n57474 & n57508 ;
  assign n57511 = ~n57474 & ~n57481 ;
  assign n57512 = ~n57510 & n57511 ;
  assign n57513 = ~n57509 & ~n57512 ;
  assign n57514 = ~n57468 & ~n57513 ;
  assign n57496 = n57468 & n57474 ;
  assign n57503 = ~n57481 & ~n57502 ;
  assign n57504 = n57481 & n57502 ;
  assign n57505 = ~n57503 & ~n57504 ;
  assign n57506 = n57487 & n57505 ;
  assign n57507 = n57496 & n57506 ;
  assign n57516 = n57504 & ~n57515 ;
  assign n57517 = ~n57481 & n57487 ;
  assign n57518 = ~n57502 & n57517 ;
  assign n57519 = ~n57516 & ~n57518 ;
  assign n57520 = ~n57474 & ~n57519 ;
  assign n57521 = ~n57507 & ~n57520 ;
  assign n57522 = ~n57514 & n57521 ;
  assign n57523 = ~n57495 & ~n57522 ;
  assign n57539 = n57474 & n57504 ;
  assign n57540 = ~n57532 & ~n57539 ;
  assign n57541 = n57487 & ~n57540 ;
  assign n57542 = n57510 & n57528 ;
  assign n57543 = ~n57541 & ~n57542 ;
  assign n57544 = ~n57468 & ~n57543 ;
  assign n57489 = n57475 & n57488 ;
  assign n57545 = ~n57487 & n57496 ;
  assign n57546 = n57503 & n57545 ;
  assign n57547 = ~n57489 & ~n57546 ;
  assign n57548 = ~n57544 & n57547 ;
  assign n57549 = ~n57523 & n57548 ;
  assign n57550 = ~n57538 & n57549 ;
  assign n57551 = ~\u0_L9_reg[31]/NET0131  & ~n57550 ;
  assign n57552 = \u0_L9_reg[31]/NET0131  & n57550 ;
  assign n57553 = ~n57551 & ~n57552 ;
  assign n57608 = decrypt_pad & ~\u0_uk_K_r9_reg[43]/NET0131  ;
  assign n57609 = ~decrypt_pad & ~\u0_uk_K_r9_reg[51]/NET0131  ;
  assign n57610 = ~n57608 & ~n57609 ;
  assign n57611 = \u0_R9_reg[24]/NET0131  & ~n57610 ;
  assign n57612 = ~\u0_R9_reg[24]/NET0131  & n57610 ;
  assign n57613 = ~n57611 & ~n57612 ;
  assign n57567 = decrypt_pad & ~\u0_uk_K_r9_reg[45]/NET0131  ;
  assign n57568 = ~decrypt_pad & ~\u0_uk_K_r9_reg[49]/NET0131  ;
  assign n57569 = ~n57567 & ~n57568 ;
  assign n57570 = \u0_R9_reg[23]/NET0131  & ~n57569 ;
  assign n57571 = ~\u0_R9_reg[23]/NET0131  & n57569 ;
  assign n57572 = ~n57570 & ~n57571 ;
  assign n57560 = decrypt_pad & ~\u0_uk_K_r9_reg[37]/NET0131  ;
  assign n57561 = ~decrypt_pad & ~\u0_uk_K_r9_reg[14]/NET0131  ;
  assign n57562 = ~n57560 & ~n57561 ;
  assign n57563 = \u0_R9_reg[21]/NET0131  & ~n57562 ;
  assign n57564 = ~\u0_R9_reg[21]/NET0131  & n57562 ;
  assign n57565 = ~n57563 & ~n57564 ;
  assign n57554 = decrypt_pad & ~\u0_uk_K_r9_reg[28]/NET0131  ;
  assign n57555 = ~decrypt_pad & ~\u0_uk_K_r9_reg[36]/NET0131  ;
  assign n57556 = ~n57554 & ~n57555 ;
  assign n57557 = \u0_R9_reg[22]/NET0131  & ~n57556 ;
  assign n57558 = ~\u0_R9_reg[22]/NET0131  & n57556 ;
  assign n57559 = ~n57557 & ~n57558 ;
  assign n57583 = decrypt_pad & ~\u0_uk_K_r9_reg[22]/NET0131  ;
  assign n57584 = ~decrypt_pad & ~\u0_uk_K_r9_reg[30]/NET0131  ;
  assign n57585 = ~n57583 & ~n57584 ;
  assign n57586 = \u0_R9_reg[20]/NET0131  & ~n57585 ;
  assign n57587 = ~\u0_R9_reg[20]/NET0131  & n57585 ;
  assign n57588 = ~n57586 & ~n57587 ;
  assign n57596 = n57559 & ~n57588 ;
  assign n57597 = n57565 & n57596 ;
  assign n57574 = decrypt_pad & ~\u0_uk_K_r9_reg[7]/NET0131  ;
  assign n57575 = ~decrypt_pad & ~\u0_uk_K_r9_reg[15]/NET0131  ;
  assign n57576 = ~n57574 & ~n57575 ;
  assign n57577 = \u0_R9_reg[25]/NET0131  & ~n57576 ;
  assign n57578 = ~\u0_R9_reg[25]/NET0131  & n57576 ;
  assign n57579 = ~n57577 & ~n57578 ;
  assign n57634 = n57559 & ~n57579 ;
  assign n57635 = n57565 & ~n57579 ;
  assign n57636 = n57588 & ~n57635 ;
  assign n57637 = ~n57565 & n57579 ;
  assign n57638 = n57636 & ~n57637 ;
  assign n57639 = ~n57634 & n57638 ;
  assign n57640 = ~n57597 & ~n57639 ;
  assign n57641 = n57572 & ~n57640 ;
  assign n57591 = n57579 & n57588 ;
  assign n57615 = n57565 & ~n57588 ;
  assign n57630 = ~n57591 & ~n57615 ;
  assign n57631 = n57559 & ~n57630 ;
  assign n57602 = n57579 & ~n57588 ;
  assign n57628 = n57565 & n57602 ;
  assign n57629 = ~n57559 & ~n57628 ;
  assign n57632 = ~n57572 & ~n57629 ;
  assign n57633 = ~n57631 & n57632 ;
  assign n57624 = ~n57559 & ~n57572 ;
  assign n57642 = n57591 & n57624 ;
  assign n57643 = ~n57565 & n57642 ;
  assign n57644 = ~n57633 & ~n57643 ;
  assign n57645 = ~n57641 & n57644 ;
  assign n57646 = n57613 & ~n57645 ;
  assign n57598 = n57565 & n57588 ;
  assign n57599 = ~n57559 & n57598 ;
  assign n57600 = ~n57597 & ~n57599 ;
  assign n57601 = ~n57572 & ~n57600 ;
  assign n57580 = ~n57559 & ~n57579 ;
  assign n57581 = ~n57565 & n57572 ;
  assign n57582 = ~n57580 & ~n57581 ;
  assign n57566 = ~n57559 & ~n57565 ;
  assign n57573 = n57566 & n57572 ;
  assign n57589 = ~n57573 & n57588 ;
  assign n57590 = ~n57582 & n57589 ;
  assign n57592 = n57559 & n57591 ;
  assign n57593 = ~n57565 & n57592 ;
  assign n57594 = ~n57559 & n57572 ;
  assign n57595 = ~n57588 & n57594 ;
  assign n57603 = n57581 & n57602 ;
  assign n57604 = ~n57595 & ~n57603 ;
  assign n57605 = ~n57593 & n57604 ;
  assign n57606 = ~n57590 & n57605 ;
  assign n57607 = ~n57601 & n57606 ;
  assign n57614 = ~n57607 & ~n57613 ;
  assign n57620 = ~n57579 & n57598 ;
  assign n57621 = ~n57572 & n57620 ;
  assign n57622 = ~n57603 & ~n57621 ;
  assign n57623 = ~n57559 & ~n57622 ;
  assign n57616 = ~n57579 & n57615 ;
  assign n57617 = ~n57559 & n57616 ;
  assign n57618 = ~n57592 & ~n57617 ;
  assign n57619 = n57572 & ~n57618 ;
  assign n57625 = ~n57579 & ~n57588 ;
  assign n57626 = n57624 & n57625 ;
  assign n57627 = ~n57565 & n57626 ;
  assign n57647 = ~n57619 & ~n57627 ;
  assign n57648 = ~n57623 & n57647 ;
  assign n57649 = ~n57614 & n57648 ;
  assign n57650 = ~n57646 & n57649 ;
  assign n57651 = ~\u0_L9_reg[11]/NET0131  & n57650 ;
  assign n57652 = \u0_L9_reg[11]/NET0131  & ~n57650 ;
  assign n57653 = ~n57651 & ~n57652 ;
  assign n57654 = decrypt_pad & ~\u0_uk_K_r9_reg[10]/NET0131  ;
  assign n57655 = ~decrypt_pad & ~\u0_uk_K_r9_reg[48]/NET0131  ;
  assign n57656 = ~n57654 & ~n57655 ;
  assign n57657 = \u0_R9_reg[12]/NET0131  & ~n57656 ;
  assign n57658 = ~\u0_R9_reg[12]/NET0131  & n57656 ;
  assign n57659 = ~n57657 & ~n57658 ;
  assign n57660 = decrypt_pad & ~\u0_uk_K_r9_reg[4]/NET0131  ;
  assign n57661 = ~decrypt_pad & ~\u0_uk_K_r9_reg[10]/NET0131  ;
  assign n57662 = ~n57660 & ~n57661 ;
  assign n57663 = \u0_R9_reg[13]/NET0131  & ~n57662 ;
  assign n57664 = ~\u0_R9_reg[13]/NET0131  & n57662 ;
  assign n57665 = ~n57663 & ~n57664 ;
  assign n57666 = ~n57659 & n57665 ;
  assign n57691 = n57659 & ~n57665 ;
  assign n57692 = ~n57666 & ~n57691 ;
  assign n57667 = decrypt_pad & ~\u0_uk_K_r9_reg[26]/NET0131  ;
  assign n57668 = ~decrypt_pad & ~\u0_uk_K_r9_reg[32]/NET0131  ;
  assign n57669 = ~n57667 & ~n57668 ;
  assign n57670 = \u0_R9_reg[17]/NET0131  & ~n57669 ;
  assign n57671 = ~\u0_R9_reg[17]/NET0131  & n57669 ;
  assign n57672 = ~n57670 & ~n57671 ;
  assign n57693 = n57659 & ~n57672 ;
  assign n57694 = ~n57659 & n57672 ;
  assign n57695 = ~n57693 & ~n57694 ;
  assign n57696 = n57692 & n57695 ;
  assign n57697 = decrypt_pad & ~\u0_uk_K_r9_reg[13]/NET0131  ;
  assign n57698 = ~decrypt_pad & ~\u0_uk_K_r9_reg[19]/NET0131  ;
  assign n57699 = ~n57697 & ~n57698 ;
  assign n57700 = \u0_R9_reg[15]/NET0131  & ~n57699 ;
  assign n57701 = ~\u0_R9_reg[15]/NET0131  & n57699 ;
  assign n57702 = ~n57700 & ~n57701 ;
  assign n57703 = ~n57696 & n57702 ;
  assign n57674 = decrypt_pad & ~\u0_uk_K_r9_reg[5]/NET0131  ;
  assign n57675 = ~decrypt_pad & ~\u0_uk_K_r9_reg[11]/NET0131  ;
  assign n57676 = ~n57674 & ~n57675 ;
  assign n57677 = \u0_R9_reg[14]/NET0131  & ~n57676 ;
  assign n57678 = ~\u0_R9_reg[14]/NET0131  & n57676 ;
  assign n57679 = ~n57677 & ~n57678 ;
  assign n57704 = n57679 & n57693 ;
  assign n57705 = ~n57665 & n57672 ;
  assign n57706 = ~n57702 & ~n57705 ;
  assign n57707 = ~n57704 & n57706 ;
  assign n57708 = ~n57703 & ~n57707 ;
  assign n57673 = n57666 & ~n57672 ;
  assign n57680 = n57673 & n57679 ;
  assign n57681 = ~n57672 & ~n57679 ;
  assign n57682 = ~n57659 & n57681 ;
  assign n57683 = ~n57665 & n57682 ;
  assign n57684 = ~n57680 & ~n57683 ;
  assign n57712 = n57659 & ~n57679 ;
  assign n57713 = ~n57665 & n57712 ;
  assign n57714 = n57672 & n57713 ;
  assign n57685 = decrypt_pad & ~\u0_uk_K_r9_reg[46]/NET0131  ;
  assign n57686 = ~decrypt_pad & ~\u0_uk_K_r9_reg[27]/P0001  ;
  assign n57687 = ~n57685 & ~n57686 ;
  assign n57688 = \u0_R9_reg[16]/NET0131  & ~n57687 ;
  assign n57689 = ~\u0_R9_reg[16]/NET0131  & n57687 ;
  assign n57690 = ~n57688 & ~n57689 ;
  assign n57709 = n57665 & n57679 ;
  assign n57710 = n57702 & n57709 ;
  assign n57711 = ~n57659 & n57710 ;
  assign n57715 = ~n57690 & ~n57711 ;
  assign n57716 = ~n57714 & n57715 ;
  assign n57717 = n57684 & n57716 ;
  assign n57718 = ~n57708 & n57717 ;
  assign n57730 = ~n57679 & ~n57702 ;
  assign n57731 = ~n57692 & n57730 ;
  assign n57723 = n57694 & n57702 ;
  assign n57724 = ~n57665 & n57723 ;
  assign n57732 = n57659 & n57672 ;
  assign n57733 = n57709 & n57732 ;
  assign n57734 = n57690 & ~n57733 ;
  assign n57735 = ~n57724 & n57734 ;
  assign n57736 = ~n57731 & n57735 ;
  assign n57719 = ~n57665 & n57679 ;
  assign n57720 = ~n57659 & n57719 ;
  assign n57721 = ~n57672 & n57720 ;
  assign n57722 = ~n57702 & n57721 ;
  assign n57725 = n57693 & n57702 ;
  assign n57726 = n57665 & n57725 ;
  assign n57727 = n57672 & ~n57679 ;
  assign n57728 = n57666 & n57727 ;
  assign n57729 = ~n57726 & ~n57728 ;
  assign n57737 = ~n57722 & n57729 ;
  assign n57738 = n57736 & n57737 ;
  assign n57739 = ~n57718 & ~n57738 ;
  assign n57740 = ~n57702 & ~n57728 ;
  assign n57741 = n57693 & n57719 ;
  assign n57742 = n57702 & ~n57741 ;
  assign n57743 = ~n57683 & n57742 ;
  assign n57744 = ~n57740 & ~n57743 ;
  assign n57745 = n57665 & ~n57679 ;
  assign n57746 = n57725 & n57745 ;
  assign n57747 = ~n57744 & ~n57746 ;
  assign n57748 = ~n57739 & n57747 ;
  assign n57749 = ~\u0_L9_reg[20]/NET0131  & ~n57748 ;
  assign n57750 = \u0_L9_reg[20]/NET0131  & n57748 ;
  assign n57751 = ~n57749 & ~n57750 ;
  assign n57752 = decrypt_pad & ~\u0_uk_K_r9_reg[52]/NET0131  ;
  assign n57753 = ~decrypt_pad & ~\u0_uk_K_r9_reg[1]/NET0131  ;
  assign n57754 = ~n57752 & ~n57753 ;
  assign n57755 = \u0_R9_reg[28]/NET0131  & ~n57754 ;
  assign n57756 = ~\u0_R9_reg[28]/NET0131  & n57754 ;
  assign n57757 = ~n57755 & ~n57756 ;
  assign n57765 = decrypt_pad & ~\u0_uk_K_r9_reg[21]/NET0131  ;
  assign n57766 = ~decrypt_pad & ~\u0_uk_K_r9_reg[29]/NET0131  ;
  assign n57767 = ~n57765 & ~n57766 ;
  assign n57768 = \u0_R9_reg[30]/NET0131  & ~n57767 ;
  assign n57769 = ~\u0_R9_reg[30]/NET0131  & n57767 ;
  assign n57770 = ~n57768 & ~n57769 ;
  assign n57758 = decrypt_pad & ~\u0_uk_K_r9_reg[51]/NET0131  ;
  assign n57759 = ~decrypt_pad & ~\u0_uk_K_r9_reg[28]/NET0131  ;
  assign n57760 = ~n57758 & ~n57759 ;
  assign n57761 = \u0_R9_reg[29]/NET0131  & ~n57760 ;
  assign n57762 = ~\u0_R9_reg[29]/NET0131  & n57760 ;
  assign n57763 = ~n57761 & ~n57762 ;
  assign n57772 = decrypt_pad & ~\u0_uk_K_r9_reg[36]/NET0131  ;
  assign n57773 = ~decrypt_pad & ~\u0_uk_K_r9_reg[44]/NET0131  ;
  assign n57774 = ~n57772 & ~n57773 ;
  assign n57775 = \u0_R9_reg[1]/NET0131  & ~n57774 ;
  assign n57776 = ~\u0_R9_reg[1]/NET0131  & n57774 ;
  assign n57777 = ~n57775 & ~n57776 ;
  assign n57797 = n57763 & ~n57777 ;
  assign n57798 = ~n57770 & n57797 ;
  assign n57782 = decrypt_pad & ~\u0_uk_K_r9_reg[9]/NET0131  ;
  assign n57783 = ~decrypt_pad & ~\u0_uk_K_r9_reg[45]/NET0131  ;
  assign n57784 = ~n57782 & ~n57783 ;
  assign n57785 = \u0_R9_reg[31]/P0001  & ~n57784 ;
  assign n57786 = ~\u0_R9_reg[31]/P0001  & n57784 ;
  assign n57787 = ~n57785 & ~n57786 ;
  assign n57794 = ~n57770 & ~n57787 ;
  assign n57795 = n57770 & n57777 ;
  assign n57796 = n57763 & n57795 ;
  assign n57799 = ~n57794 & ~n57796 ;
  assign n57800 = ~n57798 & n57799 ;
  assign n57801 = n57757 & ~n57800 ;
  assign n57764 = n57757 & ~n57763 ;
  assign n57771 = n57764 & n57770 ;
  assign n57778 = n57771 & ~n57777 ;
  assign n57779 = ~n57757 & n57777 ;
  assign n57780 = ~n57763 & n57779 ;
  assign n57781 = ~n57778 & ~n57780 ;
  assign n57788 = ~n57781 & n57787 ;
  assign n57789 = ~n57757 & n57770 ;
  assign n57790 = ~n57777 & ~n57789 ;
  assign n57791 = ~n57763 & n57777 ;
  assign n57792 = ~n57787 & ~n57791 ;
  assign n57793 = ~n57790 & n57792 ;
  assign n57802 = ~n57788 & ~n57793 ;
  assign n57803 = ~n57801 & n57802 ;
  assign n57804 = decrypt_pad & ~\u0_uk_K_r9_reg[15]/NET0131  ;
  assign n57805 = ~decrypt_pad & ~\u0_uk_K_r9_reg[23]/P0001  ;
  assign n57806 = ~n57804 & ~n57805 ;
  assign n57807 = \u0_R9_reg[32]/NET0131  & ~n57806 ;
  assign n57808 = ~\u0_R9_reg[32]/NET0131  & n57806 ;
  assign n57809 = ~n57807 & ~n57808 ;
  assign n57810 = ~n57803 & ~n57809 ;
  assign n57830 = n57757 & n57798 ;
  assign n57817 = n57757 & ~n57770 ;
  assign n57818 = ~n57797 & ~n57817 ;
  assign n57831 = n57787 & ~n57818 ;
  assign n57832 = ~n57830 & n57831 ;
  assign n57833 = ~n57757 & n57796 ;
  assign n57834 = ~n57763 & ~n57770 ;
  assign n57835 = ~n57757 & n57834 ;
  assign n57836 = ~n57787 & n57835 ;
  assign n57837 = ~n57833 & ~n57836 ;
  assign n57838 = ~n57832 & n57837 ;
  assign n57839 = n57809 & ~n57838 ;
  assign n57815 = n57757 & ~n57777 ;
  assign n57816 = n57763 & ~n57770 ;
  assign n57819 = ~n57815 & ~n57816 ;
  assign n57820 = ~n57818 & n57819 ;
  assign n57811 = ~n57763 & ~n57777 ;
  assign n57812 = ~n57757 & n57811 ;
  assign n57813 = ~n57770 & n57812 ;
  assign n57814 = n57789 & n57791 ;
  assign n57821 = ~n57813 & ~n57814 ;
  assign n57822 = ~n57820 & n57821 ;
  assign n57823 = n57787 & ~n57822 ;
  assign n57824 = n57757 & n57763 ;
  assign n57825 = ~n57777 & n57824 ;
  assign n57826 = n57794 & n57825 ;
  assign n57827 = n57770 & ~n57787 ;
  assign n57828 = n57764 & n57809 ;
  assign n57829 = n57827 & n57828 ;
  assign n57840 = ~n57826 & ~n57829 ;
  assign n57841 = ~n57823 & n57840 ;
  assign n57842 = ~n57839 & n57841 ;
  assign n57843 = ~n57810 & n57842 ;
  assign n57844 = \u0_L9_reg[5]/NET0131  & ~n57843 ;
  assign n57845 = ~\u0_L9_reg[5]/NET0131  & n57843 ;
  assign n57846 = ~n57844 & ~n57845 ;
  assign n57847 = n57702 & ~n57714 ;
  assign n57848 = ~n57728 & n57847 ;
  assign n57850 = ~n57665 & ~n57672 ;
  assign n57851 = ~n57720 & ~n57850 ;
  assign n57852 = ~n57690 & ~n57851 ;
  assign n57853 = ~n57672 & n57713 ;
  assign n57849 = n57695 & n57745 ;
  assign n57854 = ~n57702 & ~n57849 ;
  assign n57855 = ~n57853 & n57854 ;
  assign n57856 = ~n57852 & n57855 ;
  assign n57857 = ~n57848 & ~n57856 ;
  assign n57867 = ~n57659 & n57850 ;
  assign n57868 = n57702 & n57867 ;
  assign n57866 = n57665 & n57704 ;
  assign n57858 = n57666 & n57681 ;
  assign n57869 = n57690 & ~n57858 ;
  assign n57870 = ~n57866 & n57869 ;
  assign n57871 = ~n57868 & n57870 ;
  assign n57859 = ~n57665 & n57727 ;
  assign n57860 = ~n57732 & ~n57859 ;
  assign n57861 = ~n57702 & ~n57712 ;
  assign n57862 = ~n57860 & n57861 ;
  assign n57863 = n57665 & n57694 ;
  assign n57864 = ~n57723 & ~n57863 ;
  assign n57865 = n57679 & ~n57864 ;
  assign n57872 = ~n57862 & ~n57865 ;
  assign n57873 = n57871 & n57872 ;
  assign n57874 = ~n57694 & n57710 ;
  assign n57875 = ~n57690 & ~n57713 ;
  assign n57876 = ~n57874 & n57875 ;
  assign n57877 = n57729 & n57876 ;
  assign n57878 = ~n57873 & ~n57877 ;
  assign n57879 = ~n57857 & ~n57878 ;
  assign n57880 = ~\u0_L9_reg[26]/NET0131  & ~n57879 ;
  assign n57881 = \u0_L9_reg[26]/NET0131  & n57879 ;
  assign n57882 = ~n57880 & ~n57881 ;
  assign n57915 = decrypt_pad & ~\u0_uk_K_r9_reg[54]/NET0131  ;
  assign n57916 = ~decrypt_pad & ~\u0_uk_K_r9_reg[3]/NET0131  ;
  assign n57917 = ~n57915 & ~n57916 ;
  assign n57918 = \u0_R9_reg[7]/NET0131  & ~n57917 ;
  assign n57919 = ~\u0_R9_reg[7]/NET0131  & n57917 ;
  assign n57920 = ~n57918 & ~n57919 ;
  assign n57883 = decrypt_pad & ~\u0_uk_K_r9_reg[12]/NET0131  ;
  assign n57884 = ~decrypt_pad & ~\u0_uk_K_r9_reg[18]/NET0131  ;
  assign n57885 = ~n57883 & ~n57884 ;
  assign n57886 = \u0_R9_reg[5]/NET0131  & ~n57885 ;
  assign n57887 = ~\u0_R9_reg[5]/NET0131  & n57885 ;
  assign n57888 = ~n57886 & ~n57887 ;
  assign n57889 = decrypt_pad & ~\u0_uk_K_r9_reg[25]/NET0131  ;
  assign n57890 = ~decrypt_pad & ~\u0_uk_K_r9_reg[6]/NET0131  ;
  assign n57891 = ~n57889 & ~n57890 ;
  assign n57892 = \u0_R9_reg[9]/NET0131  & ~n57891 ;
  assign n57893 = ~\u0_R9_reg[9]/NET0131  & n57891 ;
  assign n57894 = ~n57892 & ~n57893 ;
  assign n57896 = decrypt_pad & ~\u0_uk_K_r9_reg[33]/NET0131  ;
  assign n57897 = ~decrypt_pad & ~\u0_uk_K_r9_reg[39]/NET0131  ;
  assign n57898 = ~n57896 & ~n57897 ;
  assign n57899 = \u0_R9_reg[4]/NET0131  & ~n57898 ;
  assign n57900 = ~\u0_R9_reg[4]/NET0131  & n57898 ;
  assign n57901 = ~n57899 & ~n57900 ;
  assign n57921 = n57894 & ~n57901 ;
  assign n57922 = n57888 & n57921 ;
  assign n57902 = decrypt_pad & ~\u0_uk_K_r9_reg[3]/NET0131  ;
  assign n57903 = ~decrypt_pad & ~\u0_uk_K_r9_reg[41]/NET0131  ;
  assign n57904 = ~n57902 & ~n57903 ;
  assign n57905 = \u0_R9_reg[6]/NET0131  & ~n57904 ;
  assign n57906 = ~\u0_R9_reg[6]/NET0131  & n57904 ;
  assign n57907 = ~n57905 & ~n57906 ;
  assign n57923 = ~n57894 & ~n57907 ;
  assign n57924 = ~n57901 & n57923 ;
  assign n57925 = ~n57922 & ~n57924 ;
  assign n57926 = n57920 & n57925 ;
  assign n57910 = ~n57888 & n57907 ;
  assign n57927 = ~n57901 & n57910 ;
  assign n57928 = ~n57920 & ~n57927 ;
  assign n57930 = n57901 & n57923 ;
  assign n57929 = ~n57888 & n57921 ;
  assign n57931 = n57888 & n57901 ;
  assign n57932 = ~n57929 & ~n57931 ;
  assign n57933 = ~n57930 & n57932 ;
  assign n57934 = n57928 & n57933 ;
  assign n57935 = ~n57926 & ~n57934 ;
  assign n57911 = n57894 & n57901 ;
  assign n57912 = ~n57894 & ~n57901 ;
  assign n57913 = ~n57911 & ~n57912 ;
  assign n57914 = n57910 & ~n57913 ;
  assign n57895 = n57888 & ~n57894 ;
  assign n57908 = n57901 & n57907 ;
  assign n57909 = n57895 & n57908 ;
  assign n57936 = decrypt_pad & ~\u0_uk_K_r9_reg[20]/NET0131  ;
  assign n57937 = ~decrypt_pad & ~\u0_uk_K_r9_reg[26]/NET0131  ;
  assign n57938 = ~n57936 & ~n57937 ;
  assign n57939 = \u0_R9_reg[8]/NET0131  & ~n57938 ;
  assign n57940 = ~\u0_R9_reg[8]/NET0131  & n57938 ;
  assign n57941 = ~n57939 & ~n57940 ;
  assign n57942 = ~n57909 & ~n57941 ;
  assign n57943 = ~n57914 & n57942 ;
  assign n57944 = ~n57935 & n57943 ;
  assign n57945 = ~n57888 & n57894 ;
  assign n57951 = ~n57895 & n57901 ;
  assign n57952 = ~n57945 & n57951 ;
  assign n57949 = n57888 & n57912 ;
  assign n57950 = n57907 & n57949 ;
  assign n57953 = n57920 & ~n57950 ;
  assign n57954 = ~n57952 & n57953 ;
  assign n57955 = ~n57909 & n57925 ;
  assign n57956 = n57928 & n57955 ;
  assign n57957 = ~n57954 & ~n57956 ;
  assign n57958 = n57907 & n57929 ;
  assign n57946 = ~n57920 & ~n57945 ;
  assign n57947 = n57901 & ~n57907 ;
  assign n57948 = ~n57946 & n57947 ;
  assign n57959 = n57941 & ~n57948 ;
  assign n57960 = ~n57958 & n57959 ;
  assign n57961 = ~n57957 & n57960 ;
  assign n57962 = ~n57944 & ~n57961 ;
  assign n57963 = ~\u0_L9_reg[28]/NET0131  & n57962 ;
  assign n57964 = \u0_L9_reg[28]/NET0131  & ~n57962 ;
  assign n57965 = ~n57963 & ~n57964 ;
  assign n57970 = ~n57566 & ~n57597 ;
  assign n57971 = ~n57579 & ~n57970 ;
  assign n57972 = ~n57638 & ~n57971 ;
  assign n57973 = n57572 & ~n57972 ;
  assign n57966 = ~n57559 & ~n57630 ;
  assign n57967 = n57598 & n57634 ;
  assign n57968 = ~n57966 & ~n57967 ;
  assign n57969 = ~n57572 & ~n57968 ;
  assign n57974 = n57596 & n57637 ;
  assign n57975 = ~n57969 & ~n57974 ;
  assign n57976 = ~n57973 & n57975 ;
  assign n57977 = ~n57613 & ~n57976 ;
  assign n57982 = n57615 & ~n57634 ;
  assign n57983 = ~n57967 & ~n57982 ;
  assign n57984 = n57572 & ~n57983 ;
  assign n57987 = n57559 & ~n57591 ;
  assign n57988 = ~n57625 & n57987 ;
  assign n57985 = ~n57565 & ~n57580 ;
  assign n57986 = n57572 & ~n57985 ;
  assign n57989 = ~n57966 & ~n57986 ;
  assign n57990 = ~n57988 & n57989 ;
  assign n57991 = ~n57984 & ~n57990 ;
  assign n57992 = n57613 & ~n57991 ;
  assign n57978 = ~n57565 & n57588 ;
  assign n57979 = n57580 & n57978 ;
  assign n57980 = n57565 & n57579 ;
  assign n57981 = n57594 & n57980 ;
  assign n57993 = ~n57979 & ~n57981 ;
  assign n57994 = ~n57992 & n57993 ;
  assign n57995 = ~n57977 & n57994 ;
  assign n57996 = \u0_L9_reg[29]/NET0131  & ~n57995 ;
  assign n57997 = ~\u0_L9_reg[29]/NET0131  & n57995 ;
  assign n57998 = ~n57996 & ~n57997 ;
  assign n58011 = n57693 & ~n57745 ;
  assign n58012 = n57740 & ~n58011 ;
  assign n58013 = ~n57673 & n57847 ;
  assign n58014 = ~n58012 & ~n58013 ;
  assign n58015 = n57672 & n57720 ;
  assign n58016 = ~n57733 & ~n58015 ;
  assign n58017 = ~n58014 & n58016 ;
  assign n58018 = n57690 & ~n58017 ;
  assign n57999 = ~n57702 & n57867 ;
  assign n58000 = n57665 & n57712 ;
  assign n58002 = n57730 & n57732 ;
  assign n58005 = ~n58000 & ~n58002 ;
  assign n58006 = ~n57999 & n58005 ;
  assign n58001 = ~n57679 & n57723 ;
  assign n58003 = n57691 & n57702 ;
  assign n58004 = ~n57727 & n58003 ;
  assign n58007 = ~n58001 & ~n58004 ;
  assign n58008 = n58006 & n58007 ;
  assign n58009 = n57684 & n58008 ;
  assign n58010 = ~n57690 & ~n58009 ;
  assign n58019 = ~n57683 & n58016 ;
  assign n58020 = ~n57702 & ~n58019 ;
  assign n58021 = ~n57711 & ~n57746 ;
  assign n58022 = ~n58020 & n58021 ;
  assign n58023 = ~n58010 & n58022 ;
  assign n58024 = ~n58018 & n58023 ;
  assign n58025 = ~\u0_L9_reg[10]/NET0131  & ~n58024 ;
  assign n58026 = \u0_L9_reg[10]/NET0131  & n58024 ;
  assign n58027 = ~n58025 & ~n58026 ;
  assign n58086 = decrypt_pad & ~\u0_uk_K_r9_reg[0]/P0001  ;
  assign n58087 = ~decrypt_pad & ~\u0_uk_K_r9_reg[8]/NET0131  ;
  assign n58088 = ~n58086 & ~n58087 ;
  assign n58089 = \u0_R9_reg[20]/NET0131  & ~n58088 ;
  assign n58090 = ~\u0_R9_reg[20]/NET0131  & n58088 ;
  assign n58091 = ~n58089 & ~n58090 ;
  assign n58056 = decrypt_pad & ~\u0_uk_K_r9_reg[16]/NET0131  ;
  assign n58057 = ~decrypt_pad & ~\u0_uk_K_r9_reg[52]/NET0131  ;
  assign n58058 = ~n58056 & ~n58057 ;
  assign n58059 = \u0_R9_reg[19]/NET0131  & ~n58058 ;
  assign n58060 = ~\u0_R9_reg[19]/NET0131  & n58058 ;
  assign n58061 = ~n58059 & ~n58060 ;
  assign n58048 = decrypt_pad & ~\u0_uk_K_r9_reg[35]/NET0131  ;
  assign n58049 = ~decrypt_pad & ~\u0_uk_K_r9_reg[43]/NET0131  ;
  assign n58050 = ~n58048 & ~n58049 ;
  assign n58051 = \u0_R9_reg[17]/NET0131  & ~n58050 ;
  assign n58052 = ~\u0_R9_reg[17]/NET0131  & n58050 ;
  assign n58053 = ~n58051 & ~n58052 ;
  assign n58034 = decrypt_pad & ~\u0_uk_K_r9_reg[44]/NET0131  ;
  assign n58035 = ~decrypt_pad & ~\u0_uk_K_r9_reg[21]/NET0131  ;
  assign n58036 = ~n58034 & ~n58035 ;
  assign n58037 = \u0_R9_reg[16]/NET0131  & ~n58036 ;
  assign n58038 = ~\u0_R9_reg[16]/NET0131  & n58036 ;
  assign n58039 = ~n58037 & ~n58038 ;
  assign n58041 = decrypt_pad & ~\u0_uk_K_r9_reg[1]/NET0131  ;
  assign n58042 = ~decrypt_pad & ~\u0_uk_K_r9_reg[9]/NET0131  ;
  assign n58043 = ~n58041 & ~n58042 ;
  assign n58044 = \u0_R9_reg[21]/NET0131  & ~n58043 ;
  assign n58045 = ~\u0_R9_reg[21]/NET0131  & n58043 ;
  assign n58046 = ~n58044 & ~n58045 ;
  assign n58093 = n58039 & ~n58046 ;
  assign n58094 = n58053 & n58093 ;
  assign n58028 = decrypt_pad & ~\u0_uk_K_r9_reg[29]/NET0131  ;
  assign n58029 = ~decrypt_pad & ~\u0_uk_K_r9_reg[37]/NET0131  ;
  assign n58030 = ~n58028 & ~n58029 ;
  assign n58031 = \u0_R9_reg[18]/NET0131  & ~n58030 ;
  assign n58032 = ~\u0_R9_reg[18]/NET0131  & n58030 ;
  assign n58033 = ~n58031 & ~n58032 ;
  assign n58054 = ~n58033 & n58053 ;
  assign n58055 = ~n58039 & n58054 ;
  assign n58040 = n58033 & n58039 ;
  assign n58095 = ~n58040 & n58046 ;
  assign n58096 = ~n58055 & n58095 ;
  assign n58097 = ~n58094 & ~n58096 ;
  assign n58098 = n58061 & ~n58097 ;
  assign n58062 = ~n58039 & ~n58046 ;
  assign n58063 = ~n58053 & n58062 ;
  assign n58075 = ~n58039 & n58046 ;
  assign n58101 = n58053 & n58075 ;
  assign n58102 = ~n58063 & ~n58101 ;
  assign n58103 = ~n58033 & ~n58061 ;
  assign n58104 = ~n58102 & n58103 ;
  assign n58072 = n58039 & n58046 ;
  assign n58073 = n58053 & n58072 ;
  assign n58105 = n58033 & ~n58061 ;
  assign n58106 = n58073 & n58105 ;
  assign n58099 = ~n58033 & n58072 ;
  assign n58100 = ~n58053 & n58099 ;
  assign n58107 = n58054 & n58093 ;
  assign n58108 = n58033 & ~n58053 ;
  assign n58109 = n58093 & n58108 ;
  assign n58110 = ~n58107 & ~n58109 ;
  assign n58111 = ~n58100 & n58110 ;
  assign n58112 = ~n58106 & n58111 ;
  assign n58113 = ~n58104 & n58112 ;
  assign n58114 = ~n58098 & n58113 ;
  assign n58115 = n58091 & ~n58114 ;
  assign n58047 = n58040 & n58046 ;
  assign n58064 = ~n58047 & n58061 ;
  assign n58065 = ~n58055 & ~n58063 ;
  assign n58066 = n58064 & n58065 ;
  assign n58076 = ~n58053 & n58075 ;
  assign n58067 = n58033 & n58053 ;
  assign n58068 = ~n58046 & n58067 ;
  assign n58077 = ~n58061 & ~n58068 ;
  assign n58078 = ~n58076 & n58077 ;
  assign n58069 = n58039 & ~n58053 ;
  assign n58070 = ~n58046 & n58069 ;
  assign n58071 = ~n58033 & n58070 ;
  assign n58074 = ~n58033 & n58073 ;
  assign n58079 = ~n58071 & ~n58074 ;
  assign n58080 = n58078 & n58079 ;
  assign n58081 = ~n58066 & ~n58080 ;
  assign n58082 = n58047 & ~n58053 ;
  assign n58083 = ~n58046 & n58055 ;
  assign n58084 = ~n58082 & ~n58083 ;
  assign n58085 = ~n58081 & n58084 ;
  assign n58092 = ~n58085 & ~n58091 ;
  assign n58116 = n58033 & n58063 ;
  assign n58117 = ~n58107 & ~n58116 ;
  assign n58118 = n58061 & ~n58117 ;
  assign n58119 = n58075 & n58108 ;
  assign n58120 = n58062 & n58067 ;
  assign n58121 = ~n58119 & ~n58120 ;
  assign n58122 = ~n58061 & ~n58121 ;
  assign n58123 = ~n58118 & ~n58122 ;
  assign n58124 = ~n58092 & n58123 ;
  assign n58125 = ~n58115 & n58124 ;
  assign n58126 = ~\u0_L9_reg[14]/NET0131  & ~n58125 ;
  assign n58127 = \u0_L9_reg[14]/NET0131  & n58125 ;
  assign n58128 = ~n58126 & ~n58127 ;
  assign n58129 = ~n57798 & ~n57824 ;
  assign n58130 = ~n57780 & n58129 ;
  assign n58131 = n57787 & ~n58130 ;
  assign n58132 = n57811 & n57817 ;
  assign n58133 = ~n58131 & ~n58132 ;
  assign n58134 = ~n57809 & ~n58133 ;
  assign n58138 = n57791 & n57827 ;
  assign n58135 = n57757 & n57816 ;
  assign n58137 = n57789 & n57797 ;
  assign n58140 = ~n58135 & ~n58137 ;
  assign n58141 = ~n58138 & n58140 ;
  assign n58136 = n57787 & n57812 ;
  assign n58139 = n57771 & n57777 ;
  assign n58142 = ~n58136 & ~n58139 ;
  assign n58143 = n58141 & n58142 ;
  assign n58144 = n57809 & ~n58143 ;
  assign n58146 = n57764 & ~n57809 ;
  assign n58145 = n57779 & n57816 ;
  assign n58148 = ~n58137 & ~n58145 ;
  assign n58149 = ~n58146 & n58148 ;
  assign n58147 = ~n57771 & ~n57787 ;
  assign n58150 = ~n57813 & n58147 ;
  assign n58151 = n58149 & n58150 ;
  assign n58152 = ~n57770 & n57780 ;
  assign n58153 = n57787 & ~n57833 ;
  assign n58154 = ~n58152 & n58153 ;
  assign n58155 = ~n58151 & ~n58154 ;
  assign n58156 = ~n58144 & ~n58155 ;
  assign n58157 = ~n58134 & n58156 ;
  assign n58158 = \u0_L9_reg[15]/P0001  & n58157 ;
  assign n58159 = ~\u0_L9_reg[15]/P0001  & ~n58157 ;
  assign n58160 = ~n58158 & ~n58159 ;
  assign n58162 = n57392 & ~n57405 ;
  assign n58163 = n57408 & n58162 ;
  assign n58161 = ~n57380 & n57409 ;
  assign n58173 = ~n57429 & ~n58161 ;
  assign n58174 = ~n58163 & n58173 ;
  assign n58172 = ~n57380 & ~n57433 ;
  assign n58175 = ~n57414 & ~n58172 ;
  assign n58176 = n58174 & n58175 ;
  assign n58164 = n57392 & n57431 ;
  assign n58165 = ~n57392 & n57409 ;
  assign n58166 = ~n58164 & ~n58165 ;
  assign n58167 = n57405 & ~n58166 ;
  assign n58168 = ~n57386 & n57406 ;
  assign n58169 = n57380 & n57444 ;
  assign n58170 = ~n58168 & ~n58169 ;
  assign n58171 = ~n57392 & ~n58170 ;
  assign n58177 = ~n58167 & ~n58171 ;
  assign n58178 = n58176 & n58177 ;
  assign n58182 = n57392 & n57399 ;
  assign n58183 = ~n57443 & ~n58182 ;
  assign n58184 = n57380 & ~n58183 ;
  assign n58181 = ~n57386 & ~n57449 ;
  assign n58180 = ~n57405 & ~n58166 ;
  assign n58179 = ~n57380 & n57445 ;
  assign n58185 = n57429 & ~n58179 ;
  assign n58186 = ~n58180 & n58185 ;
  assign n58187 = ~n58181 & n58186 ;
  assign n58188 = ~n58184 & n58187 ;
  assign n58189 = ~n58178 & ~n58188 ;
  assign n58190 = \u0_L9_reg[12]/NET0131  & n58189 ;
  assign n58191 = ~\u0_L9_reg[12]/NET0131  & ~n58189 ;
  assign n58192 = ~n58190 & ~n58191 ;
  assign n58193 = ~n57705 & ~n57713 ;
  assign n58194 = ~n57720 & n58193 ;
  assign n58195 = ~n57866 & n58194 ;
  assign n58196 = n57690 & ~n58195 ;
  assign n58197 = ~n57680 & n57702 ;
  assign n58198 = n58016 & n58197 ;
  assign n58199 = ~n58196 & n58198 ;
  assign n58200 = ~n57693 & n57745 ;
  assign n58201 = ~n57720 & ~n57863 ;
  assign n58202 = ~n58200 & n58201 ;
  assign n58203 = n57690 & ~n58202 ;
  assign n58204 = ~n57702 & ~n57721 ;
  assign n58205 = ~n57866 & n58204 ;
  assign n58206 = ~n58203 & n58205 ;
  assign n58207 = ~n58199 & ~n58206 ;
  assign n58208 = ~n57681 & ~n57705 ;
  assign n58209 = n57659 & ~n58208 ;
  assign n58210 = ~n57702 & ~n58209 ;
  assign n58211 = ~n57682 & n57742 ;
  assign n58212 = ~n58210 & ~n58211 ;
  assign n58213 = ~n57695 & n57745 ;
  assign n58214 = ~n57733 & ~n58213 ;
  assign n58215 = ~n58212 & n58214 ;
  assign n58216 = ~n57690 & ~n58215 ;
  assign n58217 = ~n58207 & ~n58216 ;
  assign n58218 = ~\u0_L9_reg[1]/NET0131  & ~n58217 ;
  assign n58219 = \u0_L9_reg[1]/NET0131  & n58217 ;
  assign n58220 = ~n58218 & ~n58219 ;
  assign n58223 = ~n57791 & n57817 ;
  assign n58224 = ~n57787 & ~n58223 ;
  assign n58225 = ~n58139 & n58224 ;
  assign n58227 = ~n57824 & ~n57834 ;
  assign n58228 = ~n58223 & ~n58227 ;
  assign n58226 = n57763 & n57779 ;
  assign n58229 = n57787 & ~n58226 ;
  assign n58230 = ~n58228 & n58229 ;
  assign n58231 = ~n58225 & ~n58230 ;
  assign n58221 = ~n57812 & ~n57825 ;
  assign n58222 = n57770 & ~n58221 ;
  assign n58232 = n57809 & ~n58152 ;
  assign n58233 = ~n58222 & n58232 ;
  assign n58234 = ~n58231 & n58233 ;
  assign n58235 = ~n57825 & ~n57835 ;
  assign n58236 = ~n57771 & n58235 ;
  assign n58237 = n57787 & ~n58236 ;
  assign n58241 = n57763 & n57789 ;
  assign n58245 = ~n57809 & ~n58241 ;
  assign n58246 = ~n57778 & n58245 ;
  assign n58242 = n57757 & n57777 ;
  assign n58243 = ~n57794 & ~n57816 ;
  assign n58244 = n58242 & ~n58243 ;
  assign n58238 = ~n57757 & ~n57787 ;
  assign n58239 = ~n57795 & ~n57797 ;
  assign n58240 = n58238 & ~n58239 ;
  assign n58247 = ~n57813 & ~n58240 ;
  assign n58248 = ~n58244 & n58247 ;
  assign n58249 = n58246 & n58248 ;
  assign n58250 = ~n58237 & n58249 ;
  assign n58251 = ~n58234 & ~n58250 ;
  assign n58252 = ~\u0_L9_reg[21]/NET0131  & n58251 ;
  assign n58253 = \u0_L9_reg[21]/NET0131  & ~n58251 ;
  assign n58254 = ~n58252 & ~n58253 ;
  assign n58258 = ~n58040 & ~n58046 ;
  assign n58259 = ~n58054 & n58258 ;
  assign n58257 = ~n58039 & ~n58053 ;
  assign n58260 = ~n58073 & ~n58257 ;
  assign n58261 = ~n58259 & n58260 ;
  assign n58262 = n58061 & ~n58261 ;
  assign n58263 = ~n58053 & n58072 ;
  assign n58264 = ~n58055 & ~n58263 ;
  assign n58265 = ~n58061 & ~n58264 ;
  assign n58255 = ~n58033 & n58046 ;
  assign n58256 = n58053 & n58255 ;
  assign n58266 = n58033 & n58094 ;
  assign n58267 = ~n58256 & ~n58266 ;
  assign n58268 = ~n58265 & n58267 ;
  assign n58269 = ~n58262 & n58268 ;
  assign n58270 = n58091 & ~n58269 ;
  assign n58278 = ~n58039 & n58067 ;
  assign n58279 = ~n58070 & ~n58278 ;
  assign n58280 = ~n58061 & ~n58279 ;
  assign n58282 = ~n58046 & n58061 ;
  assign n58283 = n58054 & n58282 ;
  assign n58277 = n58103 & n58257 ;
  assign n58281 = n58067 & n58075 ;
  assign n58284 = ~n58277 & ~n58281 ;
  assign n58285 = ~n58283 & n58284 ;
  assign n58286 = ~n58280 & n58285 ;
  assign n58287 = ~n58091 & ~n58286 ;
  assign n58271 = ~n58116 & ~n58266 ;
  assign n58272 = ~n58033 & n58075 ;
  assign n58273 = ~n58053 & n58272 ;
  assign n58274 = n58271 & ~n58273 ;
  assign n58275 = n58061 & ~n58274 ;
  assign n58276 = n58069 & n58105 ;
  assign n58288 = ~n58074 & ~n58276 ;
  assign n58289 = ~n58275 & n58288 ;
  assign n58290 = ~n58287 & n58289 ;
  assign n58291 = ~n58270 & n58290 ;
  assign n58292 = ~\u0_L9_reg[25]/NET0131  & ~n58291 ;
  assign n58293 = \u0_L9_reg[25]/NET0131  & n58291 ;
  assign n58294 = ~n58292 & ~n58293 ;
  assign n58298 = ~n57487 & ~n57505 ;
  assign n58299 = ~n57481 & n57532 ;
  assign n58300 = ~n58298 & ~n58299 ;
  assign n58301 = ~n57468 & ~n58300 ;
  assign n58302 = n57481 & n57487 ;
  assign n58303 = n57502 & n58302 ;
  assign n58304 = ~n57508 & ~n58303 ;
  assign n58305 = n57468 & ~n58304 ;
  assign n58295 = n57474 & n57487 ;
  assign n58296 = ~n57502 & n58295 ;
  assign n58297 = n57481 & n58296 ;
  assign n58306 = ~n57542 & ~n58297 ;
  assign n58307 = ~n58305 & n58306 ;
  assign n58308 = ~n58301 & n58307 ;
  assign n58309 = ~n57495 & ~n58308 ;
  assign n58311 = ~n57481 & n57502 ;
  assign n58312 = n57487 & n58311 ;
  assign n58313 = ~n57474 & ~n58312 ;
  assign n58310 = n57474 & ~n57518 ;
  assign n58314 = n57468 & ~n58310 ;
  assign n58315 = ~n58313 & n58314 ;
  assign n58318 = ~n57517 & ~n57528 ;
  assign n58319 = ~n57474 & n57481 ;
  assign n58320 = n57510 & n58319 ;
  assign n58321 = n58318 & ~n58320 ;
  assign n58322 = n57468 & ~n58321 ;
  assign n58323 = ~n57468 & ~n58319 ;
  assign n58324 = n58318 & n58323 ;
  assign n58316 = n57532 & n58302 ;
  assign n58317 = n57502 & n58295 ;
  assign n58325 = ~n58316 & ~n58317 ;
  assign n58326 = ~n58324 & n58325 ;
  assign n58327 = ~n58322 & n58326 ;
  assign n58328 = n57495 & ~n58327 ;
  assign n58329 = ~n58315 & ~n58328 ;
  assign n58330 = ~n58309 & n58329 ;
  assign n58331 = ~\u0_L9_reg[17]/NET0131  & ~n58330 ;
  assign n58332 = \u0_L9_reg[17]/NET0131  & n58330 ;
  assign n58333 = ~n58331 & ~n58332 ;
  assign n58334 = ~n57895 & ~n57929 ;
  assign n58335 = ~n57907 & ~n58334 ;
  assign n58345 = n57910 & n57920 ;
  assign n58346 = n57911 & n58345 ;
  assign n58347 = ~n58335 & ~n58346 ;
  assign n58336 = ~n57908 & ~n57945 ;
  assign n58337 = n57901 & n57945 ;
  assign n58338 = ~n57920 & ~n58337 ;
  assign n58339 = ~n58336 & n58338 ;
  assign n58340 = ~n57888 & ~n57920 ;
  assign n58341 = n57894 & ~n57907 ;
  assign n58342 = n58340 & n58341 ;
  assign n58343 = n57907 & n57922 ;
  assign n58344 = ~n58342 & ~n58343 ;
  assign n58348 = ~n58339 & n58344 ;
  assign n58349 = n58347 & n58348 ;
  assign n58350 = ~n57941 & ~n58349 ;
  assign n58351 = n57888 & ~n57907 ;
  assign n58352 = ~n57910 & ~n58351 ;
  assign n58353 = n57911 & ~n58352 ;
  assign n58354 = ~n57894 & ~n57908 ;
  assign n58355 = ~n58351 & n58354 ;
  assign n58356 = ~n58353 & ~n58355 ;
  assign n58357 = n57941 & ~n58356 ;
  assign n58358 = n57921 & n58352 ;
  assign n58359 = ~n57920 & ~n58358 ;
  assign n58360 = ~n58357 & n58359 ;
  assign n58362 = ~n57888 & n57923 ;
  assign n58363 = n57901 & n58362 ;
  assign n58364 = ~n57931 & ~n58351 ;
  assign n58365 = ~n58363 & n58364 ;
  assign n58366 = n57941 & ~n58365 ;
  assign n58367 = ~n57894 & n57910 ;
  assign n58368 = ~n57901 & n58367 ;
  assign n58361 = n57901 & n58351 ;
  assign n58369 = n57920 & ~n58361 ;
  assign n58370 = ~n58368 & n58369 ;
  assign n58371 = ~n58366 & n58370 ;
  assign n58372 = ~n58360 & ~n58371 ;
  assign n58373 = ~n58350 & ~n58372 ;
  assign n58374 = \u0_L9_reg[2]/NET0131  & n58373 ;
  assign n58375 = ~\u0_L9_reg[2]/NET0131  & ~n58373 ;
  assign n58376 = ~n58374 & ~n58375 ;
  assign n58378 = n57572 & ~n57620 ;
  assign n58377 = ~n57559 & n57602 ;
  assign n58379 = ~n57593 & ~n58377 ;
  assign n58380 = n58378 & n58379 ;
  assign n58381 = ~n57572 & ~n57616 ;
  assign n58382 = ~n57974 & n58381 ;
  assign n58383 = ~n58380 & ~n58382 ;
  assign n58384 = ~n57613 & ~n57642 ;
  assign n58385 = ~n57979 & n58384 ;
  assign n58386 = ~n58383 & n58385 ;
  assign n58388 = ~n57559 & ~n57591 ;
  assign n58387 = n57559 & ~n57980 ;
  assign n58389 = ~n57624 & ~n58387 ;
  assign n58390 = ~n58388 & n58389 ;
  assign n58391 = n57624 & ~n57636 ;
  assign n58392 = n57613 & ~n57617 ;
  assign n58393 = ~n58391 & n58392 ;
  assign n58394 = ~n58390 & n58393 ;
  assign n58395 = ~n58386 & ~n58394 ;
  assign n58399 = ~n57572 & ~n57638 ;
  assign n58396 = ~n57635 & ~n57637 ;
  assign n58397 = ~n57588 & n58396 ;
  assign n58398 = n58378 & ~n58397 ;
  assign n58400 = n57559 & ~n58398 ;
  assign n58401 = ~n58399 & n58400 ;
  assign n58402 = ~n57626 & ~n58401 ;
  assign n58403 = ~n58395 & n58402 ;
  assign n58404 = ~\u0_L9_reg[4]/NET0131  & ~n58403 ;
  assign n58405 = \u0_L9_reg[4]/NET0131  & n58403 ;
  assign n58406 = ~n58404 & ~n58405 ;
  assign n58423 = ~n57510 & ~n57518 ;
  assign n58424 = ~n57481 & ~n58423 ;
  assign n58425 = ~n57509 & ~n58424 ;
  assign n58426 = ~n57468 & ~n58425 ;
  assign n58427 = n57468 & ~n57532 ;
  assign n58428 = n57506 & n58427 ;
  assign n58429 = ~n57546 & ~n58320 ;
  assign n58430 = ~n58428 & n58429 ;
  assign n58431 = ~n58426 & n58430 ;
  assign n58432 = n57495 & ~n58431 ;
  assign n58414 = ~n57539 & ~n58302 ;
  assign n58415 = ~n57468 & ~n58414 ;
  assign n58416 = n57468 & n57518 ;
  assign n58417 = n57496 & n58311 ;
  assign n58418 = ~n57525 & ~n58317 ;
  assign n58419 = ~n58417 & n58418 ;
  assign n58420 = ~n58416 & n58419 ;
  assign n58421 = ~n58415 & n58420 ;
  assign n58422 = ~n57495 & ~n58421 ;
  assign n58407 = ~n57488 & ~n57518 ;
  assign n58408 = n57475 & ~n58407 ;
  assign n58410 = n57504 & n58295 ;
  assign n58409 = n57510 & n57511 ;
  assign n58411 = ~n58316 & ~n58409 ;
  assign n58412 = ~n58410 & n58411 ;
  assign n58413 = ~n57468 & ~n58412 ;
  assign n58433 = ~n58408 & ~n58413 ;
  assign n58434 = ~n58422 & n58433 ;
  assign n58435 = ~n58432 & n58434 ;
  assign n58436 = \u0_L9_reg[23]/NET0131  & ~n58435 ;
  assign n58437 = ~\u0_L9_reg[23]/NET0131  & n58435 ;
  assign n58438 = ~n58436 & ~n58437 ;
  assign n58442 = ~n58226 & n58235 ;
  assign n58443 = ~n57787 & ~n58442 ;
  assign n58440 = n57787 & ~n57815 ;
  assign n58441 = ~n58129 & n58440 ;
  assign n58439 = ~n57770 & n57791 ;
  assign n58444 = ~n57778 & ~n58439 ;
  assign n58445 = ~n57833 & n58444 ;
  assign n58446 = ~n58441 & n58445 ;
  assign n58447 = ~n58443 & n58446 ;
  assign n58448 = n57809 & ~n58447 ;
  assign n58452 = n57787 & ~n57798 ;
  assign n58451 = n57777 & ~n57816 ;
  assign n58453 = ~n58241 & ~n58451 ;
  assign n58454 = n58452 & n58453 ;
  assign n58450 = n57827 & n58242 ;
  assign n58449 = n57797 & n58238 ;
  assign n58455 = ~n57814 & ~n58449 ;
  assign n58456 = ~n58450 & n58455 ;
  assign n58457 = ~n58454 & n58456 ;
  assign n58458 = ~n57809 & ~n58457 ;
  assign n58461 = ~n57787 & n57820 ;
  assign n58459 = n57770 & n57787 ;
  assign n58460 = n57811 & n58459 ;
  assign n58462 = ~n57826 & ~n58460 ;
  assign n58463 = ~n58461 & n58462 ;
  assign n58464 = ~n58458 & n58463 ;
  assign n58465 = ~n58448 & n58464 ;
  assign n58466 = ~\u0_L9_reg[27]/NET0131  & ~n58465 ;
  assign n58467 = \u0_L9_reg[27]/NET0131  & n58465 ;
  assign n58468 = ~n58466 & ~n58467 ;
  assign n58469 = n57894 & n58361 ;
  assign n58470 = ~n57909 & ~n58469 ;
  assign n58471 = ~n57949 & ~n57958 ;
  assign n58472 = ~n58363 & n58471 ;
  assign n58473 = ~n57941 & ~n58472 ;
  assign n58474 = n58470 & ~n58473 ;
  assign n58475 = ~n57920 & ~n58474 ;
  assign n58480 = n57907 & n57951 ;
  assign n58478 = n57923 & n57931 ;
  assign n58479 = ~n57888 & ~n57913 ;
  assign n58481 = ~n58478 & ~n58479 ;
  assign n58482 = ~n58480 & n58481 ;
  assign n58483 = n57920 & ~n58482 ;
  assign n58476 = ~n57901 & ~n58340 ;
  assign n58477 = n58341 & n58476 ;
  assign n58484 = ~n57941 & ~n58477 ;
  assign n58485 = ~n58483 & n58484 ;
  assign n58486 = n58338 & ~n58367 ;
  assign n58487 = n57907 & n57921 ;
  assign n58488 = n57920 & ~n58362 ;
  assign n58489 = ~n58487 & n58488 ;
  assign n58490 = ~n58486 & ~n58489 ;
  assign n58491 = ~n57907 & n57949 ;
  assign n58492 = n57941 & ~n58491 ;
  assign n58493 = n58344 & n58492 ;
  assign n58494 = n58470 & n58493 ;
  assign n58495 = ~n58490 & n58494 ;
  assign n58496 = ~n58485 & ~n58495 ;
  assign n58497 = ~n58475 & ~n58496 ;
  assign n58498 = ~\u0_L9_reg[13]/NET0131  & n58497 ;
  assign n58499 = \u0_L9_reg[13]/NET0131  & ~n58497 ;
  assign n58500 = ~n58498 & ~n58499 ;
  assign n58506 = ~n57406 & ~n57444 ;
  assign n58509 = ~n57412 & n58506 ;
  assign n58510 = ~n57419 & ~n58509 ;
  assign n58507 = ~n57393 & ~n58162 ;
  assign n58508 = n58506 & n58507 ;
  assign n58511 = ~n57380 & ~n58508 ;
  assign n58512 = ~n58510 & n58511 ;
  assign n58501 = n57409 & n58162 ;
  assign n58502 = n57386 & n57406 ;
  assign n58503 = ~n57413 & ~n57440 ;
  assign n58504 = ~n58502 & n58503 ;
  assign n58505 = n57380 & ~n58504 ;
  assign n58513 = ~n58501 & ~n58505 ;
  assign n58514 = ~n58512 & n58513 ;
  assign n58515 = n57429 & ~n58514 ;
  assign n58517 = ~n57447 & ~n58168 ;
  assign n58518 = n57380 & ~n58517 ;
  assign n58523 = ~n57434 & ~n58518 ;
  assign n58519 = n57405 & n57409 ;
  assign n58520 = ~n58168 & ~n58519 ;
  assign n58521 = n57392 & ~n58520 ;
  assign n58522 = ~n58168 & n58172 ;
  assign n58524 = ~n58521 & ~n58522 ;
  assign n58525 = n58523 & n58524 ;
  assign n58526 = ~n57429 & ~n58525 ;
  assign n58516 = n57380 & n57445 ;
  assign n58527 = ~n57406 & n57438 ;
  assign n58528 = n57410 & n58527 ;
  assign n58529 = ~n58516 & ~n58528 ;
  assign n58530 = ~n58526 & n58529 ;
  assign n58531 = ~n58515 & n58530 ;
  assign n58532 = \u0_L9_reg[32]/NET0131  & n58531 ;
  assign n58533 = ~\u0_L9_reg[32]/NET0131  & ~n58531 ;
  assign n58534 = ~n58532 & ~n58533 ;
  assign n58573 = decrypt_pad & ~\u0_uk_K_r9_reg[40]/NET0131  ;
  assign n58574 = ~decrypt_pad & ~\u0_uk_K_r9_reg[46]/NET0131  ;
  assign n58575 = ~n58573 & ~n58574 ;
  assign n58576 = \u0_R9_reg[11]/P0001  & ~n58575 ;
  assign n58577 = ~\u0_R9_reg[11]/P0001  & n58575 ;
  assign n58578 = ~n58576 & ~n58577 ;
  assign n58561 = decrypt_pad & ~\u0_uk_K_r9_reg[55]/NET0131  ;
  assign n58562 = ~decrypt_pad & ~\u0_uk_K_r9_reg[4]/NET0131  ;
  assign n58563 = ~n58561 & ~n58562 ;
  assign n58564 = \u0_R9_reg[12]/NET0131  & ~n58563 ;
  assign n58565 = ~\u0_R9_reg[12]/NET0131  & n58563 ;
  assign n58566 = ~n58564 & ~n58565 ;
  assign n58535 = decrypt_pad & ~\u0_uk_K_r9_reg[11]/NET0131  ;
  assign n58536 = ~decrypt_pad & ~\u0_uk_K_r9_reg[17]/NET0131  ;
  assign n58537 = ~n58535 & ~n58536 ;
  assign n58538 = \u0_R9_reg[13]/NET0131  & ~n58537 ;
  assign n58539 = ~\u0_R9_reg[13]/NET0131  & n58537 ;
  assign n58540 = ~n58538 & ~n58539 ;
  assign n58548 = decrypt_pad & ~\u0_uk_K_r9_reg[6]/NET0131  ;
  assign n58549 = ~decrypt_pad & ~\u0_uk_K_r9_reg[12]/NET0131  ;
  assign n58550 = ~n58548 & ~n58549 ;
  assign n58551 = \u0_R9_reg[9]/NET0131  & ~n58550 ;
  assign n58552 = ~\u0_R9_reg[9]/NET0131  & n58550 ;
  assign n58553 = ~n58551 & ~n58552 ;
  assign n58570 = n58540 & ~n58553 ;
  assign n58554 = decrypt_pad & ~\u0_uk_K_r9_reg[39]/NET0131  ;
  assign n58555 = ~decrypt_pad & ~\u0_uk_K_r9_reg[20]/NET0131  ;
  assign n58556 = ~n58554 & ~n58555 ;
  assign n58557 = \u0_R9_reg[10]/NET0131  & ~n58556 ;
  assign n58558 = ~\u0_R9_reg[10]/NET0131  & n58556 ;
  assign n58559 = ~n58557 & ~n58558 ;
  assign n58541 = decrypt_pad & ~\u0_uk_K_r9_reg[34]/NET0131  ;
  assign n58542 = ~decrypt_pad & ~\u0_uk_K_r9_reg[40]/NET0131  ;
  assign n58543 = ~n58541 & ~n58542 ;
  assign n58544 = \u0_R9_reg[8]/NET0131  & ~n58543 ;
  assign n58545 = ~\u0_R9_reg[8]/NET0131  & n58543 ;
  assign n58546 = ~n58544 & ~n58545 ;
  assign n58583 = n58540 & ~n58546 ;
  assign n58603 = n58559 & n58583 ;
  assign n58569 = ~n58540 & n58553 ;
  assign n58604 = n58546 & n58569 ;
  assign n58605 = ~n58603 & ~n58604 ;
  assign n58606 = ~n58570 & n58605 ;
  assign n58607 = n58566 & ~n58606 ;
  assign n58602 = n58559 & n58570 ;
  assign n58547 = ~n58540 & ~n58546 ;
  assign n58588 = ~n58553 & ~n58559 ;
  assign n58608 = n58547 & n58588 ;
  assign n58609 = ~n58602 & ~n58608 ;
  assign n58610 = ~n58607 & n58609 ;
  assign n58611 = n58578 & ~n58610 ;
  assign n58560 = n58553 & n58559 ;
  assign n58586 = n58540 & n58546 ;
  assign n58587 = ~n58547 & ~n58586 ;
  assign n58589 = ~n58587 & ~n58588 ;
  assign n58590 = ~n58560 & n58589 ;
  assign n58584 = n58560 & n58583 ;
  assign n58585 = ~n58578 & n58584 ;
  assign n58571 = n58553 & ~n58559 ;
  assign n58593 = ~n58546 & n58578 ;
  assign n58594 = n58571 & n58593 ;
  assign n58597 = ~n58585 & ~n58594 ;
  assign n58591 = ~n58540 & n58560 ;
  assign n58592 = n58546 & n58591 ;
  assign n58595 = n58588 & ~n58593 ;
  assign n58596 = n58587 & n58595 ;
  assign n58598 = ~n58592 & ~n58596 ;
  assign n58599 = n58597 & n58598 ;
  assign n58600 = ~n58590 & n58599 ;
  assign n58601 = ~n58566 & ~n58600 ;
  assign n58567 = n58560 & n58566 ;
  assign n58568 = n58547 & n58567 ;
  assign n58572 = ~n58546 & ~n58571 ;
  assign n58579 = n58566 & ~n58578 ;
  assign n58580 = ~n58569 & ~n58570 ;
  assign n58581 = n58579 & n58580 ;
  assign n58582 = ~n58572 & n58581 ;
  assign n58612 = ~n58568 & ~n58582 ;
  assign n58613 = ~n58601 & n58612 ;
  assign n58614 = ~n58611 & n58613 ;
  assign n58615 = ~\u0_L9_reg[6]/NET0131  & ~n58614 ;
  assign n58616 = \u0_L9_reg[6]/NET0131  & n58614 ;
  assign n58617 = ~n58615 & ~n58616 ;
  assign n58618 = n57380 & ~n57429 ;
  assign n58619 = n57392 & ~n58506 ;
  assign n58620 = n57386 & n58619 ;
  assign n58621 = n57386 & ~n57446 ;
  assign n58622 = n58506 & ~n58621 ;
  assign n58623 = ~n58620 & ~n58622 ;
  assign n58624 = n58618 & ~n58623 ;
  assign n58626 = ~n57447 & ~n58619 ;
  assign n58627 = n57386 & ~n58626 ;
  assign n58628 = ~n57386 & n58509 ;
  assign n58625 = ~n57380 & n57429 ;
  assign n58629 = ~n58618 & ~n58625 ;
  assign n58630 = ~n58628 & n58629 ;
  assign n58631 = ~n58627 & n58630 ;
  assign n58632 = ~n58624 & ~n58631 ;
  assign n58633 = ~n57414 & ~n58632 ;
  assign n58634 = n57392 & ~n58502 ;
  assign n58635 = ~n57410 & ~n58634 ;
  assign n58636 = ~n58164 & n58625 ;
  assign n58637 = ~n58619 & n58636 ;
  assign n58638 = ~n58635 & n58637 ;
  assign n58639 = ~n58633 & ~n58638 ;
  assign n58640 = ~\u0_L9_reg[7]/NET0131  & n58639 ;
  assign n58641 = \u0_L9_reg[7]/NET0131  & ~n58639 ;
  assign n58642 = ~n58640 & ~n58641 ;
  assign n58655 = n58061 & ~n58071 ;
  assign n58656 = ~n58073 & n58655 ;
  assign n58657 = n58075 & ~n58108 ;
  assign n58658 = ~n58061 & ~n58263 ;
  assign n58659 = ~n58657 & n58658 ;
  assign n58660 = ~n58656 & ~n58659 ;
  assign n58661 = ~n58055 & n58271 ;
  assign n58662 = ~n58660 & n58661 ;
  assign n58663 = ~n58091 & ~n58662 ;
  assign n58643 = ~n58033 & n58063 ;
  assign n58644 = ~n58263 & ~n58643 ;
  assign n58645 = n58061 & ~n58644 ;
  assign n58646 = n58039 & n58103 ;
  assign n58647 = n58121 & ~n58646 ;
  assign n58648 = ~n58645 & n58647 ;
  assign n58649 = n58091 & ~n58648 ;
  assign n58650 = n58046 & n58055 ;
  assign n58651 = ~n58068 & ~n58119 ;
  assign n58652 = ~n58650 & n58651 ;
  assign n58653 = n58061 & ~n58652 ;
  assign n58654 = ~n58046 & n58276 ;
  assign n58664 = ~n58653 & ~n58654 ;
  assign n58665 = ~n58649 & n58664 ;
  assign n58666 = ~n58663 & n58665 ;
  assign n58667 = ~\u0_L9_reg[8]/NET0131  & ~n58666 ;
  assign n58668 = \u0_L9_reg[8]/NET0131  & n58666 ;
  assign n58669 = ~n58667 & ~n58668 ;
  assign n58672 = n57572 & ~n57599 ;
  assign n58681 = ~n57588 & ~n57635 ;
  assign n58682 = n58672 & ~n58681 ;
  assign n58679 = n57565 & n57592 ;
  assign n58680 = ~n57572 & n58397 ;
  assign n58683 = ~n58679 & ~n58680 ;
  assign n58684 = ~n58682 & n58683 ;
  assign n58685 = ~n57613 & ~n58684 ;
  assign n58673 = ~n57572 & ~n57978 ;
  assign n58674 = ~n58672 & ~n58673 ;
  assign n58670 = n57559 & n58397 ;
  assign n58671 = n58388 & ~n58396 ;
  assign n58675 = ~n57603 & ~n58671 ;
  assign n58676 = ~n58670 & n58675 ;
  assign n58677 = ~n58674 & n58676 ;
  assign n58678 = n57613 & ~n58677 ;
  assign n58686 = ~n57623 & ~n57643 ;
  assign n58687 = ~n58678 & n58686 ;
  assign n58688 = ~n58685 & n58687 ;
  assign n58689 = ~\u0_L9_reg[19]/P0001  & ~n58688 ;
  assign n58690 = \u0_L9_reg[19]/P0001  & n58688 ;
  assign n58691 = ~n58689 & ~n58690 ;
  assign n58697 = n58553 & n58586 ;
  assign n58698 = ~n58553 & ~n58586 ;
  assign n58699 = ~n58697 & ~n58698 ;
  assign n58700 = ~n58547 & ~n58699 ;
  assign n58701 = n58569 & n58593 ;
  assign n58702 = ~n58700 & ~n58701 ;
  assign n58703 = ~n58559 & ~n58702 ;
  assign n58692 = n58547 & n58559 ;
  assign n58693 = ~n58540 & ~n58559 ;
  assign n58694 = n58546 & n58693 ;
  assign n58695 = ~n58692 & ~n58694 ;
  assign n58696 = ~n58578 & ~n58695 ;
  assign n58704 = ~n58584 & ~n58696 ;
  assign n58705 = ~n58703 & n58704 ;
  assign n58706 = n58566 & ~n58705 ;
  assign n58707 = ~n58570 & ~n58693 ;
  assign n58708 = ~n58546 & ~n58707 ;
  assign n58709 = ~n58697 & ~n58708 ;
  assign n58710 = ~n58578 & ~n58709 ;
  assign n58711 = ~n58547 & n58578 ;
  assign n58712 = n58699 & n58711 ;
  assign n58713 = ~n58608 & ~n58712 ;
  assign n58714 = ~n58710 & n58713 ;
  assign n58715 = ~n58566 & ~n58714 ;
  assign n58716 = n58546 & n58559 ;
  assign n58717 = ~n58553 & n58716 ;
  assign n58718 = ~n58578 & n58717 ;
  assign n58719 = ~n58553 & n58692 ;
  assign n58720 = ~n58592 & ~n58719 ;
  assign n58721 = n58578 & ~n58720 ;
  assign n58722 = ~n58718 & ~n58721 ;
  assign n58723 = ~n58715 & n58722 ;
  assign n58724 = ~n58706 & n58723 ;
  assign n58725 = ~\u0_L9_reg[16]/NET0131  & ~n58724 ;
  assign n58726 = \u0_L9_reg[16]/NET0131  & n58724 ;
  assign n58727 = ~n58725 & ~n58726 ;
  assign n58739 = ~n58540 & n58717 ;
  assign n58740 = ~n58559 & n58583 ;
  assign n58741 = ~n58692 & ~n58740 ;
  assign n58742 = n58547 & n58553 ;
  assign n58743 = ~n58717 & ~n58742 ;
  assign n58744 = n58741 & n58743 ;
  assign n58745 = n58578 & ~n58744 ;
  assign n58746 = ~n58739 & ~n58745 ;
  assign n58747 = ~n58566 & ~n58746 ;
  assign n58731 = ~n58583 & n58588 ;
  assign n58730 = n58546 & n58560 ;
  assign n58732 = ~n58603 & ~n58730 ;
  assign n58733 = ~n58731 & n58732 ;
  assign n58734 = n58578 & ~n58733 ;
  assign n58735 = ~n58578 & n58589 ;
  assign n58736 = ~n58596 & ~n58735 ;
  assign n58737 = ~n58734 & n58736 ;
  assign n58738 = n58566 & ~n58737 ;
  assign n58748 = ~n58587 & n58588 ;
  assign n58749 = n58605 & ~n58748 ;
  assign n58750 = ~n58566 & ~n58578 ;
  assign n58751 = ~n58749 & n58750 ;
  assign n58754 = n58540 & n58594 ;
  assign n58728 = ~n58553 & n58578 ;
  assign n58729 = n58694 & n58728 ;
  assign n58752 = n58559 & ~n58578 ;
  assign n58753 = n58697 & n58752 ;
  assign n58755 = ~n58729 & ~n58753 ;
  assign n58756 = ~n58754 & n58755 ;
  assign n58757 = ~n58751 & n58756 ;
  assign n58758 = ~n58738 & n58757 ;
  assign n58759 = ~n58747 & n58758 ;
  assign n58760 = ~\u0_L9_reg[24]/NET0131  & ~n58759 ;
  assign n58761 = \u0_L9_reg[24]/NET0131  & n58759 ;
  assign n58762 = ~n58760 & ~n58761 ;
  assign n58764 = ~n58569 & ~n58716 ;
  assign n58768 = n58578 & ~n58591 ;
  assign n58769 = ~n58764 & n58768 ;
  assign n58765 = ~n58546 & ~n58553 ;
  assign n58766 = ~n58578 & ~n58765 ;
  assign n58767 = n58764 & n58766 ;
  assign n58763 = ~n58553 & n58603 ;
  assign n58770 = ~n58748 & ~n58763 ;
  assign n58771 = ~n58767 & n58770 ;
  assign n58772 = ~n58769 & n58771 ;
  assign n58773 = ~n58566 & ~n58772 ;
  assign n58774 = n58578 & ~n58741 ;
  assign n58775 = ~n58729 & ~n58774 ;
  assign n58776 = n58566 & ~n58775 ;
  assign n58777 = ~n58716 & ~n58742 ;
  assign n58778 = n58579 & ~n58777 ;
  assign n58781 = n58559 & n58586 ;
  assign n58782 = n58728 & n58781 ;
  assign n58779 = n58567 & ~n58586 ;
  assign n58780 = ~n58578 & n58591 ;
  assign n58783 = ~n58779 & ~n58780 ;
  assign n58784 = ~n58782 & n58783 ;
  assign n58785 = ~n58778 & n58784 ;
  assign n58786 = ~n58776 & n58785 ;
  assign n58787 = ~n58773 & n58786 ;
  assign n58788 = \u0_L9_reg[30]/NET0131  & ~n58787 ;
  assign n58789 = ~\u0_L9_reg[30]/NET0131  & n58787 ;
  assign n58790 = ~n58788 & ~n58789 ;
  assign n58792 = n58053 & n58062 ;
  assign n58793 = ~n58099 & ~n58792 ;
  assign n58794 = n58061 & ~n58793 ;
  assign n58791 = ~n58061 & n58101 ;
  assign n58795 = n58091 & ~n58109 ;
  assign n58796 = ~n58074 & n58795 ;
  assign n58797 = ~n58791 & n58796 ;
  assign n58798 = ~n58794 & n58797 ;
  assign n58803 = ~n58094 & ~n58272 ;
  assign n58804 = n58061 & ~n58803 ;
  assign n58800 = ~n58069 & n58255 ;
  assign n58799 = n58061 & ~n58108 ;
  assign n58801 = ~n58093 & ~n58799 ;
  assign n58802 = ~n58800 & n58801 ;
  assign n58805 = ~n58091 & ~n58802 ;
  assign n58806 = ~n58804 & n58805 ;
  assign n58807 = ~n58798 & ~n58806 ;
  assign n58808 = ~n58119 & n58655 ;
  assign n58809 = ~n58061 & ~n58107 ;
  assign n58810 = ~n58082 & n58809 ;
  assign n58811 = ~n58643 & n58810 ;
  assign n58812 = ~n58808 & ~n58811 ;
  assign n58813 = ~n58807 & ~n58812 ;
  assign n58814 = ~\u0_L9_reg[3]/NET0131  & ~n58813 ;
  assign n58815 = \u0_L9_reg[3]/NET0131  & n58813 ;
  assign n58816 = ~n58814 & ~n58815 ;
  assign n58827 = n57920 & ~n58334 ;
  assign n58828 = n57894 & n57907 ;
  assign n58829 = ~n57920 & ~n58828 ;
  assign n58830 = n57951 & n58829 ;
  assign n58831 = ~n58368 & ~n58830 ;
  assign n58832 = ~n58827 & n58831 ;
  assign n58833 = n57941 & ~n58832 ;
  assign n58818 = n57888 & n57920 ;
  assign n58821 = ~n57901 & ~n58818 ;
  assign n58822 = n58352 & n58821 ;
  assign n58819 = ~n57910 & ~n58818 ;
  assign n58820 = n57911 & ~n58819 ;
  assign n58823 = ~n57909 & ~n58362 ;
  assign n58824 = ~n58820 & n58823 ;
  assign n58825 = ~n58822 & n58824 ;
  assign n58826 = ~n57941 & ~n58825 ;
  assign n58817 = ~n57920 & n57922 ;
  assign n58834 = n57901 & n58828 ;
  assign n58835 = ~n58491 & ~n58834 ;
  assign n58836 = n57920 & ~n58835 ;
  assign n58837 = ~n58817 & ~n58836 ;
  assign n58838 = ~n58826 & n58837 ;
  assign n58839 = ~n58833 & n58838 ;
  assign n58840 = \u0_L9_reg[18]/NET0131  & n58839 ;
  assign n58841 = ~\u0_L9_reg[18]/NET0131  & ~n58839 ;
  assign n58842 = ~n58840 & ~n58841 ;
  assign n58843 = decrypt_pad & ~\u0_uk_K_r8_reg[33]/NET0131  ;
  assign n58844 = ~decrypt_pad & ~\u0_uk_K_r8_reg[11]/NET0131  ;
  assign n58845 = ~n58843 & ~n58844 ;
  assign n58846 = \u0_R8_reg[4]/NET0131  & ~n58845 ;
  assign n58847 = ~\u0_R8_reg[4]/NET0131  & n58845 ;
  assign n58848 = ~n58846 & ~n58847 ;
  assign n58862 = decrypt_pad & ~\u0_uk_K_r8_reg[10]/NET0131  ;
  assign n58863 = ~decrypt_pad & ~\u0_uk_K_r8_reg[20]/NET0131  ;
  assign n58864 = ~n58862 & ~n58863 ;
  assign n58865 = \u0_R8_reg[32]/NET0131  & ~n58864 ;
  assign n58866 = ~\u0_R8_reg[32]/NET0131  & n58864 ;
  assign n58867 = ~n58865 & ~n58866 ;
  assign n58868 = decrypt_pad & ~\u0_uk_K_r8_reg[4]/NET0131  ;
  assign n58869 = ~decrypt_pad & ~\u0_uk_K_r8_reg[39]/NET0131  ;
  assign n58870 = ~n58868 & ~n58869 ;
  assign n58871 = \u0_R8_reg[5]/NET0131  & ~n58870 ;
  assign n58872 = ~\u0_R8_reg[5]/NET0131  & n58870 ;
  assign n58873 = ~n58871 & ~n58872 ;
  assign n58875 = ~n58867 & ~n58873 ;
  assign n58849 = decrypt_pad & ~\u0_uk_K_r8_reg[55]/NET0131  ;
  assign n58850 = ~decrypt_pad & ~\u0_uk_K_r8_reg[33]/NET0131  ;
  assign n58851 = ~n58849 & ~n58850 ;
  assign n58852 = \u0_R8_reg[3]/NET0131  & ~n58851 ;
  assign n58853 = ~\u0_R8_reg[3]/NET0131  & n58851 ;
  assign n58854 = ~n58852 & ~n58853 ;
  assign n58855 = decrypt_pad & ~\u0_uk_K_r8_reg[46]/NET0131  ;
  assign n58856 = ~decrypt_pad & ~\u0_uk_K_r8_reg[24]/NET0131  ;
  assign n58857 = ~n58855 & ~n58856 ;
  assign n58858 = \u0_R8_reg[2]/NET0131  & ~n58857 ;
  assign n58859 = ~\u0_R8_reg[2]/NET0131  & n58857 ;
  assign n58860 = ~n58858 & ~n58859 ;
  assign n58885 = ~n58860 & ~n58867 ;
  assign n58906 = n58854 & n58885 ;
  assign n58876 = decrypt_pad & ~\u0_uk_K_r8_reg[6]/NET0131  ;
  assign n58877 = ~decrypt_pad & ~\u0_uk_K_r8_reg[41]/NET0131  ;
  assign n58878 = ~n58876 & ~n58877 ;
  assign n58879 = \u0_R8_reg[1]/NET0131  & ~n58878 ;
  assign n58880 = ~\u0_R8_reg[1]/NET0131  & n58878 ;
  assign n58881 = ~n58879 & ~n58880 ;
  assign n58888 = ~n58873 & ~n58881 ;
  assign n58904 = ~n58860 & n58888 ;
  assign n58905 = ~n58867 & ~n58881 ;
  assign n58907 = ~n58904 & ~n58905 ;
  assign n58908 = ~n58906 & n58907 ;
  assign n58909 = ~n58875 & ~n58908 ;
  assign n58886 = n58873 & ~n58881 ;
  assign n58910 = n58860 & n58875 ;
  assign n58911 = ~n58886 & ~n58910 ;
  assign n58912 = n58854 & ~n58911 ;
  assign n58902 = ~n58854 & n58867 ;
  assign n58903 = n58881 & n58902 ;
  assign n58913 = n58860 & n58905 ;
  assign n58914 = ~n58903 & ~n58913 ;
  assign n58915 = ~n58912 & n58914 ;
  assign n58916 = ~n58909 & n58915 ;
  assign n58917 = n58848 & ~n58916 ;
  assign n58874 = n58867 & n58873 ;
  assign n58893 = ~n58854 & n58881 ;
  assign n58894 = n58874 & ~n58893 ;
  assign n58895 = ~n58873 & n58881 ;
  assign n58896 = ~n58867 & n58895 ;
  assign n58897 = ~n58894 & ~n58896 ;
  assign n58898 = ~n58860 & ~n58897 ;
  assign n58861 = n58854 & n58860 ;
  assign n58882 = ~n58875 & n58881 ;
  assign n58883 = ~n58874 & n58882 ;
  assign n58884 = n58861 & n58883 ;
  assign n58887 = n58885 & ~n58886 ;
  assign n58889 = n58860 & n58867 ;
  assign n58890 = n58888 & n58889 ;
  assign n58891 = ~n58887 & ~n58890 ;
  assign n58892 = ~n58854 & ~n58891 ;
  assign n58899 = ~n58884 & ~n58892 ;
  assign n58900 = ~n58898 & n58899 ;
  assign n58901 = ~n58848 & ~n58900 ;
  assign n58921 = n58860 & n58873 ;
  assign n58922 = n58881 & n58921 ;
  assign n58923 = n58867 & n58922 ;
  assign n58924 = ~n58895 & ~n58921 ;
  assign n58925 = n58860 & ~n58905 ;
  assign n58926 = ~n58924 & ~n58925 ;
  assign n58927 = ~n58923 & ~n58926 ;
  assign n58928 = ~n58854 & ~n58927 ;
  assign n58918 = ~n58860 & ~n58881 ;
  assign n58919 = n58854 & n58867 ;
  assign n58920 = n58918 & n58919 ;
  assign n58929 = n58861 & ~n58881 ;
  assign n58930 = n58875 & n58929 ;
  assign n58931 = ~n58920 & ~n58930 ;
  assign n58932 = ~n58928 & n58931 ;
  assign n58933 = ~n58901 & n58932 ;
  assign n58934 = ~n58917 & n58933 ;
  assign n58935 = ~\u0_L8_reg[31]/NET0131  & ~n58934 ;
  assign n58936 = \u0_L8_reg[31]/NET0131  & n58934 ;
  assign n58937 = ~n58935 & ~n58936 ;
  assign n58938 = decrypt_pad & ~\u0_uk_K_r8_reg[2]/NET0131  ;
  assign n58939 = ~decrypt_pad & ~\u0_uk_K_r8_reg[37]/P0001  ;
  assign n58940 = ~n58938 & ~n58939 ;
  assign n58941 = \u0_R8_reg[24]/NET0131  & ~n58940 ;
  assign n58942 = ~\u0_R8_reg[24]/NET0131  & n58940 ;
  assign n58943 = ~n58941 & ~n58942 ;
  assign n58957 = decrypt_pad & ~\u0_uk_K_r8_reg[0]/NET0131  ;
  assign n58958 = ~decrypt_pad & ~\u0_uk_K_r8_reg[35]/NET0131  ;
  assign n58959 = ~n58957 & ~n58958 ;
  assign n58960 = \u0_R8_reg[23]/NET0131  & ~n58959 ;
  assign n58961 = ~\u0_R8_reg[23]/NET0131  & n58959 ;
  assign n58962 = ~n58960 & ~n58961 ;
  assign n58944 = decrypt_pad & ~\u0_uk_K_r8_reg[36]/NET0131  ;
  assign n58945 = ~decrypt_pad & ~\u0_uk_K_r8_reg[16]/NET0131  ;
  assign n58946 = ~n58944 & ~n58945 ;
  assign n58947 = \u0_R8_reg[20]/NET0131  & ~n58946 ;
  assign n58948 = ~\u0_R8_reg[20]/NET0131  & n58946 ;
  assign n58949 = ~n58947 & ~n58948 ;
  assign n58970 = decrypt_pad & ~\u0_uk_K_r8_reg[51]/NET0131  ;
  assign n58971 = ~decrypt_pad & ~\u0_uk_K_r8_reg[0]/NET0131  ;
  assign n58972 = ~n58970 & ~n58971 ;
  assign n58973 = \u0_R8_reg[21]/NET0131  & ~n58972 ;
  assign n58974 = ~\u0_R8_reg[21]/NET0131  & n58972 ;
  assign n58975 = ~n58973 & ~n58974 ;
  assign n58982 = n58949 & ~n58975 ;
  assign n58950 = decrypt_pad & ~\u0_uk_K_r8_reg[21]/NET0131  ;
  assign n58951 = ~decrypt_pad & ~\u0_uk_K_r8_reg[1]/NET0131  ;
  assign n58952 = ~n58950 & ~n58951 ;
  assign n58953 = \u0_R8_reg[25]/NET0131  & ~n58952 ;
  assign n58954 = ~\u0_R8_reg[25]/NET0131  & n58952 ;
  assign n58955 = ~n58953 & ~n58954 ;
  assign n58963 = decrypt_pad & ~\u0_uk_K_r8_reg[42]/NET0131  ;
  assign n58964 = ~decrypt_pad & ~\u0_uk_K_r8_reg[22]/NET0131  ;
  assign n58965 = ~n58963 & ~n58964 ;
  assign n58966 = \u0_R8_reg[22]/NET0131  & ~n58965 ;
  assign n58967 = ~\u0_R8_reg[22]/NET0131  & n58965 ;
  assign n58968 = ~n58966 & ~n58967 ;
  assign n59013 = ~n58955 & ~n58968 ;
  assign n59014 = n58982 & n59013 ;
  assign n58985 = ~n58949 & n58975 ;
  assign n58986 = n58968 & n58985 ;
  assign n58998 = n58949 & n58955 ;
  assign n59012 = n58975 & n58998 ;
  assign n59015 = ~n58986 & ~n59012 ;
  assign n59016 = ~n59014 & n59015 ;
  assign n59017 = n58962 & ~n59016 ;
  assign n58969 = ~n58962 & ~n58968 ;
  assign n59018 = n58969 & n58998 ;
  assign n59019 = ~n58975 & n59018 ;
  assign n59000 = ~n58968 & ~n58975 ;
  assign n59020 = ~n58986 & ~n59000 ;
  assign n59021 = ~n58962 & ~n58998 ;
  assign n59022 = ~n59013 & n59021 ;
  assign n59023 = n59020 & n59022 ;
  assign n59024 = ~n59019 & ~n59023 ;
  assign n59025 = ~n59017 & n59024 ;
  assign n59026 = n58943 & ~n59025 ;
  assign n58983 = n58968 & n58982 ;
  assign n58984 = n58955 & n58983 ;
  assign n58956 = n58949 & ~n58955 ;
  assign n58976 = ~n58968 & n58975 ;
  assign n58977 = ~n58969 & ~n58976 ;
  assign n58978 = n58956 & ~n58977 ;
  assign n58979 = ~n58949 & ~n58975 ;
  assign n58980 = n58955 & n58979 ;
  assign n58981 = n58962 & n58980 ;
  assign n58993 = ~n58978 & ~n58981 ;
  assign n58994 = ~n58984 & n58993 ;
  assign n58987 = n58949 & n58976 ;
  assign n58988 = ~n58986 & ~n58987 ;
  assign n58989 = ~n58962 & ~n58988 ;
  assign n58990 = ~n58949 & ~n58968 ;
  assign n58991 = ~n58983 & ~n58990 ;
  assign n58992 = n58962 & ~n58991 ;
  assign n58995 = ~n58989 & ~n58992 ;
  assign n58996 = n58994 & n58995 ;
  assign n58997 = ~n58943 & ~n58996 ;
  assign n59006 = n58956 & n58975 ;
  assign n59007 = ~n58962 & n59006 ;
  assign n59008 = ~n58981 & ~n59007 ;
  assign n59009 = ~n58968 & ~n59008 ;
  assign n59001 = ~n58949 & ~n58955 ;
  assign n59002 = ~n58968 & ~n59001 ;
  assign n58999 = n58968 & ~n58998 ;
  assign n59003 = n58962 & ~n59000 ;
  assign n59004 = ~n58999 & n59003 ;
  assign n59005 = ~n59002 & n59004 ;
  assign n59010 = ~n58975 & n59001 ;
  assign n59011 = n58969 & n59010 ;
  assign n59027 = ~n59005 & ~n59011 ;
  assign n59028 = ~n59009 & n59027 ;
  assign n59029 = ~n58997 & n59028 ;
  assign n59030 = ~n59026 & n59029 ;
  assign n59031 = ~\u0_L8_reg[11]/NET0131  & n59030 ;
  assign n59032 = \u0_L8_reg[11]/NET0131  & ~n59030 ;
  assign n59033 = ~n59031 & ~n59032 ;
  assign n59063 = decrypt_pad & ~\u0_uk_K_r8_reg[9]/P0001  ;
  assign n59064 = ~decrypt_pad & ~\u0_uk_K_r8_reg[44]/NET0131  ;
  assign n59065 = ~n59063 & ~n59064 ;
  assign n59066 = \u0_R8_reg[28]/NET0131  & ~n59065 ;
  assign n59067 = ~\u0_R8_reg[28]/NET0131  & n59065 ;
  assign n59068 = ~n59066 & ~n59067 ;
  assign n59049 = decrypt_pad & ~\u0_uk_K_r8_reg[22]/NET0131  ;
  assign n59050 = ~decrypt_pad & ~\u0_uk_K_r8_reg[2]/NET0131  ;
  assign n59051 = ~n59049 & ~n59050 ;
  assign n59052 = \u0_R8_reg[27]/NET0131  & ~n59051 ;
  assign n59053 = ~\u0_R8_reg[27]/NET0131  & n59051 ;
  assign n59054 = ~n59052 & ~n59053 ;
  assign n59034 = decrypt_pad & ~\u0_uk_K_r8_reg[52]/NET0131  ;
  assign n59035 = ~decrypt_pad & ~\u0_uk_K_r8_reg[28]/NET0131  ;
  assign n59036 = ~n59034 & ~n59035 ;
  assign n59037 = \u0_R8_reg[24]/NET0131  & ~n59036 ;
  assign n59038 = ~\u0_R8_reg[24]/NET0131  & n59036 ;
  assign n59039 = ~n59037 & ~n59038 ;
  assign n59055 = decrypt_pad & ~\u0_uk_K_r8_reg[28]/NET0131  ;
  assign n59056 = ~decrypt_pad & ~\u0_uk_K_r8_reg[8]/NET0131  ;
  assign n59057 = ~n59055 & ~n59056 ;
  assign n59058 = \u0_R8_reg[25]/NET0131  & ~n59057 ;
  assign n59059 = ~\u0_R8_reg[25]/NET0131  & n59057 ;
  assign n59060 = ~n59058 & ~n59059 ;
  assign n59069 = decrypt_pad & ~\u0_uk_K_r8_reg[1]/NET0131  ;
  assign n59070 = ~decrypt_pad & ~\u0_uk_K_r8_reg[36]/NET0131  ;
  assign n59071 = ~n59069 & ~n59070 ;
  assign n59072 = \u0_R8_reg[29]/NET0131  & ~n59071 ;
  assign n59073 = ~\u0_R8_reg[29]/NET0131  & n59071 ;
  assign n59074 = ~n59072 & ~n59073 ;
  assign n59077 = n59060 & ~n59074 ;
  assign n59040 = decrypt_pad & ~\u0_uk_K_r8_reg[44]/NET0131  ;
  assign n59041 = ~decrypt_pad & ~\u0_uk_K_r8_reg[52]/NET0131  ;
  assign n59042 = ~n59040 & ~n59041 ;
  assign n59043 = \u0_R8_reg[26]/NET0131  & ~n59042 ;
  assign n59044 = ~\u0_R8_reg[26]/NET0131  & n59042 ;
  assign n59045 = ~n59043 & ~n59044 ;
  assign n59078 = n59045 & n59074 ;
  assign n59079 = ~n59077 & ~n59078 ;
  assign n59080 = n59039 & ~n59079 ;
  assign n59081 = ~n59039 & ~n59060 ;
  assign n59082 = n59045 & ~n59074 ;
  assign n59083 = n59081 & n59082 ;
  assign n59084 = ~n59080 & ~n59083 ;
  assign n59085 = ~n59054 & ~n59084 ;
  assign n59088 = ~n59045 & ~n59060 ;
  assign n59086 = ~n59054 & n59074 ;
  assign n59089 = n59039 & ~n59086 ;
  assign n59090 = n59088 & n59089 ;
  assign n59046 = ~n59039 & ~n59045 ;
  assign n59047 = n59039 & n59045 ;
  assign n59048 = ~n59046 & ~n59047 ;
  assign n59075 = n59060 & n59074 ;
  assign n59076 = ~n59048 & n59075 ;
  assign n59087 = n59046 & n59086 ;
  assign n59091 = ~n59076 & ~n59087 ;
  assign n59092 = ~n59090 & n59091 ;
  assign n59093 = ~n59085 & n59092 ;
  assign n59094 = ~n59068 & ~n59093 ;
  assign n59110 = n59045 & n59060 ;
  assign n59111 = ~n59088 & ~n59110 ;
  assign n59112 = n59039 & n59054 ;
  assign n59113 = ~n59077 & n59112 ;
  assign n59114 = n59111 & n59113 ;
  assign n59103 = ~n59045 & n59074 ;
  assign n59104 = ~n59082 & ~n59103 ;
  assign n59105 = n59081 & n59104 ;
  assign n59106 = n59039 & n59060 ;
  assign n59107 = ~n59081 & ~n59106 ;
  assign n59108 = ~n59047 & n59086 ;
  assign n59109 = n59107 & n59108 ;
  assign n59115 = ~n59105 & ~n59109 ;
  assign n59116 = ~n59114 & n59115 ;
  assign n59117 = n59068 & ~n59116 ;
  assign n59061 = ~n59054 & n59060 ;
  assign n59062 = ~n59048 & n59061 ;
  assign n59095 = ~n59039 & n59045 ;
  assign n59096 = ~n59060 & n59074 ;
  assign n59097 = ~n59077 & ~n59096 ;
  assign n59098 = n59095 & ~n59097 ;
  assign n59099 = ~n59060 & ~n59074 ;
  assign n59100 = ~n59095 & n59099 ;
  assign n59101 = ~n59098 & ~n59100 ;
  assign n59102 = n59054 & ~n59101 ;
  assign n59118 = ~n59062 & ~n59102 ;
  assign n59119 = ~n59117 & n59118 ;
  assign n59120 = ~n59094 & n59119 ;
  assign n59121 = ~\u0_L8_reg[22]/NET0131  & ~n59120 ;
  assign n59122 = \u0_L8_reg[22]/NET0131  & n59120 ;
  assign n59123 = ~n59121 & ~n59122 ;
  assign n59137 = ~n58874 & ~n58875 ;
  assign n59138 = ~n58881 & ~n59137 ;
  assign n59139 = ~n58860 & n58875 ;
  assign n59140 = ~n59138 & ~n59139 ;
  assign n59141 = ~n58854 & ~n59140 ;
  assign n59142 = ~n58886 & ~n58895 ;
  assign n59143 = n58919 & n59142 ;
  assign n59136 = n58905 & n58921 ;
  assign n59144 = n58889 & n58895 ;
  assign n59145 = ~n59136 & ~n59144 ;
  assign n59146 = ~n59143 & n59145 ;
  assign n59147 = ~n59141 & n59146 ;
  assign n59148 = ~n58848 & ~n59147 ;
  assign n59126 = ~n58867 & ~n58918 ;
  assign n59127 = n58874 & n58918 ;
  assign n59128 = ~n59126 & ~n59127 ;
  assign n59129 = n58854 & ~n59128 ;
  assign n59124 = ~n58860 & n58867 ;
  assign n59130 = ~n58854 & ~n59124 ;
  assign n59131 = ~n59126 & n59130 ;
  assign n59125 = n58895 & n59124 ;
  assign n59132 = ~n58922 & ~n59125 ;
  assign n59133 = ~n59131 & n59132 ;
  assign n59134 = ~n59129 & n59133 ;
  assign n59135 = n58848 & ~n59134 ;
  assign n59149 = n58873 & n58885 ;
  assign n59150 = ~n58910 & ~n59149 ;
  assign n59151 = n58854 & n58881 ;
  assign n59152 = ~n59150 & n59151 ;
  assign n59153 = ~n59135 & ~n59152 ;
  assign n59154 = ~n59148 & n59153 ;
  assign n59155 = ~\u0_L8_reg[17]/NET0131  & ~n59154 ;
  assign n59156 = \u0_L8_reg[17]/NET0131  & n59154 ;
  assign n59157 = ~n59155 & ~n59156 ;
  assign n59164 = decrypt_pad & ~\u0_uk_K_r8_reg[18]/NET0131  ;
  assign n59165 = ~decrypt_pad & ~\u0_uk_K_r8_reg[53]/NET0131  ;
  assign n59166 = ~n59164 & ~n59165 ;
  assign n59167 = \u0_R8_reg[13]/NET0131  & ~n59166 ;
  assign n59168 = ~\u0_R8_reg[13]/NET0131  & n59166 ;
  assign n59169 = ~n59167 & ~n59168 ;
  assign n59189 = decrypt_pad & ~\u0_uk_K_r8_reg[27]/NET0131  ;
  assign n59190 = ~decrypt_pad & ~\u0_uk_K_r8_reg[5]/NET0131  ;
  assign n59191 = ~n59189 & ~n59190 ;
  assign n59192 = \u0_R8_reg[15]/NET0131  & ~n59191 ;
  assign n59193 = ~\u0_R8_reg[15]/NET0131  & n59191 ;
  assign n59194 = ~n59192 & ~n59193 ;
  assign n59158 = decrypt_pad & ~\u0_uk_K_r8_reg[40]/NET0131  ;
  assign n59159 = ~decrypt_pad & ~\u0_uk_K_r8_reg[18]/NET0131  ;
  assign n59160 = ~n59158 & ~n59159 ;
  assign n59161 = \u0_R8_reg[17]/NET0131  & ~n59160 ;
  assign n59162 = ~\u0_R8_reg[17]/NET0131  & n59160 ;
  assign n59163 = ~n59161 & ~n59162 ;
  assign n59171 = decrypt_pad & ~\u0_uk_K_r8_reg[24]/NET0131  ;
  assign n59172 = ~decrypt_pad & ~\u0_uk_K_r8_reg[34]/NET0131  ;
  assign n59173 = ~n59171 & ~n59172 ;
  assign n59174 = \u0_R8_reg[12]/NET0131  & ~n59173 ;
  assign n59175 = ~\u0_R8_reg[12]/NET0131  & n59173 ;
  assign n59176 = ~n59174 & ~n59175 ;
  assign n59203 = n59163 & ~n59176 ;
  assign n59204 = n59194 & n59203 ;
  assign n59205 = ~n59169 & n59204 ;
  assign n59217 = decrypt_pad & ~\u0_uk_K_r8_reg[3]/NET0131  ;
  assign n59218 = ~decrypt_pad & ~\u0_uk_K_r8_reg[13]/P0001  ;
  assign n59219 = ~n59217 & ~n59218 ;
  assign n59220 = \u0_R8_reg[16]/NET0131  & ~n59219 ;
  assign n59221 = ~\u0_R8_reg[16]/NET0131  & n59219 ;
  assign n59222 = ~n59220 & ~n59221 ;
  assign n59223 = ~n59205 & n59222 ;
  assign n59178 = decrypt_pad & ~\u0_uk_K_r8_reg[19]/NET0131  ;
  assign n59179 = ~decrypt_pad & ~\u0_uk_K_r8_reg[54]/NET0131  ;
  assign n59180 = ~n59178 & ~n59179 ;
  assign n59181 = \u0_R8_reg[14]/NET0131  & ~n59180 ;
  assign n59182 = ~\u0_R8_reg[14]/NET0131  & n59180 ;
  assign n59183 = ~n59181 & ~n59182 ;
  assign n59200 = ~n59183 & ~n59194 ;
  assign n59199 = n59169 & ~n59176 ;
  assign n59206 = ~n59169 & n59176 ;
  assign n59207 = ~n59199 & ~n59206 ;
  assign n59208 = n59200 & ~n59207 ;
  assign n59212 = n59163 & n59176 ;
  assign n59213 = n59183 & n59212 ;
  assign n59214 = n59169 & n59213 ;
  assign n59224 = ~n59208 & ~n59214 ;
  assign n59225 = n59223 & n59224 ;
  assign n59185 = ~n59163 & n59176 ;
  assign n59196 = n59169 & n59194 ;
  assign n59197 = n59185 & n59196 ;
  assign n59209 = n59169 & n59203 ;
  assign n59210 = ~n59183 & n59209 ;
  assign n59211 = ~n59197 & ~n59210 ;
  assign n59170 = ~n59163 & ~n59169 ;
  assign n59177 = n59170 & ~n59176 ;
  assign n59215 = n59177 & ~n59194 ;
  assign n59216 = n59183 & n59215 ;
  assign n59226 = n59211 & ~n59216 ;
  assign n59227 = n59225 & n59226 ;
  assign n59228 = n59177 & n59194 ;
  assign n59237 = n59196 & n59212 ;
  assign n59240 = ~n59222 & ~n59237 ;
  assign n59241 = ~n59228 & n59240 ;
  assign n59235 = n59183 & n59196 ;
  assign n59236 = ~n59176 & n59235 ;
  assign n59238 = ~n59169 & n59212 ;
  assign n59239 = ~n59183 & n59238 ;
  assign n59242 = ~n59236 & ~n59239 ;
  assign n59243 = n59241 & n59242 ;
  assign n59184 = n59177 & ~n59183 ;
  assign n59229 = ~n59163 & n59199 ;
  assign n59230 = n59183 & n59229 ;
  assign n59231 = ~n59184 & ~n59230 ;
  assign n59186 = n59183 & n59185 ;
  assign n59232 = n59163 & ~n59169 ;
  assign n59233 = ~n59186 & ~n59232 ;
  assign n59234 = ~n59194 & ~n59233 ;
  assign n59244 = n59231 & ~n59234 ;
  assign n59245 = n59243 & n59244 ;
  assign n59246 = ~n59227 & ~n59245 ;
  assign n59187 = ~n59169 & n59186 ;
  assign n59188 = ~n59184 & ~n59187 ;
  assign n59195 = ~n59188 & n59194 ;
  assign n59198 = ~n59183 & n59197 ;
  assign n59201 = n59163 & n59200 ;
  assign n59202 = n59199 & n59201 ;
  assign n59247 = ~n59198 & ~n59202 ;
  assign n59248 = ~n59195 & n59247 ;
  assign n59249 = ~n59246 & n59248 ;
  assign n59250 = ~\u0_L8_reg[20]/NET0131  & ~n59249 ;
  assign n59251 = \u0_L8_reg[20]/NET0131  & n59249 ;
  assign n59252 = ~n59250 & ~n59251 ;
  assign n59258 = n58956 & ~n58975 ;
  assign n59259 = ~n59012 & ~n59258 ;
  assign n59260 = ~n58955 & ~n59020 ;
  assign n59261 = n59259 & ~n59260 ;
  assign n59262 = n58962 & ~n59261 ;
  assign n59253 = n58968 & n59006 ;
  assign n59254 = ~n58956 & ~n58968 ;
  assign n59255 = ~n58979 & n59254 ;
  assign n59256 = ~n59253 & ~n59255 ;
  assign n59257 = ~n58962 & ~n59256 ;
  assign n59263 = n58968 & n58980 ;
  assign n59264 = ~n59257 & ~n59263 ;
  assign n59265 = ~n59262 & n59264 ;
  assign n59266 = ~n58943 & ~n59265 ;
  assign n59270 = ~n58955 & n58968 ;
  assign n59271 = n58985 & ~n59270 ;
  assign n59272 = ~n59253 & ~n59271 ;
  assign n59273 = n58962 & ~n59272 ;
  assign n59276 = n58999 & ~n59001 ;
  assign n59274 = ~n58975 & ~n59013 ;
  assign n59275 = n58962 & ~n59274 ;
  assign n59277 = ~n59255 & ~n59275 ;
  assign n59278 = ~n59276 & n59277 ;
  assign n59279 = ~n59273 & ~n59278 ;
  assign n59280 = n58943 & ~n59279 ;
  assign n59267 = n58962 & ~n58968 ;
  assign n59268 = n58955 & n58975 ;
  assign n59269 = n59267 & n59268 ;
  assign n59281 = ~n59014 & ~n59269 ;
  assign n59282 = ~n59280 & n59281 ;
  assign n59283 = ~n59266 & n59282 ;
  assign n59284 = \u0_L8_reg[29]/NET0131  & ~n59283 ;
  assign n59285 = ~\u0_L8_reg[29]/NET0131  & n59283 ;
  assign n59286 = ~n59284 & ~n59285 ;
  assign n59310 = decrypt_pad & ~\u0_uk_K_r8_reg[11]/NET0131  ;
  assign n59311 = ~decrypt_pad & ~\u0_uk_K_r8_reg[46]/NET0131  ;
  assign n59312 = ~n59310 & ~n59311 ;
  assign n59313 = \u0_R8_reg[7]/NET0131  & ~n59312 ;
  assign n59314 = ~\u0_R8_reg[7]/NET0131  & n59312 ;
  assign n59315 = ~n59313 & ~n59314 ;
  assign n59287 = decrypt_pad & ~\u0_uk_K_r8_reg[39]/NET0131  ;
  assign n59288 = ~decrypt_pad & ~\u0_uk_K_r8_reg[17]/NET0131  ;
  assign n59289 = ~n59287 & ~n59288 ;
  assign n59290 = \u0_R8_reg[9]/NET0131  & ~n59289 ;
  assign n59291 = ~\u0_R8_reg[9]/NET0131  & n59289 ;
  assign n59292 = ~n59290 & ~n59291 ;
  assign n59293 = decrypt_pad & ~\u0_uk_K_r8_reg[47]/NET0131  ;
  assign n59294 = ~decrypt_pad & ~\u0_uk_K_r8_reg[25]/NET0131  ;
  assign n59295 = ~n59293 & ~n59294 ;
  assign n59296 = \u0_R8_reg[4]/NET0131  & ~n59295 ;
  assign n59297 = ~\u0_R8_reg[4]/NET0131  & n59295 ;
  assign n59298 = ~n59296 & ~n59297 ;
  assign n59332 = n59292 & ~n59298 ;
  assign n59300 = decrypt_pad & ~\u0_uk_K_r8_reg[26]/NET0131  ;
  assign n59301 = ~decrypt_pad & ~\u0_uk_K_r8_reg[4]/NET0131  ;
  assign n59302 = ~n59300 & ~n59301 ;
  assign n59303 = \u0_R8_reg[5]/NET0131  & ~n59302 ;
  assign n59304 = ~\u0_R8_reg[5]/NET0131  & n59302 ;
  assign n59305 = ~n59303 & ~n59304 ;
  assign n59318 = decrypt_pad & ~\u0_uk_K_r8_reg[17]/NET0131  ;
  assign n59319 = ~decrypt_pad & ~\u0_uk_K_r8_reg[27]/NET0131  ;
  assign n59320 = ~n59318 & ~n59319 ;
  assign n59321 = \u0_R8_reg[6]/NET0131  & ~n59320 ;
  assign n59322 = ~\u0_R8_reg[6]/NET0131  & n59320 ;
  assign n59323 = ~n59321 & ~n59322 ;
  assign n59345 = n59305 & n59323 ;
  assign n59346 = ~n59305 & ~n59323 ;
  assign n59347 = ~n59345 & ~n59346 ;
  assign n59348 = n59332 & ~n59347 ;
  assign n59338 = decrypt_pad & ~\u0_uk_K_r8_reg[34]/NET0131  ;
  assign n59339 = ~decrypt_pad & ~\u0_uk_K_r8_reg[12]/NET0131  ;
  assign n59340 = ~n59338 & ~n59339 ;
  assign n59341 = \u0_R8_reg[8]/NET0131  & ~n59340 ;
  assign n59342 = ~\u0_R8_reg[8]/NET0131  & n59340 ;
  assign n59343 = ~n59341 & ~n59342 ;
  assign n59349 = ~n59305 & n59332 ;
  assign n59299 = ~n59292 & n59298 ;
  assign n59330 = n59298 & n59305 ;
  assign n59331 = ~n59299 & ~n59330 ;
  assign n59350 = n59323 & ~n59331 ;
  assign n59351 = ~n59349 & ~n59350 ;
  assign n59352 = ~n59343 & ~n59351 ;
  assign n59353 = ~n59348 & ~n59352 ;
  assign n59354 = ~n59315 & ~n59353 ;
  assign n59306 = n59299 & ~n59305 ;
  assign n59307 = n59292 & n59298 ;
  assign n59308 = n59305 & n59307 ;
  assign n59309 = ~n59306 & ~n59308 ;
  assign n59316 = n59305 & n59315 ;
  assign n59317 = n59309 & ~n59316 ;
  assign n59324 = ~n59317 & ~n59323 ;
  assign n59325 = ~n59305 & ~n59315 ;
  assign n59326 = ~n59298 & ~n59325 ;
  assign n59327 = ~n59292 & ~n59298 ;
  assign n59328 = ~n59316 & ~n59327 ;
  assign n59329 = ~n59326 & ~n59328 ;
  assign n59333 = ~n59315 & n59323 ;
  assign n59334 = ~n59332 & n59333 ;
  assign n59335 = n59331 & n59334 ;
  assign n59336 = ~n59329 & ~n59335 ;
  assign n59337 = ~n59324 & n59336 ;
  assign n59344 = ~n59337 & n59343 ;
  assign n59355 = ~n59292 & n59305 ;
  assign n59356 = ~n59349 & ~n59355 ;
  assign n59357 = ~n59323 & ~n59356 ;
  assign n59358 = n59292 & ~n59323 ;
  assign n59359 = n59325 & n59358 ;
  assign n59360 = n59323 & n59332 ;
  assign n59361 = n59305 & n59360 ;
  assign n59362 = ~n59359 & ~n59361 ;
  assign n59363 = ~n59357 & n59362 ;
  assign n59364 = ~n59343 & ~n59363 ;
  assign n59365 = n59307 & n59323 ;
  assign n59366 = ~n59305 & n59365 ;
  assign n59367 = ~n59343 & n59366 ;
  assign n59368 = ~n59323 & n59330 ;
  assign n59369 = ~n59305 & n59323 ;
  assign n59370 = ~n59292 & n59369 ;
  assign n59371 = ~n59298 & n59370 ;
  assign n59372 = ~n59368 & ~n59371 ;
  assign n59373 = ~n59367 & n59372 ;
  assign n59374 = n59315 & ~n59373 ;
  assign n59375 = ~n59364 & ~n59374 ;
  assign n59376 = ~n59344 & n59375 ;
  assign n59377 = ~n59354 & n59376 ;
  assign n59378 = \u0_L8_reg[2]/NET0131  & n59377 ;
  assign n59379 = ~\u0_L8_reg[2]/NET0131  & ~n59377 ;
  assign n59380 = ~n59378 & ~n59379 ;
  assign n59381 = n58955 & ~n58991 ;
  assign n59382 = ~n59006 & ~n59381 ;
  assign n59383 = n58962 & ~n59382 ;
  assign n59384 = n58975 & n59001 ;
  assign n59385 = ~n59263 & ~n59384 ;
  assign n59386 = ~n58962 & ~n59385 ;
  assign n59387 = ~n59014 & ~n59018 ;
  assign n59388 = ~n59386 & n59387 ;
  assign n59389 = ~n59383 & n59388 ;
  assign n59390 = ~n58943 & ~n59389 ;
  assign n59392 = n58975 & n59013 ;
  assign n59393 = ~n58990 & ~n59392 ;
  assign n59394 = ~n58962 & ~n59393 ;
  assign n59391 = n58998 & n59267 ;
  assign n59395 = n58975 & ~n59270 ;
  assign n59396 = ~n59002 & n59395 ;
  assign n59397 = ~n59391 & ~n59396 ;
  assign n59398 = ~n59394 & n59397 ;
  assign n59399 = n58943 & ~n59398 ;
  assign n59400 = n58968 & n59259 ;
  assign n59401 = ~n58962 & ~n59002 ;
  assign n59402 = ~n59400 & n59401 ;
  assign n59403 = n58955 & n58985 ;
  assign n59404 = ~n59010 & ~n59403 ;
  assign n59405 = ~n59006 & n59404 ;
  assign n59406 = n58962 & n58968 ;
  assign n59407 = ~n59405 & n59406 ;
  assign n59408 = ~n59402 & ~n59407 ;
  assign n59409 = ~n59399 & n59408 ;
  assign n59410 = ~n59390 & n59409 ;
  assign n59411 = ~\u0_L8_reg[4]/NET0131  & ~n59410 ;
  assign n59412 = \u0_L8_reg[4]/NET0131  & n59410 ;
  assign n59413 = ~n59411 & ~n59412 ;
  assign n59414 = decrypt_pad & ~\u0_uk_K_r8_reg[29]/NET0131  ;
  assign n59415 = ~decrypt_pad & ~\u0_uk_K_r8_reg[9]/P0001  ;
  assign n59416 = ~n59414 & ~n59415 ;
  assign n59417 = \u0_R8_reg[32]/NET0131  & ~n59416 ;
  assign n59418 = ~\u0_R8_reg[32]/NET0131  & n59416 ;
  assign n59419 = ~n59417 & ~n59418 ;
  assign n59439 = decrypt_pad & ~\u0_uk_K_r8_reg[50]/NET0131  ;
  assign n59440 = ~decrypt_pad & ~\u0_uk_K_r8_reg[30]/NET0131  ;
  assign n59441 = ~n59439 & ~n59440 ;
  assign n59442 = \u0_R8_reg[1]/NET0131  & ~n59441 ;
  assign n59443 = ~\u0_R8_reg[1]/NET0131  & n59441 ;
  assign n59444 = ~n59442 & ~n59443 ;
  assign n59420 = decrypt_pad & ~\u0_uk_K_r8_reg[35]/NET0131  ;
  assign n59421 = ~decrypt_pad & ~\u0_uk_K_r8_reg[15]/NET0131  ;
  assign n59422 = ~n59420 & ~n59421 ;
  assign n59423 = \u0_R8_reg[30]/NET0131  & ~n59422 ;
  assign n59424 = ~\u0_R8_reg[30]/NET0131  & n59422 ;
  assign n59425 = ~n59423 & ~n59424 ;
  assign n59426 = decrypt_pad & ~\u0_uk_K_r8_reg[38]/NET0131  ;
  assign n59427 = ~decrypt_pad & ~\u0_uk_K_r8_reg[14]/NET0131  ;
  assign n59428 = ~n59426 & ~n59427 ;
  assign n59429 = \u0_R8_reg[29]/NET0131  & ~n59428 ;
  assign n59430 = ~\u0_R8_reg[29]/NET0131  & n59428 ;
  assign n59431 = ~n59429 & ~n59430 ;
  assign n59432 = decrypt_pad & ~\u0_uk_K_r8_reg[7]/NET0131  ;
  assign n59433 = ~decrypt_pad & ~\u0_uk_K_r8_reg[42]/NET0131  ;
  assign n59434 = ~n59432 & ~n59433 ;
  assign n59435 = \u0_R8_reg[28]/NET0131  & ~n59434 ;
  assign n59436 = ~\u0_R8_reg[28]/NET0131  & n59434 ;
  assign n59437 = ~n59435 & ~n59436 ;
  assign n59447 = ~n59431 & n59437 ;
  assign n59448 = n59425 & n59447 ;
  assign n59449 = ~n59444 & n59448 ;
  assign n59450 = ~n59437 & n59444 ;
  assign n59451 = ~n59431 & n59450 ;
  assign n59452 = ~n59449 & ~n59451 ;
  assign n59453 = decrypt_pad & ~\u0_uk_K_r8_reg[23]/NET0131  ;
  assign n59454 = ~decrypt_pad & ~\u0_uk_K_r8_reg[31]/NET0131  ;
  assign n59455 = ~n59453 & ~n59454 ;
  assign n59456 = \u0_R8_reg[31]/P0001  & ~n59455 ;
  assign n59457 = ~\u0_R8_reg[31]/P0001  & n59455 ;
  assign n59458 = ~n59456 & ~n59457 ;
  assign n59459 = ~n59452 & n59458 ;
  assign n59464 = n59425 & ~n59437 ;
  assign n59465 = ~n59444 & ~n59464 ;
  assign n59466 = ~n59431 & n59444 ;
  assign n59467 = ~n59458 & ~n59466 ;
  assign n59468 = ~n59465 & n59467 ;
  assign n59438 = n59431 & n59437 ;
  assign n59445 = n59438 & n59444 ;
  assign n59446 = n59425 & n59445 ;
  assign n59460 = ~n59425 & n59437 ;
  assign n59461 = ~n59458 & n59460 ;
  assign n59462 = n59431 & ~n59444 ;
  assign n59463 = n59460 & n59462 ;
  assign n59469 = ~n59461 & ~n59463 ;
  assign n59470 = ~n59446 & n59469 ;
  assign n59471 = ~n59468 & n59470 ;
  assign n59472 = ~n59459 & n59471 ;
  assign n59473 = ~n59419 & ~n59472 ;
  assign n59494 = n59425 & n59451 ;
  assign n59489 = ~n59431 & ~n59444 ;
  assign n59490 = ~n59437 & n59489 ;
  assign n59491 = ~n59425 & n59490 ;
  assign n59479 = ~n59460 & ~n59462 ;
  assign n59492 = ~n59464 & ~n59466 ;
  assign n59493 = ~n59479 & ~n59492 ;
  assign n59495 = ~n59491 & ~n59493 ;
  assign n59496 = ~n59494 & n59495 ;
  assign n59497 = n59458 & ~n59496 ;
  assign n59480 = n59458 & ~n59463 ;
  assign n59481 = ~n59479 & n59480 ;
  assign n59474 = n59431 & n59450 ;
  assign n59475 = n59425 & n59474 ;
  assign n59476 = ~n59425 & ~n59431 ;
  assign n59477 = ~n59437 & n59476 ;
  assign n59478 = ~n59458 & n59477 ;
  assign n59482 = ~n59475 & ~n59478 ;
  assign n59483 = ~n59481 & n59482 ;
  assign n59484 = n59419 & ~n59483 ;
  assign n59485 = ~n59458 & n59463 ;
  assign n59486 = n59425 & ~n59458 ;
  assign n59487 = n59419 & n59447 ;
  assign n59488 = n59486 & n59487 ;
  assign n59498 = ~n59485 & ~n59488 ;
  assign n59499 = ~n59484 & n59498 ;
  assign n59500 = ~n59497 & n59499 ;
  assign n59501 = ~n59473 & n59500 ;
  assign n59502 = \u0_L8_reg[5]/NET0131  & ~n59501 ;
  assign n59503 = ~\u0_L8_reg[5]/NET0131  & n59501 ;
  assign n59504 = ~n59502 & ~n59503 ;
  assign n59505 = n59299 & n59345 ;
  assign n59506 = n59292 & n59368 ;
  assign n59507 = ~n59505 & ~n59506 ;
  assign n59509 = ~n59305 & n59360 ;
  assign n59508 = n59305 & n59327 ;
  assign n59510 = n59299 & n59346 ;
  assign n59511 = ~n59508 & ~n59510 ;
  assign n59512 = ~n59509 & n59511 ;
  assign n59513 = ~n59343 & ~n59512 ;
  assign n59514 = n59507 & ~n59513 ;
  assign n59515 = ~n59315 & ~n59514 ;
  assign n59516 = ~n59299 & ~n59305 ;
  assign n59517 = ~n59332 & n59516 ;
  assign n59518 = n59299 & ~n59323 ;
  assign n59519 = n59305 & n59518 ;
  assign n59520 = ~n59517 & ~n59519 ;
  assign n59521 = n59315 & ~n59520 ;
  assign n59525 = n59326 & n59358 ;
  assign n59522 = n59298 & n59315 ;
  assign n59523 = n59323 & ~n59355 ;
  assign n59524 = n59522 & n59523 ;
  assign n59526 = ~n59343 & ~n59524 ;
  assign n59527 = ~n59525 & n59526 ;
  assign n59528 = ~n59521 & n59527 ;
  assign n59529 = ~n59292 & n59346 ;
  assign n59530 = n59315 & ~n59360 ;
  assign n59531 = ~n59529 & n59530 ;
  assign n59532 = ~n59305 & n59307 ;
  assign n59533 = ~n59315 & ~n59370 ;
  assign n59534 = ~n59532 & n59533 ;
  assign n59535 = ~n59531 & ~n59534 ;
  assign n59536 = ~n59323 & n59327 ;
  assign n59537 = n59305 & n59536 ;
  assign n59538 = n59343 & ~n59537 ;
  assign n59539 = n59362 & n59538 ;
  assign n59540 = n59507 & n59539 ;
  assign n59541 = ~n59535 & n59540 ;
  assign n59542 = ~n59528 & ~n59541 ;
  assign n59543 = ~n59515 & ~n59542 ;
  assign n59544 = ~\u0_L8_reg[13]/NET0131  & n59543 ;
  assign n59545 = \u0_L8_reg[13]/NET0131  & ~n59543 ;
  assign n59546 = ~n59544 & ~n59545 ;
  assign n59567 = decrypt_pad & ~\u0_uk_K_r8_reg[43]/NET0131  ;
  assign n59568 = ~decrypt_pad & ~\u0_uk_K_r8_reg[23]/NET0131  ;
  assign n59569 = ~n59567 & ~n59568 ;
  assign n59570 = \u0_R8_reg[18]/NET0131  & ~n59569 ;
  assign n59571 = ~\u0_R8_reg[18]/NET0131  & n59569 ;
  assign n59572 = ~n59570 & ~n59571 ;
  assign n59574 = decrypt_pad & ~\u0_uk_K_r8_reg[30]/NET0131  ;
  assign n59575 = ~decrypt_pad & ~\u0_uk_K_r8_reg[38]/NET0131  ;
  assign n59576 = ~n59574 & ~n59575 ;
  assign n59577 = \u0_R8_reg[19]/NET0131  & ~n59576 ;
  assign n59578 = ~\u0_R8_reg[19]/NET0131  & n59576 ;
  assign n59579 = ~n59577 & ~n59578 ;
  assign n59580 = ~n59572 & ~n59579 ;
  assign n59553 = decrypt_pad & ~\u0_uk_K_r8_reg[49]/NET0131  ;
  assign n59554 = ~decrypt_pad & ~\u0_uk_K_r8_reg[29]/NET0131  ;
  assign n59555 = ~n59553 & ~n59554 ;
  assign n59556 = \u0_R8_reg[17]/NET0131  & ~n59555 ;
  assign n59557 = ~\u0_R8_reg[17]/NET0131  & n59555 ;
  assign n59558 = ~n59556 & ~n59557 ;
  assign n59547 = decrypt_pad & ~\u0_uk_K_r8_reg[15]/NET0131  ;
  assign n59548 = ~decrypt_pad & ~\u0_uk_K_r8_reg[50]/NET0131  ;
  assign n59549 = ~n59547 & ~n59548 ;
  assign n59550 = \u0_R8_reg[21]/NET0131  & ~n59549 ;
  assign n59551 = ~\u0_R8_reg[21]/NET0131  & n59549 ;
  assign n59552 = ~n59550 & ~n59551 ;
  assign n59560 = decrypt_pad & ~\u0_uk_K_r8_reg[31]/NET0131  ;
  assign n59561 = ~decrypt_pad & ~\u0_uk_K_r8_reg[7]/NET0131  ;
  assign n59562 = ~n59560 & ~n59561 ;
  assign n59563 = \u0_R8_reg[16]/NET0131  & ~n59562 ;
  assign n59564 = ~\u0_R8_reg[16]/NET0131  & n59562 ;
  assign n59565 = ~n59563 & ~n59564 ;
  assign n59581 = n59552 & ~n59565 ;
  assign n59582 = n59558 & n59581 ;
  assign n59583 = ~n59552 & ~n59565 ;
  assign n59584 = ~n59558 & n59583 ;
  assign n59585 = ~n59582 & ~n59584 ;
  assign n59586 = n59580 & ~n59585 ;
  assign n59559 = ~n59552 & n59558 ;
  assign n59566 = n59559 & n59565 ;
  assign n59573 = n59566 & ~n59572 ;
  assign n59607 = n59572 & ~n59579 ;
  assign n59608 = n59558 & ~n59607 ;
  assign n59606 = n59552 & n59565 ;
  assign n59609 = ~n59558 & n59572 ;
  assign n59610 = n59606 & ~n59609 ;
  assign n59611 = ~n59608 & n59610 ;
  assign n59612 = ~n59573 & ~n59611 ;
  assign n59613 = ~n59586 & n59612 ;
  assign n59587 = n59558 & ~n59572 ;
  assign n59588 = ~n59565 & n59587 ;
  assign n59589 = n59552 & n59572 ;
  assign n59590 = n59565 & n59589 ;
  assign n59591 = ~n59588 & ~n59590 ;
  assign n59592 = ~n59552 & ~n59558 ;
  assign n59593 = n59579 & ~n59583 ;
  assign n59594 = ~n59592 & n59593 ;
  assign n59595 = n59591 & n59594 ;
  assign n59596 = ~n59558 & n59565 ;
  assign n59597 = ~n59552 & n59596 ;
  assign n59598 = n59572 & n59597 ;
  assign n59599 = decrypt_pad & ~\u0_uk_K_r8_reg[14]/NET0131  ;
  assign n59600 = ~decrypt_pad & ~\u0_uk_K_r8_reg[49]/NET0131  ;
  assign n59601 = ~n59599 & ~n59600 ;
  assign n59602 = \u0_R8_reg[20]/NET0131  & ~n59601 ;
  assign n59603 = ~\u0_R8_reg[20]/NET0131  & n59601 ;
  assign n59604 = ~n59602 & ~n59603 ;
  assign n59605 = ~n59598 & n59604 ;
  assign n59614 = ~n59595 & n59605 ;
  assign n59615 = n59613 & n59614 ;
  assign n59622 = ~n59558 & ~n59565 ;
  assign n59623 = n59552 & n59622 ;
  assign n59620 = n59558 & n59572 ;
  assign n59621 = ~n59552 & n59620 ;
  assign n59624 = ~n59579 & ~n59621 ;
  assign n59625 = ~n59623 & n59624 ;
  assign n59617 = n59558 & n59606 ;
  assign n59618 = ~n59572 & n59617 ;
  assign n59619 = ~n59572 & n59597 ;
  assign n59626 = ~n59618 & ~n59619 ;
  assign n59627 = n59625 & n59626 ;
  assign n59628 = n59579 & ~n59584 ;
  assign n59629 = n59591 & n59628 ;
  assign n59630 = ~n59627 & ~n59629 ;
  assign n59631 = ~n59552 & n59588 ;
  assign n59616 = n59589 & n59596 ;
  assign n59632 = ~n59604 & ~n59616 ;
  assign n59633 = ~n59631 & n59632 ;
  assign n59634 = ~n59630 & n59633 ;
  assign n59635 = ~n59615 & ~n59634 ;
  assign n59636 = n59572 & n59583 ;
  assign n59637 = ~n59558 & n59636 ;
  assign n59638 = ~n59573 & ~n59637 ;
  assign n59639 = n59579 & ~n59638 ;
  assign n59640 = n59589 & n59622 ;
  assign n59641 = n59583 & n59620 ;
  assign n59642 = ~n59640 & ~n59641 ;
  assign n59643 = ~n59579 & ~n59642 ;
  assign n59644 = ~n59639 & ~n59643 ;
  assign n59645 = ~n59635 & n59644 ;
  assign n59646 = ~\u0_L8_reg[14]/NET0131  & ~n59645 ;
  assign n59647 = \u0_L8_reg[14]/NET0131  & n59645 ;
  assign n59648 = ~n59646 & ~n59647 ;
  assign n59670 = ~n59176 & ~n59183 ;
  assign n59671 = ~n59163 & n59670 ;
  assign n59672 = ~n59187 & ~n59671 ;
  assign n59673 = n59194 & ~n59672 ;
  assign n59674 = ~n59183 & n59185 ;
  assign n59675 = ~n59238 & ~n59674 ;
  assign n59676 = ~n59194 & ~n59675 ;
  assign n59661 = n59169 & ~n59183 ;
  assign n59668 = ~n59185 & ~n59203 ;
  assign n59669 = n59661 & ~n59668 ;
  assign n59677 = ~n59214 & ~n59669 ;
  assign n59678 = ~n59676 & n59677 ;
  assign n59679 = ~n59673 & n59678 ;
  assign n59680 = ~n59222 & ~n59679 ;
  assign n59662 = ~n59185 & n59661 ;
  assign n59663 = ~n59209 & ~n59662 ;
  assign n59664 = ~n59194 & ~n59663 ;
  assign n59649 = ~n59169 & n59183 ;
  assign n59650 = ~n59176 & n59649 ;
  assign n59659 = n59169 & n59186 ;
  assign n59665 = ~n59650 & ~n59659 ;
  assign n59666 = ~n59664 & n59665 ;
  assign n59667 = n59222 & ~n59666 ;
  assign n59651 = n59163 & n59650 ;
  assign n59652 = ~n59214 & ~n59651 ;
  assign n59653 = ~n59230 & n59652 ;
  assign n59654 = n59194 & ~n59653 ;
  assign n59660 = ~n59194 & n59659 ;
  assign n59655 = ~n59183 & n59206 ;
  assign n59656 = ~n59232 & ~n59655 ;
  assign n59657 = n59194 & n59222 ;
  assign n59658 = ~n59656 & n59657 ;
  assign n59681 = ~n59216 & ~n59658 ;
  assign n59682 = ~n59660 & n59681 ;
  assign n59683 = ~n59654 & n59682 ;
  assign n59684 = ~n59667 & n59683 ;
  assign n59685 = ~n59680 & n59684 ;
  assign n59686 = ~\u0_L8_reg[1]/NET0131  & ~n59685 ;
  assign n59687 = \u0_L8_reg[1]/NET0131  & n59685 ;
  assign n59688 = ~n59686 & ~n59687 ;
  assign n59701 = n59185 & ~n59661 ;
  assign n59702 = ~n59210 & ~n59701 ;
  assign n59703 = ~n59194 & ~n59702 ;
  assign n59699 = ~n59229 & ~n59239 ;
  assign n59700 = n59194 & ~n59699 ;
  assign n59704 = n59652 & ~n59700 ;
  assign n59705 = ~n59703 & n59704 ;
  assign n59706 = n59222 & ~n59705 ;
  assign n59690 = ~n59170 & ~n59649 ;
  assign n59691 = n59194 & ~n59690 ;
  assign n59692 = ~n59201 & ~n59661 ;
  assign n59693 = ~n59691 & n59692 ;
  assign n59694 = n59176 & ~n59693 ;
  assign n59689 = ~n59183 & n59204 ;
  assign n59695 = ~n59215 & ~n59689 ;
  assign n59696 = n59231 & n59695 ;
  assign n59697 = ~n59694 & n59696 ;
  assign n59698 = ~n59222 & ~n59697 ;
  assign n59707 = ~n59184 & n59652 ;
  assign n59708 = ~n59194 & ~n59707 ;
  assign n59709 = ~n59198 & ~n59236 ;
  assign n59710 = ~n59708 & n59709 ;
  assign n59711 = ~n59698 & n59710 ;
  assign n59712 = ~n59706 & n59711 ;
  assign n59713 = ~\u0_L8_reg[10]/NET0131  & ~n59712 ;
  assign n59714 = \u0_L8_reg[10]/NET0131  & n59712 ;
  assign n59715 = ~n59713 & ~n59714 ;
  assign n59716 = n59054 & ~n59095 ;
  assign n59717 = ~n59096 & n59716 ;
  assign n59718 = ~n59107 & n59717 ;
  assign n59720 = n59078 & n59081 ;
  assign n59721 = ~n59054 & n59720 ;
  assign n59719 = ~n59104 & n59107 ;
  assign n59722 = n59068 & ~n59719 ;
  assign n59723 = ~n59721 & n59722 ;
  assign n59724 = ~n59718 & n59723 ;
  assign n59727 = ~n59039 & n59074 ;
  assign n59731 = n59039 & ~n59074 ;
  assign n59733 = ~n59727 & ~n59731 ;
  assign n59734 = ~n59106 & n59111 ;
  assign n59735 = n59733 & n59734 ;
  assign n59725 = ~n59047 & ~n59097 ;
  assign n59726 = ~n59054 & ~n59725 ;
  assign n59728 = n59054 & ~n59060 ;
  assign n59729 = ~n59110 & ~n59728 ;
  assign n59730 = n59727 & ~n59729 ;
  assign n59732 = n59088 & n59731 ;
  assign n59736 = ~n59068 & ~n59732 ;
  assign n59737 = ~n59730 & n59736 ;
  assign n59738 = ~n59726 & n59737 ;
  assign n59739 = ~n59735 & n59738 ;
  assign n59740 = ~n59724 & ~n59739 ;
  assign n59741 = \u0_L8_reg[12]/NET0131  & n59740 ;
  assign n59742 = ~\u0_L8_reg[12]/NET0131  & ~n59740 ;
  assign n59743 = ~n59741 & ~n59742 ;
  assign n59744 = n59458 & n59477 ;
  assign n59745 = ~n59419 & ~n59744 ;
  assign n59752 = ~n59474 & ~n59477 ;
  assign n59751 = n59425 & n59438 ;
  assign n59750 = n59444 & n59476 ;
  assign n59753 = n59458 & ~n59750 ;
  assign n59754 = ~n59751 & n59753 ;
  assign n59755 = n59752 & n59754 ;
  assign n59757 = n59444 & n59448 ;
  assign n59756 = ~n59444 & n59460 ;
  assign n59758 = ~n59458 & ~n59756 ;
  assign n59759 = ~n59757 & n59758 ;
  assign n59760 = ~n59755 & ~n59759 ;
  assign n59746 = n59450 & n59476 ;
  assign n59747 = n59437 & n59462 ;
  assign n59748 = ~n59490 & ~n59747 ;
  assign n59749 = n59425 & ~n59748 ;
  assign n59761 = ~n59746 & ~n59749 ;
  assign n59762 = ~n59760 & n59761 ;
  assign n59763 = ~n59745 & ~n59762 ;
  assign n59764 = n59444 & n59461 ;
  assign n59765 = n59431 & n59764 ;
  assign n59778 = ~n59449 & ~n59491 ;
  assign n59779 = ~n59764 & n59778 ;
  assign n59769 = ~n59448 & ~n59747 ;
  assign n59770 = n59458 & ~n59769 ;
  assign n59766 = n59437 & n59444 ;
  assign n59767 = ~n59425 & n59431 ;
  assign n59768 = n59766 & n59767 ;
  assign n59771 = n59431 & n59464 ;
  assign n59775 = ~n59768 & ~n59771 ;
  assign n59772 = n59450 & n59486 ;
  assign n59773 = ~n59437 & ~n59458 ;
  assign n59774 = n59462 & n59773 ;
  assign n59776 = ~n59772 & ~n59774 ;
  assign n59777 = n59775 & n59776 ;
  assign n59780 = ~n59770 & n59777 ;
  assign n59781 = n59779 & n59780 ;
  assign n59782 = ~n59419 & ~n59781 ;
  assign n59783 = ~n59765 & ~n59782 ;
  assign n59784 = ~n59763 & n59783 ;
  assign n59785 = ~\u0_L8_reg[21]/NET0131  & ~n59784 ;
  assign n59786 = \u0_L8_reg[21]/NET0131  & n59784 ;
  assign n59787 = ~n59785 & ~n59786 ;
  assign n59788 = ~n59444 & n59767 ;
  assign n59789 = ~n59438 & ~n59451 ;
  assign n59790 = ~n59788 & n59789 ;
  assign n59791 = n59458 & ~n59790 ;
  assign n59792 = n59460 & n59489 ;
  assign n59793 = ~n59791 & ~n59792 ;
  assign n59794 = ~n59419 & ~n59793 ;
  assign n59798 = n59466 & n59486 ;
  assign n59795 = n59431 & n59460 ;
  assign n59797 = n59462 & n59464 ;
  assign n59799 = ~n59795 & ~n59797 ;
  assign n59800 = ~n59798 & n59799 ;
  assign n59796 = n59458 & n59490 ;
  assign n59801 = ~n59757 & ~n59796 ;
  assign n59802 = n59800 & n59801 ;
  assign n59803 = n59419 & ~n59802 ;
  assign n59805 = ~n59419 & n59447 ;
  assign n59804 = n59450 & n59767 ;
  assign n59807 = ~n59797 & ~n59804 ;
  assign n59808 = ~n59805 & n59807 ;
  assign n59806 = ~n59448 & ~n59458 ;
  assign n59809 = ~n59491 & n59806 ;
  assign n59810 = n59808 & n59809 ;
  assign n59811 = n59458 & ~n59746 ;
  assign n59812 = ~n59475 & n59811 ;
  assign n59813 = ~n59810 & ~n59812 ;
  assign n59814 = ~n59803 & ~n59813 ;
  assign n59815 = ~n59794 & n59814 ;
  assign n59816 = \u0_L8_reg[15]/P0001  & n59815 ;
  assign n59817 = ~\u0_L8_reg[15]/P0001  & ~n59815 ;
  assign n59818 = ~n59816 & ~n59817 ;
  assign n59831 = n58949 & ~n58976 ;
  assign n59832 = ~n59384 & ~n59831 ;
  assign n59833 = n58962 & ~n59832 ;
  assign n59829 = n58968 & n59012 ;
  assign n59830 = ~n58962 & ~n59404 ;
  assign n59834 = ~n59829 & ~n59830 ;
  assign n59835 = ~n59833 & n59834 ;
  assign n59836 = ~n58943 & ~n59835 ;
  assign n59822 = ~n58980 & ~n58987 ;
  assign n59823 = n58962 & ~n59822 ;
  assign n59819 = n58968 & ~n59404 ;
  assign n59820 = ~n58968 & n58980 ;
  assign n59821 = ~n58962 & n58982 ;
  assign n59824 = ~n59392 & ~n59821 ;
  assign n59825 = ~n59820 & n59824 ;
  assign n59826 = ~n59819 & n59825 ;
  assign n59827 = ~n59823 & n59826 ;
  assign n59828 = n58943 & ~n59827 ;
  assign n59837 = ~n59009 & ~n59019 ;
  assign n59838 = ~n59828 & n59837 ;
  assign n59839 = ~n59836 & n59838 ;
  assign n59840 = ~\u0_L8_reg[19]/NET0131  & ~n59839 ;
  assign n59841 = \u0_L8_reg[19]/NET0131  & n59839 ;
  assign n59842 = ~n59840 & ~n59841 ;
  assign n59843 = n58885 & n58886 ;
  assign n59844 = ~n59125 & ~n59843 ;
  assign n59845 = ~n58854 & ~n59844 ;
  assign n59846 = n58854 & ~n58905 ;
  assign n59847 = ~n58882 & n59846 ;
  assign n59848 = ~n58923 & ~n59847 ;
  assign n59849 = ~n59845 & n59848 ;
  assign n59850 = ~n58861 & ~n59849 ;
  assign n59851 = n58883 & ~n59124 ;
  assign n59852 = n58854 & ~n59851 ;
  assign n59853 = ~n58867 & ~n59142 ;
  assign n59854 = ~n58854 & ~n58890 ;
  assign n59855 = ~n59853 & n59854 ;
  assign n59856 = ~n59852 & ~n59855 ;
  assign n59857 = n58848 & ~n59127 ;
  assign n59858 = ~n58930 & n59857 ;
  assign n59859 = ~n59856 & n59858 ;
  assign n59864 = ~n58848 & ~n58904 ;
  assign n59865 = ~n58922 & n59864 ;
  assign n59860 = ~n58888 & n58902 ;
  assign n59861 = ~n58918 & n59860 ;
  assign n59862 = n58854 & ~n58867 ;
  assign n59863 = ~n58924 & n59862 ;
  assign n59866 = ~n59861 & ~n59863 ;
  assign n59867 = n59865 & n59866 ;
  assign n59868 = ~n59859 & ~n59867 ;
  assign n59869 = ~n59850 & ~n59868 ;
  assign n59870 = \u0_L8_reg[23]/NET0131  & ~n59869 ;
  assign n59871 = ~\u0_L8_reg[23]/NET0131  & n59869 ;
  assign n59872 = ~n59870 & ~n59871 ;
  assign n59876 = ~n59170 & ~n59650 ;
  assign n59877 = ~n59222 & ~n59876 ;
  assign n59873 = n59169 & ~n59668 ;
  assign n59874 = ~n59661 & ~n59674 ;
  assign n59875 = ~n59873 & ~n59874 ;
  assign n59878 = ~n59194 & ~n59875 ;
  assign n59879 = ~n59877 & n59878 ;
  assign n59880 = n59194 & ~n59210 ;
  assign n59881 = ~n59239 & n59880 ;
  assign n59882 = ~n59879 & ~n59881 ;
  assign n59883 = ~n59186 & ~n59671 ;
  assign n59884 = n59169 & ~n59883 ;
  assign n59890 = n59222 & ~n59228 ;
  assign n59891 = ~n59884 & n59890 ;
  assign n59885 = n59232 & n59670 ;
  assign n59886 = ~n59213 & ~n59885 ;
  assign n59887 = ~n59194 & ~n59886 ;
  assign n59888 = ~n59204 & ~n59209 ;
  assign n59889 = n59183 & ~n59888 ;
  assign n59892 = ~n59887 & ~n59889 ;
  assign n59893 = n59891 & n59892 ;
  assign n59894 = ~n59203 & n59235 ;
  assign n59895 = ~n59222 & ~n59655 ;
  assign n59896 = ~n59894 & n59895 ;
  assign n59897 = n59211 & n59896 ;
  assign n59898 = ~n59893 & ~n59897 ;
  assign n59899 = ~n59882 & ~n59898 ;
  assign n59900 = ~\u0_L8_reg[26]/NET0131  & ~n59899 ;
  assign n59901 = \u0_L8_reg[26]/NET0131  & n59899 ;
  assign n59902 = ~n59900 & ~n59901 ;
  assign n59920 = n59327 & n59345 ;
  assign n59921 = n59309 & ~n59920 ;
  assign n59922 = n59315 & ~n59921 ;
  assign n59904 = n59305 & n59332 ;
  assign n59905 = ~n59536 & ~n59904 ;
  assign n59919 = ~n59315 & ~n59905 ;
  assign n59917 = ~n59522 & ~n59532 ;
  assign n59918 = ~n59323 & ~n59917 ;
  assign n59923 = ~n59509 & ~n59918 ;
  assign n59924 = ~n59919 & n59923 ;
  assign n59925 = ~n59922 & n59924 ;
  assign n59926 = n59343 & ~n59925 ;
  assign n59907 = ~n59330 & ~n59349 ;
  assign n59908 = ~n59518 & n59907 ;
  assign n59909 = ~n59315 & ~n59908 ;
  assign n59906 = n59315 & ~n59905 ;
  assign n59903 = n59323 & n59517 ;
  assign n59910 = ~n59505 & ~n59903 ;
  assign n59911 = ~n59906 & n59910 ;
  assign n59912 = ~n59909 & n59911 ;
  assign n59913 = ~n59343 & ~n59912 ;
  assign n59914 = ~n59298 & n59369 ;
  assign n59915 = ~n59505 & ~n59914 ;
  assign n59916 = ~n59315 & ~n59915 ;
  assign n59927 = ~n59913 & ~n59916 ;
  assign n59928 = ~n59926 & n59927 ;
  assign n59929 = ~\u0_L8_reg[28]/NET0131  & ~n59928 ;
  assign n59930 = \u0_L8_reg[28]/NET0131  & n59928 ;
  assign n59931 = ~n59929 & ~n59930 ;
  assign n59932 = ~n59617 & ~n59619 ;
  assign n59933 = n59579 & ~n59932 ;
  assign n59938 = n59566 & n59572 ;
  assign n59939 = ~n59637 & ~n59938 ;
  assign n59934 = n59581 & ~n59609 ;
  assign n59935 = ~n59558 & n59606 ;
  assign n59936 = ~n59934 & ~n59935 ;
  assign n59937 = ~n59579 & ~n59936 ;
  assign n59940 = ~n59588 & ~n59937 ;
  assign n59941 = n59939 & n59940 ;
  assign n59942 = ~n59933 & n59941 ;
  assign n59943 = ~n59604 & ~n59942 ;
  assign n59944 = ~n59572 & n59592 ;
  assign n59945 = ~n59565 & n59944 ;
  assign n59946 = ~n59935 & ~n59945 ;
  assign n59947 = n59579 & ~n59946 ;
  assign n59948 = n59565 & n59580 ;
  assign n59949 = n59642 & ~n59948 ;
  assign n59950 = ~n59947 & n59949 ;
  assign n59951 = n59604 & ~n59950 ;
  assign n59952 = ~n59579 & n59598 ;
  assign n59953 = ~n59587 & ~n59609 ;
  assign n59954 = n59581 & ~n59953 ;
  assign n59955 = ~n59621 & ~n59954 ;
  assign n59956 = n59579 & ~n59955 ;
  assign n59957 = ~n59952 & ~n59956 ;
  assign n59958 = ~n59951 & n59957 ;
  assign n59959 = ~n59943 & n59958 ;
  assign n59960 = ~\u0_L8_reg[8]/NET0131  & ~n59959 ;
  assign n59961 = \u0_L8_reg[8]/NET0131  & n59959 ;
  assign n59962 = ~n59960 & ~n59961 ;
  assign n59978 = ~n59747 & n59752 ;
  assign n59979 = ~n59458 & ~n59978 ;
  assign n59975 = ~n59437 & n59788 ;
  assign n59976 = ~n59445 & ~n59975 ;
  assign n59977 = n59458 & ~n59976 ;
  assign n59980 = ~n59449 & ~n59750 ;
  assign n59981 = ~n59475 & n59980 ;
  assign n59982 = ~n59977 & n59981 ;
  assign n59983 = ~n59979 & n59982 ;
  assign n59984 = n59419 & ~n59983 ;
  assign n59965 = n59458 & ~n59771 ;
  assign n59964 = n59444 & ~n59767 ;
  assign n59966 = ~n59788 & ~n59964 ;
  assign n59967 = n59965 & n59966 ;
  assign n59963 = n59486 & n59766 ;
  assign n59968 = ~n59774 & ~n59963 ;
  assign n59969 = ~n59494 & n59968 ;
  assign n59970 = ~n59967 & n59969 ;
  assign n59971 = ~n59419 & ~n59970 ;
  assign n59974 = ~n59458 & n59493 ;
  assign n59972 = n59425 & n59458 ;
  assign n59973 = n59489 & n59972 ;
  assign n59985 = ~n59485 & ~n59973 ;
  assign n59986 = ~n59974 & n59985 ;
  assign n59987 = ~n59971 & n59986 ;
  assign n59988 = ~n59984 & n59987 ;
  assign n59989 = ~\u0_L8_reg[27]/NET0131  & ~n59988 ;
  assign n59990 = \u0_L8_reg[27]/NET0131  & n59988 ;
  assign n59991 = ~n59989 & ~n59990 ;
  assign n59993 = n59088 & ~n59733 ;
  assign n59995 = ~n59039 & n59077 ;
  assign n59994 = n59047 & n59096 ;
  assign n59996 = ~n59054 & ~n59994 ;
  assign n59997 = ~n59995 & n59996 ;
  assign n59998 = ~n59993 & n59997 ;
  assign n59999 = ~n59045 & n59731 ;
  assign n60000 = ~n59078 & ~n59999 ;
  assign n60001 = ~n59725 & n60000 ;
  assign n60002 = n59054 & ~n59720 ;
  assign n60003 = ~n60001 & n60002 ;
  assign n60004 = ~n59998 & ~n60003 ;
  assign n59992 = n59110 & n59731 ;
  assign n60005 = n59068 & ~n59992 ;
  assign n60006 = ~n60004 & n60005 ;
  assign n60010 = n59104 & n59106 ;
  assign n60013 = ~n59068 & ~n59098 ;
  assign n60014 = ~n60010 & n60013 ;
  assign n60007 = n59039 & n59096 ;
  assign n60008 = ~n59999 & ~n60007 ;
  assign n60009 = n59054 & ~n60008 ;
  assign n60011 = ~n59054 & n59097 ;
  assign n60012 = ~n59999 & n60011 ;
  assign n60015 = ~n60009 & ~n60012 ;
  assign n60016 = n60014 & n60015 ;
  assign n60017 = ~n60006 & ~n60016 ;
  assign n60018 = n59061 & ~n59731 ;
  assign n60019 = n59048 & n60018 ;
  assign n60020 = ~n60017 & ~n60019 ;
  assign n60021 = \u0_L8_reg[32]/NET0131  & n60020 ;
  assign n60022 = ~\u0_L8_reg[32]/NET0131  & ~n60020 ;
  assign n60023 = ~n60021 & ~n60022 ;
  assign n60027 = n59579 & ~n59609 ;
  assign n60028 = ~n59583 & ~n59589 ;
  assign n60029 = ~n59935 & n60028 ;
  assign n60030 = ~n60027 & ~n60029 ;
  assign n60024 = ~n59572 & n59581 ;
  assign n60025 = ~n59566 & ~n60024 ;
  assign n60026 = n59579 & ~n60025 ;
  assign n60031 = ~n59604 & ~n60026 ;
  assign n60032 = ~n60030 & n60031 ;
  assign n60033 = ~n59572 & n59606 ;
  assign n60034 = n59559 & ~n59565 ;
  assign n60035 = ~n60033 & ~n60034 ;
  assign n60036 = n59579 & ~n60035 ;
  assign n60037 = ~n59579 & n59582 ;
  assign n60038 = ~n59618 & ~n60037 ;
  assign n60039 = n59605 & n60038 ;
  assign n60040 = ~n60036 & n60039 ;
  assign n60041 = ~n60032 & ~n60040 ;
  assign n60042 = ~n59579 & ~n59616 ;
  assign n60043 = ~n59573 & n60042 ;
  assign n60044 = ~n59945 & n60043 ;
  assign n60045 = n59579 & ~n59640 ;
  assign n60046 = ~n59619 & n60045 ;
  assign n60047 = ~n60044 & ~n60046 ;
  assign n60048 = ~n60041 & ~n60047 ;
  assign n60049 = ~\u0_L8_reg[3]/NET0131  & ~n60048 ;
  assign n60050 = \u0_L8_reg[3]/NET0131  & n60048 ;
  assign n60051 = ~n60049 & ~n60050 ;
  assign n60058 = decrypt_pad & ~\u0_uk_K_r8_reg[54]/NET0131  ;
  assign n60059 = ~decrypt_pad & ~\u0_uk_K_r8_reg[32]/NET0131  ;
  assign n60060 = ~n60058 & ~n60059 ;
  assign n60061 = \u0_R8_reg[11]/NET0131  & ~n60060 ;
  assign n60062 = ~\u0_R8_reg[11]/NET0131  & n60060 ;
  assign n60063 = ~n60061 & ~n60062 ;
  assign n60052 = decrypt_pad & ~\u0_uk_K_r8_reg[12]/NET0131  ;
  assign n60053 = ~decrypt_pad & ~\u0_uk_K_r8_reg[47]/NET0131  ;
  assign n60054 = ~n60052 & ~n60053 ;
  assign n60055 = \u0_R8_reg[12]/NET0131  & ~n60054 ;
  assign n60056 = ~\u0_R8_reg[12]/NET0131  & n60054 ;
  assign n60057 = ~n60055 & ~n60056 ;
  assign n60064 = decrypt_pad & ~\u0_uk_K_r8_reg[25]/NET0131  ;
  assign n60065 = ~decrypt_pad & ~\u0_uk_K_r8_reg[3]/NET0131  ;
  assign n60066 = ~n60064 & ~n60065 ;
  assign n60067 = \u0_R8_reg[13]/NET0131  & ~n60066 ;
  assign n60068 = ~\u0_R8_reg[13]/NET0131  & n60066 ;
  assign n60069 = ~n60067 & ~n60068 ;
  assign n60077 = decrypt_pad & ~\u0_uk_K_r8_reg[20]/NET0131  ;
  assign n60078 = ~decrypt_pad & ~\u0_uk_K_r8_reg[55]/NET0131  ;
  assign n60079 = ~n60077 & ~n60078 ;
  assign n60080 = \u0_R8_reg[9]/NET0131  & ~n60079 ;
  assign n60081 = ~\u0_R8_reg[9]/NET0131  & n60079 ;
  assign n60082 = ~n60080 & ~n60081 ;
  assign n60122 = n60069 & ~n60082 ;
  assign n60070 = decrypt_pad & ~\u0_uk_K_r8_reg[48]/NET0131  ;
  assign n60071 = ~decrypt_pad & ~\u0_uk_K_r8_reg[26]/NET0131  ;
  assign n60072 = ~n60070 & ~n60071 ;
  assign n60073 = \u0_R8_reg[8]/NET0131  & ~n60072 ;
  assign n60074 = ~\u0_R8_reg[8]/NET0131  & n60072 ;
  assign n60075 = ~n60073 & ~n60074 ;
  assign n60102 = ~n60069 & n60082 ;
  assign n60103 = n60075 & n60102 ;
  assign n60076 = n60069 & ~n60075 ;
  assign n60084 = decrypt_pad & ~\u0_uk_K_r8_reg[53]/NET0131  ;
  assign n60085 = ~decrypt_pad & ~\u0_uk_K_r8_reg[6]/NET0131  ;
  assign n60086 = ~n60084 & ~n60085 ;
  assign n60087 = \u0_R8_reg[10]/NET0131  & ~n60086 ;
  assign n60088 = ~\u0_R8_reg[10]/NET0131  & n60086 ;
  assign n60089 = ~n60087 & ~n60088 ;
  assign n60124 = n60076 & n60089 ;
  assign n60125 = ~n60103 & ~n60124 ;
  assign n60126 = ~n60122 & n60125 ;
  assign n60127 = n60057 & ~n60126 ;
  assign n60123 = n60089 & n60122 ;
  assign n60094 = ~n60069 & ~n60075 ;
  assign n60128 = ~n60089 & n60094 ;
  assign n60129 = ~n60082 & n60128 ;
  assign n60130 = ~n60123 & ~n60129 ;
  assign n60131 = ~n60127 & n60130 ;
  assign n60132 = n60063 & ~n60131 ;
  assign n60095 = n60069 & n60075 ;
  assign n60096 = ~n60094 & ~n60095 ;
  assign n60093 = ~n60082 & ~n60089 ;
  assign n60099 = n60063 & ~n60075 ;
  assign n60105 = n60093 & ~n60099 ;
  assign n60106 = n60096 & n60105 ;
  assign n60100 = n60082 & ~n60089 ;
  assign n60101 = n60099 & n60100 ;
  assign n60104 = n60089 & n60103 ;
  assign n60107 = ~n60101 & ~n60104 ;
  assign n60108 = ~n60106 & n60107 ;
  assign n60083 = n60076 & n60082 ;
  assign n60090 = n60083 & n60089 ;
  assign n60091 = ~n60063 & n60090 ;
  assign n60092 = n60082 & n60089 ;
  assign n60097 = ~n60093 & ~n60096 ;
  assign n60098 = ~n60092 & n60097 ;
  assign n60109 = ~n60091 & ~n60098 ;
  assign n60110 = n60108 & n60109 ;
  assign n60111 = ~n60057 & ~n60110 ;
  assign n60112 = n60057 & n60092 ;
  assign n60113 = n60094 & n60112 ;
  assign n60114 = n60069 & n60100 ;
  assign n60115 = n60075 & ~n60082 ;
  assign n60116 = ~n60069 & n60115 ;
  assign n60117 = n60082 & n60095 ;
  assign n60118 = ~n60116 & ~n60117 ;
  assign n60119 = ~n60114 & n60118 ;
  assign n60120 = n60057 & ~n60063 ;
  assign n60121 = ~n60119 & n60120 ;
  assign n60133 = ~n60113 & ~n60121 ;
  assign n60134 = ~n60111 & n60133 ;
  assign n60135 = ~n60132 & n60134 ;
  assign n60136 = ~\u0_L8_reg[6]/NET0131  & ~n60135 ;
  assign n60137 = \u0_L8_reg[6]/NET0131  & n60135 ;
  assign n60138 = ~n60136 & ~n60137 ;
  assign n60139 = n59054 & ~n59068 ;
  assign n60141 = ~n59045 & n59733 ;
  assign n60140 = n59110 & ~n59733 ;
  assign n60142 = ~n60007 & ~n60140 ;
  assign n60143 = ~n60141 & n60142 ;
  assign n60144 = n60139 & ~n60143 ;
  assign n60146 = ~n59099 & n60141 ;
  assign n60145 = ~n59054 & n59068 ;
  assign n60147 = ~n60139 & ~n60145 ;
  assign n60148 = ~n59994 & n60147 ;
  assign n60149 = ~n60140 & n60148 ;
  assign n60150 = ~n60146 & n60149 ;
  assign n60151 = ~n60144 & ~n60150 ;
  assign n60152 = ~n59083 & ~n60151 ;
  assign n60155 = n59060 & ~n59733 ;
  assign n60154 = ~n59039 & ~n59111 ;
  assign n60153 = n59047 & ~n59075 ;
  assign n60156 = n60145 & ~n60153 ;
  assign n60157 = ~n60154 & n60156 ;
  assign n60158 = ~n60155 & n60157 ;
  assign n60159 = ~n60152 & ~n60158 ;
  assign n60160 = ~\u0_L8_reg[7]/NET0131  & n60159 ;
  assign n60161 = \u0_L8_reg[7]/NET0131  & ~n60159 ;
  assign n60162 = ~n60160 & ~n60161 ;
  assign n60179 = n58860 & ~n58883 ;
  assign n60180 = ~n59138 & n60179 ;
  assign n60166 = ~n58874 & n59142 ;
  assign n60177 = n58854 & ~n58860 ;
  assign n60178 = n60166 & n60177 ;
  assign n60181 = ~n59125 & ~n60178 ;
  assign n60182 = ~n60180 & n60181 ;
  assign n60183 = n58848 & ~n60182 ;
  assign n60163 = n58881 & n59124 ;
  assign n60164 = n58854 & ~n59142 ;
  assign n60165 = ~n60163 & n60164 ;
  assign n60169 = n58873 & n60163 ;
  assign n60170 = ~n60165 & ~n60169 ;
  assign n60167 = ~n58854 & n60166 ;
  assign n60168 = n58860 & n59138 ;
  assign n60171 = ~n60167 & ~n60168 ;
  assign n60172 = n60170 & n60171 ;
  assign n60173 = ~n58848 & ~n60172 ;
  assign n60174 = ~n58867 & n58922 ;
  assign n60175 = ~n60169 & ~n60174 ;
  assign n60176 = ~n58854 & ~n60175 ;
  assign n60184 = ~n60173 & ~n60176 ;
  assign n60185 = ~n60183 & n60184 ;
  assign n60186 = ~\u0_L8_reg[9]/NET0131  & ~n60185 ;
  assign n60187 = \u0_L8_reg[9]/NET0131  & n60185 ;
  assign n60188 = ~n60186 & ~n60187 ;
  assign n60189 = n60076 & ~n60082 ;
  assign n60206 = n60099 & n60102 ;
  assign n60207 = ~n60189 & ~n60206 ;
  assign n60208 = n60118 & n60207 ;
  assign n60209 = ~n60089 & ~n60208 ;
  assign n60200 = n60089 & n60094 ;
  assign n60210 = n60075 & ~n60089 ;
  assign n60211 = ~n60069 & n60210 ;
  assign n60212 = ~n60200 & ~n60211 ;
  assign n60213 = ~n60063 & ~n60212 ;
  assign n60214 = ~n60090 & ~n60213 ;
  assign n60215 = ~n60209 & n60214 ;
  assign n60216 = n60057 & ~n60215 ;
  assign n60190 = ~n60117 & ~n60128 ;
  assign n60191 = ~n60189 & n60190 ;
  assign n60192 = ~n60063 & ~n60191 ;
  assign n60193 = ~n60082 & ~n60095 ;
  assign n60194 = n60063 & ~n60094 ;
  assign n60195 = ~n60117 & n60194 ;
  assign n60196 = ~n60193 & n60195 ;
  assign n60197 = ~n60129 & ~n60196 ;
  assign n60198 = ~n60192 & n60197 ;
  assign n60199 = ~n60057 & ~n60198 ;
  assign n60201 = ~n60082 & n60200 ;
  assign n60202 = ~n60104 & ~n60201 ;
  assign n60203 = n60063 & ~n60202 ;
  assign n60204 = ~n60063 & n60089 ;
  assign n60205 = n60115 & n60204 ;
  assign n60217 = ~n60203 & ~n60205 ;
  assign n60218 = ~n60199 & n60217 ;
  assign n60219 = ~n60216 & n60218 ;
  assign n60220 = ~\u0_L8_reg[16]/NET0131  & ~n60219 ;
  assign n60221 = \u0_L8_reg[16]/NET0131  & n60219 ;
  assign n60222 = ~n60220 & ~n60221 ;
  assign n60239 = ~n60063 & n60097 ;
  assign n60233 = n60075 & n60092 ;
  assign n60234 = ~n60124 & ~n60233 ;
  assign n60235 = n60063 & ~n60234 ;
  assign n60236 = n60063 & ~n60089 ;
  assign n60237 = ~n60076 & ~n60082 ;
  assign n60238 = n60236 & n60237 ;
  assign n60240 = ~n60106 & ~n60238 ;
  assign n60241 = ~n60235 & n60240 ;
  assign n60242 = ~n60239 & n60241 ;
  assign n60243 = n60057 & ~n60242 ;
  assign n60223 = n60076 & ~n60089 ;
  assign n60224 = ~n60200 & ~n60223 ;
  assign n60225 = n60082 & n60094 ;
  assign n60226 = n60089 & n60115 ;
  assign n60227 = ~n60225 & ~n60226 ;
  assign n60228 = n60224 & n60227 ;
  assign n60229 = n60063 & ~n60228 ;
  assign n60230 = n60089 & n60116 ;
  assign n60231 = ~n60229 & ~n60230 ;
  assign n60232 = ~n60057 & ~n60231 ;
  assign n60247 = n60093 & ~n60096 ;
  assign n60248 = n60125 & ~n60247 ;
  assign n60249 = ~n60057 & ~n60063 ;
  assign n60250 = ~n60248 & n60249 ;
  assign n60244 = n60117 & n60204 ;
  assign n60245 = ~n60083 & ~n60116 ;
  assign n60246 = n60236 & ~n60245 ;
  assign n60251 = ~n60244 & ~n60246 ;
  assign n60252 = ~n60250 & n60251 ;
  assign n60253 = ~n60232 & n60252 ;
  assign n60254 = ~n60243 & n60253 ;
  assign n60255 = ~\u0_L8_reg[24]/NET0131  & ~n60254 ;
  assign n60256 = \u0_L8_reg[24]/NET0131  & n60254 ;
  assign n60257 = ~n60255 & ~n60256 ;
  assign n60263 = n60089 & n60189 ;
  assign n60267 = ~n60057 & ~n60247 ;
  assign n60268 = ~n60263 & n60267 ;
  assign n60258 = n60075 & n60089 ;
  assign n60259 = ~n60102 & n60258 ;
  assign n60260 = ~n60069 & n60100 ;
  assign n60261 = ~n60259 & ~n60260 ;
  assign n60262 = n60063 & ~n60261 ;
  assign n60264 = ~n60102 & n60210 ;
  assign n60265 = ~n60083 & ~n60264 ;
  assign n60266 = ~n60063 & ~n60265 ;
  assign n60269 = ~n60262 & ~n60266 ;
  assign n60270 = n60268 & n60269 ;
  assign n60273 = ~n60089 & n60116 ;
  assign n60274 = n60224 & ~n60273 ;
  assign n60275 = n60063 & ~n60274 ;
  assign n60271 = ~n60225 & ~n60258 ;
  assign n60272 = ~n60063 & ~n60271 ;
  assign n60276 = n60057 & ~n60272 ;
  assign n60277 = ~n60275 & n60276 ;
  assign n60278 = ~n60270 & ~n60277 ;
  assign n60281 = n60063 & n60122 ;
  assign n60282 = n60258 & n60281 ;
  assign n60279 = ~n60095 & n60112 ;
  assign n60280 = n60102 & n60204 ;
  assign n60283 = ~n60279 & ~n60280 ;
  assign n60284 = ~n60282 & n60283 ;
  assign n60285 = ~n60278 & n60284 ;
  assign n60286 = \u0_L8_reg[30]/NET0131  & ~n60285 ;
  assign n60287 = ~\u0_L8_reg[30]/NET0131  & n60285 ;
  assign n60288 = ~n60286 & ~n60287 ;
  assign n60293 = n59315 & ~n59356 ;
  assign n60290 = n59298 & n59358 ;
  assign n60291 = ~n59306 & ~n60290 ;
  assign n60292 = ~n59315 & ~n60291 ;
  assign n60294 = ~n59371 & ~n60292 ;
  assign n60295 = ~n60293 & n60294 ;
  assign n60296 = n59343 & ~n60295 ;
  assign n60297 = n59307 & n59316 ;
  assign n60300 = ~n59505 & ~n59529 ;
  assign n60301 = ~n60297 & n60300 ;
  assign n60298 = ~n59298 & ~n59316 ;
  assign n60299 = ~n59347 & n60298 ;
  assign n60302 = ~n59366 & ~n60299 ;
  assign n60303 = n60301 & n60302 ;
  assign n60304 = ~n59343 & ~n60303 ;
  assign n60289 = ~n59315 & n59904 ;
  assign n60305 = ~n59365 & ~n59537 ;
  assign n60306 = n59315 & ~n60305 ;
  assign n60307 = ~n60289 & ~n60306 ;
  assign n60308 = ~n60304 & n60307 ;
  assign n60309 = ~n60296 & n60308 ;
  assign n60310 = \u0_L8_reg[18]/NET0131  & n60309 ;
  assign n60311 = ~\u0_L8_reg[18]/NET0131  & ~n60309 ;
  assign n60312 = ~n60310 & ~n60311 ;
  assign n60313 = decrypt_pad & ~\u0_uk_K_r7_reg[23]/P0001  ;
  assign n60314 = ~decrypt_pad & ~\u0_uk_K_r7_reg[30]/P0001  ;
  assign n60315 = ~n60313 & ~n60314 ;
  assign n60316 = \u0_R7_reg[28]/NET0131  & ~n60315 ;
  assign n60317 = ~\u0_R7_reg[28]/NET0131  & n60315 ;
  assign n60318 = ~n60316 & ~n60317 ;
  assign n60348 = decrypt_pad & ~\u0_uk_K_r7_reg[36]/NET0131  ;
  assign n60349 = ~decrypt_pad & ~\u0_uk_K_r7_reg[43]/NET0131  ;
  assign n60350 = ~n60348 & ~n60349 ;
  assign n60351 = \u0_R7_reg[27]/NET0131  & ~n60350 ;
  assign n60352 = ~\u0_R7_reg[27]/NET0131  & n60350 ;
  assign n60353 = ~n60351 & ~n60352 ;
  assign n60319 = decrypt_pad & ~\u0_uk_K_r7_reg[31]/NET0131  ;
  assign n60320 = ~decrypt_pad & ~\u0_uk_K_r7_reg[38]/NET0131  ;
  assign n60321 = ~n60319 & ~n60320 ;
  assign n60322 = \u0_R7_reg[26]/NET0131  & ~n60321 ;
  assign n60323 = ~\u0_R7_reg[26]/NET0131  & n60321 ;
  assign n60324 = ~n60322 & ~n60323 ;
  assign n60325 = decrypt_pad & ~\u0_uk_K_r7_reg[7]/NET0131  ;
  assign n60326 = ~decrypt_pad & ~\u0_uk_K_r7_reg[14]/NET0131  ;
  assign n60327 = ~n60325 & ~n60326 ;
  assign n60328 = \u0_R7_reg[24]/NET0131  & ~n60327 ;
  assign n60329 = ~\u0_R7_reg[24]/NET0131  & n60327 ;
  assign n60330 = ~n60328 & ~n60329 ;
  assign n60331 = n60324 & ~n60330 ;
  assign n60332 = ~n60324 & n60330 ;
  assign n60333 = ~n60331 & ~n60332 ;
  assign n60334 = decrypt_pad & ~\u0_uk_K_r7_reg[15]/NET0131  ;
  assign n60335 = ~decrypt_pad & ~\u0_uk_K_r7_reg[22]/NET0131  ;
  assign n60336 = ~n60334 & ~n60335 ;
  assign n60337 = \u0_R7_reg[29]/NET0131  & ~n60336 ;
  assign n60338 = ~\u0_R7_reg[29]/NET0131  & n60336 ;
  assign n60339 = ~n60337 & ~n60338 ;
  assign n60357 = n60333 & n60339 ;
  assign n60340 = decrypt_pad & ~\u0_uk_K_r7_reg[42]/NET0131  ;
  assign n60341 = ~decrypt_pad & ~\u0_uk_K_r7_reg[49]/NET0131  ;
  assign n60342 = ~n60340 & ~n60341 ;
  assign n60343 = \u0_R7_reg[25]/NET0131  & ~n60342 ;
  assign n60344 = ~\u0_R7_reg[25]/NET0131  & n60342 ;
  assign n60345 = ~n60343 & ~n60344 ;
  assign n60354 = n60324 & ~n60345 ;
  assign n60355 = n60330 & ~n60339 ;
  assign n60356 = ~n60354 & n60355 ;
  assign n60358 = ~n60339 & ~n60345 ;
  assign n60359 = n60331 & n60358 ;
  assign n60360 = ~n60356 & ~n60359 ;
  assign n60361 = ~n60357 & n60360 ;
  assign n60362 = ~n60353 & ~n60361 ;
  assign n60346 = n60339 & n60345 ;
  assign n60347 = n60333 & n60346 ;
  assign n60363 = n60332 & ~n60345 ;
  assign n60364 = n60353 & n60363 ;
  assign n60365 = ~n60347 & ~n60364 ;
  assign n60366 = ~n60362 & n60365 ;
  assign n60367 = ~n60318 & ~n60366 ;
  assign n60368 = ~n60332 & ~n60345 ;
  assign n60369 = n60330 & n60345 ;
  assign n60370 = n60318 & n60339 ;
  assign n60371 = ~n60369 & n60370 ;
  assign n60372 = ~n60333 & ~n60371 ;
  assign n60373 = ~n60368 & ~n60372 ;
  assign n60374 = ~n60353 & ~n60373 ;
  assign n60375 = ~n60330 & ~n60339 ;
  assign n60376 = n60324 & n60345 ;
  assign n60377 = n60375 & n60376 ;
  assign n60381 = n60353 & ~n60377 ;
  assign n60378 = ~n60330 & n60339 ;
  assign n60379 = n60354 & n60378 ;
  assign n60380 = ~n60331 & n60358 ;
  assign n60382 = ~n60379 & ~n60380 ;
  assign n60383 = n60381 & n60382 ;
  assign n60384 = ~n60374 & ~n60383 ;
  assign n60387 = ~n60324 & n60346 ;
  assign n60388 = ~n60354 & ~n60387 ;
  assign n60389 = n60330 & n60353 ;
  assign n60390 = ~n60388 & n60389 ;
  assign n60385 = ~n60324 & ~n60345 ;
  assign n60386 = n60375 & n60385 ;
  assign n60391 = ~n60379 & ~n60386 ;
  assign n60392 = ~n60390 & n60391 ;
  assign n60393 = n60318 & ~n60392 ;
  assign n60394 = ~n60384 & ~n60393 ;
  assign n60395 = ~n60367 & n60394 ;
  assign n60396 = ~\u0_L7_reg[22]/NET0131  & ~n60395 ;
  assign n60397 = \u0_L7_reg[22]/NET0131  & n60395 ;
  assign n60398 = ~n60396 & ~n60397 ;
  assign n60412 = decrypt_pad & ~\u0_uk_K_r7_reg[24]/NET0131  ;
  assign n60413 = ~decrypt_pad & ~\u0_uk_K_r7_reg[6]/NET0131  ;
  assign n60414 = ~n60412 & ~n60413 ;
  assign n60415 = \u0_R7_reg[32]/NET0131  & ~n60414 ;
  assign n60416 = ~\u0_R7_reg[32]/NET0131  & n60414 ;
  assign n60417 = ~n60415 & ~n60416 ;
  assign n60426 = decrypt_pad & ~\u0_uk_K_r7_reg[18]/NET0131  ;
  assign n60427 = ~decrypt_pad & ~\u0_uk_K_r7_reg[25]/NET0131  ;
  assign n60428 = ~n60426 & ~n60427 ;
  assign n60429 = \u0_R7_reg[5]/NET0131  & ~n60428 ;
  assign n60430 = ~\u0_R7_reg[5]/NET0131  & n60428 ;
  assign n60431 = ~n60429 & ~n60430 ;
  assign n60435 = ~n60417 & n60431 ;
  assign n60399 = decrypt_pad & ~\u0_uk_K_r7_reg[12]/NET0131  ;
  assign n60400 = ~decrypt_pad & ~\u0_uk_K_r7_reg[19]/NET0131  ;
  assign n60401 = ~n60399 & ~n60400 ;
  assign n60402 = \u0_R7_reg[3]/NET0131  & ~n60401 ;
  assign n60403 = ~\u0_R7_reg[3]/NET0131  & n60401 ;
  assign n60404 = ~n60402 & ~n60403 ;
  assign n60405 = decrypt_pad & ~\u0_uk_K_r7_reg[3]/NET0131  ;
  assign n60406 = ~decrypt_pad & ~\u0_uk_K_r7_reg[10]/NET0131  ;
  assign n60407 = ~n60405 & ~n60406 ;
  assign n60408 = \u0_R7_reg[2]/NET0131  & ~n60407 ;
  assign n60409 = ~\u0_R7_reg[2]/NET0131  & n60407 ;
  assign n60410 = ~n60408 & ~n60409 ;
  assign n60411 = n60404 & ~n60410 ;
  assign n60418 = decrypt_pad & ~\u0_uk_K_r7_reg[20]/NET0131  ;
  assign n60419 = ~decrypt_pad & ~\u0_uk_K_r7_reg[27]/NET0131  ;
  assign n60420 = ~n60418 & ~n60419 ;
  assign n60421 = \u0_R7_reg[1]/NET0131  & ~n60420 ;
  assign n60422 = ~\u0_R7_reg[1]/NET0131  & n60420 ;
  assign n60423 = ~n60421 & ~n60422 ;
  assign n60461 = ~n60411 & n60423 ;
  assign n60462 = n60435 & ~n60461 ;
  assign n60440 = decrypt_pad & ~\u0_uk_K_r7_reg[47]/NET0131  ;
  assign n60441 = ~decrypt_pad & ~\u0_uk_K_r7_reg[54]/NET0131  ;
  assign n60442 = ~n60440 & ~n60441 ;
  assign n60443 = \u0_R7_reg[4]/NET0131  & ~n60442 ;
  assign n60444 = ~\u0_R7_reg[4]/NET0131  & n60442 ;
  assign n60445 = ~n60443 & ~n60444 ;
  assign n60448 = ~n60410 & n60417 ;
  assign n60457 = ~n60423 & ~n60431 ;
  assign n60467 = n60448 & n60457 ;
  assign n60472 = n60445 & ~n60467 ;
  assign n60473 = ~n60462 & n60472 ;
  assign n60447 = n60410 & ~n60417 ;
  assign n60463 = ~n60431 & ~n60447 ;
  assign n60464 = n60423 & n60431 ;
  assign n60465 = n60404 & ~n60464 ;
  assign n60466 = ~n60463 & n60465 ;
  assign n60468 = ~n60417 & n60423 ;
  assign n60469 = ~n60404 & n60423 ;
  assign n60470 = ~n60447 & ~n60469 ;
  assign n60471 = ~n60468 & ~n60470 ;
  assign n60474 = ~n60466 & ~n60471 ;
  assign n60475 = n60473 & n60474 ;
  assign n60432 = n60417 & n60431 ;
  assign n60480 = n60432 & ~n60469 ;
  assign n60476 = ~n60417 & ~n60431 ;
  assign n60481 = n60423 & n60476 ;
  assign n60482 = ~n60480 & ~n60481 ;
  assign n60483 = ~n60410 & ~n60482 ;
  assign n60477 = ~n60432 & ~n60476 ;
  assign n60433 = n60410 & n60423 ;
  assign n60478 = n60404 & n60433 ;
  assign n60479 = n60477 & n60478 ;
  assign n60484 = ~n60445 & ~n60479 ;
  assign n60485 = ~n60483 & n60484 ;
  assign n60486 = ~n60475 & ~n60485 ;
  assign n60449 = ~n60447 & ~n60448 ;
  assign n60446 = ~n60423 & n60431 ;
  assign n60450 = ~n60433 & ~n60445 ;
  assign n60451 = ~n60446 & n60450 ;
  assign n60452 = n60449 & n60451 ;
  assign n60436 = n60410 & n60435 ;
  assign n60437 = ~n60423 & n60436 ;
  assign n60434 = n60432 & n60433 ;
  assign n60438 = ~n60410 & n60423 ;
  assign n60439 = ~n60431 & n60438 ;
  assign n60453 = ~n60434 & ~n60439 ;
  assign n60454 = ~n60437 & n60453 ;
  assign n60455 = ~n60452 & n60454 ;
  assign n60456 = ~n60404 & ~n60455 ;
  assign n60424 = n60417 & ~n60423 ;
  assign n60425 = n60411 & n60424 ;
  assign n60458 = n60410 & n60457 ;
  assign n60459 = n60404 & ~n60417 ;
  assign n60460 = n60458 & n60459 ;
  assign n60487 = ~n60425 & ~n60460 ;
  assign n60488 = ~n60456 & n60487 ;
  assign n60489 = ~n60486 & n60488 ;
  assign n60490 = ~\u0_L7_reg[31]/NET0131  & ~n60489 ;
  assign n60491 = \u0_L7_reg[31]/NET0131  & n60489 ;
  assign n60492 = ~n60490 & ~n60491 ;
  assign n60499 = decrypt_pad & ~\u0_uk_K_r7_reg[14]/NET0131  ;
  assign n60500 = ~decrypt_pad & ~\u0_uk_K_r7_reg[21]/NET0131  ;
  assign n60501 = ~n60499 & ~n60500 ;
  assign n60502 = \u0_R7_reg[23]/NET0131  & ~n60501 ;
  assign n60503 = ~\u0_R7_reg[23]/NET0131  & n60501 ;
  assign n60504 = ~n60502 & ~n60503 ;
  assign n60505 = decrypt_pad & ~\u0_uk_K_r7_reg[35]/NET0131  ;
  assign n60506 = ~decrypt_pad & ~\u0_uk_K_r7_reg[42]/NET0131  ;
  assign n60507 = ~n60505 & ~n60506 ;
  assign n60508 = \u0_R7_reg[25]/NET0131  & ~n60507 ;
  assign n60509 = ~\u0_R7_reg[25]/NET0131  & n60507 ;
  assign n60510 = ~n60508 & ~n60509 ;
  assign n60511 = decrypt_pad & ~\u0_uk_K_r7_reg[50]/NET0131  ;
  assign n60512 = ~decrypt_pad & ~\u0_uk_K_r7_reg[2]/NET0131  ;
  assign n60513 = ~n60511 & ~n60512 ;
  assign n60514 = \u0_R7_reg[20]/NET0131  & ~n60513 ;
  assign n60515 = ~\u0_R7_reg[20]/NET0131  & n60513 ;
  assign n60516 = ~n60514 & ~n60515 ;
  assign n60517 = n60510 & n60516 ;
  assign n60526 = decrypt_pad & ~\u0_uk_K_r7_reg[1]/NET0131  ;
  assign n60527 = ~decrypt_pad & ~\u0_uk_K_r7_reg[8]/NET0131  ;
  assign n60528 = ~n60526 & ~n60527 ;
  assign n60529 = \u0_R7_reg[22]/NET0131  & ~n60528 ;
  assign n60530 = ~\u0_R7_reg[22]/NET0131  & n60528 ;
  assign n60531 = ~n60529 & ~n60530 ;
  assign n60562 = n60517 & n60531 ;
  assign n60518 = decrypt_pad & ~\u0_uk_K_r7_reg[38]/NET0131  ;
  assign n60519 = ~decrypt_pad & ~\u0_uk_K_r7_reg[45]/NET0131  ;
  assign n60520 = ~n60518 & ~n60519 ;
  assign n60521 = \u0_R7_reg[21]/NET0131  & ~n60520 ;
  assign n60522 = ~\u0_R7_reg[21]/NET0131  & n60520 ;
  assign n60523 = ~n60521 & ~n60522 ;
  assign n60569 = ~n60516 & ~n60523 ;
  assign n60572 = n60510 & n60569 ;
  assign n60573 = ~n60516 & ~n60531 ;
  assign n60574 = ~n60572 & ~n60573 ;
  assign n60493 = decrypt_pad & ~\u0_uk_K_r7_reg[16]/NET0131  ;
  assign n60494 = ~decrypt_pad & ~\u0_uk_K_r7_reg[23]/P0001  ;
  assign n60495 = ~n60493 & ~n60494 ;
  assign n60496 = \u0_R7_reg[24]/NET0131  & ~n60495 ;
  assign n60497 = ~\u0_R7_reg[24]/NET0131  & n60495 ;
  assign n60498 = ~n60496 & ~n60497 ;
  assign n60575 = ~n60510 & n60573 ;
  assign n60576 = n60523 & n60575 ;
  assign n60577 = n60498 & ~n60576 ;
  assign n60578 = ~n60574 & ~n60577 ;
  assign n60579 = ~n60562 & ~n60578 ;
  assign n60580 = n60504 & ~n60579 ;
  assign n60533 = ~n60510 & n60516 ;
  assign n60534 = ~n60523 & n60533 ;
  assign n60535 = ~n60531 & n60534 ;
  assign n60524 = n60517 & n60523 ;
  assign n60525 = ~n60516 & n60523 ;
  assign n60532 = n60525 & n60531 ;
  assign n60536 = ~n60524 & ~n60532 ;
  assign n60537 = ~n60535 & n60536 ;
  assign n60538 = n60504 & ~n60537 ;
  assign n60542 = n60510 & n60523 ;
  assign n60543 = ~n60531 & ~n60542 ;
  assign n60544 = ~n60504 & ~n60517 ;
  assign n60545 = ~n60532 & n60544 ;
  assign n60546 = ~n60543 & n60545 ;
  assign n60539 = n60517 & ~n60531 ;
  assign n60540 = ~n60504 & ~n60523 ;
  assign n60541 = n60539 & n60540 ;
  assign n60547 = n60498 & ~n60541 ;
  assign n60548 = ~n60546 & n60547 ;
  assign n60549 = ~n60538 & n60548 ;
  assign n60550 = n60523 & ~n60531 ;
  assign n60551 = n60516 & n60550 ;
  assign n60552 = ~n60532 & ~n60551 ;
  assign n60553 = ~n60504 & ~n60552 ;
  assign n60565 = ~n60498 & ~n60553 ;
  assign n60554 = n60504 & n60531 ;
  assign n60555 = ~n60523 & n60554 ;
  assign n60556 = ~n60510 & n60523 ;
  assign n60557 = ~n60531 & n60556 ;
  assign n60558 = ~n60555 & ~n60557 ;
  assign n60559 = n60516 & ~n60558 ;
  assign n60560 = ~n60504 & ~n60531 ;
  assign n60561 = n60533 & n60560 ;
  assign n60563 = ~n60523 & n60562 ;
  assign n60564 = ~n60561 & ~n60563 ;
  assign n60566 = ~n60559 & n60564 ;
  assign n60567 = n60565 & n60566 ;
  assign n60568 = ~n60549 & ~n60567 ;
  assign n60570 = ~n60510 & n60569 ;
  assign n60571 = n60560 & n60570 ;
  assign n60581 = n60516 & n60556 ;
  assign n60582 = ~n60504 & ~n60581 ;
  assign n60583 = ~n60531 & n60572 ;
  assign n60584 = ~n60560 & ~n60583 ;
  assign n60585 = ~n60582 & ~n60584 ;
  assign n60586 = ~n60571 & ~n60585 ;
  assign n60587 = ~n60568 & n60586 ;
  assign n60588 = ~n60580 & n60587 ;
  assign n60589 = \u0_L7_reg[11]/NET0131  & ~n60588 ;
  assign n60590 = ~\u0_L7_reg[11]/NET0131  & n60588 ;
  assign n60591 = ~n60589 & ~n60590 ;
  assign n60592 = decrypt_pad & ~\u0_uk_K_r7_reg[37]/NET0131  ;
  assign n60593 = ~decrypt_pad & ~\u0_uk_K_r7_reg[44]/NET0131  ;
  assign n60594 = ~n60592 & ~n60593 ;
  assign n60595 = \u0_R7_reg[31]/P0001  & ~n60594 ;
  assign n60596 = ~\u0_R7_reg[31]/P0001  & n60594 ;
  assign n60597 = ~n60595 & ~n60596 ;
  assign n60598 = decrypt_pad & ~\u0_uk_K_r7_reg[21]/NET0131  ;
  assign n60599 = ~decrypt_pad & ~\u0_uk_K_r7_reg[28]/NET0131  ;
  assign n60600 = ~n60598 & ~n60599 ;
  assign n60601 = \u0_R7_reg[28]/NET0131  & ~n60600 ;
  assign n60602 = ~\u0_R7_reg[28]/NET0131  & n60600 ;
  assign n60603 = ~n60601 & ~n60602 ;
  assign n60611 = decrypt_pad & ~\u0_uk_K_r7_reg[49]/NET0131  ;
  assign n60612 = ~decrypt_pad & ~\u0_uk_K_r7_reg[1]/NET0131  ;
  assign n60613 = ~n60611 & ~n60612 ;
  assign n60614 = \u0_R7_reg[30]/NET0131  & ~n60613 ;
  assign n60615 = ~\u0_R7_reg[30]/NET0131  & n60613 ;
  assign n60616 = ~n60614 & ~n60615 ;
  assign n60625 = n60603 & ~n60616 ;
  assign n60604 = decrypt_pad & ~\u0_uk_K_r7_reg[9]/NET0131  ;
  assign n60605 = ~decrypt_pad & ~\u0_uk_K_r7_reg[16]/NET0131  ;
  assign n60606 = ~n60604 & ~n60605 ;
  assign n60607 = \u0_R7_reg[1]/NET0131  & ~n60606 ;
  assign n60608 = ~\u0_R7_reg[1]/NET0131  & n60606 ;
  assign n60609 = ~n60607 & ~n60608 ;
  assign n60617 = decrypt_pad & ~\u0_uk_K_r7_reg[52]/NET0131  ;
  assign n60618 = ~decrypt_pad & ~\u0_uk_K_r7_reg[0]/NET0131  ;
  assign n60619 = ~n60617 & ~n60618 ;
  assign n60620 = \u0_R7_reg[29]/NET0131  & ~n60619 ;
  assign n60621 = ~\u0_R7_reg[29]/NET0131  & n60619 ;
  assign n60622 = ~n60620 & ~n60621 ;
  assign n60626 = ~n60609 & n60622 ;
  assign n60627 = ~n60625 & ~n60626 ;
  assign n60610 = n60603 & ~n60609 ;
  assign n60623 = ~n60616 & n60622 ;
  assign n60624 = n60610 & n60623 ;
  assign n60628 = decrypt_pad & ~\u0_uk_K_r7_reg[43]/NET0131  ;
  assign n60629 = ~decrypt_pad & ~\u0_uk_K_r7_reg[50]/NET0131  ;
  assign n60630 = ~n60628 & ~n60629 ;
  assign n60631 = \u0_R7_reg[32]/NET0131  & ~n60630 ;
  assign n60632 = ~\u0_R7_reg[32]/NET0131  & n60630 ;
  assign n60633 = ~n60631 & ~n60632 ;
  assign n60634 = ~n60624 & n60633 ;
  assign n60635 = ~n60627 & n60634 ;
  assign n60641 = ~n60603 & ~n60616 ;
  assign n60642 = ~n60622 & n60641 ;
  assign n60643 = ~n60609 & n60642 ;
  assign n60636 = n60609 & ~n60622 ;
  assign n60637 = ~n60603 & n60616 ;
  assign n60638 = n60636 & n60637 ;
  assign n60639 = ~n60610 & ~n60623 ;
  assign n60640 = ~n60627 & n60639 ;
  assign n60644 = ~n60638 & ~n60640 ;
  assign n60645 = ~n60643 & n60644 ;
  assign n60646 = ~n60635 & n60645 ;
  assign n60647 = n60597 & ~n60646 ;
  assign n60652 = n60597 & ~n60624 ;
  assign n60648 = ~n60609 & ~n60622 ;
  assign n60649 = n60603 & n60616 ;
  assign n60650 = n60648 & n60649 ;
  assign n60651 = ~n60603 & n60636 ;
  assign n60653 = ~n60650 & ~n60651 ;
  assign n60654 = n60652 & n60653 ;
  assign n60655 = ~n60609 & ~n60616 ;
  assign n60656 = ~n60610 & ~n60636 ;
  assign n60657 = ~n60655 & n60656 ;
  assign n60658 = ~n60597 & ~n60625 ;
  assign n60659 = ~n60657 & n60658 ;
  assign n60660 = ~n60654 & ~n60659 ;
  assign n60661 = n60622 & n60649 ;
  assign n60662 = n60609 & n60661 ;
  assign n60663 = ~n60633 & ~n60662 ;
  assign n60664 = ~n60660 & n60663 ;
  assign n60668 = ~n60622 & n60649 ;
  assign n60669 = ~n60642 & ~n60668 ;
  assign n60670 = ~n60624 & n60669 ;
  assign n60671 = ~n60597 & ~n60670 ;
  assign n60665 = ~n60603 & n60609 ;
  assign n60666 = n60622 & n60665 ;
  assign n60667 = n60616 & n60666 ;
  assign n60672 = n60633 & ~n60667 ;
  assign n60673 = ~n60671 & n60672 ;
  assign n60674 = ~n60664 & ~n60673 ;
  assign n60675 = ~n60647 & ~n60674 ;
  assign n60676 = \u0_L7_reg[5]/NET0131  & ~n60675 ;
  assign n60677 = ~\u0_L7_reg[5]/NET0131  & n60675 ;
  assign n60678 = ~n60676 & ~n60677 ;
  assign n60680 = n60597 & ~n60603 ;
  assign n60681 = n60616 & n60636 ;
  assign n60682 = ~n60680 & n60681 ;
  assign n60679 = n60622 & n60625 ;
  assign n60685 = n60633 & ~n60679 ;
  assign n60683 = n60626 & n60637 ;
  assign n60684 = n60648 & n60680 ;
  assign n60686 = ~n60683 & ~n60684 ;
  assign n60687 = n60685 & n60686 ;
  assign n60688 = ~n60682 & n60687 ;
  assign n60691 = n60597 & ~n60666 ;
  assign n60692 = n60622 & ~n60637 ;
  assign n60693 = ~n60665 & ~n60692 ;
  assign n60694 = n60691 & ~n60693 ;
  assign n60689 = n60603 & ~n60622 ;
  assign n60690 = n60655 & n60689 ;
  assign n60695 = ~n60633 & ~n60690 ;
  assign n60696 = ~n60694 & n60695 ;
  assign n60697 = ~n60688 & ~n60696 ;
  assign n60698 = ~n60616 & n60651 ;
  assign n60699 = n60597 & ~n60667 ;
  assign n60700 = ~n60698 & n60699 ;
  assign n60704 = ~n60597 & ~n60683 ;
  assign n60701 = ~n60616 & n60633 ;
  assign n60702 = n60689 & ~n60701 ;
  assign n60703 = n60623 & n60665 ;
  assign n60705 = ~n60702 & ~n60703 ;
  assign n60706 = n60704 & n60705 ;
  assign n60707 = ~n60643 & n60706 ;
  assign n60708 = ~n60700 & ~n60707 ;
  assign n60709 = ~n60697 & ~n60708 ;
  assign n60710 = \u0_L7_reg[15]/P0001  & n60709 ;
  assign n60711 = ~\u0_L7_reg[15]/P0001  & ~n60709 ;
  assign n60712 = ~n60710 & ~n60711 ;
  assign n60748 = decrypt_pad & ~\u0_uk_K_r7_reg[54]/NET0131  ;
  assign n60749 = ~decrypt_pad & ~\u0_uk_K_r7_reg[4]/NET0131  ;
  assign n60750 = ~n60748 & ~n60749 ;
  assign n60751 = \u0_R7_reg[17]/NET0131  & ~n60750 ;
  assign n60752 = ~\u0_R7_reg[17]/NET0131  & n60750 ;
  assign n60753 = ~n60751 & ~n60752 ;
  assign n60725 = decrypt_pad & ~\u0_uk_K_r7_reg[33]/NET0131  ;
  assign n60726 = ~decrypt_pad & ~\u0_uk_K_r7_reg[40]/NET0131  ;
  assign n60727 = ~n60725 & ~n60726 ;
  assign n60728 = \u0_R7_reg[14]/NET0131  & ~n60727 ;
  assign n60729 = ~\u0_R7_reg[14]/NET0131  & n60727 ;
  assign n60730 = ~n60728 & ~n60729 ;
  assign n60732 = decrypt_pad & ~\u0_uk_K_r7_reg[32]/NET0131  ;
  assign n60733 = ~decrypt_pad & ~\u0_uk_K_r7_reg[39]/NET0131  ;
  assign n60734 = ~n60732 & ~n60733 ;
  assign n60735 = \u0_R7_reg[13]/NET0131  & ~n60734 ;
  assign n60736 = ~\u0_R7_reg[13]/NET0131  & n60734 ;
  assign n60737 = ~n60735 & ~n60736 ;
  assign n60771 = ~n60730 & n60737 ;
  assign n60719 = decrypt_pad & ~\u0_uk_K_r7_reg[13]/NET0131  ;
  assign n60720 = ~decrypt_pad & ~\u0_uk_K_r7_reg[20]/NET0131  ;
  assign n60721 = ~n60719 & ~n60720 ;
  assign n60722 = \u0_R7_reg[12]/NET0131  & ~n60721 ;
  assign n60723 = ~\u0_R7_reg[12]/NET0131  & n60721 ;
  assign n60724 = ~n60722 & ~n60723 ;
  assign n60739 = ~n60724 & n60730 ;
  assign n60741 = decrypt_pad & ~\u0_uk_K_r7_reg[41]/NET0131  ;
  assign n60742 = ~decrypt_pad & ~\u0_uk_K_r7_reg[48]/NET0131  ;
  assign n60743 = ~n60741 & ~n60742 ;
  assign n60744 = \u0_R7_reg[15]/NET0131  & ~n60743 ;
  assign n60745 = ~\u0_R7_reg[15]/NET0131  & n60743 ;
  assign n60746 = ~n60744 & ~n60745 ;
  assign n60777 = ~n60739 & n60746 ;
  assign n60778 = ~n60771 & ~n60777 ;
  assign n60779 = n60753 & ~n60778 ;
  assign n60781 = n60737 & n60753 ;
  assign n60780 = ~n60737 & n60746 ;
  assign n60782 = n60739 & ~n60780 ;
  assign n60783 = ~n60781 & n60782 ;
  assign n60784 = n60724 & n60780 ;
  assign n60754 = ~n60737 & ~n60753 ;
  assign n60755 = ~n60746 & n60754 ;
  assign n60713 = decrypt_pad & ~\u0_uk_K_r7_reg[17]/NET0131  ;
  assign n60714 = ~decrypt_pad & ~\u0_uk_K_r7_reg[24]/NET0131  ;
  assign n60715 = ~n60713 & ~n60714 ;
  assign n60716 = \u0_R7_reg[16]/NET0131  & ~n60715 ;
  assign n60717 = ~\u0_R7_reg[16]/NET0131  & n60715 ;
  assign n60718 = ~n60716 & ~n60717 ;
  assign n60731 = n60724 & ~n60730 ;
  assign n60785 = n60718 & ~n60731 ;
  assign n60786 = ~n60755 & n60785 ;
  assign n60787 = ~n60784 & n60786 ;
  assign n60788 = ~n60783 & n60787 ;
  assign n60789 = ~n60779 & n60788 ;
  assign n60740 = ~n60737 & n60739 ;
  assign n60747 = n60740 & ~n60746 ;
  assign n60738 = n60731 & ~n60737 ;
  assign n60766 = ~n60738 & ~n60755 ;
  assign n60767 = ~n60747 & n60766 ;
  assign n60756 = n60724 & ~n60753 ;
  assign n60757 = n60737 & n60746 ;
  assign n60758 = n60756 & n60757 ;
  assign n60759 = ~n60724 & n60737 ;
  assign n60760 = ~n60730 & n60753 ;
  assign n60761 = n60759 & n60760 ;
  assign n60762 = ~n60758 & ~n60761 ;
  assign n60763 = ~n60724 & n60753 ;
  assign n60764 = n60730 & n60757 ;
  assign n60765 = ~n60763 & n60764 ;
  assign n60768 = n60762 & ~n60765 ;
  assign n60769 = n60767 & n60768 ;
  assign n60770 = ~n60718 & ~n60769 ;
  assign n60772 = ~n60756 & ~n60763 ;
  assign n60773 = n60771 & n60772 ;
  assign n60774 = n60731 & n60754 ;
  assign n60775 = ~n60773 & ~n60774 ;
  assign n60776 = ~n60746 & ~n60775 ;
  assign n60790 = ~n60724 & n60771 ;
  assign n60791 = ~n60738 & ~n60790 ;
  assign n60792 = n60746 & n60753 ;
  assign n60793 = ~n60791 & n60792 ;
  assign n60794 = ~n60776 & ~n60793 ;
  assign n60795 = ~n60770 & n60794 ;
  assign n60796 = ~n60789 & n60795 ;
  assign n60797 = ~\u0_L7_reg[26]/NET0131  & ~n60796 ;
  assign n60798 = \u0_L7_reg[26]/NET0131  & n60796 ;
  assign n60799 = ~n60797 & ~n60798 ;
  assign n60810 = n60516 & ~n60556 ;
  assign n60811 = n60560 & ~n60810 ;
  assign n60808 = n60504 & ~n60531 ;
  assign n60809 = n60517 & n60808 ;
  assign n60812 = n60531 & n60542 ;
  assign n60813 = ~n60809 & ~n60812 ;
  assign n60814 = ~n60811 & n60813 ;
  assign n60815 = n60577 & n60814 ;
  assign n60816 = n60531 & n60572 ;
  assign n60817 = ~n60504 & ~n60816 ;
  assign n60818 = ~n60510 & n60525 ;
  assign n60819 = ~n60539 & ~n60818 ;
  assign n60820 = n60817 & n60819 ;
  assign n60821 = n60510 & n60573 ;
  assign n60822 = n60504 & ~n60581 ;
  assign n60823 = ~n60821 & n60822 ;
  assign n60824 = ~n60563 & n60823 ;
  assign n60825 = ~n60820 & ~n60824 ;
  assign n60826 = ~n60498 & ~n60535 ;
  assign n60827 = ~n60825 & n60826 ;
  assign n60828 = ~n60815 & ~n60827 ;
  assign n60800 = n60510 & n60525 ;
  assign n60801 = ~n60570 & ~n60800 ;
  assign n60802 = ~n60581 & n60801 ;
  assign n60803 = n60554 & ~n60802 ;
  assign n60804 = ~n60524 & ~n60534 ;
  assign n60805 = n60531 & ~n60804 ;
  assign n60806 = ~n60575 & ~n60805 ;
  assign n60807 = ~n60504 & ~n60806 ;
  assign n60829 = ~n60803 & ~n60807 ;
  assign n60830 = ~n60828 & n60829 ;
  assign n60831 = ~\u0_L7_reg[4]/NET0131  & ~n60830 ;
  assign n60832 = \u0_L7_reg[4]/NET0131  & n60830 ;
  assign n60833 = ~n60831 & ~n60832 ;
  assign n60834 = n60730 & ~n60753 ;
  assign n60857 = n60724 & ~n60781 ;
  assign n60858 = ~n60834 & n60857 ;
  assign n60859 = ~n60746 & ~n60858 ;
  assign n60846 = n60730 & n60756 ;
  assign n60861 = ~n60737 & n60846 ;
  assign n60842 = ~n60724 & ~n60753 ;
  assign n60860 = ~n60730 & n60842 ;
  assign n60862 = n60746 & ~n60860 ;
  assign n60863 = ~n60861 & n60862 ;
  assign n60864 = ~n60859 & ~n60863 ;
  assign n60836 = n60724 & n60781 ;
  assign n60837 = n60730 & n60836 ;
  assign n60865 = n60771 & ~n60772 ;
  assign n60866 = ~n60837 & ~n60865 ;
  assign n60867 = ~n60864 & n60866 ;
  assign n60868 = ~n60718 & ~n60867 ;
  assign n60850 = ~n60753 & ~n60790 ;
  assign n60851 = ~n60759 & ~n60771 ;
  assign n60852 = ~n60746 & ~n60851 ;
  assign n60853 = ~n60850 & n60852 ;
  assign n60847 = n60737 & n60846 ;
  assign n60854 = ~n60740 & ~n60847 ;
  assign n60855 = ~n60853 & n60854 ;
  assign n60856 = n60718 & ~n60855 ;
  assign n60835 = n60759 & n60834 ;
  assign n60838 = n60740 & n60753 ;
  assign n60839 = ~n60837 & ~n60838 ;
  assign n60840 = ~n60835 & n60839 ;
  assign n60841 = n60746 & ~n60840 ;
  assign n60848 = ~n60746 & n60847 ;
  assign n60843 = n60718 & n60780 ;
  assign n60844 = ~n60834 & ~n60842 ;
  assign n60845 = n60843 & n60844 ;
  assign n60849 = n60739 & n60755 ;
  assign n60869 = ~n60845 & ~n60849 ;
  assign n60870 = ~n60848 & n60869 ;
  assign n60871 = ~n60841 & n60870 ;
  assign n60872 = ~n60856 & n60871 ;
  assign n60873 = ~n60868 & n60872 ;
  assign n60874 = ~\u0_L7_reg[1]/NET0131  & ~n60873 ;
  assign n60875 = \u0_L7_reg[1]/NET0131  & n60873 ;
  assign n60876 = ~n60874 & ~n60875 ;
  assign n60898 = ~n60410 & n60476 ;
  assign n60899 = n60423 & ~n60898 ;
  assign n60900 = ~n60404 & ~n60477 ;
  assign n60901 = ~n60899 & n60900 ;
  assign n60894 = ~n60457 & ~n60464 ;
  assign n60895 = n60417 & ~n60894 ;
  assign n60896 = n60404 & n60895 ;
  assign n60890 = ~n60431 & n60433 ;
  assign n60897 = n60417 & n60890 ;
  assign n60902 = ~n60437 & ~n60897 ;
  assign n60903 = ~n60896 & n60902 ;
  assign n60904 = ~n60901 & n60903 ;
  assign n60905 = ~n60445 & ~n60904 ;
  assign n60878 = ~n60410 & ~n60423 ;
  assign n60879 = ~n60417 & ~n60878 ;
  assign n60880 = n60432 & n60878 ;
  assign n60881 = ~n60879 & ~n60880 ;
  assign n60882 = n60404 & ~n60881 ;
  assign n60884 = ~n60404 & ~n60468 ;
  assign n60885 = n60449 & n60884 ;
  assign n60877 = n60431 & n60433 ;
  assign n60883 = n60417 & n60439 ;
  assign n60886 = ~n60877 & ~n60883 ;
  assign n60887 = ~n60885 & n60886 ;
  assign n60888 = ~n60882 & n60887 ;
  assign n60889 = n60445 & ~n60888 ;
  assign n60891 = n60431 & n60438 ;
  assign n60892 = ~n60890 & ~n60891 ;
  assign n60893 = n60459 & ~n60892 ;
  assign n60906 = ~n60889 & ~n60893 ;
  assign n60907 = ~n60905 & n60906 ;
  assign n60908 = ~\u0_L7_reg[17]/NET0131  & ~n60907 ;
  assign n60909 = \u0_L7_reg[17]/NET0131  & n60907 ;
  assign n60910 = ~n60908 & ~n60909 ;
  assign n60911 = decrypt_pad & ~\u0_uk_K_r7_reg[48]/NET0131  ;
  assign n60912 = ~decrypt_pad & ~\u0_uk_K_r7_reg[55]/P0001  ;
  assign n60913 = ~n60911 & ~n60912 ;
  assign n60914 = \u0_R7_reg[8]/NET0131  & ~n60913 ;
  assign n60915 = ~\u0_R7_reg[8]/NET0131  & n60913 ;
  assign n60916 = ~n60914 & ~n60915 ;
  assign n60917 = decrypt_pad & ~\u0_uk_K_r7_reg[6]/NET0131  ;
  assign n60918 = ~decrypt_pad & ~\u0_uk_K_r7_reg[13]/NET0131  ;
  assign n60919 = ~n60917 & ~n60918 ;
  assign n60920 = \u0_R7_reg[6]/NET0131  & ~n60919 ;
  assign n60921 = ~\u0_R7_reg[6]/NET0131  & n60919 ;
  assign n60922 = ~n60920 & ~n60921 ;
  assign n60923 = decrypt_pad & ~\u0_uk_K_r7_reg[53]/NET0131  ;
  assign n60924 = ~decrypt_pad & ~\u0_uk_K_r7_reg[3]/NET0131  ;
  assign n60925 = ~n60923 & ~n60924 ;
  assign n60926 = \u0_R7_reg[9]/NET0131  & ~n60925 ;
  assign n60927 = ~\u0_R7_reg[9]/NET0131  & n60925 ;
  assign n60928 = ~n60926 & ~n60927 ;
  assign n60929 = ~n60922 & n60928 ;
  assign n60930 = decrypt_pad & ~\u0_uk_K_r7_reg[40]/NET0131  ;
  assign n60931 = ~decrypt_pad & ~\u0_uk_K_r7_reg[47]/NET0131  ;
  assign n60932 = ~n60930 & ~n60931 ;
  assign n60933 = \u0_R7_reg[5]/NET0131  & ~n60932 ;
  assign n60934 = ~\u0_R7_reg[5]/NET0131  & n60932 ;
  assign n60935 = ~n60933 & ~n60934 ;
  assign n60936 = decrypt_pad & ~\u0_uk_K_r7_reg[25]/NET0131  ;
  assign n60937 = ~decrypt_pad & ~\u0_uk_K_r7_reg[32]/NET0131  ;
  assign n60938 = ~n60936 & ~n60937 ;
  assign n60939 = \u0_R7_reg[7]/NET0131  & ~n60938 ;
  assign n60940 = ~\u0_R7_reg[7]/NET0131  & n60938 ;
  assign n60941 = ~n60939 & ~n60940 ;
  assign n60942 = ~n60935 & ~n60941 ;
  assign n60943 = n60929 & n60942 ;
  assign n60944 = decrypt_pad & ~\u0_uk_K_r7_reg[4]/NET0131  ;
  assign n60945 = ~decrypt_pad & ~\u0_uk_K_r7_reg[11]/NET0131  ;
  assign n60946 = ~n60944 & ~n60945 ;
  assign n60947 = \u0_R7_reg[4]/NET0131  & ~n60946 ;
  assign n60948 = ~\u0_R7_reg[4]/NET0131  & n60946 ;
  assign n60949 = ~n60947 & ~n60948 ;
  assign n60950 = n60928 & ~n60949 ;
  assign n60951 = n60935 & n60950 ;
  assign n60952 = n60922 & n60951 ;
  assign n60953 = ~n60943 & ~n60952 ;
  assign n60955 = n60928 & ~n60935 ;
  assign n60960 = n60922 & n60949 ;
  assign n60961 = n60955 & n60960 ;
  assign n60962 = n60941 & n60961 ;
  assign n60967 = n60953 & ~n60962 ;
  assign n60954 = n60928 & n60949 ;
  assign n60956 = ~n60928 & n60935 ;
  assign n60957 = ~n60955 & ~n60956 ;
  assign n60958 = ~n60954 & ~n60957 ;
  assign n60959 = ~n60922 & n60958 ;
  assign n60963 = ~n60935 & n60954 ;
  assign n60964 = ~n60941 & ~n60963 ;
  assign n60965 = ~n60955 & ~n60960 ;
  assign n60966 = n60964 & ~n60965 ;
  assign n60968 = ~n60959 & ~n60966 ;
  assign n60969 = n60967 & n60968 ;
  assign n60970 = ~n60916 & ~n60969 ;
  assign n60972 = ~n60928 & ~n60949 ;
  assign n60989 = ~n60961 & ~n60972 ;
  assign n60990 = n60916 & ~n60989 ;
  assign n60971 = n60922 & ~n60935 ;
  assign n60991 = n60950 & ~n60971 ;
  assign n60992 = ~n60990 & ~n60991 ;
  assign n60988 = ~n60922 & n60935 ;
  assign n60993 = ~n60941 & ~n60988 ;
  assign n60994 = ~n60992 & n60993 ;
  assign n60973 = n60971 & n60972 ;
  assign n60974 = n60935 & n60949 ;
  assign n60975 = ~n60922 & n60974 ;
  assign n60976 = ~n60973 & ~n60975 ;
  assign n60977 = n60941 & ~n60976 ;
  assign n60978 = ~n60928 & ~n60935 ;
  assign n60979 = ~n60922 & n60978 ;
  assign n60980 = n60949 & n60979 ;
  assign n60981 = n60922 & ~n60949 ;
  assign n60982 = n60935 & n60941 ;
  assign n60983 = ~n60981 & n60982 ;
  assign n60984 = n60929 & n60974 ;
  assign n60985 = ~n60983 & ~n60984 ;
  assign n60986 = ~n60980 & n60985 ;
  assign n60987 = n60916 & ~n60986 ;
  assign n60995 = ~n60977 & ~n60987 ;
  assign n60996 = ~n60994 & n60995 ;
  assign n60997 = ~n60970 & n60996 ;
  assign n60998 = \u0_L7_reg[2]/NET0131  & n60997 ;
  assign n60999 = ~\u0_L7_reg[2]/NET0131  & ~n60997 ;
  assign n61000 = ~n60998 & ~n60999 ;
  assign n61007 = ~n60655 & ~n60681 ;
  assign n61008 = n60603 & ~n61007 ;
  assign n61009 = ~n60597 & ~n61008 ;
  assign n61010 = ~n60616 & n60636 ;
  assign n61011 = ~n60661 & ~n61010 ;
  assign n61012 = n60691 & n61011 ;
  assign n61013 = ~n61009 & ~n61012 ;
  assign n61004 = ~n60610 & ~n60648 ;
  assign n61005 = n60616 & ~n60689 ;
  assign n61006 = ~n61004 & n61005 ;
  assign n61014 = n60633 & ~n60698 ;
  assign n61015 = ~n61006 & n61014 ;
  assign n61016 = ~n61013 & n61015 ;
  assign n61023 = n60597 & ~n60622 ;
  assign n61026 = n60609 & n60625 ;
  assign n61027 = ~n61023 & n61026 ;
  assign n61024 = n60637 & ~n60648 ;
  assign n61025 = ~n61023 & n61024 ;
  assign n61021 = ~n60597 & ~n60603 ;
  assign n61022 = n60626 & n61021 ;
  assign n61028 = ~n60633 & ~n61022 ;
  assign n61029 = ~n61025 & n61028 ;
  assign n61030 = ~n61027 & n61029 ;
  assign n61017 = ~n60609 & ~n60669 ;
  assign n61018 = n60603 & n60626 ;
  assign n61019 = ~n60668 & ~n61018 ;
  assign n61020 = n60597 & ~n61019 ;
  assign n61031 = ~n61017 & ~n61020 ;
  assign n61032 = n61030 & n61031 ;
  assign n61033 = ~n61016 & ~n61032 ;
  assign n61001 = ~n60597 & n60609 ;
  assign n61002 = n60679 & n61001 ;
  assign n61003 = n60597 & n60642 ;
  assign n61034 = ~n61002 & ~n61003 ;
  assign n61035 = ~n61033 & n61034 ;
  assign n61036 = ~\u0_L7_reg[21]/NET0131  & ~n61035 ;
  assign n61037 = \u0_L7_reg[21]/NET0131  & n61035 ;
  assign n61038 = ~n61036 & ~n61037 ;
  assign n61039 = n60531 & n60533 ;
  assign n61040 = ~n60573 & ~n61039 ;
  assign n61041 = n60523 & ~n61040 ;
  assign n61042 = ~n60800 & ~n61041 ;
  assign n61043 = n60504 & ~n61042 ;
  assign n61044 = ~n60510 & ~n60550 ;
  assign n61045 = ~n60516 & n61044 ;
  assign n61046 = ~n60562 & ~n61045 ;
  assign n61047 = ~n60504 & ~n61046 ;
  assign n61048 = n60531 & n60570 ;
  assign n61049 = ~n60583 & ~n61048 ;
  assign n61050 = n60564 & n61049 ;
  assign n61051 = ~n61047 & n61050 ;
  assign n61052 = ~n61043 & n61051 ;
  assign n61053 = n60498 & ~n61052 ;
  assign n61058 = ~n60525 & n60531 ;
  assign n61059 = n61044 & ~n61058 ;
  assign n61060 = n60804 & ~n60816 ;
  assign n61061 = ~n61059 & n61060 ;
  assign n61062 = ~n60498 & ~n60817 ;
  assign n61063 = ~n61061 & n61062 ;
  assign n61055 = ~n60539 & ~n61041 ;
  assign n61056 = ~n60498 & ~n60504 ;
  assign n61057 = ~n61055 & n61056 ;
  assign n61054 = n60542 & n60808 ;
  assign n61064 = ~n60535 & ~n61054 ;
  assign n61065 = ~n61057 & n61064 ;
  assign n61066 = ~n61063 & n61065 ;
  assign n61067 = ~n61053 & n61066 ;
  assign n61068 = \u0_L7_reg[29]/NET0131  & ~n61067 ;
  assign n61069 = ~\u0_L7_reg[29]/NET0131  & n61067 ;
  assign n61070 = ~n61068 & ~n61069 ;
  assign n61129 = decrypt_pad & ~\u0_uk_K_r7_reg[28]/NET0131  ;
  assign n61130 = ~decrypt_pad & ~\u0_uk_K_r7_reg[35]/NET0131  ;
  assign n61131 = ~n61129 & ~n61130 ;
  assign n61132 = \u0_R7_reg[20]/NET0131  & ~n61131 ;
  assign n61133 = ~\u0_R7_reg[20]/NET0131  & n61131 ;
  assign n61134 = ~n61132 & ~n61133 ;
  assign n61099 = decrypt_pad & ~\u0_uk_K_r7_reg[44]/NET0131  ;
  assign n61100 = ~decrypt_pad & ~\u0_uk_K_r7_reg[51]/NET0131  ;
  assign n61101 = ~n61099 & ~n61100 ;
  assign n61102 = \u0_R7_reg[19]/NET0131  & ~n61101 ;
  assign n61103 = ~\u0_R7_reg[19]/NET0131  & n61101 ;
  assign n61104 = ~n61102 & ~n61103 ;
  assign n61091 = decrypt_pad & ~\u0_uk_K_r7_reg[8]/NET0131  ;
  assign n61092 = ~decrypt_pad & ~\u0_uk_K_r7_reg[15]/NET0131  ;
  assign n61093 = ~n61091 & ~n61092 ;
  assign n61094 = \u0_R7_reg[17]/NET0131  & ~n61093 ;
  assign n61095 = ~\u0_R7_reg[17]/NET0131  & n61093 ;
  assign n61096 = ~n61094 & ~n61095 ;
  assign n61077 = decrypt_pad & ~\u0_uk_K_r7_reg[45]/NET0131  ;
  assign n61078 = ~decrypt_pad & ~\u0_uk_K_r7_reg[52]/NET0131  ;
  assign n61079 = ~n61077 & ~n61078 ;
  assign n61080 = \u0_R7_reg[16]/NET0131  & ~n61079 ;
  assign n61081 = ~\u0_R7_reg[16]/NET0131  & n61079 ;
  assign n61082 = ~n61080 & ~n61081 ;
  assign n61084 = decrypt_pad & ~\u0_uk_K_r7_reg[29]/NET0131  ;
  assign n61085 = ~decrypt_pad & ~\u0_uk_K_r7_reg[36]/NET0131  ;
  assign n61086 = ~n61084 & ~n61085 ;
  assign n61087 = \u0_R7_reg[21]/NET0131  & ~n61086 ;
  assign n61088 = ~\u0_R7_reg[21]/NET0131  & n61086 ;
  assign n61089 = ~n61087 & ~n61088 ;
  assign n61136 = n61082 & ~n61089 ;
  assign n61137 = n61096 & n61136 ;
  assign n61071 = decrypt_pad & ~\u0_uk_K_r7_reg[2]/NET0131  ;
  assign n61072 = ~decrypt_pad & ~\u0_uk_K_r7_reg[9]/NET0131  ;
  assign n61073 = ~n61071 & ~n61072 ;
  assign n61074 = \u0_R7_reg[18]/NET0131  & ~n61073 ;
  assign n61075 = ~\u0_R7_reg[18]/NET0131  & n61073 ;
  assign n61076 = ~n61074 & ~n61075 ;
  assign n61097 = ~n61076 & n61096 ;
  assign n61098 = ~n61082 & n61097 ;
  assign n61083 = n61076 & n61082 ;
  assign n61138 = ~n61083 & n61089 ;
  assign n61139 = ~n61098 & n61138 ;
  assign n61140 = ~n61137 & ~n61139 ;
  assign n61141 = n61104 & ~n61140 ;
  assign n61105 = ~n61082 & ~n61089 ;
  assign n61106 = ~n61096 & n61105 ;
  assign n61118 = ~n61082 & n61089 ;
  assign n61144 = n61096 & n61118 ;
  assign n61145 = ~n61106 & ~n61144 ;
  assign n61146 = ~n61076 & ~n61104 ;
  assign n61147 = ~n61145 & n61146 ;
  assign n61115 = n61082 & n61089 ;
  assign n61116 = n61096 & n61115 ;
  assign n61148 = n61076 & ~n61104 ;
  assign n61149 = n61116 & n61148 ;
  assign n61142 = ~n61076 & n61115 ;
  assign n61143 = ~n61096 & n61142 ;
  assign n61150 = n61097 & n61136 ;
  assign n61151 = n61076 & ~n61096 ;
  assign n61152 = n61136 & n61151 ;
  assign n61153 = ~n61150 & ~n61152 ;
  assign n61154 = ~n61143 & n61153 ;
  assign n61155 = ~n61149 & n61154 ;
  assign n61156 = ~n61147 & n61155 ;
  assign n61157 = ~n61141 & n61156 ;
  assign n61158 = n61134 & ~n61157 ;
  assign n61090 = n61083 & n61089 ;
  assign n61107 = ~n61090 & n61104 ;
  assign n61108 = ~n61098 & ~n61106 ;
  assign n61109 = n61107 & n61108 ;
  assign n61119 = ~n61096 & n61118 ;
  assign n61110 = n61076 & n61096 ;
  assign n61111 = ~n61089 & n61110 ;
  assign n61120 = ~n61104 & ~n61111 ;
  assign n61121 = ~n61119 & n61120 ;
  assign n61112 = n61082 & ~n61096 ;
  assign n61113 = ~n61089 & n61112 ;
  assign n61114 = ~n61076 & n61113 ;
  assign n61117 = ~n61076 & n61116 ;
  assign n61122 = ~n61114 & ~n61117 ;
  assign n61123 = n61121 & n61122 ;
  assign n61124 = ~n61109 & ~n61123 ;
  assign n61125 = n61090 & ~n61096 ;
  assign n61126 = ~n61089 & n61098 ;
  assign n61127 = ~n61125 & ~n61126 ;
  assign n61128 = ~n61124 & n61127 ;
  assign n61135 = ~n61128 & ~n61134 ;
  assign n61159 = n61076 & n61106 ;
  assign n61160 = ~n61150 & ~n61159 ;
  assign n61161 = n61104 & ~n61160 ;
  assign n61162 = n61118 & n61151 ;
  assign n61163 = n61105 & n61110 ;
  assign n61164 = ~n61162 & ~n61163 ;
  assign n61165 = ~n61104 & ~n61164 ;
  assign n61166 = ~n61161 & ~n61165 ;
  assign n61167 = ~n61135 & n61166 ;
  assign n61168 = ~n61158 & n61167 ;
  assign n61169 = ~\u0_L7_reg[14]/NET0131  & ~n61168 ;
  assign n61170 = \u0_L7_reg[14]/NET0131  & n61168 ;
  assign n61171 = ~n61169 & ~n61170 ;
  assign n61175 = ~n60922 & n60972 ;
  assign n61176 = ~n60951 & ~n61175 ;
  assign n61177 = n60941 & n61176 ;
  assign n61181 = ~n60935 & n60981 ;
  assign n61182 = ~n60941 & ~n61181 ;
  assign n61179 = ~n60928 & n60949 ;
  assign n61180 = ~n60922 & n61179 ;
  assign n61178 = ~n60935 & n60950 ;
  assign n61183 = ~n60974 & ~n61178 ;
  assign n61184 = ~n61180 & n61183 ;
  assign n61185 = n61182 & n61184 ;
  assign n61186 = ~n61177 & ~n61185 ;
  assign n61173 = ~n60954 & ~n60972 ;
  assign n61174 = n60971 & ~n61173 ;
  assign n61172 = n60956 & n60960 ;
  assign n61187 = ~n60916 & ~n61172 ;
  assign n61188 = ~n61174 & n61187 ;
  assign n61189 = ~n61186 & n61188 ;
  assign n61195 = n60949 & n60957 ;
  assign n61194 = n60956 & n60981 ;
  assign n61196 = n60941 & ~n61194 ;
  assign n61197 = ~n61195 & n61196 ;
  assign n61198 = ~n61172 & n61176 ;
  assign n61199 = n61182 & n61198 ;
  assign n61200 = ~n61197 & ~n61199 ;
  assign n61190 = n60941 & n60949 ;
  assign n61191 = ~n60963 & ~n61190 ;
  assign n61192 = ~n60922 & ~n61191 ;
  assign n61193 = n60950 & n60971 ;
  assign n61201 = n60916 & ~n61193 ;
  assign n61202 = ~n61192 & n61201 ;
  assign n61203 = ~n61200 & n61202 ;
  assign n61204 = ~n61189 & ~n61203 ;
  assign n61205 = ~\u0_L7_reg[28]/NET0131  & n61204 ;
  assign n61206 = \u0_L7_reg[28]/NET0131  & ~n61204 ;
  assign n61207 = ~n61205 & ~n61206 ;
  assign n61219 = ~n60345 & ~n60353 ;
  assign n61218 = ~n60324 & n60345 ;
  assign n61220 = n60378 & ~n61218 ;
  assign n61221 = ~n61219 & n61220 ;
  assign n61216 = n60330 & n60339 ;
  assign n61217 = n60354 & n61216 ;
  assign n61222 = ~n60318 & ~n60359 ;
  assign n61223 = ~n61217 & n61222 ;
  assign n61224 = ~n61221 & n61223 ;
  assign n61208 = n60345 & n60375 ;
  assign n61209 = n60330 & n60358 ;
  assign n61210 = ~n61208 & ~n61209 ;
  assign n61211 = ~n60324 & ~n61210 ;
  assign n61212 = n60324 & n60330 ;
  assign n61213 = ~n60346 & ~n61212 ;
  assign n61214 = ~n60358 & n61213 ;
  assign n61215 = ~n60353 & ~n61214 ;
  assign n61225 = ~n61211 & ~n61215 ;
  assign n61226 = n61224 & n61225 ;
  assign n61227 = ~n60369 & ~n60386 ;
  assign n61228 = n60353 & ~n61227 ;
  assign n61229 = ~n60353 & n60379 ;
  assign n61233 = n60318 & ~n61229 ;
  assign n61230 = ~n60376 & ~n61216 ;
  assign n61231 = n61213 & ~n61230 ;
  assign n61232 = ~n61213 & n61230 ;
  assign n61234 = ~n61231 & ~n61232 ;
  assign n61235 = n61233 & n61234 ;
  assign n61236 = ~n61228 & n61235 ;
  assign n61237 = ~n61226 & ~n61236 ;
  assign n61238 = \u0_L7_reg[12]/NET0131  & n61237 ;
  assign n61239 = ~\u0_L7_reg[12]/NET0131  & ~n61237 ;
  assign n61240 = ~n61238 & ~n61239 ;
  assign n61257 = n60730 & n60746 ;
  assign n61252 = ~n60737 & n60842 ;
  assign n61258 = n60746 & n60763 ;
  assign n61259 = ~n61252 & ~n61258 ;
  assign n61260 = ~n61257 & ~n61259 ;
  assign n61262 = n60731 & ~n60754 ;
  assign n61263 = ~n60780 & n61262 ;
  assign n61261 = ~n60760 & n60784 ;
  assign n61264 = ~n60835 & ~n61261 ;
  assign n61265 = ~n61263 & n61264 ;
  assign n61266 = ~n61260 & n61265 ;
  assign n61267 = ~n60718 & ~n61266 ;
  assign n61246 = n60756 & ~n60771 ;
  assign n61247 = ~n60761 & ~n61246 ;
  assign n61248 = ~n60746 & ~n61247 ;
  assign n61241 = ~n60737 & n60753 ;
  assign n61242 = n60731 & n61241 ;
  assign n61243 = ~n60753 & n60759 ;
  assign n61244 = ~n61242 & ~n61243 ;
  assign n61245 = n60746 & ~n61244 ;
  assign n61249 = n60839 & ~n61245 ;
  assign n61250 = ~n61248 & n61249 ;
  assign n61251 = n60718 & ~n61250 ;
  assign n61253 = ~n60730 & n61252 ;
  assign n61254 = n60839 & ~n61253 ;
  assign n61255 = ~n60746 & ~n61254 ;
  assign n61256 = ~n60730 & n60758 ;
  assign n61268 = n60739 & n60757 ;
  assign n61269 = ~n61256 & ~n61268 ;
  assign n61270 = ~n61255 & n61269 ;
  assign n61271 = ~n61251 & n61270 ;
  assign n61272 = ~n61267 & n61271 ;
  assign n61273 = ~\u0_L7_reg[10]/NET0131  & ~n61272 ;
  assign n61274 = \u0_L7_reg[10]/NET0131  & n61272 ;
  assign n61275 = ~n61273 & ~n61274 ;
  assign n61279 = ~n61083 & ~n61089 ;
  assign n61280 = ~n61097 & n61279 ;
  assign n61278 = ~n61082 & ~n61096 ;
  assign n61281 = ~n61116 & ~n61278 ;
  assign n61282 = ~n61280 & n61281 ;
  assign n61283 = n61104 & ~n61282 ;
  assign n61284 = ~n61096 & n61115 ;
  assign n61285 = ~n61098 & ~n61284 ;
  assign n61286 = ~n61104 & ~n61285 ;
  assign n61276 = ~n61076 & n61089 ;
  assign n61277 = n61096 & n61276 ;
  assign n61287 = n61076 & n61137 ;
  assign n61288 = ~n61277 & ~n61287 ;
  assign n61289 = ~n61286 & n61288 ;
  assign n61290 = ~n61283 & n61289 ;
  assign n61291 = n61134 & ~n61290 ;
  assign n61299 = ~n61082 & n61110 ;
  assign n61300 = ~n61113 & ~n61299 ;
  assign n61301 = ~n61104 & ~n61300 ;
  assign n61303 = ~n61089 & n61104 ;
  assign n61304 = n61097 & n61303 ;
  assign n61298 = n61146 & n61278 ;
  assign n61302 = n61110 & n61118 ;
  assign n61305 = ~n61298 & ~n61302 ;
  assign n61306 = ~n61304 & n61305 ;
  assign n61307 = ~n61301 & n61306 ;
  assign n61308 = ~n61134 & ~n61307 ;
  assign n61292 = ~n61159 & ~n61287 ;
  assign n61293 = ~n61076 & n61118 ;
  assign n61294 = ~n61096 & n61293 ;
  assign n61295 = n61292 & ~n61294 ;
  assign n61296 = n61104 & ~n61295 ;
  assign n61297 = n61112 & n61148 ;
  assign n61309 = ~n61117 & ~n61297 ;
  assign n61310 = ~n61296 & n61309 ;
  assign n61311 = ~n61308 & n61310 ;
  assign n61312 = ~n61291 & n61311 ;
  assign n61313 = ~\u0_L7_reg[25]/NET0131  & ~n61312 ;
  assign n61314 = \u0_L7_reg[25]/NET0131  & n61312 ;
  assign n61315 = ~n61313 & ~n61314 ;
  assign n61320 = ~n60504 & ~n60801 ;
  assign n61316 = n60516 & ~n60550 ;
  assign n61317 = ~n60818 & ~n61316 ;
  assign n61318 = n60504 & ~n61317 ;
  assign n61319 = n60524 & n60531 ;
  assign n61321 = ~n60498 & ~n61319 ;
  assign n61322 = ~n61318 & n61321 ;
  assign n61323 = ~n61320 & n61322 ;
  assign n61324 = n60516 & n60540 ;
  assign n61328 = n60498 & ~n60557 ;
  assign n61329 = ~n61324 & n61328 ;
  assign n61330 = ~n60583 & n61329 ;
  assign n61325 = ~n60551 & ~n60572 ;
  assign n61326 = n60504 & ~n61325 ;
  assign n61327 = n60531 & ~n60801 ;
  assign n61331 = ~n61326 & ~n61327 ;
  assign n61332 = n61330 & n61331 ;
  assign n61333 = ~n61323 & ~n61332 ;
  assign n61334 = ~n60541 & ~n60585 ;
  assign n61335 = ~n61333 & n61334 ;
  assign n61336 = ~\u0_L7_reg[19]/NET0131  & ~n61335 ;
  assign n61337 = \u0_L7_reg[19]/NET0131  & n61335 ;
  assign n61338 = ~n61336 & ~n61337 ;
  assign n61354 = ~n60639 & ~n60655 ;
  assign n61355 = ~n60648 & ~n61354 ;
  assign n61356 = n60597 & ~n61355 ;
  assign n61357 = n60649 & n61001 ;
  assign n61358 = ~n60638 & ~n61022 ;
  assign n61359 = ~n61357 & n61358 ;
  assign n61360 = ~n61356 & n61359 ;
  assign n61361 = ~n60633 & ~n61360 ;
  assign n61339 = ~n60610 & ~n60665 ;
  assign n61340 = n60692 & n61339 ;
  assign n61341 = n60597 & ~n61340 ;
  assign n61342 = n60622 & ~n61339 ;
  assign n61343 = ~n60597 & ~n60642 ;
  assign n61344 = ~n61342 & n61343 ;
  assign n61345 = ~n61341 & ~n61344 ;
  assign n61346 = ~n60650 & ~n61010 ;
  assign n61347 = ~n60667 & n61346 ;
  assign n61348 = ~n61345 & n61347 ;
  assign n61349 = n60633 & ~n61348 ;
  assign n61350 = n60597 & n60616 ;
  assign n61351 = n60648 & n61350 ;
  assign n61352 = ~n60624 & ~n60640 ;
  assign n61353 = ~n60597 & ~n61352 ;
  assign n61362 = ~n61351 & ~n61353 ;
  assign n61363 = ~n61349 & n61362 ;
  assign n61364 = ~n61361 & n61363 ;
  assign n61365 = ~\u0_L7_reg[27]/NET0131  & ~n61364 ;
  assign n61366 = \u0_L7_reg[27]/NET0131  & n61364 ;
  assign n61367 = ~n61365 & ~n61366 ;
  assign n61371 = ~n60330 & ~n60354 ;
  assign n61372 = ~n61218 & n61371 ;
  assign n61368 = ~n60339 & n61212 ;
  assign n61369 = ~n60355 & ~n60378 ;
  assign n61370 = n60345 & ~n61369 ;
  assign n61373 = ~n61368 & ~n61370 ;
  assign n61374 = ~n61372 & n61373 ;
  assign n61375 = ~n60353 & ~n61374 ;
  assign n61379 = n60324 & n61370 ;
  assign n61380 = ~n61217 & ~n61379 ;
  assign n61376 = ~n60324 & n61369 ;
  assign n61377 = ~n60358 & n61376 ;
  assign n61378 = n60353 & n61377 ;
  assign n61381 = n60318 & ~n61378 ;
  assign n61382 = n61380 & n61381 ;
  assign n61383 = ~n61375 & n61382 ;
  assign n61384 = ~n60345 & n61216 ;
  assign n61385 = n60353 & ~n61384 ;
  assign n61386 = ~n61376 & n61385 ;
  assign n61387 = ~n61379 & n61386 ;
  assign n61388 = ~n60318 & ~n61387 ;
  assign n61389 = ~n61383 & ~n61388 ;
  assign n61390 = ~n60353 & ~n61380 ;
  assign n61391 = ~n60353 & n61377 ;
  assign n61392 = ~n60359 & ~n61391 ;
  assign n61393 = n60318 & ~n60353 ;
  assign n61394 = ~n61392 & ~n61393 ;
  assign n61395 = ~n61390 & ~n61394 ;
  assign n61396 = ~n61389 & n61395 ;
  assign n61397 = ~\u0_L7_reg[7]/NET0131  & ~n61396 ;
  assign n61398 = \u0_L7_reg[7]/NET0131  & n61396 ;
  assign n61399 = ~n61397 & ~n61398 ;
  assign n61412 = n61104 & ~n61114 ;
  assign n61413 = ~n61116 & n61412 ;
  assign n61414 = n61118 & ~n61151 ;
  assign n61415 = ~n61104 & ~n61284 ;
  assign n61416 = ~n61414 & n61415 ;
  assign n61417 = ~n61413 & ~n61416 ;
  assign n61418 = ~n61098 & n61292 ;
  assign n61419 = ~n61417 & n61418 ;
  assign n61420 = ~n61134 & ~n61419 ;
  assign n61400 = ~n61076 & n61106 ;
  assign n61401 = ~n61284 & ~n61400 ;
  assign n61402 = n61104 & ~n61401 ;
  assign n61403 = n61082 & n61146 ;
  assign n61404 = n61164 & ~n61403 ;
  assign n61405 = ~n61402 & n61404 ;
  assign n61406 = n61134 & ~n61405 ;
  assign n61407 = n61089 & n61098 ;
  assign n61408 = ~n61111 & ~n61162 ;
  assign n61409 = ~n61407 & n61408 ;
  assign n61410 = n61104 & ~n61409 ;
  assign n61411 = ~n61089 & n61297 ;
  assign n61421 = ~n61410 & ~n61411 ;
  assign n61422 = ~n61406 & n61421 ;
  assign n61423 = ~n61420 & n61422 ;
  assign n61424 = ~\u0_L7_reg[8]/NET0131  & ~n61423 ;
  assign n61425 = \u0_L7_reg[8]/NET0131  & n61423 ;
  assign n61426 = ~n61424 & ~n61425 ;
  assign n61428 = n60353 & ~n60387 ;
  assign n61427 = ~n60330 & n60358 ;
  assign n61429 = ~n61368 & ~n61427 ;
  assign n61430 = n61428 & n61429 ;
  assign n61431 = n60385 & ~n61369 ;
  assign n61432 = ~n60353 & ~n61208 ;
  assign n61433 = ~n61217 & n61432 ;
  assign n61434 = ~n61431 & n61433 ;
  assign n61435 = ~n61430 & ~n61434 ;
  assign n61436 = n60324 & ~n60339 ;
  assign n61437 = n60369 & n61436 ;
  assign n61438 = ~n61435 & ~n61437 ;
  assign n61439 = n60318 & ~n61438 ;
  assign n61446 = n60345 & ~n60355 ;
  assign n61447 = ~n60333 & n61446 ;
  assign n61448 = ~n60346 & ~n60358 ;
  assign n61449 = ~n60318 & ~n60363 ;
  assign n61450 = ~n61448 & n61449 ;
  assign n61451 = ~n61447 & ~n61450 ;
  assign n61452 = ~n60353 & ~n61451 ;
  assign n61440 = n60379 & ~n61393 ;
  assign n61441 = n60330 & ~n61219 ;
  assign n61442 = ~n61436 & n61441 ;
  assign n61443 = ~n60387 & n61442 ;
  assign n61444 = ~n60377 & ~n61443 ;
  assign n61445 = ~n60318 & ~n61444 ;
  assign n61453 = ~n61440 & ~n61445 ;
  assign n61454 = ~n61452 & n61453 ;
  assign n61455 = ~n61439 & n61454 ;
  assign n61456 = \u0_L7_reg[32]/NET0131  & n61455 ;
  assign n61457 = ~\u0_L7_reg[32]/NET0131  & ~n61455 ;
  assign n61458 = ~n61456 & ~n61457 ;
  assign n61459 = ~n60433 & ~n60878 ;
  assign n61460 = ~n60894 & ~n61459 ;
  assign n61461 = ~n60445 & ~n61460 ;
  assign n61462 = n60417 & ~n60457 ;
  assign n61463 = ~n60878 & n61462 ;
  assign n61464 = n61461 & ~n61463 ;
  assign n61466 = ~n60460 & ~n60880 ;
  assign n61467 = n60417 & n60458 ;
  assign n61465 = ~n60417 & n60894 ;
  assign n61468 = n60445 & ~n61465 ;
  assign n61469 = ~n61467 & n61468 ;
  assign n61470 = n61466 & n61469 ;
  assign n61471 = ~n61464 & ~n61470 ;
  assign n61472 = n60431 & n60449 ;
  assign n61473 = ~n61459 & n61472 ;
  assign n61474 = ~n60404 & ~n60883 ;
  assign n61475 = ~n61473 & n61474 ;
  assign n61476 = ~n61471 & n61475 ;
  assign n61479 = n60423 & n60435 ;
  assign n61480 = n60445 & ~n61479 ;
  assign n61481 = ~n60897 & n61480 ;
  assign n61482 = n61466 & n61481 ;
  assign n61483 = ~n60436 & ~n60481 ;
  assign n61484 = n61461 & n61483 ;
  assign n61485 = ~n61482 & ~n61484 ;
  assign n61477 = ~n60424 & ~n60481 ;
  assign n61478 = ~n60410 & ~n61477 ;
  assign n61486 = n60404 & ~n61478 ;
  assign n61487 = ~n61485 & n61486 ;
  assign n61488 = ~n61476 & ~n61487 ;
  assign n61489 = \u0_L7_reg[23]/NET0131  & n61488 ;
  assign n61490 = ~\u0_L7_reg[23]/NET0131  & ~n61488 ;
  assign n61491 = ~n61489 & ~n61490 ;
  assign n61492 = ~n60984 & ~n61172 ;
  assign n61493 = ~n60949 & n60956 ;
  assign n61494 = ~n61193 & ~n61493 ;
  assign n61495 = ~n60980 & n61494 ;
  assign n61496 = ~n60916 & ~n61495 ;
  assign n61497 = n61492 & ~n61496 ;
  assign n61498 = ~n60941 & ~n61497 ;
  assign n61504 = ~n60935 & n61173 ;
  assign n61503 = n60935 & ~n61180 ;
  assign n61505 = n60941 & ~n61503 ;
  assign n61506 = ~n61504 & n61505 ;
  assign n61501 = ~n60922 & ~n60942 ;
  assign n61502 = n60950 & n61501 ;
  assign n61499 = n60922 & ~n60956 ;
  assign n61500 = n61190 & n61499 ;
  assign n61507 = ~n60916 & ~n61500 ;
  assign n61508 = ~n61502 & n61507 ;
  assign n61509 = ~n61506 & n61508 ;
  assign n61510 = ~n60928 & n60971 ;
  assign n61511 = n60964 & ~n61510 ;
  assign n61512 = n60922 & n60950 ;
  assign n61513 = n60941 & ~n60979 ;
  assign n61514 = ~n61512 & n61513 ;
  assign n61515 = ~n61511 & ~n61514 ;
  assign n61516 = ~n60922 & n61493 ;
  assign n61517 = n60916 & n61492 ;
  assign n61518 = ~n61516 & n61517 ;
  assign n61519 = n60953 & n61518 ;
  assign n61520 = ~n61515 & n61519 ;
  assign n61521 = ~n61509 & ~n61520 ;
  assign n61522 = ~n61498 & ~n61521 ;
  assign n61523 = ~\u0_L7_reg[13]/NET0131  & n61522 ;
  assign n61524 = \u0_L7_reg[13]/NET0131  & ~n61522 ;
  assign n61525 = ~n61523 & ~n61524 ;
  assign n61560 = decrypt_pad & ~\u0_uk_K_r7_reg[11]/NET0131  ;
  assign n61561 = ~decrypt_pad & ~\u0_uk_K_r7_reg[18]/NET0131  ;
  assign n61562 = ~n61560 & ~n61561 ;
  assign n61563 = \u0_R7_reg[11]/P0001  & ~n61562 ;
  assign n61564 = ~\u0_R7_reg[11]/P0001  & n61562 ;
  assign n61565 = ~n61563 & ~n61564 ;
  assign n61552 = decrypt_pad & ~\u0_uk_K_r7_reg[26]/P0001  ;
  assign n61553 = ~decrypt_pad & ~\u0_uk_K_r7_reg[33]/NET0131  ;
  assign n61554 = ~n61552 & ~n61553 ;
  assign n61555 = \u0_R7_reg[12]/NET0131  & ~n61554 ;
  assign n61556 = ~\u0_R7_reg[12]/NET0131  & n61554 ;
  assign n61557 = ~n61555 & ~n61556 ;
  assign n61526 = decrypt_pad & ~\u0_uk_K_r7_reg[39]/NET0131  ;
  assign n61527 = ~decrypt_pad & ~\u0_uk_K_r7_reg[46]/NET0131  ;
  assign n61528 = ~n61526 & ~n61527 ;
  assign n61529 = \u0_R7_reg[13]/NET0131  & ~n61528 ;
  assign n61530 = ~\u0_R7_reg[13]/NET0131  & n61528 ;
  assign n61531 = ~n61529 & ~n61530 ;
  assign n61539 = decrypt_pad & ~\u0_uk_K_r7_reg[34]/NET0131  ;
  assign n61540 = ~decrypt_pad & ~\u0_uk_K_r7_reg[41]/NET0131  ;
  assign n61541 = ~n61539 & ~n61540 ;
  assign n61542 = \u0_R7_reg[9]/NET0131  & ~n61541 ;
  assign n61543 = ~\u0_R7_reg[9]/NET0131  & n61541 ;
  assign n61544 = ~n61542 & ~n61543 ;
  assign n61566 = n61531 & ~n61544 ;
  assign n61545 = decrypt_pad & ~\u0_uk_K_r7_reg[10]/NET0131  ;
  assign n61546 = ~decrypt_pad & ~\u0_uk_K_r7_reg[17]/NET0131  ;
  assign n61547 = ~n61545 & ~n61546 ;
  assign n61548 = \u0_R7_reg[10]/NET0131  & ~n61547 ;
  assign n61549 = ~\u0_R7_reg[10]/NET0131  & n61547 ;
  assign n61550 = ~n61548 & ~n61549 ;
  assign n61532 = decrypt_pad & ~\u0_uk_K_r7_reg[5]/NET0131  ;
  assign n61533 = ~decrypt_pad & ~\u0_uk_K_r7_reg[12]/NET0131  ;
  assign n61534 = ~n61532 & ~n61533 ;
  assign n61535 = \u0_R7_reg[8]/NET0131  & ~n61534 ;
  assign n61536 = ~\u0_R7_reg[8]/NET0131  & n61534 ;
  assign n61537 = ~n61535 & ~n61536 ;
  assign n61568 = n61531 & ~n61537 ;
  assign n61569 = n61550 & n61568 ;
  assign n61570 = ~n61531 & n61544 ;
  assign n61571 = n61537 & n61570 ;
  assign n61572 = ~n61569 & ~n61571 ;
  assign n61573 = ~n61566 & n61572 ;
  assign n61574 = n61557 & ~n61573 ;
  assign n61567 = n61550 & n61566 ;
  assign n61538 = ~n61531 & ~n61537 ;
  assign n61575 = n61538 & ~n61550 ;
  assign n61576 = ~n61544 & n61575 ;
  assign n61577 = ~n61567 & ~n61576 ;
  assign n61578 = ~n61574 & n61577 ;
  assign n61579 = n61565 & ~n61578 ;
  assign n61551 = n61544 & n61550 ;
  assign n61586 = ~n61544 & ~n61550 ;
  assign n61587 = ~n61551 & ~n61586 ;
  assign n61588 = n61531 & n61537 ;
  assign n61589 = ~n61538 & ~n61588 ;
  assign n61590 = ~n61537 & n61565 ;
  assign n61594 = n61589 & ~n61590 ;
  assign n61595 = ~n61587 & ~n61594 ;
  assign n61591 = n61544 & n61590 ;
  assign n61592 = n61587 & n61589 ;
  assign n61593 = ~n61591 & n61592 ;
  assign n61596 = ~n61557 & ~n61593 ;
  assign n61597 = ~n61595 & n61596 ;
  assign n61558 = n61551 & n61557 ;
  assign n61559 = n61538 & n61558 ;
  assign n61580 = n61544 & ~n61550 ;
  assign n61581 = ~n61537 & ~n61580 ;
  assign n61582 = n61557 & ~n61565 ;
  assign n61583 = ~n61566 & n61582 ;
  assign n61584 = ~n61570 & n61583 ;
  assign n61585 = ~n61581 & n61584 ;
  assign n61598 = ~n61559 & ~n61585 ;
  assign n61599 = ~n61597 & n61598 ;
  assign n61600 = ~n61579 & n61599 ;
  assign n61601 = ~\u0_L7_reg[6]/NET0131  & ~n61600 ;
  assign n61602 = \u0_L7_reg[6]/NET0131  & n61600 ;
  assign n61603 = ~n61601 & ~n61602 ;
  assign n61619 = ~n61565 & n61586 ;
  assign n61621 = ~n61568 & n61586 ;
  assign n61622 = ~n61565 & ~n61589 ;
  assign n61623 = ~n61621 & ~n61622 ;
  assign n61624 = ~n61619 & ~n61623 ;
  assign n61616 = n61537 & n61551 ;
  assign n61617 = ~n61569 & ~n61616 ;
  assign n61618 = n61565 & ~n61617 ;
  assign n61620 = n61568 & n61619 ;
  assign n61625 = n61537 & ~n61550 ;
  assign n61626 = ~n61531 & n61625 ;
  assign n61627 = ~n61544 & n61626 ;
  assign n61628 = ~n61620 & ~n61627 ;
  assign n61629 = ~n61618 & n61628 ;
  assign n61630 = ~n61624 & n61629 ;
  assign n61631 = n61557 & ~n61630 ;
  assign n61604 = n61537 & n61550 ;
  assign n61605 = ~n61544 & n61604 ;
  assign n61606 = ~n61531 & n61605 ;
  assign n61607 = n61538 & n61550 ;
  assign n61608 = ~n61550 & n61568 ;
  assign n61609 = ~n61607 & ~n61608 ;
  assign n61610 = n61538 & n61544 ;
  assign n61611 = ~n61605 & ~n61610 ;
  assign n61612 = n61609 & n61611 ;
  assign n61613 = n61565 & ~n61612 ;
  assign n61614 = ~n61606 & ~n61613 ;
  assign n61615 = ~n61557 & ~n61614 ;
  assign n61638 = n61586 & ~n61589 ;
  assign n61639 = n61572 & ~n61638 ;
  assign n61640 = ~n61557 & ~n61565 ;
  assign n61641 = ~n61639 & n61640 ;
  assign n61632 = n61544 & n61608 ;
  assign n61633 = ~n61627 & ~n61632 ;
  assign n61634 = n61565 & ~n61633 ;
  assign n61635 = n61550 & ~n61565 ;
  assign n61636 = n61544 & n61588 ;
  assign n61637 = n61635 & n61636 ;
  assign n61642 = ~n61634 & ~n61637 ;
  assign n61643 = ~n61641 & n61642 ;
  assign n61644 = ~n61615 & n61643 ;
  assign n61645 = ~n61631 & n61644 ;
  assign n61646 = ~\u0_L7_reg[24]/NET0131  & ~n61645 ;
  assign n61647 = \u0_L7_reg[24]/NET0131  & n61645 ;
  assign n61648 = ~n61646 & ~n61647 ;
  assign n61649 = ~n60446 & ~n60481 ;
  assign n61650 = ~n60890 & n61649 ;
  assign n61651 = n60404 & ~n61650 ;
  assign n61654 = ~n60435 & ~n60463 ;
  assign n61655 = n61459 & n61654 ;
  assign n61652 = ~n60432 & ~n60894 ;
  assign n61653 = ~n60404 & n61652 ;
  assign n61656 = ~n60445 & ~n61653 ;
  assign n61657 = ~n61655 & n61656 ;
  assign n61658 = ~n61651 & n61657 ;
  assign n61660 = ~n60895 & ~n61465 ;
  assign n61661 = n60410 & ~n61660 ;
  assign n61659 = n60411 & n61652 ;
  assign n61662 = n60445 & ~n60883 ;
  assign n61663 = ~n61659 & n61662 ;
  assign n61664 = ~n61661 & n61663 ;
  assign n61665 = ~n61658 & ~n61664 ;
  assign n61666 = ~n60404 & n60464 ;
  assign n61667 = ~n60449 & n61666 ;
  assign n61668 = ~n61665 & ~n61667 ;
  assign n61669 = ~\u0_L7_reg[9]/NET0131  & ~n61668 ;
  assign n61670 = \u0_L7_reg[9]/NET0131  & n61668 ;
  assign n61671 = ~n61669 & ~n61670 ;
  assign n61672 = n61565 & n61609 ;
  assign n61673 = ~n61627 & n61672 ;
  assign n61674 = ~n61565 & ~n61604 ;
  assign n61675 = ~n61610 & n61674 ;
  assign n61676 = ~n61673 & ~n61675 ;
  assign n61677 = n61557 & ~n61676 ;
  assign n61681 = ~n61531 & n61580 ;
  assign n61680 = ~n61570 & n61604 ;
  assign n61682 = n61565 & ~n61680 ;
  assign n61683 = ~n61681 & n61682 ;
  assign n61685 = ~n61570 & n61625 ;
  assign n61684 = n61544 & n61568 ;
  assign n61686 = ~n61565 & ~n61684 ;
  assign n61687 = ~n61685 & n61686 ;
  assign n61688 = ~n61683 & ~n61687 ;
  assign n61678 = ~n61544 & n61568 ;
  assign n61679 = n61550 & n61678 ;
  assign n61689 = ~n61557 & ~n61638 ;
  assign n61690 = ~n61679 & n61689 ;
  assign n61691 = ~n61688 & n61690 ;
  assign n61692 = ~n61677 & ~n61691 ;
  assign n61695 = n61531 & n61565 ;
  assign n61696 = n61605 & n61695 ;
  assign n61693 = n61558 & ~n61588 ;
  assign n61694 = n61570 & n61635 ;
  assign n61697 = ~n61693 & ~n61694 ;
  assign n61698 = ~n61696 & n61697 ;
  assign n61699 = ~n61692 & n61698 ;
  assign n61700 = \u0_L7_reg[30]/NET0131  & ~n61699 ;
  assign n61701 = ~\u0_L7_reg[30]/NET0131  & n61699 ;
  assign n61702 = ~n61700 & ~n61701 ;
  assign n61704 = n61096 & n61105 ;
  assign n61705 = ~n61142 & ~n61704 ;
  assign n61706 = n61104 & ~n61705 ;
  assign n61703 = ~n61104 & n61144 ;
  assign n61707 = n61134 & ~n61152 ;
  assign n61708 = ~n61117 & n61707 ;
  assign n61709 = ~n61703 & n61708 ;
  assign n61710 = ~n61706 & n61709 ;
  assign n61715 = ~n61137 & ~n61293 ;
  assign n61716 = n61104 & ~n61715 ;
  assign n61712 = ~n61112 & n61276 ;
  assign n61711 = n61104 & ~n61151 ;
  assign n61713 = ~n61136 & ~n61711 ;
  assign n61714 = ~n61712 & n61713 ;
  assign n61717 = ~n61134 & ~n61714 ;
  assign n61718 = ~n61716 & n61717 ;
  assign n61719 = ~n61710 & ~n61718 ;
  assign n61720 = ~n61162 & n61412 ;
  assign n61721 = ~n61104 & ~n61150 ;
  assign n61722 = ~n61125 & n61721 ;
  assign n61723 = ~n61400 & n61722 ;
  assign n61724 = ~n61720 & ~n61723 ;
  assign n61725 = ~n61719 & ~n61724 ;
  assign n61726 = ~\u0_L7_reg[3]/NET0131  & ~n61725 ;
  assign n61727 = \u0_L7_reg[3]/NET0131  & n61725 ;
  assign n61728 = ~n61726 & ~n61727 ;
  assign n61730 = ~n61544 & ~n61588 ;
  assign n61731 = ~n61636 & ~n61730 ;
  assign n61732 = ~n61538 & ~n61731 ;
  assign n61733 = ~n61531 & n61591 ;
  assign n61734 = ~n61732 & ~n61733 ;
  assign n61735 = ~n61550 & ~n61734 ;
  assign n61729 = n61550 & n61684 ;
  assign n61736 = ~n61607 & ~n61626 ;
  assign n61737 = ~n61565 & ~n61736 ;
  assign n61738 = ~n61729 & ~n61737 ;
  assign n61739 = ~n61735 & n61738 ;
  assign n61740 = n61557 & ~n61739 ;
  assign n61741 = ~n61575 & ~n61636 ;
  assign n61742 = ~n61678 & n61741 ;
  assign n61743 = ~n61565 & ~n61742 ;
  assign n61744 = ~n61538 & n61565 ;
  assign n61745 = n61731 & n61744 ;
  assign n61746 = ~n61576 & ~n61745 ;
  assign n61747 = ~n61743 & n61746 ;
  assign n61748 = ~n61557 & ~n61747 ;
  assign n61749 = ~n61544 & n61607 ;
  assign n61750 = n61550 & n61571 ;
  assign n61751 = ~n61749 & ~n61750 ;
  assign n61752 = n61565 & ~n61751 ;
  assign n61753 = ~n61565 & n61605 ;
  assign n61754 = ~n61752 & ~n61753 ;
  assign n61755 = ~n61748 & n61754 ;
  assign n61756 = ~n61740 & n61755 ;
  assign n61757 = ~\u0_L7_reg[16]/NET0131  & ~n61756 ;
  assign n61758 = \u0_L7_reg[16]/NET0131  & n61756 ;
  assign n61759 = ~n61757 & ~n61758 ;
  assign n61772 = ~n60971 & ~n60982 ;
  assign n61774 = n60954 & ~n61772 ;
  assign n61768 = ~n60949 & ~n60988 ;
  assign n61773 = n61768 & n61772 ;
  assign n61775 = ~n60979 & ~n61172 ;
  assign n61776 = ~n61773 & n61775 ;
  assign n61777 = ~n61774 & n61776 ;
  assign n61778 = ~n60916 & ~n61777 ;
  assign n61765 = n60941 & n60958 ;
  assign n61766 = ~n60973 & ~n61765 ;
  assign n61767 = n60916 & ~n61766 ;
  assign n61760 = ~n60929 & ~n60978 ;
  assign n61761 = n60916 & n60949 ;
  assign n61762 = ~n61760 & n61761 ;
  assign n61763 = ~n60951 & ~n61762 ;
  assign n61764 = ~n60941 & ~n61763 ;
  assign n61769 = ~n60929 & n60941 ;
  assign n61770 = ~n61179 & n61769 ;
  assign n61771 = ~n61768 & n61770 ;
  assign n61779 = ~n61764 & ~n61771 ;
  assign n61780 = ~n61767 & n61779 ;
  assign n61781 = ~n61778 & n61780 ;
  assign n61782 = \u0_L7_reg[18]/NET0131  & n61781 ;
  assign n61783 = ~\u0_L7_reg[18]/NET0131  & ~n61781 ;
  assign n61784 = ~n61782 & ~n61783 ;
  assign n61819 = decrypt_pad & ~\u0_uk_K_r6_reg[54]/NET0131  ;
  assign n61820 = ~decrypt_pad & ~\u0_uk_K_r6_reg[47]/NET0131  ;
  assign n61821 = ~n61819 & ~n61820 ;
  assign n61822 = \u0_R6_reg[4]/NET0131  & ~n61821 ;
  assign n61823 = ~\u0_R6_reg[4]/NET0131  & n61821 ;
  assign n61824 = ~n61822 & ~n61823 ;
  assign n61798 = decrypt_pad & ~\u0_uk_K_r6_reg[19]/NET0131  ;
  assign n61799 = ~decrypt_pad & ~\u0_uk_K_r6_reg[12]/NET0131  ;
  assign n61800 = ~n61798 & ~n61799 ;
  assign n61801 = \u0_R6_reg[3]/NET0131  & ~n61800 ;
  assign n61802 = ~\u0_R6_reg[3]/NET0131  & n61800 ;
  assign n61803 = ~n61801 & ~n61802 ;
  assign n61785 = decrypt_pad & ~\u0_uk_K_r6_reg[25]/NET0131  ;
  assign n61786 = ~decrypt_pad & ~\u0_uk_K_r6_reg[18]/NET0131  ;
  assign n61787 = ~n61785 & ~n61786 ;
  assign n61788 = \u0_R6_reg[5]/NET0131  & ~n61787 ;
  assign n61789 = ~\u0_R6_reg[5]/NET0131  & n61787 ;
  assign n61790 = ~n61788 & ~n61789 ;
  assign n61791 = decrypt_pad & ~\u0_uk_K_r6_reg[27]/NET0131  ;
  assign n61792 = ~decrypt_pad & ~\u0_uk_K_r6_reg[20]/NET0131  ;
  assign n61793 = ~n61791 & ~n61792 ;
  assign n61794 = \u0_R6_reg[1]/NET0131  & ~n61793 ;
  assign n61795 = ~\u0_R6_reg[1]/NET0131  & n61793 ;
  assign n61796 = ~n61794 & ~n61795 ;
  assign n61827 = n61790 & ~n61796 ;
  assign n61804 = decrypt_pad & ~\u0_uk_K_r6_reg[6]/NET0131  ;
  assign n61805 = ~decrypt_pad & ~\u0_uk_K_r6_reg[24]/NET0131  ;
  assign n61806 = ~n61804 & ~n61805 ;
  assign n61807 = \u0_R6_reg[32]/NET0131  & ~n61806 ;
  assign n61808 = ~\u0_R6_reg[32]/NET0131  & n61806 ;
  assign n61809 = ~n61807 & ~n61808 ;
  assign n61811 = decrypt_pad & ~\u0_uk_K_r6_reg[10]/NET0131  ;
  assign n61812 = ~decrypt_pad & ~\u0_uk_K_r6_reg[3]/NET0131  ;
  assign n61813 = ~n61811 & ~n61812 ;
  assign n61814 = \u0_R6_reg[2]/NET0131  & ~n61813 ;
  assign n61815 = ~\u0_R6_reg[2]/NET0131  & n61813 ;
  assign n61816 = ~n61814 & ~n61815 ;
  assign n61828 = ~n61809 & n61816 ;
  assign n61829 = ~n61790 & n61828 ;
  assign n61830 = ~n61827 & ~n61829 ;
  assign n61831 = n61803 & ~n61830 ;
  assign n61836 = n61796 & ~n61809 ;
  assign n61837 = n61796 & ~n61803 ;
  assign n61838 = ~n61828 & ~n61837 ;
  assign n61839 = ~n61836 & ~n61838 ;
  assign n61797 = ~n61790 & ~n61796 ;
  assign n61825 = n61809 & ~n61816 ;
  assign n61826 = n61797 & n61825 ;
  assign n61832 = n61790 & ~n61809 ;
  assign n61833 = n61803 & ~n61816 ;
  assign n61834 = n61796 & ~n61833 ;
  assign n61835 = n61832 & ~n61834 ;
  assign n61840 = ~n61826 & ~n61835 ;
  assign n61841 = ~n61839 & n61840 ;
  assign n61842 = ~n61831 & n61841 ;
  assign n61843 = n61824 & ~n61842 ;
  assign n61845 = n61790 & n61809 ;
  assign n61859 = ~n61837 & n61845 ;
  assign n61860 = ~n61790 & n61836 ;
  assign n61861 = ~n61859 & ~n61860 ;
  assign n61862 = ~n61816 & ~n61861 ;
  assign n61863 = ~n61790 & ~n61809 ;
  assign n61864 = ~n61845 & ~n61863 ;
  assign n61865 = n61796 & n61864 ;
  assign n61866 = n61803 & n61816 ;
  assign n61867 = n61865 & n61866 ;
  assign n61868 = ~n61862 & ~n61867 ;
  assign n61869 = ~n61824 & ~n61868 ;
  assign n61851 = ~n61825 & ~n61828 ;
  assign n61850 = n61796 & n61816 ;
  assign n61852 = ~n61824 & ~n61827 ;
  assign n61853 = ~n61850 & n61852 ;
  assign n61854 = n61851 & n61853 ;
  assign n61846 = n61796 & n61845 ;
  assign n61847 = n61816 & n61846 ;
  assign n61844 = n61827 & n61828 ;
  assign n61848 = n61796 & ~n61816 ;
  assign n61849 = ~n61790 & n61848 ;
  assign n61855 = ~n61844 & ~n61849 ;
  assign n61856 = ~n61847 & n61855 ;
  assign n61857 = ~n61854 & n61856 ;
  assign n61858 = ~n61803 & ~n61857 ;
  assign n61810 = n61803 & ~n61809 ;
  assign n61817 = n61810 & n61816 ;
  assign n61818 = n61797 & n61817 ;
  assign n61870 = ~n61796 & n61809 ;
  assign n61871 = n61833 & n61870 ;
  assign n61872 = ~n61818 & ~n61871 ;
  assign n61873 = ~n61858 & n61872 ;
  assign n61874 = ~n61869 & n61873 ;
  assign n61875 = ~n61843 & n61874 ;
  assign n61876 = ~\u0_L6_reg[31]/NET0131  & ~n61875 ;
  assign n61877 = \u0_L6_reg[31]/NET0131  & n61875 ;
  assign n61878 = ~n61876 & ~n61877 ;
  assign n61879 = decrypt_pad & ~\u0_uk_K_r6_reg[23]/P0001  ;
  assign n61880 = ~decrypt_pad & ~\u0_uk_K_r6_reg[16]/NET0131  ;
  assign n61881 = ~n61879 & ~n61880 ;
  assign n61882 = \u0_R6_reg[24]/NET0131  & ~n61881 ;
  assign n61883 = ~\u0_R6_reg[24]/NET0131  & n61881 ;
  assign n61884 = ~n61882 & ~n61883 ;
  assign n61913 = decrypt_pad & ~\u0_uk_K_r6_reg[21]/NET0131  ;
  assign n61914 = ~decrypt_pad & ~\u0_uk_K_r6_reg[14]/NET0131  ;
  assign n61915 = ~n61913 & ~n61914 ;
  assign n61916 = \u0_R6_reg[23]/NET0131  & ~n61915 ;
  assign n61917 = ~\u0_R6_reg[23]/NET0131  & n61915 ;
  assign n61918 = ~n61916 & ~n61917 ;
  assign n61885 = decrypt_pad & ~\u0_uk_K_r6_reg[45]/NET0131  ;
  assign n61886 = ~decrypt_pad & ~\u0_uk_K_r6_reg[38]/NET0131  ;
  assign n61887 = ~n61885 & ~n61886 ;
  assign n61888 = \u0_R6_reg[21]/NET0131  & ~n61887 ;
  assign n61889 = ~\u0_R6_reg[21]/NET0131  & n61887 ;
  assign n61890 = ~n61888 & ~n61889 ;
  assign n61891 = decrypt_pad & ~\u0_uk_K_r6_reg[2]/NET0131  ;
  assign n61892 = ~decrypt_pad & ~\u0_uk_K_r6_reg[50]/NET0131  ;
  assign n61893 = ~n61891 & ~n61892 ;
  assign n61894 = \u0_R6_reg[20]/NET0131  & ~n61893 ;
  assign n61895 = ~\u0_R6_reg[20]/NET0131  & n61893 ;
  assign n61896 = ~n61894 & ~n61895 ;
  assign n61897 = ~n61890 & n61896 ;
  assign n61898 = decrypt_pad & ~\u0_uk_K_r6_reg[8]/NET0131  ;
  assign n61899 = ~decrypt_pad & ~\u0_uk_K_r6_reg[1]/NET0131  ;
  assign n61900 = ~n61898 & ~n61899 ;
  assign n61901 = \u0_R6_reg[22]/NET0131  & ~n61900 ;
  assign n61902 = ~\u0_R6_reg[22]/NET0131  & n61900 ;
  assign n61903 = ~n61901 & ~n61902 ;
  assign n61905 = decrypt_pad & ~\u0_uk_K_r6_reg[42]/NET0131  ;
  assign n61906 = ~decrypt_pad & ~\u0_uk_K_r6_reg[35]/NET0131  ;
  assign n61907 = ~n61905 & ~n61906 ;
  assign n61908 = \u0_R6_reg[25]/NET0131  & ~n61907 ;
  assign n61909 = ~\u0_R6_reg[25]/NET0131  & n61907 ;
  assign n61910 = ~n61908 & ~n61909 ;
  assign n61952 = ~n61903 & ~n61910 ;
  assign n61953 = n61897 & n61952 ;
  assign n61926 = n61890 & ~n61896 ;
  assign n61927 = n61903 & n61926 ;
  assign n61941 = n61896 & n61910 ;
  assign n61951 = n61890 & n61941 ;
  assign n61954 = ~n61927 & ~n61951 ;
  assign n61955 = ~n61953 & n61954 ;
  assign n61956 = n61918 & ~n61955 ;
  assign n61919 = ~n61903 & ~n61918 ;
  assign n61957 = n61919 & n61941 ;
  assign n61958 = ~n61890 & n61957 ;
  assign n61920 = n61890 & ~n61903 ;
  assign n61959 = n61903 & ~n61926 ;
  assign n61960 = ~n61920 & ~n61959 ;
  assign n61961 = ~n61918 & ~n61941 ;
  assign n61962 = ~n61952 & n61961 ;
  assign n61963 = ~n61960 & n61962 ;
  assign n61964 = ~n61958 & ~n61963 ;
  assign n61965 = ~n61956 & n61964 ;
  assign n61966 = n61884 & ~n61965 ;
  assign n61923 = ~n61890 & ~n61896 ;
  assign n61924 = n61910 & n61923 ;
  assign n61925 = n61918 & n61924 ;
  assign n61904 = n61897 & n61903 ;
  assign n61911 = n61904 & n61910 ;
  assign n61912 = n61896 & ~n61910 ;
  assign n61921 = ~n61919 & ~n61920 ;
  assign n61922 = n61912 & ~n61921 ;
  assign n61934 = ~n61911 & ~n61922 ;
  assign n61935 = ~n61925 & n61934 ;
  assign n61928 = n61896 & n61920 ;
  assign n61929 = ~n61927 & ~n61928 ;
  assign n61930 = ~n61918 & ~n61929 ;
  assign n61931 = ~n61896 & ~n61903 ;
  assign n61932 = ~n61904 & ~n61931 ;
  assign n61933 = n61918 & ~n61932 ;
  assign n61936 = ~n61930 & ~n61933 ;
  assign n61937 = n61935 & n61936 ;
  assign n61938 = ~n61884 & ~n61937 ;
  assign n61945 = n61890 & n61912 ;
  assign n61946 = ~n61918 & n61945 ;
  assign n61947 = ~n61925 & ~n61946 ;
  assign n61948 = ~n61903 & ~n61947 ;
  assign n61942 = ~n61920 & ~n61941 ;
  assign n61939 = ~n61896 & ~n61910 ;
  assign n61940 = ~n61903 & ~n61939 ;
  assign n61943 = n61918 & ~n61940 ;
  assign n61944 = ~n61942 & n61943 ;
  assign n61949 = ~n61890 & n61939 ;
  assign n61950 = n61919 & n61949 ;
  assign n61967 = ~n61944 & ~n61950 ;
  assign n61968 = ~n61948 & n61967 ;
  assign n61969 = ~n61938 & n61968 ;
  assign n61970 = ~n61966 & n61969 ;
  assign n61971 = ~\u0_L6_reg[11]/NET0131  & n61970 ;
  assign n61972 = \u0_L6_reg[11]/NET0131  & ~n61970 ;
  assign n61973 = ~n61971 & ~n61972 ;
  assign n61974 = decrypt_pad & ~\u0_uk_K_r6_reg[38]/NET0131  ;
  assign n61975 = ~decrypt_pad & ~\u0_uk_K_r6_reg[31]/NET0131  ;
  assign n61976 = ~n61974 & ~n61975 ;
  assign n61977 = \u0_R6_reg[26]/NET0131  & ~n61976 ;
  assign n61978 = ~\u0_R6_reg[26]/NET0131  & n61976 ;
  assign n61979 = ~n61977 & ~n61978 ;
  assign n61980 = decrypt_pad & ~\u0_uk_K_r6_reg[49]/NET0131  ;
  assign n61981 = ~decrypt_pad & ~\u0_uk_K_r6_reg[42]/NET0131  ;
  assign n61982 = ~n61980 & ~n61981 ;
  assign n61983 = \u0_R6_reg[25]/NET0131  & ~n61982 ;
  assign n61984 = ~\u0_R6_reg[25]/NET0131  & n61982 ;
  assign n61985 = ~n61983 & ~n61984 ;
  assign n61986 = n61979 & ~n61985 ;
  assign n61987 = decrypt_pad & ~\u0_uk_K_r6_reg[14]/NET0131  ;
  assign n61988 = ~decrypt_pad & ~\u0_uk_K_r6_reg[7]/NET0131  ;
  assign n61989 = ~n61987 & ~n61988 ;
  assign n61990 = \u0_R6_reg[24]/NET0131  & ~n61989 ;
  assign n61991 = ~\u0_R6_reg[24]/NET0131  & n61989 ;
  assign n61992 = ~n61990 & ~n61991 ;
  assign n61993 = decrypt_pad & ~\u0_uk_K_r6_reg[22]/NET0131  ;
  assign n61994 = ~decrypt_pad & ~\u0_uk_K_r6_reg[15]/NET0131  ;
  assign n61995 = ~n61993 & ~n61994 ;
  assign n61996 = \u0_R6_reg[29]/NET0131  & ~n61995 ;
  assign n61997 = ~\u0_R6_reg[29]/NET0131  & n61995 ;
  assign n61998 = ~n61996 & ~n61997 ;
  assign n61999 = ~n61992 & n61998 ;
  assign n62000 = n61986 & n61999 ;
  assign n62001 = n61979 & n61985 ;
  assign n62002 = ~n61992 & n62001 ;
  assign n62003 = ~n61998 & n62002 ;
  assign n62004 = ~n62000 & ~n62003 ;
  assign n62005 = ~n61985 & ~n61998 ;
  assign n62006 = n61985 & n61998 ;
  assign n62007 = ~n61979 & n62006 ;
  assign n62008 = ~n61986 & ~n62007 ;
  assign n62009 = decrypt_pad & ~\u0_uk_K_r6_reg[30]/P0001  ;
  assign n62010 = ~decrypt_pad & ~\u0_uk_K_r6_reg[23]/P0001  ;
  assign n62011 = ~n62009 & ~n62010 ;
  assign n62012 = \u0_R6_reg[28]/NET0131  & ~n62011 ;
  assign n62013 = ~\u0_R6_reg[28]/NET0131  & n62011 ;
  assign n62014 = ~n62012 & ~n62013 ;
  assign n62015 = ~n62008 & n62014 ;
  assign n62016 = ~n62005 & ~n62015 ;
  assign n62017 = n61992 & ~n62016 ;
  assign n62018 = n62004 & ~n62017 ;
  assign n62019 = decrypt_pad & ~\u0_uk_K_r6_reg[43]/NET0131  ;
  assign n62020 = ~decrypt_pad & ~\u0_uk_K_r6_reg[36]/NET0131  ;
  assign n62021 = ~n62019 & ~n62020 ;
  assign n62022 = \u0_R6_reg[27]/NET0131  & ~n62021 ;
  assign n62023 = ~\u0_R6_reg[27]/NET0131  & n62021 ;
  assign n62024 = ~n62022 & ~n62023 ;
  assign n62025 = ~n62018 & n62024 ;
  assign n62026 = ~n61985 & n62024 ;
  assign n62027 = ~n61979 & n62026 ;
  assign n62028 = ~n61979 & n61998 ;
  assign n62029 = ~n61986 & ~n62024 ;
  assign n62030 = ~n62028 & n62029 ;
  assign n62031 = ~n62027 & ~n62030 ;
  assign n62032 = n61992 & ~n62031 ;
  assign n62033 = ~n61992 & n62005 ;
  assign n62034 = n61979 & n62033 ;
  assign n62035 = ~n62024 & n62034 ;
  assign n62036 = ~n61979 & ~n61992 ;
  assign n62037 = n61979 & n61992 ;
  assign n62038 = ~n62036 & ~n62037 ;
  assign n62039 = n61998 & ~n62026 ;
  assign n62040 = ~n62038 & n62039 ;
  assign n62041 = ~n62035 & ~n62040 ;
  assign n62042 = ~n62032 & n62041 ;
  assign n62043 = ~n62014 & ~n62042 ;
  assign n62047 = ~n61985 & n61992 ;
  assign n62048 = n62028 & n62047 ;
  assign n62049 = n61985 & n61999 ;
  assign n62050 = ~n62048 & ~n62049 ;
  assign n62051 = ~n62024 & ~n62050 ;
  assign n62052 = n62005 & n62036 ;
  assign n62053 = ~n62000 & ~n62052 ;
  assign n62054 = ~n62051 & n62053 ;
  assign n62055 = n62014 & ~n62054 ;
  assign n62044 = n61985 & ~n62024 ;
  assign n62045 = ~n62038 & n62044 ;
  assign n62046 = ~n61998 & n62027 ;
  assign n62056 = ~n62045 & ~n62046 ;
  assign n62057 = ~n62055 & n62056 ;
  assign n62058 = ~n62043 & n62057 ;
  assign n62059 = ~n62025 & n62058 ;
  assign n62060 = ~\u0_L6_reg[22]/NET0131  & ~n62059 ;
  assign n62061 = \u0_L6_reg[22]/NET0131  & n62059 ;
  assign n62062 = ~n62060 & ~n62061 ;
  assign n62063 = decrypt_pad & ~\u0_uk_K_r6_reg[48]/NET0131  ;
  assign n62064 = ~decrypt_pad & ~\u0_uk_K_r6_reg[41]/NET0131  ;
  assign n62065 = ~n62063 & ~n62064 ;
  assign n62066 = \u0_R6_reg[15]/NET0131  & ~n62065 ;
  assign n62067 = ~\u0_R6_reg[15]/NET0131  & n62065 ;
  assign n62068 = ~n62066 & ~n62067 ;
  assign n62089 = decrypt_pad & ~\u0_uk_K_r6_reg[39]/NET0131  ;
  assign n62090 = ~decrypt_pad & ~\u0_uk_K_r6_reg[32]/NET0131  ;
  assign n62091 = ~n62089 & ~n62090 ;
  assign n62092 = \u0_R6_reg[13]/NET0131  & ~n62091 ;
  assign n62093 = ~\u0_R6_reg[13]/NET0131  & n62091 ;
  assign n62094 = ~n62092 & ~n62093 ;
  assign n62076 = decrypt_pad & ~\u0_uk_K_r6_reg[20]/NET0131  ;
  assign n62077 = ~decrypt_pad & ~\u0_uk_K_r6_reg[13]/NET0131  ;
  assign n62078 = ~n62076 & ~n62077 ;
  assign n62079 = \u0_R6_reg[12]/NET0131  & ~n62078 ;
  assign n62080 = ~\u0_R6_reg[12]/NET0131  & n62078 ;
  assign n62081 = ~n62079 & ~n62080 ;
  assign n62069 = decrypt_pad & ~\u0_uk_K_r6_reg[40]/NET0131  ;
  assign n62070 = ~decrypt_pad & ~\u0_uk_K_r6_reg[33]/NET0131  ;
  assign n62071 = ~n62069 & ~n62070 ;
  assign n62072 = \u0_R6_reg[14]/NET0131  & ~n62071 ;
  assign n62073 = ~\u0_R6_reg[14]/NET0131  & n62071 ;
  assign n62074 = ~n62072 & ~n62073 ;
  assign n62082 = decrypt_pad & ~\u0_uk_K_r6_reg[4]/NET0131  ;
  assign n62083 = ~decrypt_pad & ~\u0_uk_K_r6_reg[54]/NET0131  ;
  assign n62084 = ~n62082 & ~n62083 ;
  assign n62085 = \u0_R6_reg[17]/NET0131  & ~n62084 ;
  assign n62086 = ~\u0_R6_reg[17]/NET0131  & n62084 ;
  assign n62087 = ~n62085 & ~n62086 ;
  assign n62107 = ~n62074 & ~n62087 ;
  assign n62108 = ~n62081 & n62107 ;
  assign n62109 = ~n62094 & n62108 ;
  assign n62110 = ~n62068 & ~n62109 ;
  assign n62111 = ~n62087 & ~n62094 ;
  assign n62112 = ~n62081 & n62111 ;
  assign n62113 = n62081 & n62087 ;
  assign n62114 = n62094 & n62113 ;
  assign n62115 = ~n62112 & ~n62114 ;
  assign n62116 = ~n62110 & ~n62115 ;
  assign n62117 = ~n62081 & n62094 ;
  assign n62118 = ~n62087 & n62117 ;
  assign n62119 = n62074 & n62118 ;
  assign n62120 = decrypt_pad & ~\u0_uk_K_r6_reg[24]/NET0131  ;
  assign n62121 = ~decrypt_pad & ~\u0_uk_K_r6_reg[17]/NET0131  ;
  assign n62122 = ~n62120 & ~n62121 ;
  assign n62123 = \u0_R6_reg[16]/NET0131  & ~n62122 ;
  assign n62124 = ~\u0_R6_reg[16]/NET0131  & n62122 ;
  assign n62125 = ~n62123 & ~n62124 ;
  assign n62126 = ~n62119 & ~n62125 ;
  assign n62097 = n62087 & ~n62094 ;
  assign n62100 = n62081 & ~n62087 ;
  assign n62101 = n62074 & n62100 ;
  assign n62102 = ~n62097 & ~n62101 ;
  assign n62103 = ~n62068 & ~n62102 ;
  assign n62098 = ~n62074 & n62097 ;
  assign n62099 = n62081 & n62098 ;
  assign n62104 = n62068 & n62074 ;
  assign n62105 = n62094 & n62104 ;
  assign n62106 = ~n62081 & n62105 ;
  assign n62127 = ~n62099 & ~n62106 ;
  assign n62128 = ~n62103 & n62127 ;
  assign n62129 = n62126 & n62128 ;
  assign n62130 = ~n62116 & n62129 ;
  assign n62088 = ~n62081 & n62087 ;
  assign n62131 = n62068 & n62088 ;
  assign n62132 = ~n62094 & n62131 ;
  assign n62133 = ~n62074 & n62087 ;
  assign n62134 = n62117 & n62133 ;
  assign n62144 = n62125 & ~n62134 ;
  assign n62145 = ~n62132 & n62144 ;
  assign n62135 = n62074 & ~n62081 ;
  assign n62136 = ~n62068 & n62111 ;
  assign n62137 = n62135 & n62136 ;
  assign n62075 = ~n62068 & ~n62074 ;
  assign n62138 = n62081 & ~n62094 ;
  assign n62139 = ~n62117 & ~n62138 ;
  assign n62140 = n62075 & ~n62139 ;
  assign n62146 = ~n62137 & ~n62140 ;
  assign n62141 = n62074 & n62114 ;
  assign n62142 = n62094 & n62100 ;
  assign n62143 = n62068 & n62142 ;
  assign n62147 = ~n62141 & ~n62143 ;
  assign n62148 = n62146 & n62147 ;
  assign n62149 = n62145 & n62148 ;
  assign n62150 = ~n62130 & ~n62149 ;
  assign n62095 = n62088 & n62094 ;
  assign n62096 = n62075 & n62095 ;
  assign n62153 = ~n62094 & n62101 ;
  assign n62151 = ~n62074 & n62094 ;
  assign n62152 = n62100 & n62151 ;
  assign n62154 = ~n62109 & ~n62152 ;
  assign n62155 = ~n62153 & n62154 ;
  assign n62156 = n62068 & ~n62155 ;
  assign n62157 = ~n62096 & ~n62156 ;
  assign n62158 = ~n62150 & n62157 ;
  assign n62159 = ~\u0_L6_reg[20]/NET0131  & ~n62158 ;
  assign n62160 = \u0_L6_reg[20]/NET0131  & n62158 ;
  assign n62161 = ~n62159 & ~n62160 ;
  assign n62205 = decrypt_pad & ~\u0_uk_K_r6_reg[44]/NET0131  ;
  assign n62206 = ~decrypt_pad & ~\u0_uk_K_r6_reg[37]/NET0131  ;
  assign n62207 = ~n62205 & ~n62206 ;
  assign n62208 = \u0_R6_reg[31]/P0001  & ~n62207 ;
  assign n62209 = ~\u0_R6_reg[31]/P0001  & n62207 ;
  assign n62210 = ~n62208 & ~n62209 ;
  assign n62168 = decrypt_pad & ~\u0_uk_K_r6_reg[1]/NET0131  ;
  assign n62169 = ~decrypt_pad & ~\u0_uk_K_r6_reg[49]/NET0131  ;
  assign n62170 = ~n62168 & ~n62169 ;
  assign n62171 = \u0_R6_reg[30]/NET0131  & ~n62170 ;
  assign n62172 = ~\u0_R6_reg[30]/NET0131  & n62170 ;
  assign n62173 = ~n62171 & ~n62172 ;
  assign n62174 = decrypt_pad & ~\u0_uk_K_r6_reg[28]/NET0131  ;
  assign n62175 = ~decrypt_pad & ~\u0_uk_K_r6_reg[21]/NET0131  ;
  assign n62176 = ~n62174 & ~n62175 ;
  assign n62177 = \u0_R6_reg[28]/NET0131  & ~n62176 ;
  assign n62178 = ~\u0_R6_reg[28]/NET0131  & n62176 ;
  assign n62179 = ~n62177 & ~n62178 ;
  assign n62181 = decrypt_pad & ~\u0_uk_K_r6_reg[0]/NET0131  ;
  assign n62182 = ~decrypt_pad & ~\u0_uk_K_r6_reg[52]/NET0131  ;
  assign n62183 = ~n62181 & ~n62182 ;
  assign n62184 = \u0_R6_reg[29]/NET0131  & ~n62183 ;
  assign n62185 = ~\u0_R6_reg[29]/NET0131  & n62183 ;
  assign n62186 = ~n62184 & ~n62185 ;
  assign n62188 = decrypt_pad & ~\u0_uk_K_r6_reg[16]/NET0131  ;
  assign n62189 = ~decrypt_pad & ~\u0_uk_K_r6_reg[9]/NET0131  ;
  assign n62190 = ~n62188 & ~n62189 ;
  assign n62191 = \u0_R6_reg[1]/NET0131  & ~n62190 ;
  assign n62192 = ~\u0_R6_reg[1]/NET0131  & n62190 ;
  assign n62193 = ~n62191 & ~n62192 ;
  assign n62217 = n62186 & ~n62193 ;
  assign n62228 = n62179 & n62217 ;
  assign n62229 = ~n62173 & n62228 ;
  assign n62162 = decrypt_pad & ~\u0_uk_K_r6_reg[50]/NET0131  ;
  assign n62163 = ~decrypt_pad & ~\u0_uk_K_r6_reg[43]/NET0131  ;
  assign n62164 = ~n62162 & ~n62163 ;
  assign n62165 = \u0_R6_reg[32]/NET0131  & ~n62164 ;
  assign n62166 = ~\u0_R6_reg[32]/NET0131  & n62164 ;
  assign n62167 = ~n62165 & ~n62166 ;
  assign n62216 = ~n62173 & n62179 ;
  assign n62232 = ~n62216 & ~n62217 ;
  assign n62233 = n62167 & ~n62232 ;
  assign n62234 = ~n62229 & n62233 ;
  assign n62239 = ~n62179 & ~n62193 ;
  assign n62240 = ~n62186 & n62239 ;
  assign n62241 = ~n62173 & n62240 ;
  assign n62199 = n62173 & ~n62186 ;
  assign n62235 = ~n62179 & n62193 ;
  assign n62236 = n62199 & n62235 ;
  assign n62180 = n62173 & ~n62179 ;
  assign n62202 = ~n62186 & n62193 ;
  assign n62237 = ~n62180 & ~n62202 ;
  assign n62238 = ~n62232 & ~n62237 ;
  assign n62242 = ~n62236 & ~n62238 ;
  assign n62243 = ~n62241 & n62242 ;
  assign n62244 = ~n62234 & n62243 ;
  assign n62245 = n62210 & ~n62244 ;
  assign n62200 = n62179 & n62199 ;
  assign n62201 = ~n62193 & n62200 ;
  assign n62203 = ~n62179 & n62202 ;
  assign n62204 = ~n62201 & ~n62203 ;
  assign n62211 = ~n62204 & n62210 ;
  assign n62212 = n62186 & n62193 ;
  assign n62213 = n62180 & ~n62193 ;
  assign n62214 = ~n62212 & ~n62213 ;
  assign n62215 = ~n62210 & ~n62214 ;
  assign n62196 = n62179 & n62186 ;
  assign n62197 = n62173 & n62196 ;
  assign n62198 = n62193 & n62197 ;
  assign n62218 = n62210 & ~n62217 ;
  assign n62219 = n62216 & ~n62218 ;
  assign n62220 = ~n62198 & ~n62219 ;
  assign n62221 = ~n62215 & n62220 ;
  assign n62222 = ~n62211 & n62221 ;
  assign n62223 = ~n62167 & ~n62222 ;
  assign n62187 = n62180 & n62186 ;
  assign n62194 = n62187 & n62193 ;
  assign n62195 = n62167 & n62194 ;
  assign n62224 = ~n62173 & ~n62186 ;
  assign n62225 = ~n62179 & n62224 ;
  assign n62226 = ~n62200 & ~n62225 ;
  assign n62227 = n62167 & ~n62226 ;
  assign n62230 = ~n62227 & ~n62229 ;
  assign n62231 = ~n62210 & ~n62230 ;
  assign n62246 = ~n62195 & ~n62231 ;
  assign n62247 = ~n62223 & n62246 ;
  assign n62248 = ~n62245 & n62247 ;
  assign n62249 = \u0_L6_reg[5]/NET0131  & ~n62248 ;
  assign n62250 = ~\u0_L6_reg[5]/NET0131  & n62248 ;
  assign n62251 = ~n62249 & ~n62250 ;
  assign n62252 = decrypt_pad & ~\u0_uk_K_r6_reg[55]/P0001  ;
  assign n62253 = ~decrypt_pad & ~\u0_uk_K_r6_reg[48]/NET0131  ;
  assign n62254 = ~n62252 & ~n62253 ;
  assign n62255 = \u0_R6_reg[8]/NET0131  & ~n62254 ;
  assign n62256 = ~\u0_R6_reg[8]/NET0131  & n62254 ;
  assign n62257 = ~n62255 & ~n62256 ;
  assign n62258 = decrypt_pad & ~\u0_uk_K_r6_reg[13]/NET0131  ;
  assign n62259 = ~decrypt_pad & ~\u0_uk_K_r6_reg[6]/NET0131  ;
  assign n62260 = ~n62258 & ~n62259 ;
  assign n62261 = \u0_R6_reg[6]/NET0131  & ~n62260 ;
  assign n62262 = ~\u0_R6_reg[6]/NET0131  & n62260 ;
  assign n62263 = ~n62261 & ~n62262 ;
  assign n62264 = decrypt_pad & ~\u0_uk_K_r6_reg[3]/NET0131  ;
  assign n62265 = ~decrypt_pad & ~\u0_uk_K_r6_reg[53]/NET0131  ;
  assign n62266 = ~n62264 & ~n62265 ;
  assign n62267 = \u0_R6_reg[9]/NET0131  & ~n62266 ;
  assign n62268 = ~\u0_R6_reg[9]/NET0131  & n62266 ;
  assign n62269 = ~n62267 & ~n62268 ;
  assign n62270 = ~n62263 & n62269 ;
  assign n62271 = decrypt_pad & ~\u0_uk_K_r6_reg[47]/NET0131  ;
  assign n62272 = ~decrypt_pad & ~\u0_uk_K_r6_reg[40]/NET0131  ;
  assign n62273 = ~n62271 & ~n62272 ;
  assign n62274 = \u0_R6_reg[5]/NET0131  & ~n62273 ;
  assign n62275 = ~\u0_R6_reg[5]/NET0131  & n62273 ;
  assign n62276 = ~n62274 & ~n62275 ;
  assign n62277 = decrypt_pad & ~\u0_uk_K_r6_reg[32]/NET0131  ;
  assign n62278 = ~decrypt_pad & ~\u0_uk_K_r6_reg[25]/NET0131  ;
  assign n62279 = ~n62277 & ~n62278 ;
  assign n62280 = \u0_R6_reg[7]/NET0131  & ~n62279 ;
  assign n62281 = ~\u0_R6_reg[7]/NET0131  & n62279 ;
  assign n62282 = ~n62280 & ~n62281 ;
  assign n62283 = ~n62276 & ~n62282 ;
  assign n62284 = n62270 & n62283 ;
  assign n62285 = decrypt_pad & ~\u0_uk_K_r6_reg[11]/NET0131  ;
  assign n62286 = ~decrypt_pad & ~\u0_uk_K_r6_reg[4]/NET0131  ;
  assign n62287 = ~n62285 & ~n62286 ;
  assign n62288 = \u0_R6_reg[4]/NET0131  & ~n62287 ;
  assign n62289 = ~\u0_R6_reg[4]/NET0131  & n62287 ;
  assign n62290 = ~n62288 & ~n62289 ;
  assign n62291 = n62269 & ~n62290 ;
  assign n62292 = n62276 & n62291 ;
  assign n62293 = n62263 & n62292 ;
  assign n62294 = ~n62284 & ~n62293 ;
  assign n62296 = n62269 & ~n62276 ;
  assign n62301 = n62263 & n62290 ;
  assign n62302 = n62296 & n62301 ;
  assign n62303 = n62282 & n62302 ;
  assign n62308 = n62294 & ~n62303 ;
  assign n62295 = n62269 & n62290 ;
  assign n62297 = ~n62269 & n62276 ;
  assign n62298 = ~n62296 & ~n62297 ;
  assign n62299 = ~n62295 & ~n62298 ;
  assign n62300 = ~n62263 & n62299 ;
  assign n62304 = ~n62276 & n62295 ;
  assign n62305 = ~n62282 & ~n62304 ;
  assign n62306 = ~n62296 & ~n62301 ;
  assign n62307 = n62305 & ~n62306 ;
  assign n62309 = ~n62300 & ~n62307 ;
  assign n62310 = n62308 & n62309 ;
  assign n62311 = ~n62257 & ~n62310 ;
  assign n62313 = ~n62269 & ~n62290 ;
  assign n62330 = ~n62302 & ~n62313 ;
  assign n62331 = n62257 & ~n62330 ;
  assign n62312 = n62263 & ~n62276 ;
  assign n62332 = n62291 & ~n62312 ;
  assign n62333 = ~n62331 & ~n62332 ;
  assign n62329 = ~n62263 & n62276 ;
  assign n62334 = ~n62282 & ~n62329 ;
  assign n62335 = ~n62333 & n62334 ;
  assign n62314 = n62312 & n62313 ;
  assign n62315 = n62276 & n62290 ;
  assign n62316 = ~n62263 & n62315 ;
  assign n62317 = ~n62314 & ~n62316 ;
  assign n62318 = n62282 & ~n62317 ;
  assign n62319 = ~n62269 & ~n62276 ;
  assign n62320 = ~n62263 & n62319 ;
  assign n62321 = n62290 & n62320 ;
  assign n62322 = n62263 & ~n62290 ;
  assign n62323 = n62276 & n62282 ;
  assign n62324 = ~n62322 & n62323 ;
  assign n62325 = n62270 & n62315 ;
  assign n62326 = ~n62324 & ~n62325 ;
  assign n62327 = ~n62321 & n62326 ;
  assign n62328 = n62257 & ~n62327 ;
  assign n62336 = ~n62318 & ~n62328 ;
  assign n62337 = ~n62335 & n62336 ;
  assign n62338 = ~n62311 & n62337 ;
  assign n62339 = \u0_L6_reg[2]/NET0131  & n62338 ;
  assign n62340 = ~\u0_L6_reg[2]/NET0131  & ~n62338 ;
  assign n62341 = ~n62339 & ~n62340 ;
  assign n62363 = ~n61890 & n61912 ;
  assign n62364 = ~n61951 & ~n62363 ;
  assign n62365 = ~n61910 & n61960 ;
  assign n62366 = n62364 & ~n62365 ;
  assign n62367 = n61918 & ~n62366 ;
  assign n62343 = n61903 & n61945 ;
  assign n62350 = ~n61903 & ~n61912 ;
  assign n62351 = ~n61923 & n62350 ;
  assign n62361 = ~n62343 & ~n62351 ;
  assign n62362 = ~n61918 & ~n62361 ;
  assign n62368 = n61903 & n61924 ;
  assign n62369 = ~n62362 & ~n62368 ;
  assign n62370 = ~n62367 & n62369 ;
  assign n62371 = ~n61884 & ~n62370 ;
  assign n62342 = n61910 & n61926 ;
  assign n62344 = n61890 & n61931 ;
  assign n62345 = ~n62342 & ~n62344 ;
  assign n62346 = ~n62343 & n62345 ;
  assign n62347 = n61918 & ~n62346 ;
  assign n62352 = n61903 & ~n61939 ;
  assign n62353 = ~n61941 & n62352 ;
  assign n62348 = ~n61890 & ~n61952 ;
  assign n62349 = n61918 & ~n62348 ;
  assign n62354 = ~n62349 & ~n62351 ;
  assign n62355 = ~n62353 & n62354 ;
  assign n62356 = ~n62347 & ~n62355 ;
  assign n62357 = n61884 & ~n62356 ;
  assign n62358 = n61890 & n61910 ;
  assign n62359 = ~n61903 & n61918 ;
  assign n62360 = n62358 & n62359 ;
  assign n62372 = ~n61953 & ~n62360 ;
  assign n62373 = ~n62357 & n62372 ;
  assign n62374 = ~n62371 & n62373 ;
  assign n62375 = \u0_L6_reg[29]/NET0131  & ~n62374 ;
  assign n62376 = ~\u0_L6_reg[29]/NET0131  & n62374 ;
  assign n62377 = ~n62375 & ~n62376 ;
  assign n62380 = ~n61796 & ~n61864 ;
  assign n62382 = n61816 & ~n62380 ;
  assign n62381 = ~n61863 & ~n62380 ;
  assign n62383 = ~n61803 & ~n62381 ;
  assign n62384 = ~n62382 & n62383 ;
  assign n62385 = ~n61790 & n61870 ;
  assign n62386 = ~n61846 & ~n62385 ;
  assign n62387 = n61803 & ~n62386 ;
  assign n62378 = ~n61790 & n61850 ;
  assign n62379 = n61809 & n62378 ;
  assign n62388 = ~n61844 & ~n62379 ;
  assign n62389 = ~n62387 & n62388 ;
  assign n62390 = ~n62384 & n62389 ;
  assign n62391 = ~n61824 & ~n62390 ;
  assign n62392 = n61790 & n61848 ;
  assign n62393 = ~n62378 & ~n62392 ;
  assign n62394 = n61810 & ~n62393 ;
  assign n62399 = ~n61796 & ~n61816 ;
  assign n62401 = n61809 & ~n62399 ;
  assign n62400 = ~n61845 & n62399 ;
  assign n62402 = n61803 & ~n62400 ;
  assign n62403 = ~n62401 & n62402 ;
  assign n62398 = n61809 & n61849 ;
  assign n62395 = n61790 & n61850 ;
  assign n62396 = ~n61803 & ~n61836 ;
  assign n62397 = n61851 & n62396 ;
  assign n62404 = ~n62395 & ~n62397 ;
  assign n62405 = ~n62398 & n62404 ;
  assign n62406 = ~n62403 & n62405 ;
  assign n62407 = n61824 & ~n62406 ;
  assign n62408 = ~n62394 & ~n62407 ;
  assign n62409 = ~n62391 & n62408 ;
  assign n62410 = ~\u0_L6_reg[17]/NET0131  & ~n62409 ;
  assign n62411 = \u0_L6_reg[17]/NET0131  & n62409 ;
  assign n62412 = ~n62410 & ~n62411 ;
  assign n62415 = n61890 & n61952 ;
  assign n62416 = ~n61931 & ~n62415 ;
  assign n62417 = ~n61918 & ~n62416 ;
  assign n62413 = n61890 & n61939 ;
  assign n62414 = ~n61903 & n62413 ;
  assign n62419 = n61903 & n62358 ;
  assign n62418 = n61941 & n62359 ;
  assign n62420 = n61884 & ~n62418 ;
  assign n62421 = ~n62419 & n62420 ;
  assign n62422 = ~n62414 & n62421 ;
  assign n62423 = ~n62417 & n62422 ;
  assign n62426 = n61910 & ~n61932 ;
  assign n62427 = ~n61945 & ~n62426 ;
  assign n62428 = n61918 & ~n62427 ;
  assign n62424 = ~n62368 & ~n62413 ;
  assign n62425 = ~n61918 & ~n62424 ;
  assign n62429 = ~n61884 & ~n61953 ;
  assign n62430 = ~n61957 & n62429 ;
  assign n62431 = ~n62425 & n62430 ;
  assign n62432 = ~n62428 & n62431 ;
  assign n62433 = ~n62423 & ~n62432 ;
  assign n62434 = n61903 & n62364 ;
  assign n62435 = ~n61918 & ~n61940 ;
  assign n62436 = ~n62434 & n62435 ;
  assign n62437 = ~n61949 & ~n62342 ;
  assign n62438 = ~n61945 & n62437 ;
  assign n62439 = n61903 & n61918 ;
  assign n62440 = ~n62438 & n62439 ;
  assign n62441 = ~n62436 & ~n62440 ;
  assign n62442 = ~n62433 & n62441 ;
  assign n62443 = ~\u0_L6_reg[4]/NET0131  & ~n62442 ;
  assign n62444 = \u0_L6_reg[4]/NET0131  & n62442 ;
  assign n62445 = ~n62443 & ~n62444 ;
  assign n62452 = n61985 & n61992 ;
  assign n62453 = ~n62052 & ~n62452 ;
  assign n62454 = n62024 & ~n62453 ;
  assign n62455 = n62014 & ~n62048 ;
  assign n62456 = ~n62003 & n62455 ;
  assign n62447 = n61992 & ~n61998 ;
  assign n62448 = ~n61999 & ~n62447 ;
  assign n62446 = ~n61992 & n62024 ;
  assign n62449 = n61986 & ~n62446 ;
  assign n62450 = ~n62448 & n62449 ;
  assign n62451 = ~n61992 & n62007 ;
  assign n62457 = ~n62450 & ~n62451 ;
  assign n62458 = n62456 & n62457 ;
  assign n62459 = ~n62454 & n62458 ;
  assign n62464 = ~n61985 & n62036 ;
  assign n62465 = n61979 & ~n61998 ;
  assign n62466 = n61992 & n62465 ;
  assign n62467 = ~n62464 & ~n62466 ;
  assign n62463 = n61985 & ~n62036 ;
  assign n62468 = n61998 & ~n62037 ;
  assign n62469 = ~n62463 & ~n62468 ;
  assign n62470 = n62467 & n62469 ;
  assign n62471 = ~n62005 & ~n62006 ;
  assign n62472 = ~n62024 & ~n62471 ;
  assign n62461 = ~n62001 & ~n62026 ;
  assign n62462 = n61999 & ~n62461 ;
  assign n62460 = ~n62024 & n62037 ;
  assign n62473 = ~n62014 & ~n62460 ;
  assign n62474 = ~n62462 & n62473 ;
  assign n62475 = ~n62472 & n62474 ;
  assign n62476 = ~n62470 & n62475 ;
  assign n62477 = ~n62459 & ~n62476 ;
  assign n62478 = \u0_L6_reg[12]/NET0131  & n62477 ;
  assign n62479 = ~\u0_L6_reg[12]/NET0131  & ~n62477 ;
  assign n62480 = ~n62478 & ~n62479 ;
  assign n62493 = n61896 & ~n61920 ;
  assign n62494 = ~n62413 & ~n62493 ;
  assign n62495 = n61918 & ~n62494 ;
  assign n62491 = n61903 & n61951 ;
  assign n62492 = ~n61918 & ~n62437 ;
  assign n62496 = ~n62491 & ~n62492 ;
  assign n62497 = ~n62495 & n62496 ;
  assign n62498 = ~n61884 & ~n62497 ;
  assign n62485 = n61903 & ~n62437 ;
  assign n62481 = ~n61924 & ~n61928 ;
  assign n62482 = n61918 & ~n62481 ;
  assign n62483 = ~n61903 & n61924 ;
  assign n62484 = n61897 & ~n61918 ;
  assign n62486 = ~n62415 & ~n62484 ;
  assign n62487 = ~n62483 & n62486 ;
  assign n62488 = ~n62482 & n62487 ;
  assign n62489 = ~n62485 & n62488 ;
  assign n62490 = n61884 & ~n62489 ;
  assign n62499 = ~n61948 & ~n61958 ;
  assign n62500 = ~n62490 & n62499 ;
  assign n62501 = ~n62498 & n62500 ;
  assign n62502 = ~\u0_L6_reg[19]/P0001  & ~n62501 ;
  assign n62503 = \u0_L6_reg[19]/P0001  & n62501 ;
  assign n62504 = ~n62502 & ~n62503 ;
  assign n62539 = decrypt_pad & ~\u0_uk_K_r6_reg[35]/NET0131  ;
  assign n62540 = ~decrypt_pad & ~\u0_uk_K_r6_reg[28]/NET0131  ;
  assign n62541 = ~n62539 & ~n62540 ;
  assign n62542 = \u0_R6_reg[20]/NET0131  & ~n62541 ;
  assign n62543 = ~\u0_R6_reg[20]/NET0131  & n62541 ;
  assign n62544 = ~n62542 & ~n62543 ;
  assign n62505 = decrypt_pad & ~\u0_uk_K_r6_reg[15]/NET0131  ;
  assign n62506 = ~decrypt_pad & ~\u0_uk_K_r6_reg[8]/NET0131  ;
  assign n62507 = ~n62505 & ~n62506 ;
  assign n62508 = \u0_R6_reg[17]/NET0131  & ~n62507 ;
  assign n62509 = ~\u0_R6_reg[17]/NET0131  & n62507 ;
  assign n62510 = ~n62508 & ~n62509 ;
  assign n62511 = decrypt_pad & ~\u0_uk_K_r6_reg[52]/NET0131  ;
  assign n62512 = ~decrypt_pad & ~\u0_uk_K_r6_reg[45]/NET0131  ;
  assign n62513 = ~n62511 & ~n62512 ;
  assign n62514 = \u0_R6_reg[16]/NET0131  & ~n62513 ;
  assign n62515 = ~\u0_R6_reg[16]/NET0131  & n62513 ;
  assign n62516 = ~n62514 & ~n62515 ;
  assign n62518 = decrypt_pad & ~\u0_uk_K_r6_reg[36]/NET0131  ;
  assign n62519 = ~decrypt_pad & ~\u0_uk_K_r6_reg[29]/NET0131  ;
  assign n62520 = ~n62518 & ~n62519 ;
  assign n62521 = \u0_R6_reg[21]/NET0131  & ~n62520 ;
  assign n62522 = ~\u0_R6_reg[21]/NET0131  & n62520 ;
  assign n62523 = ~n62521 & ~n62522 ;
  assign n62551 = n62516 & n62523 ;
  assign n62572 = n62510 & n62551 ;
  assign n62525 = decrypt_pad & ~\u0_uk_K_r6_reg[51]/NET0131  ;
  assign n62526 = ~decrypt_pad & ~\u0_uk_K_r6_reg[44]/NET0131  ;
  assign n62527 = ~n62525 & ~n62526 ;
  assign n62528 = \u0_R6_reg[19]/NET0131  & ~n62527 ;
  assign n62529 = ~\u0_R6_reg[19]/NET0131  & n62527 ;
  assign n62530 = ~n62528 & ~n62529 ;
  assign n62517 = ~n62510 & n62516 ;
  assign n62531 = decrypt_pad & ~\u0_uk_K_r6_reg[9]/NET0131  ;
  assign n62532 = ~decrypt_pad & ~\u0_uk_K_r6_reg[2]/NET0131  ;
  assign n62533 = ~n62531 & ~n62532 ;
  assign n62534 = \u0_R6_reg[18]/NET0131  & ~n62533 ;
  assign n62535 = ~\u0_R6_reg[18]/NET0131  & n62533 ;
  assign n62536 = ~n62534 & ~n62535 ;
  assign n62553 = ~n62523 & ~n62536 ;
  assign n62573 = n62517 & n62553 ;
  assign n62574 = n62530 & ~n62573 ;
  assign n62575 = ~n62572 & n62574 ;
  assign n62545 = ~n62516 & n62523 ;
  assign n62564 = ~n62510 & n62536 ;
  assign n62576 = n62545 & ~n62564 ;
  assign n62552 = ~n62510 & n62551 ;
  assign n62577 = ~n62530 & ~n62552 ;
  assign n62578 = ~n62576 & n62577 ;
  assign n62579 = ~n62575 & ~n62578 ;
  assign n62566 = n62510 & ~n62536 ;
  assign n62567 = ~n62516 & n62566 ;
  assign n62547 = n62510 & ~n62523 ;
  assign n62580 = n62516 & n62547 ;
  assign n62581 = ~n62516 & ~n62523 ;
  assign n62582 = ~n62510 & n62581 ;
  assign n62583 = ~n62580 & ~n62582 ;
  assign n62584 = n62536 & ~n62583 ;
  assign n62585 = ~n62567 & ~n62584 ;
  assign n62586 = ~n62579 & n62585 ;
  assign n62587 = ~n62544 & ~n62586 ;
  assign n62554 = ~n62510 & ~n62516 ;
  assign n62555 = n62553 & n62554 ;
  assign n62556 = ~n62552 & ~n62555 ;
  assign n62557 = n62530 & ~n62556 ;
  assign n62546 = ~n62510 & n62545 ;
  assign n62548 = ~n62516 & n62547 ;
  assign n62549 = ~n62546 & ~n62548 ;
  assign n62550 = n62536 & ~n62549 ;
  assign n62558 = ~n62530 & ~n62536 ;
  assign n62559 = n62516 & n62558 ;
  assign n62560 = ~n62550 & ~n62559 ;
  assign n62561 = ~n62557 & n62560 ;
  assign n62562 = n62544 & ~n62561 ;
  assign n62524 = n62517 & ~n62523 ;
  assign n62537 = ~n62530 & n62536 ;
  assign n62538 = n62524 & n62537 ;
  assign n62568 = n62523 & n62567 ;
  assign n62563 = n62536 & n62547 ;
  assign n62565 = n62545 & n62564 ;
  assign n62569 = ~n62563 & ~n62565 ;
  assign n62570 = ~n62568 & n62569 ;
  assign n62571 = n62530 & ~n62570 ;
  assign n62588 = ~n62538 & ~n62571 ;
  assign n62589 = ~n62562 & n62588 ;
  assign n62590 = ~n62587 & n62589 ;
  assign n62591 = ~\u0_L6_reg[8]/NET0131  & ~n62590 ;
  assign n62592 = \u0_L6_reg[8]/NET0131  & n62590 ;
  assign n62593 = ~n62591 & ~n62592 ;
  assign n62600 = n62179 & ~n62212 ;
  assign n62601 = ~n62224 & n62600 ;
  assign n62602 = ~n62225 & ~n62601 ;
  assign n62603 = n62210 & ~n62602 ;
  assign n62597 = ~n62193 & ~n62226 ;
  assign n62598 = ~n62179 & ~n62210 ;
  assign n62599 = n62217 & n62598 ;
  assign n62606 = ~n62167 & ~n62187 ;
  assign n62607 = ~n62599 & n62606 ;
  assign n62594 = n62193 & ~n62210 ;
  assign n62595 = n62173 & n62594 ;
  assign n62596 = ~n62179 & n62595 ;
  assign n62604 = ~n62212 & ~n62594 ;
  assign n62605 = n62216 & ~n62604 ;
  assign n62608 = ~n62596 & ~n62605 ;
  assign n62609 = n62607 & n62608 ;
  assign n62610 = ~n62597 & n62609 ;
  assign n62611 = ~n62603 & n62610 ;
  assign n62615 = n62193 & n62200 ;
  assign n62616 = ~n62202 & n62216 ;
  assign n62617 = ~n62210 & ~n62616 ;
  assign n62618 = ~n62615 & n62617 ;
  assign n62619 = ~n62179 & ~n62199 ;
  assign n62620 = ~n62217 & n62619 ;
  assign n62621 = ~n62173 & n62202 ;
  assign n62622 = ~n62197 & n62210 ;
  assign n62623 = ~n62621 & n62622 ;
  assign n62624 = ~n62620 & n62623 ;
  assign n62625 = ~n62618 & ~n62624 ;
  assign n62613 = ~n62228 & ~n62240 ;
  assign n62614 = n62173 & ~n62613 ;
  assign n62612 = ~n62173 & n62203 ;
  assign n62626 = n62167 & ~n62612 ;
  assign n62627 = ~n62614 & n62626 ;
  assign n62628 = ~n62625 & n62627 ;
  assign n62629 = ~n62611 & ~n62628 ;
  assign n62630 = ~\u0_L6_reg[21]/NET0131  & n62629 ;
  assign n62631 = \u0_L6_reg[21]/NET0131  & ~n62629 ;
  assign n62632 = ~n62630 & ~n62631 ;
  assign n62633 = ~n61827 & ~n61860 ;
  assign n62634 = ~n61809 & ~n62633 ;
  assign n62635 = n61816 & n62385 ;
  assign n62636 = ~n62634 & ~n62635 ;
  assign n62637 = ~n61803 & ~n62636 ;
  assign n62639 = n61803 & ~n61825 ;
  assign n62640 = n61865 & n62639 ;
  assign n62638 = n61845 & n62399 ;
  assign n62641 = ~n61818 & ~n62638 ;
  assign n62642 = ~n62640 & n62641 ;
  assign n62643 = ~n62637 & n62642 ;
  assign n62644 = n61824 & ~n62643 ;
  assign n62646 = ~n61817 & ~n61850 ;
  assign n62647 = n61790 & ~n62646 ;
  assign n62650 = n61803 & n61860 ;
  assign n62645 = ~n61790 & n62399 ;
  assign n62648 = ~n61797 & ~n61803 ;
  assign n62649 = n62401 & n62648 ;
  assign n62651 = ~n62645 & ~n62649 ;
  assign n62652 = ~n62650 & n62651 ;
  assign n62653 = ~n62647 & n62652 ;
  assign n62654 = ~n61824 & ~n62653 ;
  assign n62655 = ~n61860 & ~n61870 ;
  assign n62656 = n61833 & ~n62655 ;
  assign n62657 = n61832 & n62399 ;
  assign n62658 = ~n61847 & ~n62657 ;
  assign n62659 = ~n62398 & n62658 ;
  assign n62660 = ~n61803 & ~n62659 ;
  assign n62661 = ~n62656 & ~n62660 ;
  assign n62662 = ~n62654 & n62661 ;
  assign n62663 = ~n62644 & n62662 ;
  assign n62664 = \u0_L6_reg[23]/NET0131  & ~n62663 ;
  assign n62665 = ~\u0_L6_reg[23]/NET0131  & n62663 ;
  assign n62666 = ~n62664 & ~n62665 ;
  assign n62670 = ~n62263 & n62313 ;
  assign n62671 = ~n62292 & ~n62670 ;
  assign n62672 = n62282 & n62671 ;
  assign n62676 = ~n62276 & n62322 ;
  assign n62677 = ~n62282 & ~n62676 ;
  assign n62674 = ~n62269 & n62290 ;
  assign n62675 = ~n62263 & n62674 ;
  assign n62673 = ~n62276 & n62291 ;
  assign n62678 = ~n62315 & ~n62673 ;
  assign n62679 = ~n62675 & n62678 ;
  assign n62680 = n62677 & n62679 ;
  assign n62681 = ~n62672 & ~n62680 ;
  assign n62668 = ~n62295 & ~n62313 ;
  assign n62669 = n62312 & ~n62668 ;
  assign n62667 = n62297 & n62301 ;
  assign n62682 = ~n62257 & ~n62667 ;
  assign n62683 = ~n62669 & n62682 ;
  assign n62684 = ~n62681 & n62683 ;
  assign n62690 = n62290 & n62298 ;
  assign n62689 = n62297 & n62322 ;
  assign n62691 = n62282 & ~n62689 ;
  assign n62692 = ~n62690 & n62691 ;
  assign n62693 = ~n62667 & n62671 ;
  assign n62694 = n62677 & n62693 ;
  assign n62695 = ~n62692 & ~n62694 ;
  assign n62685 = n62282 & n62290 ;
  assign n62686 = ~n62304 & ~n62685 ;
  assign n62687 = ~n62263 & ~n62686 ;
  assign n62688 = n62291 & n62312 ;
  assign n62696 = n62257 & ~n62688 ;
  assign n62697 = ~n62687 & n62696 ;
  assign n62698 = ~n62695 & n62697 ;
  assign n62699 = ~n62684 & ~n62698 ;
  assign n62700 = ~\u0_L6_reg[28]/NET0131  & n62699 ;
  assign n62701 = \u0_L6_reg[28]/NET0131  & ~n62699 ;
  assign n62702 = ~n62700 & ~n62701 ;
  assign n62728 = ~n62536 & n62551 ;
  assign n62727 = n62545 & ~n62566 ;
  assign n62729 = ~n62580 & ~n62727 ;
  assign n62730 = ~n62728 & n62729 ;
  assign n62731 = n62530 & ~n62730 ;
  assign n62720 = n62510 & n62545 ;
  assign n62721 = ~n62582 & ~n62720 ;
  assign n62722 = n62558 & ~n62721 ;
  assign n62713 = n62523 & n62536 ;
  assign n62725 = n62517 & ~n62553 ;
  assign n62726 = ~n62713 & n62725 ;
  assign n62723 = ~n62536 & n62580 ;
  assign n62724 = n62537 & n62572 ;
  assign n62732 = ~n62723 & ~n62724 ;
  assign n62733 = ~n62726 & n62732 ;
  assign n62734 = ~n62722 & n62733 ;
  assign n62735 = ~n62731 & n62734 ;
  assign n62736 = n62544 & ~n62735 ;
  assign n62707 = ~n62536 & n62572 ;
  assign n62708 = ~n62546 & ~n62563 ;
  assign n62709 = ~n62573 & n62708 ;
  assign n62710 = ~n62707 & n62709 ;
  assign n62711 = ~n62530 & ~n62710 ;
  assign n62703 = n62536 & n62551 ;
  assign n62704 = ~n62567 & ~n62582 ;
  assign n62705 = ~n62703 & n62704 ;
  assign n62706 = n62530 & ~n62705 ;
  assign n62714 = ~n62581 & ~n62713 ;
  assign n62712 = n62510 & n62536 ;
  assign n62715 = ~n62554 & ~n62712 ;
  assign n62716 = ~n62714 & n62715 ;
  assign n62717 = ~n62706 & ~n62716 ;
  assign n62718 = ~n62711 & n62717 ;
  assign n62719 = ~n62544 & ~n62718 ;
  assign n62737 = ~n62530 & ~n62550 ;
  assign n62738 = n62536 & n62582 ;
  assign n62739 = n62530 & ~n62723 ;
  assign n62740 = ~n62738 & n62739 ;
  assign n62741 = ~n62737 & ~n62740 ;
  assign n62742 = ~n62719 & ~n62741 ;
  assign n62743 = ~n62736 & n62742 ;
  assign n62744 = ~\u0_L6_reg[14]/NET0131  & ~n62743 ;
  assign n62745 = \u0_L6_reg[14]/NET0131  & n62743 ;
  assign n62746 = ~n62744 & ~n62745 ;
  assign n62771 = ~n62213 & ~n62216 ;
  assign n62772 = n62186 & ~n62771 ;
  assign n62768 = n62210 & n62239 ;
  assign n62769 = ~n62595 & ~n62768 ;
  assign n62770 = ~n62186 & ~n62769 ;
  assign n62773 = ~n62615 & ~n62770 ;
  assign n62774 = ~n62772 & n62773 ;
  assign n62775 = n62167 & ~n62774 ;
  assign n62747 = ~n62173 & n62186 ;
  assign n62748 = ~n62193 & n62747 ;
  assign n62749 = ~n62196 & ~n62203 ;
  assign n62750 = ~n62748 & n62749 ;
  assign n62751 = n62210 & ~n62750 ;
  assign n62752 = ~n62186 & ~n62193 ;
  assign n62753 = n62216 & n62752 ;
  assign n62754 = ~n62751 & ~n62753 ;
  assign n62755 = ~n62167 & ~n62754 ;
  assign n62763 = ~n62193 & ~n62747 ;
  assign n62764 = n62619 & n62763 ;
  assign n62762 = n62235 & n62747 ;
  assign n62765 = ~n62200 & ~n62762 ;
  assign n62766 = ~n62764 & n62765 ;
  assign n62767 = ~n62210 & ~n62766 ;
  assign n62756 = ~n62167 & n62179 ;
  assign n62757 = ~n62186 & ~n62210 ;
  assign n62758 = n62756 & n62757 ;
  assign n62759 = n62193 & ~n62747 ;
  assign n62760 = n62210 & n62619 ;
  assign n62761 = n62759 & n62760 ;
  assign n62776 = ~n62758 & ~n62761 ;
  assign n62777 = ~n62767 & n62776 ;
  assign n62778 = ~n62755 & n62777 ;
  assign n62779 = ~n62775 & n62778 ;
  assign n62780 = \u0_L6_reg[15]/P0001  & n62779 ;
  assign n62781 = ~\u0_L6_reg[15]/P0001  & ~n62779 ;
  assign n62782 = ~n62780 & ~n62781 ;
  assign n62783 = ~n62325 & ~n62667 ;
  assign n62784 = ~n62290 & n62297 ;
  assign n62785 = ~n62688 & ~n62784 ;
  assign n62786 = ~n62321 & n62785 ;
  assign n62787 = ~n62257 & ~n62786 ;
  assign n62788 = n62783 & ~n62787 ;
  assign n62789 = ~n62282 & ~n62788 ;
  assign n62795 = ~n62276 & n62668 ;
  assign n62794 = n62276 & ~n62675 ;
  assign n62796 = n62282 & ~n62794 ;
  assign n62797 = ~n62795 & n62796 ;
  assign n62792 = ~n62263 & ~n62283 ;
  assign n62793 = n62291 & n62792 ;
  assign n62790 = n62263 & ~n62297 ;
  assign n62791 = n62685 & n62790 ;
  assign n62798 = ~n62257 & ~n62791 ;
  assign n62799 = ~n62793 & n62798 ;
  assign n62800 = ~n62797 & n62799 ;
  assign n62801 = ~n62269 & n62312 ;
  assign n62802 = n62305 & ~n62801 ;
  assign n62803 = n62263 & n62291 ;
  assign n62804 = n62282 & ~n62320 ;
  assign n62805 = ~n62803 & n62804 ;
  assign n62806 = ~n62802 & ~n62805 ;
  assign n62807 = ~n62263 & n62784 ;
  assign n62808 = n62257 & n62783 ;
  assign n62809 = ~n62807 & n62808 ;
  assign n62810 = n62294 & n62809 ;
  assign n62811 = ~n62806 & n62810 ;
  assign n62812 = ~n62800 & ~n62811 ;
  assign n62813 = ~n62789 & ~n62812 ;
  assign n62814 = ~\u0_L6_reg[13]/NET0131  & n62813 ;
  assign n62815 = \u0_L6_reg[13]/NET0131  & ~n62813 ;
  assign n62816 = ~n62814 & ~n62815 ;
  assign n62819 = ~n62112 & ~n62131 ;
  assign n62820 = ~n62104 & ~n62819 ;
  assign n62822 = n62068 & ~n62133 ;
  assign n62823 = n62138 & n62822 ;
  assign n62817 = ~n62074 & n62081 ;
  assign n62818 = n62094 & n62817 ;
  assign n62821 = n62075 & n62113 ;
  assign n62824 = ~n62818 & ~n62821 ;
  assign n62825 = ~n62823 & n62824 ;
  assign n62826 = n62126 & n62825 ;
  assign n62827 = ~n62820 & n62826 ;
  assign n62831 = ~n62099 & ~n62118 ;
  assign n62832 = n62068 & ~n62831 ;
  assign n62833 = ~n62094 & n62135 ;
  assign n62834 = n62087 & n62833 ;
  assign n62835 = ~n62141 & ~n62834 ;
  assign n62828 = n62100 & ~n62151 ;
  assign n62829 = ~n62134 & ~n62828 ;
  assign n62830 = ~n62068 & ~n62829 ;
  assign n62836 = n62125 & ~n62830 ;
  assign n62837 = n62835 & n62836 ;
  assign n62838 = ~n62832 & n62837 ;
  assign n62839 = ~n62827 & ~n62838 ;
  assign n62840 = n62068 & ~n62152 ;
  assign n62841 = n62110 & n62835 ;
  assign n62842 = ~n62840 & ~n62841 ;
  assign n62843 = ~n62106 & ~n62842 ;
  assign n62844 = ~n62839 & n62843 ;
  assign n62845 = ~\u0_L6_reg[10]/NET0131  & ~n62844 ;
  assign n62846 = \u0_L6_reg[10]/NET0131  & n62844 ;
  assign n62847 = ~n62845 & ~n62846 ;
  assign n62848 = ~n62087 & ~n62139 ;
  assign n62849 = ~n62114 & ~n62848 ;
  assign n62850 = ~n62074 & ~n62849 ;
  assign n62851 = ~n62111 & ~n62833 ;
  assign n62852 = ~n62125 & ~n62851 ;
  assign n62853 = ~n62068 & ~n62852 ;
  assign n62854 = ~n62850 & n62853 ;
  assign n62855 = n62068 & ~n62134 ;
  assign n62856 = ~n62099 & n62855 ;
  assign n62857 = ~n62854 & ~n62856 ;
  assign n62859 = ~n62074 & ~n62118 ;
  assign n62860 = ~n62095 & ~n62142 ;
  assign n62861 = n62074 & ~n62131 ;
  assign n62862 = n62860 & n62861 ;
  assign n62863 = ~n62859 & ~n62862 ;
  assign n62864 = ~n62098 & ~n62113 ;
  assign n62865 = ~n62068 & ~n62817 ;
  assign n62866 = ~n62864 & n62865 ;
  assign n62858 = n62068 & n62112 ;
  assign n62867 = n62125 & ~n62858 ;
  assign n62868 = ~n62866 & n62867 ;
  assign n62869 = ~n62863 & n62868 ;
  assign n62871 = ~n62094 & n62817 ;
  assign n62872 = ~n62125 & ~n62134 ;
  assign n62873 = ~n62871 & n62872 ;
  assign n62870 = ~n62088 & n62105 ;
  assign n62874 = ~n62143 & ~n62870 ;
  assign n62875 = n62873 & n62874 ;
  assign n62876 = ~n62869 & ~n62875 ;
  assign n62877 = ~n62857 & ~n62876 ;
  assign n62878 = ~\u0_L6_reg[26]/NET0131  & ~n62877 ;
  assign n62879 = \u0_L6_reg[26]/NET0131  & n62877 ;
  assign n62880 = ~n62878 & ~n62879 ;
  assign n62881 = ~n62553 & ~n62581 ;
  assign n62882 = ~n62554 & n62881 ;
  assign n62883 = ~n62566 & ~n62882 ;
  assign n62884 = ~n62572 & ~n62883 ;
  assign n62885 = n62530 & ~n62884 ;
  assign n62886 = ~n62552 & ~n62567 ;
  assign n62887 = ~n62530 & ~n62886 ;
  assign n62888 = n62510 & ~n62713 ;
  assign n62889 = n62881 & n62888 ;
  assign n62890 = ~n62887 & ~n62889 ;
  assign n62891 = ~n62885 & n62890 ;
  assign n62892 = n62544 & ~n62891 ;
  assign n62896 = ~n62523 & n62530 ;
  assign n62897 = ~n62516 & n62712 ;
  assign n62898 = ~n62524 & ~n62897 ;
  assign n62899 = ~n62896 & ~n62898 ;
  assign n62901 = n62530 & ~n62547 ;
  assign n62900 = ~n62530 & ~n62554 ;
  assign n62902 = ~n62536 & ~n62900 ;
  assign n62903 = ~n62901 & n62902 ;
  assign n62904 = ~n62899 & ~n62903 ;
  assign n62905 = ~n62544 & ~n62904 ;
  assign n62893 = ~n62536 & n62546 ;
  assign n62894 = ~n62584 & ~n62893 ;
  assign n62895 = n62530 & ~n62894 ;
  assign n62906 = n62517 & n62537 ;
  assign n62907 = ~n62707 & ~n62906 ;
  assign n62908 = ~n62895 & n62907 ;
  assign n62909 = ~n62905 & n62908 ;
  assign n62910 = ~n62892 & n62909 ;
  assign n62911 = ~\u0_L6_reg[25]/NET0131  & ~n62910 ;
  assign n62912 = \u0_L6_reg[25]/NET0131  & n62910 ;
  assign n62913 = ~n62911 & ~n62912 ;
  assign n62927 = ~n62097 & ~n62107 ;
  assign n62928 = n62081 & ~n62927 ;
  assign n62929 = ~n62068 & ~n62928 ;
  assign n62930 = n62068 & ~n62108 ;
  assign n62931 = ~n62153 & n62930 ;
  assign n62932 = ~n62929 & ~n62931 ;
  assign n62933 = ~n62074 & ~n62860 ;
  assign n62934 = ~n62141 & ~n62933 ;
  assign n62935 = ~n62932 & n62934 ;
  assign n62936 = ~n62125 & ~n62935 ;
  assign n62921 = ~n62100 & n62151 ;
  assign n62922 = ~n62095 & ~n62921 ;
  assign n62923 = ~n62068 & ~n62922 ;
  assign n62919 = n62074 & n62142 ;
  assign n62924 = ~n62833 & ~n62919 ;
  assign n62925 = ~n62923 & n62924 ;
  assign n62926 = n62125 & ~n62925 ;
  assign n62914 = ~n62119 & n62835 ;
  assign n62915 = n62068 & ~n62914 ;
  assign n62920 = ~n62068 & n62919 ;
  assign n62916 = ~n62097 & ~n62871 ;
  assign n62917 = n62068 & n62125 ;
  assign n62918 = ~n62916 & n62917 ;
  assign n62937 = ~n62137 & ~n62918 ;
  assign n62938 = ~n62920 & n62937 ;
  assign n62939 = ~n62915 & n62938 ;
  assign n62940 = ~n62926 & n62939 ;
  assign n62941 = ~n62936 & n62940 ;
  assign n62942 = ~\u0_L6_reg[1]/NET0131  & ~n62941 ;
  assign n62943 = \u0_L6_reg[1]/NET0131  & n62941 ;
  assign n62944 = ~n62942 & ~n62943 ;
  assign n62951 = ~n62028 & n62471 ;
  assign n62952 = n62448 & ~n62951 ;
  assign n62950 = n61985 & ~n62448 ;
  assign n62949 = n61979 & ~n62448 ;
  assign n62953 = ~n62024 & ~n62949 ;
  assign n62954 = ~n62950 & n62953 ;
  assign n62955 = ~n62952 & n62954 ;
  assign n62945 = ~n61985 & ~n62024 ;
  assign n62946 = n62466 & ~n62945 ;
  assign n62947 = ~n62007 & ~n62033 ;
  assign n62948 = n62024 & ~n62947 ;
  assign n62956 = ~n62946 & ~n62948 ;
  assign n62957 = ~n62955 & n62956 ;
  assign n62958 = n62014 & ~n62957 ;
  assign n62962 = n61992 & ~n62465 ;
  assign n62963 = ~n62945 & n62962 ;
  assign n62964 = ~n62007 & n62963 ;
  assign n62960 = ~n61979 & n62447 ;
  assign n62961 = n62472 & ~n62960 ;
  assign n62965 = n62004 & ~n62961 ;
  assign n62966 = ~n62964 & n62965 ;
  assign n62967 = ~n62014 & ~n62966 ;
  assign n62959 = n62000 & n62024 ;
  assign n62968 = n62044 & ~n62447 ;
  assign n62969 = n62038 & n62968 ;
  assign n62970 = ~n62959 & ~n62969 ;
  assign n62971 = ~n62967 & n62970 ;
  assign n62972 = ~n62958 & n62971 ;
  assign n62973 = \u0_L6_reg[32]/NET0131  & n62972 ;
  assign n62974 = ~\u0_L6_reg[32]/NET0131  & ~n62972 ;
  assign n62975 = ~n62973 & ~n62974 ;
  assign n62991 = ~n62228 & ~n62620 ;
  assign n62992 = ~n62210 & ~n62991 ;
  assign n62988 = ~n62179 & ~n62748 ;
  assign n62989 = n62210 & ~n62600 ;
  assign n62990 = ~n62988 & n62989 ;
  assign n62993 = ~n62194 & ~n62621 ;
  assign n62994 = ~n62201 & n62993 ;
  assign n62995 = ~n62990 & n62994 ;
  assign n62996 = ~n62992 & n62995 ;
  assign n62997 = n62167 & ~n62996 ;
  assign n62979 = ~n62187 & n62210 ;
  assign n62980 = ~n62748 & ~n62759 ;
  assign n62981 = n62979 & n62980 ;
  assign n62978 = n62179 & n62595 ;
  assign n62982 = ~n62236 & ~n62599 ;
  assign n62983 = ~n62978 & n62982 ;
  assign n62984 = ~n62981 & n62983 ;
  assign n62985 = ~n62167 & ~n62984 ;
  assign n62976 = ~n62229 & ~n62238 ;
  assign n62977 = ~n62210 & ~n62976 ;
  assign n62986 = ~n62193 & n62210 ;
  assign n62987 = n62199 & n62986 ;
  assign n62998 = ~n62977 & ~n62987 ;
  assign n62999 = ~n62985 & n62998 ;
  assign n63000 = ~n62997 & n62999 ;
  assign n63001 = ~\u0_L6_reg[27]/NET0131  & ~n63000 ;
  assign n63002 = \u0_L6_reg[27]/NET0131  & n63000 ;
  assign n63003 = ~n63001 & ~n63002 ;
  assign n63010 = decrypt_pad & ~\u0_uk_K_r6_reg[12]/NET0131  ;
  assign n63011 = ~decrypt_pad & ~\u0_uk_K_r6_reg[5]/NET0131  ;
  assign n63012 = ~n63010 & ~n63011 ;
  assign n63013 = \u0_R6_reg[8]/NET0131  & ~n63012 ;
  assign n63014 = ~\u0_R6_reg[8]/NET0131  & n63012 ;
  assign n63015 = ~n63013 & ~n63014 ;
  assign n63016 = decrypt_pad & ~\u0_uk_K_r6_reg[46]/NET0131  ;
  assign n63017 = ~decrypt_pad & ~\u0_uk_K_r6_reg[39]/NET0131  ;
  assign n63018 = ~n63016 & ~n63017 ;
  assign n63019 = \u0_R6_reg[13]/NET0131  & ~n63018 ;
  assign n63020 = ~\u0_R6_reg[13]/NET0131  & n63018 ;
  assign n63021 = ~n63019 & ~n63020 ;
  assign n63040 = ~n63015 & ~n63021 ;
  assign n63041 = n63015 & n63021 ;
  assign n63042 = ~n63040 & ~n63041 ;
  assign n63004 = decrypt_pad & ~\u0_uk_K_r6_reg[18]/NET0131  ;
  assign n63005 = ~decrypt_pad & ~\u0_uk_K_r6_reg[11]/NET0131  ;
  assign n63006 = ~n63004 & ~n63005 ;
  assign n63007 = \u0_R6_reg[11]/NET0131  & ~n63006 ;
  assign n63008 = ~\u0_R6_reg[11]/NET0131  & n63006 ;
  assign n63009 = ~n63007 & ~n63008 ;
  assign n63038 = n63009 & ~n63015 ;
  assign n63023 = decrypt_pad & ~\u0_uk_K_r6_reg[17]/NET0131  ;
  assign n63024 = ~decrypt_pad & ~\u0_uk_K_r6_reg[10]/NET0131  ;
  assign n63025 = ~n63023 & ~n63024 ;
  assign n63026 = \u0_R6_reg[10]/NET0131  & ~n63025 ;
  assign n63027 = ~\u0_R6_reg[10]/NET0131  & n63025 ;
  assign n63028 = ~n63026 & ~n63027 ;
  assign n63030 = decrypt_pad & ~\u0_uk_K_r6_reg[41]/NET0131  ;
  assign n63031 = ~decrypt_pad & ~\u0_uk_K_r6_reg[34]/NET0131  ;
  assign n63032 = ~n63030 & ~n63031 ;
  assign n63033 = \u0_R6_reg[9]/NET0131  & ~n63032 ;
  assign n63034 = ~\u0_R6_reg[9]/NET0131  & n63032 ;
  assign n63035 = ~n63033 & ~n63034 ;
  assign n63039 = ~n63028 & ~n63035 ;
  assign n63043 = ~n63038 & n63039 ;
  assign n63044 = n63042 & n63043 ;
  assign n63051 = n63028 & n63035 ;
  assign n63056 = n63015 & ~n63021 ;
  assign n63057 = n63051 & n63056 ;
  assign n63045 = decrypt_pad & ~\u0_uk_K_r6_reg[33]/NET0131  ;
  assign n63046 = ~decrypt_pad & ~\u0_uk_K_r6_reg[26]/P0001  ;
  assign n63047 = ~n63045 & ~n63046 ;
  assign n63048 = \u0_R6_reg[12]/NET0131  & ~n63047 ;
  assign n63049 = ~\u0_R6_reg[12]/NET0131  & n63047 ;
  assign n63050 = ~n63048 & ~n63049 ;
  assign n63054 = ~n63028 & n63035 ;
  assign n63055 = n63038 & n63054 ;
  assign n63058 = ~n63050 & ~n63055 ;
  assign n63059 = ~n63057 & n63058 ;
  assign n63060 = ~n63044 & n63059 ;
  assign n63022 = ~n63015 & n63021 ;
  assign n63029 = n63022 & n63028 ;
  assign n63036 = n63029 & n63035 ;
  assign n63037 = ~n63009 & n63036 ;
  assign n63052 = ~n63039 & ~n63042 ;
  assign n63053 = ~n63051 & n63052 ;
  assign n63061 = ~n63037 & ~n63053 ;
  assign n63062 = n63060 & n63061 ;
  assign n63067 = ~n63015 & ~n63054 ;
  assign n63066 = n63021 & ~n63035 ;
  assign n63065 = ~n63021 & n63035 ;
  assign n63068 = ~n63009 & ~n63065 ;
  assign n63069 = ~n63066 & n63068 ;
  assign n63070 = ~n63067 & n63069 ;
  assign n63063 = n63028 & n63040 ;
  assign n63064 = n63035 & n63063 ;
  assign n63071 = n63050 & ~n63064 ;
  assign n63072 = ~n63070 & n63071 ;
  assign n63073 = ~n63062 & ~n63072 ;
  assign n63075 = n63035 & n63056 ;
  assign n63076 = ~n63029 & ~n63075 ;
  assign n63077 = ~n63066 & n63076 ;
  assign n63078 = n63050 & ~n63077 ;
  assign n63074 = n63028 & n63066 ;
  assign n63079 = ~n63028 & n63040 ;
  assign n63080 = ~n63035 & n63079 ;
  assign n63081 = ~n63074 & ~n63080 ;
  assign n63082 = ~n63078 & n63081 ;
  assign n63083 = n63009 & ~n63082 ;
  assign n63084 = ~n63073 & ~n63083 ;
  assign n63085 = ~\u0_L6_reg[6]/NET0131  & ~n63084 ;
  assign n63086 = \u0_L6_reg[6]/NET0131  & n63084 ;
  assign n63087 = ~n63085 & ~n63086 ;
  assign n63088 = ~n62565 & n62574 ;
  assign n63089 = ~n62558 & ~n62577 ;
  assign n63090 = ~n62536 & ~n62583 ;
  assign n63091 = ~n63089 & ~n63090 ;
  assign n63092 = ~n63088 & ~n63091 ;
  assign n63096 = ~n62536 & n62545 ;
  assign n63097 = ~n62580 & ~n63096 ;
  assign n63098 = n62530 & ~n63097 ;
  assign n63093 = n62530 & ~n62564 ;
  assign n63094 = ~n62552 & n62714 ;
  assign n63095 = ~n63093 & ~n63094 ;
  assign n63099 = ~n62544 & ~n63095 ;
  assign n63100 = ~n63098 & n63099 ;
  assign n63102 = ~n62548 & ~n62728 ;
  assign n63103 = n62530 & ~n63102 ;
  assign n63105 = n62544 & ~n62707 ;
  assign n63101 = ~n62530 & n62720 ;
  assign n63104 = n62524 & n62536 ;
  assign n63106 = ~n63101 & ~n63104 ;
  assign n63107 = n63105 & n63106 ;
  assign n63108 = ~n63103 & n63107 ;
  assign n63109 = ~n63100 & ~n63108 ;
  assign n63110 = ~n63092 & ~n63109 ;
  assign n63111 = ~\u0_L6_reg[3]/NET0131  & ~n63110 ;
  assign n63112 = \u0_L6_reg[3]/NET0131  & n63110 ;
  assign n63113 = ~n63111 & ~n63112 ;
  assign n63114 = ~n62014 & n62024 ;
  assign n63115 = n61979 & ~n62047 ;
  assign n63116 = n62448 & ~n63115 ;
  assign n63117 = n62001 & ~n62448 ;
  assign n63118 = ~n63116 & ~n63117 ;
  assign n63119 = n63114 & ~n63118 ;
  assign n63121 = ~n62001 & ~n62005 ;
  assign n63122 = n62448 & n63121 ;
  assign n63120 = n62014 & ~n62024 ;
  assign n63123 = ~n63114 & ~n63120 ;
  assign n63124 = ~n63117 & n63123 ;
  assign n63125 = ~n63122 & n63124 ;
  assign n63126 = ~n63119 & ~n63125 ;
  assign n63127 = ~n62034 & ~n63126 ;
  assign n63128 = n61979 & n61998 ;
  assign n63129 = n62047 & n63128 ;
  assign n63130 = ~n62002 & n63120 ;
  assign n63131 = ~n63129 & n63130 ;
  assign n63132 = n62467 & ~n62950 ;
  assign n63133 = n63131 & n63132 ;
  assign n63134 = ~n63127 & ~n63133 ;
  assign n63135 = ~\u0_L6_reg[7]/NET0131  & n63134 ;
  assign n63136 = \u0_L6_reg[7]/NET0131  & ~n63134 ;
  assign n63137 = ~n63135 & ~n63136 ;
  assign n63149 = ~n61865 & n62382 ;
  assign n63142 = n61790 & n61836 ;
  assign n63147 = ~n61797 & ~n63142 ;
  assign n63148 = n61833 & ~n63147 ;
  assign n63150 = ~n62398 & ~n63148 ;
  assign n63151 = ~n63149 & n63150 ;
  assign n63152 = n61824 & ~n63151 ;
  assign n63138 = ~n61816 & ~n61846 ;
  assign n63139 = ~n62382 & ~n63138 ;
  assign n63140 = n61803 & ~n62378 ;
  assign n63141 = n62633 & n63140 ;
  assign n63143 = n62648 & ~n63142 ;
  assign n63144 = ~n63141 & ~n63143 ;
  assign n63145 = ~n63139 & ~n63144 ;
  assign n63146 = ~n61824 & ~n63145 ;
  assign n63153 = n61790 & n61837 ;
  assign n63154 = ~n61851 & n63153 ;
  assign n63155 = ~n63146 & ~n63154 ;
  assign n63156 = ~n63152 & n63155 ;
  assign n63157 = ~\u0_L6_reg[9]/NET0131  & ~n63156 ;
  assign n63158 = \u0_L6_reg[9]/NET0131  & n63156 ;
  assign n63159 = ~n63157 & ~n63158 ;
  assign n63172 = ~n62312 & ~n62323 ;
  assign n63174 = n62295 & ~n63172 ;
  assign n63168 = ~n62290 & ~n62329 ;
  assign n63173 = n63168 & n63172 ;
  assign n63175 = ~n62320 & ~n62667 ;
  assign n63176 = ~n63173 & n63175 ;
  assign n63177 = ~n63174 & n63176 ;
  assign n63178 = ~n62257 & ~n63177 ;
  assign n63165 = n62282 & n62299 ;
  assign n63166 = ~n62314 & ~n63165 ;
  assign n63167 = n62257 & ~n63166 ;
  assign n63160 = ~n62270 & ~n62319 ;
  assign n63161 = n62257 & n62290 ;
  assign n63162 = ~n63160 & n63161 ;
  assign n63163 = ~n62292 & ~n63162 ;
  assign n63164 = ~n62282 & ~n63163 ;
  assign n63169 = ~n62270 & n62282 ;
  assign n63170 = ~n62674 & n63169 ;
  assign n63171 = ~n63168 & n63170 ;
  assign n63179 = ~n63164 & ~n63171 ;
  assign n63180 = ~n63167 & n63179 ;
  assign n63181 = ~n63178 & n63180 ;
  assign n63182 = \u0_L6_reg[18]/NET0131  & n63181 ;
  assign n63183 = ~\u0_L6_reg[18]/NET0131  & ~n63181 ;
  assign n63184 = ~n63182 & ~n63183 ;
  assign n63188 = n63035 & n63041 ;
  assign n63189 = ~n63035 & ~n63041 ;
  assign n63190 = ~n63188 & ~n63189 ;
  assign n63191 = ~n63040 & ~n63190 ;
  assign n63192 = n63038 & n63065 ;
  assign n63193 = ~n63191 & ~n63192 ;
  assign n63194 = ~n63028 & ~n63193 ;
  assign n63185 = ~n63028 & n63056 ;
  assign n63186 = ~n63063 & ~n63185 ;
  assign n63187 = ~n63009 & ~n63186 ;
  assign n63195 = ~n63036 & ~n63187 ;
  assign n63196 = ~n63194 & n63195 ;
  assign n63197 = n63050 & ~n63196 ;
  assign n63198 = n63009 & ~n63080 ;
  assign n63199 = ~n63015 & ~n63035 ;
  assign n63200 = n63021 & n63199 ;
  assign n63201 = ~n63079 & ~n63188 ;
  assign n63202 = ~n63200 & n63201 ;
  assign n63203 = ~n63198 & ~n63202 ;
  assign n63204 = n63009 & ~n63040 ;
  assign n63205 = n63190 & n63204 ;
  assign n63206 = ~n63203 & ~n63205 ;
  assign n63207 = ~n63050 & ~n63206 ;
  assign n63208 = ~n63035 & n63063 ;
  assign n63209 = ~n63057 & ~n63208 ;
  assign n63210 = n63009 & ~n63209 ;
  assign n63211 = n63015 & n63028 ;
  assign n63212 = ~n63035 & n63211 ;
  assign n63213 = ~n63009 & n63212 ;
  assign n63214 = ~n63210 & ~n63213 ;
  assign n63215 = ~n63207 & n63214 ;
  assign n63216 = ~n63197 & n63215 ;
  assign n63217 = ~\u0_L6_reg[16]/NET0131  & ~n63216 ;
  assign n63218 = \u0_L6_reg[16]/NET0131  & n63216 ;
  assign n63219 = ~n63217 & ~n63218 ;
  assign n63220 = ~n63009 & ~n63211 ;
  assign n63221 = n63035 & n63040 ;
  assign n63222 = n63220 & ~n63221 ;
  assign n63223 = n63022 & ~n63028 ;
  assign n63224 = n63009 & ~n63063 ;
  assign n63225 = ~n63223 & n63224 ;
  assign n63226 = n63039 & n63056 ;
  assign n63227 = n63225 & ~n63226 ;
  assign n63228 = ~n63222 & ~n63227 ;
  assign n63229 = n63050 & ~n63228 ;
  assign n63234 = ~n63065 & n63211 ;
  assign n63235 = ~n63021 & n63054 ;
  assign n63236 = ~n63234 & ~n63235 ;
  assign n63237 = n63009 & ~n63236 ;
  assign n63230 = ~n63015 & n63074 ;
  assign n63238 = ~n63050 & ~n63230 ;
  assign n63231 = n63039 & ~n63042 ;
  assign n63232 = ~n63065 & ~n63199 ;
  assign n63233 = n63220 & n63232 ;
  assign n63239 = ~n63231 & ~n63233 ;
  assign n63240 = n63238 & n63239 ;
  assign n63241 = ~n63237 & n63240 ;
  assign n63242 = ~n63229 & ~n63241 ;
  assign n63247 = n63009 & n63015 ;
  assign n63248 = n63074 & n63247 ;
  assign n63243 = ~n63009 & n63028 ;
  assign n63244 = n63065 & n63243 ;
  assign n63245 = ~n63041 & n63050 ;
  assign n63246 = n63051 & n63245 ;
  assign n63249 = ~n63244 & ~n63246 ;
  assign n63250 = ~n63248 & n63249 ;
  assign n63251 = ~n63242 & n63250 ;
  assign n63252 = \u0_L6_reg[30]/NET0131  & ~n63251 ;
  assign n63253 = ~\u0_L6_reg[30]/NET0131  & n63251 ;
  assign n63254 = ~n63252 & ~n63253 ;
  assign n63256 = ~n63009 & n63076 ;
  assign n63255 = ~n63021 & n63212 ;
  assign n63257 = ~n63231 & ~n63255 ;
  assign n63258 = n63256 & n63257 ;
  assign n63259 = ~n63212 & ~n63221 ;
  assign n63260 = n63225 & n63259 ;
  assign n63261 = ~n63258 & ~n63260 ;
  assign n63262 = ~n63050 & ~n63261 ;
  assign n63264 = n63009 & ~n63028 ;
  assign n63265 = ~n63022 & ~n63035 ;
  assign n63266 = n63264 & n63265 ;
  assign n63270 = ~n63044 & n63050 ;
  assign n63271 = ~n63266 & n63270 ;
  assign n63263 = ~n63009 & n63052 ;
  assign n63267 = n63035 & n63211 ;
  assign n63268 = ~n63029 & ~n63267 ;
  assign n63269 = n63009 & ~n63268 ;
  assign n63272 = ~n63263 & ~n63269 ;
  assign n63273 = n63271 & n63272 ;
  assign n63274 = ~n63262 & ~n63273 ;
  assign n63275 = n63188 & n63243 ;
  assign n63276 = ~n63041 & n63264 ;
  assign n63277 = n63232 & n63276 ;
  assign n63278 = ~n63275 & ~n63277 ;
  assign n63279 = ~n63274 & n63278 ;
  assign n63280 = ~\u0_L6_reg[24]/NET0131  & ~n63279 ;
  assign n63281 = \u0_L6_reg[24]/NET0131  & n63279 ;
  assign n63282 = ~n63280 & ~n63281 ;
  assign n63283 = decrypt_pad & ~\u0_uk_K_r5_reg[44]/NET0131  ;
  assign n63284 = ~decrypt_pad & ~\u0_uk_K_r5_reg[9]/NET0131  ;
  assign n63285 = ~n63283 & ~n63284 ;
  assign n63286 = \u0_R5_reg[28]/NET0131  & ~n63285 ;
  assign n63287 = ~\u0_R5_reg[28]/NET0131  & n63285 ;
  assign n63288 = ~n63286 & ~n63287 ;
  assign n63319 = decrypt_pad & ~\u0_uk_K_r5_reg[2]/NET0131  ;
  assign n63320 = ~decrypt_pad & ~\u0_uk_K_r5_reg[22]/NET0131  ;
  assign n63321 = ~n63319 & ~n63320 ;
  assign n63322 = \u0_R5_reg[27]/NET0131  & ~n63321 ;
  assign n63323 = ~\u0_R5_reg[27]/NET0131  & n63321 ;
  assign n63324 = ~n63322 & ~n63323 ;
  assign n63289 = decrypt_pad & ~\u0_uk_K_r5_reg[28]/NET0131  ;
  assign n63290 = ~decrypt_pad & ~\u0_uk_K_r5_reg[52]/NET0131  ;
  assign n63291 = ~n63289 & ~n63290 ;
  assign n63292 = \u0_R5_reg[24]/NET0131  & ~n63291 ;
  assign n63293 = ~\u0_R5_reg[24]/NET0131  & n63291 ;
  assign n63294 = ~n63292 & ~n63293 ;
  assign n63295 = decrypt_pad & ~\u0_uk_K_r5_reg[52]/NET0131  ;
  assign n63296 = ~decrypt_pad & ~\u0_uk_K_r5_reg[44]/NET0131  ;
  assign n63297 = ~n63295 & ~n63296 ;
  assign n63298 = \u0_R5_reg[26]/NET0131  & ~n63297 ;
  assign n63299 = ~\u0_R5_reg[26]/NET0131  & n63297 ;
  assign n63300 = ~n63298 & ~n63299 ;
  assign n63302 = decrypt_pad & ~\u0_uk_K_r5_reg[36]/NET0131  ;
  assign n63303 = ~decrypt_pad & ~\u0_uk_K_r5_reg[1]/NET0131  ;
  assign n63304 = ~n63302 & ~n63303 ;
  assign n63305 = \u0_R5_reg[29]/NET0131  & ~n63304 ;
  assign n63306 = ~\u0_R5_reg[29]/NET0131  & n63304 ;
  assign n63307 = ~n63305 & ~n63306 ;
  assign n63308 = decrypt_pad & ~\u0_uk_K_r5_reg[8]/NET0131  ;
  assign n63309 = ~decrypt_pad & ~\u0_uk_K_r5_reg[28]/NET0131  ;
  assign n63310 = ~n63308 & ~n63309 ;
  assign n63311 = \u0_R5_reg[25]/NET0131  & ~n63310 ;
  assign n63312 = ~\u0_R5_reg[25]/NET0131  & n63310 ;
  assign n63313 = ~n63311 & ~n63312 ;
  assign n63314 = ~n63307 & ~n63313 ;
  assign n63357 = n63300 & n63314 ;
  assign n63358 = ~n63294 & n63357 ;
  assign n63355 = n63294 & n63313 ;
  assign n63356 = ~n63307 & n63355 ;
  assign n63325 = n63294 & n63307 ;
  assign n63359 = n63300 & n63325 ;
  assign n63360 = ~n63356 & ~n63359 ;
  assign n63361 = ~n63358 & n63360 ;
  assign n63362 = ~n63324 & ~n63361 ;
  assign n63326 = ~n63300 & ~n63313 ;
  assign n63332 = n63294 & n63324 ;
  assign n63366 = n63294 & ~n63307 ;
  assign n63367 = ~n63332 & ~n63366 ;
  assign n63368 = n63326 & ~n63367 ;
  assign n63317 = ~n63294 & n63307 ;
  assign n63363 = ~n63300 & ~n63324 ;
  assign n63364 = n63317 & n63363 ;
  assign n63328 = n63307 & n63313 ;
  assign n63301 = ~n63294 & ~n63300 ;
  assign n63344 = n63294 & n63300 ;
  assign n63345 = ~n63301 & ~n63344 ;
  assign n63365 = n63328 & ~n63345 ;
  assign n63369 = ~n63364 & ~n63365 ;
  assign n63370 = ~n63368 & n63369 ;
  assign n63371 = ~n63362 & n63370 ;
  assign n63372 = ~n63288 & ~n63371 ;
  assign n63327 = n63325 & n63326 ;
  assign n63329 = ~n63294 & n63328 ;
  assign n63330 = ~n63327 & ~n63329 ;
  assign n63331 = ~n63324 & ~n63330 ;
  assign n63333 = n63300 & n63313 ;
  assign n63334 = ~n63326 & ~n63333 ;
  assign n63335 = ~n63300 & ~n63307 ;
  assign n63336 = n63332 & ~n63335 ;
  assign n63337 = n63334 & n63336 ;
  assign n63315 = n63301 & n63314 ;
  assign n63316 = n63300 & ~n63313 ;
  assign n63318 = n63316 & n63317 ;
  assign n63338 = ~n63315 & ~n63318 ;
  assign n63339 = ~n63337 & n63338 ;
  assign n63340 = ~n63331 & n63339 ;
  assign n63341 = n63288 & ~n63340 ;
  assign n63349 = ~n63294 & ~n63307 ;
  assign n63350 = n63313 & n63349 ;
  assign n63351 = n63300 & n63350 ;
  assign n63348 = n63294 & n63314 ;
  assign n63352 = ~n63318 & ~n63348 ;
  assign n63353 = ~n63351 & n63352 ;
  assign n63354 = n63324 & ~n63353 ;
  assign n63342 = ~n63313 & n63324 ;
  assign n63343 = n63335 & n63342 ;
  assign n63346 = n63313 & ~n63324 ;
  assign n63347 = ~n63345 & n63346 ;
  assign n63373 = ~n63343 & ~n63347 ;
  assign n63374 = ~n63354 & n63373 ;
  assign n63375 = ~n63341 & n63374 ;
  assign n63376 = ~n63372 & n63375 ;
  assign n63377 = ~\u0_L5_reg[22]/NET0131  & ~n63376 ;
  assign n63378 = \u0_L5_reg[22]/NET0131  & n63376 ;
  assign n63379 = ~n63377 & ~n63378 ;
  assign n63414 = decrypt_pad & ~\u0_uk_K_r5_reg[11]/NET0131  ;
  assign n63415 = ~decrypt_pad & ~\u0_uk_K_r5_reg[33]/NET0131  ;
  assign n63416 = ~n63414 & ~n63415 ;
  assign n63417 = \u0_R5_reg[4]/NET0131  & ~n63416 ;
  assign n63418 = ~\u0_R5_reg[4]/NET0131  & n63416 ;
  assign n63419 = ~n63417 & ~n63418 ;
  assign n63405 = decrypt_pad & ~\u0_uk_K_r5_reg[20]/NET0131  ;
  assign n63406 = ~decrypt_pad & ~\u0_uk_K_r5_reg[10]/NET0131  ;
  assign n63407 = ~n63405 & ~n63406 ;
  assign n63408 = \u0_R5_reg[32]/NET0131  & ~n63407 ;
  assign n63409 = ~\u0_R5_reg[32]/NET0131  & n63407 ;
  assign n63410 = ~n63408 & ~n63409 ;
  assign n63380 = decrypt_pad & ~\u0_uk_K_r5_reg[41]/NET0131  ;
  assign n63381 = ~decrypt_pad & ~\u0_uk_K_r5_reg[6]/NET0131  ;
  assign n63382 = ~n63380 & ~n63381 ;
  assign n63383 = \u0_R5_reg[1]/NET0131  & ~n63382 ;
  assign n63384 = ~\u0_R5_reg[1]/NET0131  & n63382 ;
  assign n63385 = ~n63383 & ~n63384 ;
  assign n63392 = decrypt_pad & ~\u0_uk_K_r5_reg[24]/NET0131  ;
  assign n63393 = ~decrypt_pad & ~\u0_uk_K_r5_reg[46]/NET0131  ;
  assign n63394 = ~n63392 & ~n63393 ;
  assign n63395 = \u0_R5_reg[2]/NET0131  & ~n63394 ;
  assign n63396 = ~\u0_R5_reg[2]/NET0131  & n63394 ;
  assign n63397 = ~n63395 & ~n63396 ;
  assign n63399 = decrypt_pad & ~\u0_uk_K_r5_reg[39]/NET0131  ;
  assign n63400 = ~decrypt_pad & ~\u0_uk_K_r5_reg[4]/NET0131  ;
  assign n63401 = ~n63399 & ~n63400 ;
  assign n63402 = \u0_R5_reg[5]/NET0131  & ~n63401 ;
  assign n63403 = ~\u0_R5_reg[5]/NET0131  & n63401 ;
  assign n63404 = ~n63402 & ~n63403 ;
  assign n63450 = ~n63397 & ~n63404 ;
  assign n63451 = ~n63385 & n63450 ;
  assign n63452 = n63410 & ~n63451 ;
  assign n63411 = ~n63404 & ~n63410 ;
  assign n63386 = decrypt_pad & ~\u0_uk_K_r5_reg[33]/NET0131  ;
  assign n63387 = ~decrypt_pad & ~\u0_uk_K_r5_reg[55]/NET0131  ;
  assign n63388 = ~n63386 & ~n63387 ;
  assign n63389 = \u0_R5_reg[3]/NET0131  & ~n63388 ;
  assign n63390 = ~\u0_R5_reg[3]/NET0131  & n63388 ;
  assign n63391 = ~n63389 & ~n63390 ;
  assign n63448 = n63391 & ~n63397 ;
  assign n63449 = n63385 & ~n63448 ;
  assign n63453 = ~n63411 & ~n63449 ;
  assign n63454 = ~n63452 & n63453 ;
  assign n63427 = ~n63385 & n63404 ;
  assign n63441 = n63397 & ~n63410 ;
  assign n63442 = ~n63404 & n63441 ;
  assign n63443 = ~n63427 & ~n63442 ;
  assign n63444 = n63391 & ~n63443 ;
  assign n63445 = n63385 & ~n63410 ;
  assign n63432 = n63385 & ~n63391 ;
  assign n63446 = ~n63432 & ~n63441 ;
  assign n63447 = ~n63445 & ~n63446 ;
  assign n63455 = ~n63444 & ~n63447 ;
  assign n63456 = ~n63454 & n63455 ;
  assign n63457 = n63419 & ~n63456 ;
  assign n63424 = ~n63385 & n63410 ;
  assign n63425 = ~n63404 & n63424 ;
  assign n63426 = n63397 & n63425 ;
  assign n63428 = ~n63397 & ~n63410 ;
  assign n63429 = ~n63427 & n63428 ;
  assign n63430 = ~n63426 & ~n63429 ;
  assign n63431 = ~n63391 & ~n63430 ;
  assign n63398 = n63391 & n63397 ;
  assign n63420 = n63404 & n63410 ;
  assign n63421 = ~n63411 & ~n63420 ;
  assign n63422 = n63385 & n63421 ;
  assign n63423 = n63398 & n63422 ;
  assign n63433 = n63420 & ~n63432 ;
  assign n63434 = n63385 & ~n63404 ;
  assign n63435 = ~n63410 & n63434 ;
  assign n63436 = ~n63433 & ~n63435 ;
  assign n63437 = ~n63397 & ~n63436 ;
  assign n63438 = ~n63423 & ~n63437 ;
  assign n63439 = ~n63431 & n63438 ;
  assign n63440 = ~n63419 & ~n63439 ;
  assign n63459 = n63385 & n63420 ;
  assign n63460 = n63397 & n63459 ;
  assign n63461 = n63427 & n63441 ;
  assign n63462 = ~n63397 & n63434 ;
  assign n63463 = ~n63461 & ~n63462 ;
  assign n63464 = ~n63460 & n63463 ;
  assign n63465 = ~n63391 & ~n63464 ;
  assign n63412 = ~n63385 & n63398 ;
  assign n63413 = n63411 & n63412 ;
  assign n63458 = n63424 & n63448 ;
  assign n63466 = ~n63413 & ~n63458 ;
  assign n63467 = ~n63465 & n63466 ;
  assign n63468 = ~n63440 & n63467 ;
  assign n63469 = ~n63457 & n63468 ;
  assign n63470 = ~\u0_L5_reg[31]/NET0131  & ~n63469 ;
  assign n63471 = \u0_L5_reg[31]/NET0131  & n63469 ;
  assign n63472 = ~n63470 & ~n63471 ;
  assign n63521 = decrypt_pad & ~\u0_uk_K_r5_reg[37]/P0001  ;
  assign n63522 = ~decrypt_pad & ~\u0_uk_K_r5_reg[2]/NET0131  ;
  assign n63523 = ~n63521 & ~n63522 ;
  assign n63524 = \u0_R5_reg[24]/NET0131  & ~n63523 ;
  assign n63525 = ~\u0_R5_reg[24]/NET0131  & n63523 ;
  assign n63526 = ~n63524 & ~n63525 ;
  assign n63486 = decrypt_pad & ~\u0_uk_K_r5_reg[22]/NET0131  ;
  assign n63487 = ~decrypt_pad & ~\u0_uk_K_r5_reg[42]/NET0131  ;
  assign n63488 = ~n63486 & ~n63487 ;
  assign n63489 = \u0_R5_reg[22]/NET0131  & ~n63488 ;
  assign n63490 = ~\u0_R5_reg[22]/NET0131  & n63488 ;
  assign n63491 = ~n63489 & ~n63490 ;
  assign n63473 = decrypt_pad & ~\u0_uk_K_r5_reg[1]/NET0131  ;
  assign n63474 = ~decrypt_pad & ~\u0_uk_K_r5_reg[21]/NET0131  ;
  assign n63475 = ~n63473 & ~n63474 ;
  assign n63476 = \u0_R5_reg[25]/NET0131  & ~n63475 ;
  assign n63477 = ~\u0_R5_reg[25]/NET0131  & n63475 ;
  assign n63478 = ~n63476 & ~n63477 ;
  assign n63479 = decrypt_pad & ~\u0_uk_K_r5_reg[16]/NET0131  ;
  assign n63480 = ~decrypt_pad & ~\u0_uk_K_r5_reg[36]/NET0131  ;
  assign n63481 = ~n63479 & ~n63480 ;
  assign n63482 = \u0_R5_reg[20]/NET0131  & ~n63481 ;
  assign n63483 = ~\u0_R5_reg[20]/NET0131  & n63481 ;
  assign n63484 = ~n63482 & ~n63483 ;
  assign n63485 = n63478 & n63484 ;
  assign n63493 = decrypt_pad & ~\u0_uk_K_r5_reg[0]/NET0131  ;
  assign n63494 = ~decrypt_pad & ~\u0_uk_K_r5_reg[51]/NET0131  ;
  assign n63495 = ~n63493 & ~n63494 ;
  assign n63496 = \u0_R5_reg[21]/NET0131  & ~n63495 ;
  assign n63497 = ~\u0_R5_reg[21]/NET0131  & n63495 ;
  assign n63498 = ~n63496 & ~n63497 ;
  assign n63499 = ~n63484 & n63498 ;
  assign n63558 = ~n63485 & ~n63499 ;
  assign n63559 = n63491 & ~n63558 ;
  assign n63503 = decrypt_pad & ~\u0_uk_K_r5_reg[35]/NET0131  ;
  assign n63504 = ~decrypt_pad & ~\u0_uk_K_r5_reg[0]/NET0131  ;
  assign n63505 = ~n63503 & ~n63504 ;
  assign n63506 = \u0_R5_reg[23]/NET0131  & ~n63505 ;
  assign n63507 = ~\u0_R5_reg[23]/NET0131  & n63505 ;
  assign n63508 = ~n63506 & ~n63507 ;
  assign n63555 = n63478 & n63498 ;
  assign n63556 = ~n63484 & n63555 ;
  assign n63557 = ~n63491 & ~n63556 ;
  assign n63560 = ~n63508 & ~n63557 ;
  assign n63561 = ~n63559 & n63560 ;
  assign n63516 = ~n63478 & n63484 ;
  assign n63547 = ~n63498 & n63516 ;
  assign n63548 = ~n63491 & n63547 ;
  assign n63527 = n63491 & n63499 ;
  assign n63549 = n63485 & n63498 ;
  assign n63550 = ~n63527 & ~n63549 ;
  assign n63551 = ~n63548 & n63550 ;
  assign n63552 = n63508 & ~n63551 ;
  assign n63510 = ~n63491 & ~n63508 ;
  assign n63553 = n63485 & n63510 ;
  assign n63554 = ~n63498 & n63553 ;
  assign n63562 = ~n63552 & ~n63554 ;
  assign n63563 = ~n63561 & n63562 ;
  assign n63564 = n63526 & ~n63563 ;
  assign n63528 = ~n63491 & n63498 ;
  assign n63529 = n63484 & n63528 ;
  assign n63530 = ~n63527 & ~n63529 ;
  assign n63531 = ~n63508 & ~n63530 ;
  assign n63533 = n63484 & ~n63498 ;
  assign n63534 = n63491 & n63508 ;
  assign n63535 = n63533 & n63534 ;
  assign n63536 = n63516 & n63528 ;
  assign n63540 = ~n63535 & ~n63536 ;
  assign n63537 = n63510 & n63516 ;
  assign n63538 = ~n63484 & ~n63491 ;
  assign n63539 = n63508 & n63538 ;
  assign n63541 = ~n63537 & ~n63539 ;
  assign n63542 = n63540 & n63541 ;
  assign n63511 = ~n63484 & ~n63498 ;
  assign n63514 = n63478 & n63511 ;
  assign n63515 = n63508 & n63514 ;
  assign n63492 = n63485 & n63491 ;
  assign n63532 = n63492 & ~n63498 ;
  assign n63543 = ~n63515 & ~n63532 ;
  assign n63544 = n63542 & n63543 ;
  assign n63545 = ~n63531 & n63544 ;
  assign n63546 = ~n63526 & ~n63545 ;
  assign n63517 = n63498 & n63516 ;
  assign n63518 = ~n63508 & n63517 ;
  assign n63519 = ~n63515 & ~n63518 ;
  assign n63520 = ~n63491 & ~n63519 ;
  assign n63500 = ~n63478 & n63499 ;
  assign n63501 = ~n63491 & n63500 ;
  assign n63502 = ~n63492 & ~n63501 ;
  assign n63509 = ~n63502 & n63508 ;
  assign n63512 = ~n63478 & n63511 ;
  assign n63513 = n63510 & n63512 ;
  assign n63565 = ~n63509 & ~n63513 ;
  assign n63566 = ~n63520 & n63565 ;
  assign n63567 = ~n63546 & n63566 ;
  assign n63568 = ~n63564 & n63567 ;
  assign n63569 = \u0_L5_reg[11]/NET0131  & ~n63568 ;
  assign n63570 = ~\u0_L5_reg[11]/NET0131  & n63568 ;
  assign n63571 = ~n63569 & ~n63570 ;
  assign n63578 = decrypt_pad & ~\u0_uk_K_r5_reg[54]/NET0131  ;
  assign n63579 = ~decrypt_pad & ~\u0_uk_K_r5_reg[19]/NET0131  ;
  assign n63580 = ~n63578 & ~n63579 ;
  assign n63581 = \u0_R5_reg[14]/NET0131  & ~n63580 ;
  assign n63582 = ~\u0_R5_reg[14]/NET0131  & n63580 ;
  assign n63583 = ~n63581 & ~n63582 ;
  assign n63585 = decrypt_pad & ~\u0_uk_K_r5_reg[53]/NET0131  ;
  assign n63586 = ~decrypt_pad & ~\u0_uk_K_r5_reg[18]/NET0131  ;
  assign n63587 = ~n63585 & ~n63586 ;
  assign n63588 = \u0_R5_reg[13]/NET0131  & ~n63587 ;
  assign n63589 = ~\u0_R5_reg[13]/NET0131  & n63587 ;
  assign n63590 = ~n63588 & ~n63589 ;
  assign n63591 = decrypt_pad & ~\u0_uk_K_r5_reg[34]/NET0131  ;
  assign n63592 = ~decrypt_pad & ~\u0_uk_K_r5_reg[24]/NET0131  ;
  assign n63593 = ~n63591 & ~n63592 ;
  assign n63594 = \u0_R5_reg[12]/NET0131  & ~n63593 ;
  assign n63595 = ~\u0_R5_reg[12]/NET0131  & n63593 ;
  assign n63596 = ~n63594 & ~n63595 ;
  assign n63601 = decrypt_pad & ~\u0_uk_K_r5_reg[18]/NET0131  ;
  assign n63602 = ~decrypt_pad & ~\u0_uk_K_r5_reg[40]/NET0131  ;
  assign n63603 = ~n63601 & ~n63602 ;
  assign n63604 = \u0_R5_reg[17]/NET0131  & ~n63603 ;
  assign n63605 = ~\u0_R5_reg[17]/NET0131  & n63603 ;
  assign n63606 = ~n63604 & ~n63605 ;
  assign n63626 = n63596 & n63606 ;
  assign n63627 = n63590 & n63626 ;
  assign n63628 = n63583 & n63627 ;
  assign n63572 = decrypt_pad & ~\u0_uk_K_r5_reg[5]/NET0131  ;
  assign n63573 = ~decrypt_pad & ~\u0_uk_K_r5_reg[27]/NET0131  ;
  assign n63574 = ~n63572 & ~n63573 ;
  assign n63575 = \u0_R5_reg[15]/NET0131  & ~n63574 ;
  assign n63576 = ~\u0_R5_reg[15]/NET0131  & n63574 ;
  assign n63577 = ~n63575 & ~n63576 ;
  assign n63607 = ~n63596 & n63606 ;
  assign n63608 = n63577 & n63607 ;
  assign n63609 = ~n63590 & n63608 ;
  assign n63620 = n63577 & n63590 ;
  assign n63621 = n63596 & ~n63606 ;
  assign n63622 = n63620 & n63621 ;
  assign n63623 = ~n63583 & n63590 ;
  assign n63624 = n63607 & n63623 ;
  assign n63625 = ~n63622 & ~n63624 ;
  assign n63630 = ~n63609 & n63625 ;
  assign n63631 = ~n63628 & n63630 ;
  assign n63616 = ~n63590 & ~n63606 ;
  assign n63617 = ~n63596 & n63616 ;
  assign n63618 = ~n63577 & n63617 ;
  assign n63619 = n63583 & n63618 ;
  assign n63584 = ~n63577 & ~n63583 ;
  assign n63597 = n63590 & ~n63596 ;
  assign n63598 = ~n63590 & n63596 ;
  assign n63599 = ~n63597 & ~n63598 ;
  assign n63600 = n63584 & ~n63599 ;
  assign n63610 = decrypt_pad & ~\u0_uk_K_r5_reg[13]/P0001  ;
  assign n63611 = ~decrypt_pad & ~\u0_uk_K_r5_reg[3]/NET0131  ;
  assign n63612 = ~n63610 & ~n63611 ;
  assign n63613 = \u0_R5_reg[16]/NET0131  & ~n63612 ;
  assign n63614 = ~\u0_R5_reg[16]/NET0131  & n63612 ;
  assign n63615 = ~n63613 & ~n63614 ;
  assign n63629 = ~n63600 & n63615 ;
  assign n63632 = ~n63619 & n63629 ;
  assign n63633 = n63631 & n63632 ;
  assign n63636 = n63577 & ~n63617 ;
  assign n63637 = ~n63627 & n63636 ;
  assign n63639 = n63583 & n63621 ;
  assign n63638 = ~n63590 & n63606 ;
  assign n63640 = ~n63577 & ~n63638 ;
  assign n63641 = ~n63639 & n63640 ;
  assign n63642 = ~n63637 & ~n63641 ;
  assign n63643 = ~n63583 & n63598 ;
  assign n63644 = n63606 & n63643 ;
  assign n63634 = ~n63583 & ~n63596 ;
  assign n63635 = n63616 & n63634 ;
  assign n63649 = ~n63615 & ~n63635 ;
  assign n63650 = ~n63644 & n63649 ;
  assign n63645 = n63583 & n63620 ;
  assign n63646 = ~n63596 & n63645 ;
  assign n63647 = n63597 & ~n63606 ;
  assign n63648 = n63583 & n63647 ;
  assign n63651 = ~n63646 & ~n63648 ;
  assign n63652 = n63650 & n63651 ;
  assign n63653 = ~n63642 & n63652 ;
  assign n63654 = ~n63633 & ~n63653 ;
  assign n63655 = ~n63577 & ~n63624 ;
  assign n63656 = n63583 & ~n63590 ;
  assign n63657 = n63621 & n63656 ;
  assign n63658 = n63577 & ~n63657 ;
  assign n63659 = ~n63635 & n63658 ;
  assign n63660 = ~n63655 & ~n63659 ;
  assign n63661 = ~n63583 & n63622 ;
  assign n63662 = ~n63660 & ~n63661 ;
  assign n63663 = ~n63654 & n63662 ;
  assign n63664 = ~\u0_L5_reg[20]/NET0131  & ~n63663 ;
  assign n63665 = \u0_L5_reg[20]/NET0131  & n63663 ;
  assign n63666 = ~n63664 & ~n63665 ;
  assign n63667 = decrypt_pad & ~\u0_uk_K_r5_reg[42]/NET0131  ;
  assign n63668 = ~decrypt_pad & ~\u0_uk_K_r5_reg[7]/NET0131  ;
  assign n63669 = ~n63667 & ~n63668 ;
  assign n63670 = \u0_R5_reg[28]/NET0131  & ~n63669 ;
  assign n63671 = ~\u0_R5_reg[28]/NET0131  & n63669 ;
  assign n63672 = ~n63670 & ~n63671 ;
  assign n63680 = decrypt_pad & ~\u0_uk_K_r5_reg[15]/NET0131  ;
  assign n63681 = ~decrypt_pad & ~\u0_uk_K_r5_reg[35]/NET0131  ;
  assign n63682 = ~n63680 & ~n63681 ;
  assign n63683 = \u0_R5_reg[30]/NET0131  & ~n63682 ;
  assign n63684 = ~\u0_R5_reg[30]/NET0131  & n63682 ;
  assign n63685 = ~n63683 & ~n63684 ;
  assign n63673 = decrypt_pad & ~\u0_uk_K_r5_reg[14]/NET0131  ;
  assign n63674 = ~decrypt_pad & ~\u0_uk_K_r5_reg[38]/NET0131  ;
  assign n63675 = ~n63673 & ~n63674 ;
  assign n63676 = \u0_R5_reg[29]/NET0131  & ~n63675 ;
  assign n63677 = ~\u0_R5_reg[29]/NET0131  & n63675 ;
  assign n63678 = ~n63676 & ~n63677 ;
  assign n63687 = decrypt_pad & ~\u0_uk_K_r5_reg[30]/NET0131  ;
  assign n63688 = ~decrypt_pad & ~\u0_uk_K_r5_reg[50]/NET0131  ;
  assign n63689 = ~n63687 & ~n63688 ;
  assign n63690 = \u0_R5_reg[1]/NET0131  & ~n63689 ;
  assign n63691 = ~\u0_R5_reg[1]/NET0131  & n63689 ;
  assign n63692 = ~n63690 & ~n63691 ;
  assign n63712 = n63678 & ~n63692 ;
  assign n63713 = ~n63685 & n63712 ;
  assign n63697 = decrypt_pad & ~\u0_uk_K_r5_reg[31]/NET0131  ;
  assign n63698 = ~decrypt_pad & ~\u0_uk_K_r5_reg[23]/NET0131  ;
  assign n63699 = ~n63697 & ~n63698 ;
  assign n63700 = \u0_R5_reg[31]/P0001  & ~n63699 ;
  assign n63701 = ~\u0_R5_reg[31]/P0001  & n63699 ;
  assign n63702 = ~n63700 & ~n63701 ;
  assign n63709 = ~n63685 & ~n63702 ;
  assign n63710 = n63685 & n63692 ;
  assign n63711 = n63678 & n63710 ;
  assign n63714 = ~n63709 & ~n63711 ;
  assign n63715 = ~n63713 & n63714 ;
  assign n63716 = n63672 & ~n63715 ;
  assign n63679 = n63672 & ~n63678 ;
  assign n63686 = n63679 & n63685 ;
  assign n63693 = n63686 & ~n63692 ;
  assign n63694 = ~n63672 & n63692 ;
  assign n63695 = ~n63678 & n63694 ;
  assign n63696 = ~n63693 & ~n63695 ;
  assign n63703 = ~n63696 & n63702 ;
  assign n63704 = ~n63672 & n63685 ;
  assign n63705 = ~n63692 & ~n63704 ;
  assign n63706 = ~n63678 & n63692 ;
  assign n63707 = ~n63702 & ~n63706 ;
  assign n63708 = ~n63705 & n63707 ;
  assign n63717 = ~n63703 & ~n63708 ;
  assign n63718 = ~n63716 & n63717 ;
  assign n63719 = decrypt_pad & ~\u0_uk_K_r5_reg[9]/NET0131  ;
  assign n63720 = ~decrypt_pad & ~\u0_uk_K_r5_reg[29]/NET0131  ;
  assign n63721 = ~n63719 & ~n63720 ;
  assign n63722 = \u0_R5_reg[32]/NET0131  & ~n63721 ;
  assign n63723 = ~\u0_R5_reg[32]/NET0131  & n63721 ;
  assign n63724 = ~n63722 & ~n63723 ;
  assign n63725 = ~n63718 & ~n63724 ;
  assign n63745 = n63672 & n63713 ;
  assign n63732 = n63672 & ~n63685 ;
  assign n63733 = ~n63712 & ~n63732 ;
  assign n63746 = n63702 & ~n63733 ;
  assign n63747 = ~n63745 & n63746 ;
  assign n63748 = ~n63672 & n63711 ;
  assign n63749 = ~n63678 & ~n63685 ;
  assign n63750 = ~n63672 & n63749 ;
  assign n63751 = ~n63702 & n63750 ;
  assign n63752 = ~n63748 & ~n63751 ;
  assign n63753 = ~n63747 & n63752 ;
  assign n63754 = n63724 & ~n63753 ;
  assign n63730 = n63672 & ~n63692 ;
  assign n63731 = n63678 & ~n63685 ;
  assign n63734 = ~n63730 & ~n63731 ;
  assign n63735 = ~n63733 & n63734 ;
  assign n63726 = ~n63678 & ~n63692 ;
  assign n63727 = ~n63672 & n63726 ;
  assign n63728 = ~n63685 & n63727 ;
  assign n63729 = n63704 & n63706 ;
  assign n63736 = ~n63728 & ~n63729 ;
  assign n63737 = ~n63735 & n63736 ;
  assign n63738 = n63702 & ~n63737 ;
  assign n63739 = n63672 & n63678 ;
  assign n63740 = ~n63692 & n63739 ;
  assign n63741 = n63709 & n63740 ;
  assign n63742 = n63685 & ~n63702 ;
  assign n63743 = n63679 & n63724 ;
  assign n63744 = n63742 & n63743 ;
  assign n63755 = ~n63741 & ~n63744 ;
  assign n63756 = ~n63738 & n63755 ;
  assign n63757 = ~n63754 & n63756 ;
  assign n63758 = ~n63725 & n63757 ;
  assign n63759 = \u0_L5_reg[5]/NET0131  & ~n63758 ;
  assign n63760 = ~\u0_L5_reg[5]/NET0131  & n63758 ;
  assign n63761 = ~n63759 & ~n63760 ;
  assign n63762 = n63391 & ~n63425 ;
  assign n63763 = ~n63459 & n63762 ;
  assign n63764 = ~n63385 & ~n63421 ;
  assign n63765 = ~n63404 & n63428 ;
  assign n63766 = ~n63391 & ~n63765 ;
  assign n63767 = ~n63764 & n63766 ;
  assign n63768 = ~n63763 & ~n63767 ;
  assign n63769 = n63397 & n63434 ;
  assign n63770 = n63410 & n63769 ;
  assign n63771 = ~n63419 & ~n63461 ;
  assign n63772 = ~n63770 & n63771 ;
  assign n63773 = ~n63768 & n63772 ;
  assign n63774 = ~n63441 & ~n63445 ;
  assign n63775 = ~n63397 & n63410 ;
  assign n63780 = n63427 & n63775 ;
  assign n63781 = n63774 & ~n63780 ;
  assign n63782 = n63391 & ~n63781 ;
  assign n63783 = n63410 & n63462 ;
  assign n63776 = ~n63391 & ~n63775 ;
  assign n63777 = n63774 & n63776 ;
  assign n63778 = n63397 & n63404 ;
  assign n63779 = n63385 & n63778 ;
  assign n63784 = n63419 & ~n63779 ;
  assign n63785 = ~n63777 & n63784 ;
  assign n63786 = ~n63783 & n63785 ;
  assign n63787 = ~n63782 & n63786 ;
  assign n63788 = ~n63773 & ~n63787 ;
  assign n63789 = n63391 & n63445 ;
  assign n63790 = ~n63450 & ~n63778 ;
  assign n63791 = n63789 & n63790 ;
  assign n63792 = ~n63788 & ~n63791 ;
  assign n63793 = ~\u0_L5_reg[17]/NET0131  & ~n63792 ;
  assign n63794 = \u0_L5_reg[17]/NET0131  & n63792 ;
  assign n63795 = ~n63793 & ~n63794 ;
  assign n63818 = ~n63547 & ~n63549 ;
  assign n63801 = ~n63478 & ~n63528 ;
  assign n63819 = n63491 & ~n63499 ;
  assign n63820 = n63801 & ~n63819 ;
  assign n63821 = n63818 & ~n63820 ;
  assign n63822 = n63508 & ~n63821 ;
  assign n63796 = n63491 & n63517 ;
  assign n63815 = ~n63491 & ~n63558 ;
  assign n63816 = ~n63796 & ~n63815 ;
  assign n63817 = ~n63508 & ~n63816 ;
  assign n63823 = n63491 & n63514 ;
  assign n63824 = ~n63817 & ~n63823 ;
  assign n63825 = ~n63822 & n63824 ;
  assign n63826 = ~n63526 & ~n63825 ;
  assign n63802 = ~n63484 & n63801 ;
  assign n63803 = ~n63492 & ~n63802 ;
  assign n63804 = ~n63508 & ~n63803 ;
  assign n63797 = ~n63478 & n63491 ;
  assign n63798 = n63499 & ~n63797 ;
  assign n63799 = ~n63796 & ~n63798 ;
  assign n63800 = n63508 & ~n63799 ;
  assign n63805 = n63478 & ~n63491 ;
  assign n63806 = ~n63797 & ~n63805 ;
  assign n63807 = n63511 & ~n63806 ;
  assign n63808 = ~n63532 & ~n63537 ;
  assign n63809 = ~n63807 & n63808 ;
  assign n63810 = ~n63800 & n63809 ;
  assign n63811 = ~n63804 & n63810 ;
  assign n63812 = n63526 & ~n63811 ;
  assign n63813 = ~n63491 & n63508 ;
  assign n63814 = n63555 & n63813 ;
  assign n63827 = ~n63548 & ~n63814 ;
  assign n63828 = ~n63812 & n63827 ;
  assign n63829 = ~n63826 & n63828 ;
  assign n63830 = \u0_L5_reg[29]/NET0131  & ~n63829 ;
  assign n63831 = ~\u0_L5_reg[29]/NET0131  & n63829 ;
  assign n63832 = ~n63830 & ~n63831 ;
  assign n63833 = decrypt_pad & ~\u0_uk_K_r5_reg[12]/NET0131  ;
  assign n63834 = ~decrypt_pad & ~\u0_uk_K_r5_reg[34]/NET0131  ;
  assign n63835 = ~n63833 & ~n63834 ;
  assign n63836 = \u0_R5_reg[8]/NET0131  & ~n63835 ;
  assign n63837 = ~\u0_R5_reg[8]/NET0131  & n63835 ;
  assign n63838 = ~n63836 & ~n63837 ;
  assign n63839 = decrypt_pad & ~\u0_uk_K_r5_reg[46]/NET0131  ;
  assign n63840 = ~decrypt_pad & ~\u0_uk_K_r5_reg[11]/NET0131  ;
  assign n63841 = ~n63839 & ~n63840 ;
  assign n63842 = \u0_R5_reg[7]/NET0131  & ~n63841 ;
  assign n63843 = ~\u0_R5_reg[7]/NET0131  & n63841 ;
  assign n63844 = ~n63842 & ~n63843 ;
  assign n63858 = decrypt_pad & ~\u0_uk_K_r5_reg[4]/NET0131  ;
  assign n63859 = ~decrypt_pad & ~\u0_uk_K_r5_reg[26]/NET0131  ;
  assign n63860 = ~n63858 & ~n63859 ;
  assign n63861 = \u0_R5_reg[5]/NET0131  & ~n63860 ;
  assign n63862 = ~\u0_R5_reg[5]/NET0131  & n63860 ;
  assign n63863 = ~n63861 & ~n63862 ;
  assign n63845 = decrypt_pad & ~\u0_uk_K_r5_reg[25]/NET0131  ;
  assign n63846 = ~decrypt_pad & ~\u0_uk_K_r5_reg[47]/NET0131  ;
  assign n63847 = ~n63845 & ~n63846 ;
  assign n63848 = \u0_R5_reg[4]/NET0131  & ~n63847 ;
  assign n63849 = ~\u0_R5_reg[4]/NET0131  & n63847 ;
  assign n63850 = ~n63848 & ~n63849 ;
  assign n63851 = decrypt_pad & ~\u0_uk_K_r5_reg[17]/NET0131  ;
  assign n63852 = ~decrypt_pad & ~\u0_uk_K_r5_reg[39]/NET0131  ;
  assign n63853 = ~n63851 & ~n63852 ;
  assign n63854 = \u0_R5_reg[9]/NET0131  & ~n63853 ;
  assign n63855 = ~\u0_R5_reg[9]/NET0131  & n63853 ;
  assign n63856 = ~n63854 & ~n63855 ;
  assign n63873 = ~n63850 & n63856 ;
  assign n63874 = ~n63863 & n63873 ;
  assign n63865 = decrypt_pad & ~\u0_uk_K_r5_reg[27]/NET0131  ;
  assign n63866 = ~decrypt_pad & ~\u0_uk_K_r5_reg[17]/NET0131  ;
  assign n63867 = ~n63865 & ~n63866 ;
  assign n63868 = \u0_R5_reg[6]/NET0131  & ~n63867 ;
  assign n63869 = ~\u0_R5_reg[6]/NET0131  & n63867 ;
  assign n63870 = ~n63868 & ~n63869 ;
  assign n63875 = n63850 & n63863 ;
  assign n63876 = n63850 & ~n63856 ;
  assign n63877 = ~n63875 & ~n63876 ;
  assign n63878 = n63870 & ~n63877 ;
  assign n63879 = ~n63874 & ~n63878 ;
  assign n63880 = ~n63844 & ~n63879 ;
  assign n63881 = ~n63856 & n63863 ;
  assign n63882 = ~n63874 & ~n63881 ;
  assign n63883 = ~n63870 & ~n63882 ;
  assign n63857 = n63850 & n63856 ;
  assign n63864 = n63857 & ~n63863 ;
  assign n63871 = n63864 & n63870 ;
  assign n63872 = n63844 & n63871 ;
  assign n63884 = ~n63844 & ~n63863 ;
  assign n63885 = n63856 & ~n63870 ;
  assign n63886 = n63884 & n63885 ;
  assign n63887 = n63863 & n63870 ;
  assign n63888 = n63873 & n63887 ;
  assign n63889 = ~n63886 & ~n63888 ;
  assign n63890 = ~n63872 & n63889 ;
  assign n63891 = ~n63883 & n63890 ;
  assign n63892 = ~n63880 & n63891 ;
  assign n63893 = ~n63838 & ~n63892 ;
  assign n63899 = ~n63863 & n63876 ;
  assign n63900 = ~n63870 & n63899 ;
  assign n63894 = ~n63850 & ~n63856 ;
  assign n63895 = n63884 & n63894 ;
  assign n63896 = ~n63850 & n63870 ;
  assign n63897 = n63844 & n63863 ;
  assign n63898 = ~n63896 & n63897 ;
  assign n63906 = ~n63895 & ~n63898 ;
  assign n63907 = ~n63900 & n63906 ;
  assign n63901 = n63857 & n63863 ;
  assign n63902 = ~n63870 & n63901 ;
  assign n63903 = ~n63844 & n63870 ;
  assign n63904 = ~n63873 & n63903 ;
  assign n63905 = n63877 & n63904 ;
  assign n63908 = ~n63902 & ~n63905 ;
  assign n63909 = n63907 & n63908 ;
  assign n63910 = n63838 & ~n63909 ;
  assign n63911 = ~n63863 & ~n63870 ;
  assign n63912 = ~n63887 & ~n63911 ;
  assign n63913 = n63873 & ~n63912 ;
  assign n63914 = ~n63844 & ~n63913 ;
  assign n63916 = ~n63863 & n63870 ;
  assign n63917 = ~n63856 & n63916 ;
  assign n63918 = ~n63850 & n63917 ;
  assign n63915 = ~n63870 & n63875 ;
  assign n63919 = n63844 & ~n63915 ;
  assign n63920 = ~n63918 & n63919 ;
  assign n63921 = ~n63914 & ~n63920 ;
  assign n63922 = ~n63910 & ~n63921 ;
  assign n63923 = ~n63893 & n63922 ;
  assign n63924 = \u0_L5_reg[2]/NET0131  & n63923 ;
  assign n63925 = ~\u0_L5_reg[2]/NET0131  & ~n63923 ;
  assign n63926 = ~n63924 & ~n63925 ;
  assign n63927 = n63577 & ~n63644 ;
  assign n63928 = ~n63647 & n63927 ;
  assign n63929 = n63621 & ~n63623 ;
  assign n63930 = n63655 & ~n63929 ;
  assign n63931 = ~n63928 & ~n63930 ;
  assign n63932 = n63607 & n63656 ;
  assign n63933 = ~n63628 & ~n63932 ;
  assign n63934 = ~n63931 & n63933 ;
  assign n63935 = n63615 & ~n63934 ;
  assign n63936 = n63599 & ~n63638 ;
  assign n63937 = ~n63608 & ~n63936 ;
  assign n63938 = ~n63583 & ~n63937 ;
  assign n63942 = n63584 & n63626 ;
  assign n63943 = ~n63618 & ~n63942 ;
  assign n63939 = ~n63616 & ~n63656 ;
  assign n63940 = n63577 & n63596 ;
  assign n63941 = ~n63939 & n63940 ;
  assign n63944 = ~n63648 & ~n63941 ;
  assign n63945 = n63943 & n63944 ;
  assign n63946 = ~n63938 & n63945 ;
  assign n63947 = ~n63615 & ~n63946 ;
  assign n63948 = ~n63635 & n63933 ;
  assign n63949 = ~n63577 & ~n63948 ;
  assign n63950 = ~n63646 & ~n63661 ;
  assign n63951 = ~n63949 & n63950 ;
  assign n63952 = ~n63947 & n63951 ;
  assign n63953 = ~n63935 & n63952 ;
  assign n63954 = ~\u0_L5_reg[10]/NET0131  & ~n63953 ;
  assign n63955 = \u0_L5_reg[10]/NET0131  & n63953 ;
  assign n63956 = ~n63954 & ~n63955 ;
  assign n63962 = ~n63317 & ~n63366 ;
  assign n63963 = n63316 & n63962 ;
  assign n63957 = ~n63333 & ~n63342 ;
  assign n63958 = n63317 & ~n63957 ;
  assign n63966 = ~n63288 & ~n63958 ;
  assign n63967 = ~n63963 & n63966 ;
  assign n63959 = ~n63328 & ~n63344 ;
  assign n63960 = ~n63314 & n63959 ;
  assign n63961 = ~n63324 & ~n63960 ;
  assign n63964 = ~n63348 & ~n63350 ;
  assign n63965 = ~n63300 & ~n63964 ;
  assign n63968 = ~n63961 & ~n63965 ;
  assign n63969 = n63967 & n63968 ;
  assign n63974 = ~n63315 & ~n63355 ;
  assign n63975 = n63324 & ~n63974 ;
  assign n63970 = n63318 & ~n63324 ;
  assign n63976 = n63288 & ~n63970 ;
  assign n63971 = ~n63325 & ~n63333 ;
  assign n63972 = n63959 & ~n63971 ;
  assign n63973 = ~n63959 & n63971 ;
  assign n63977 = ~n63972 & ~n63973 ;
  assign n63978 = n63976 & n63977 ;
  assign n63979 = ~n63975 & n63978 ;
  assign n63980 = ~n63969 & ~n63979 ;
  assign n63981 = \u0_L5_reg[12]/NET0131  & n63980 ;
  assign n63982 = ~\u0_L5_reg[12]/NET0131  & ~n63980 ;
  assign n63983 = ~n63981 & ~n63982 ;
  assign n63984 = decrypt_pad & ~\u0_uk_K_r5_reg[49]/NET0131  ;
  assign n63985 = ~decrypt_pad & ~\u0_uk_K_r5_reg[14]/NET0131  ;
  assign n63986 = ~n63984 & ~n63985 ;
  assign n63987 = \u0_R5_reg[20]/NET0131  & ~n63986 ;
  assign n63988 = ~\u0_R5_reg[20]/NET0131  & n63986 ;
  assign n63989 = ~n63987 & ~n63988 ;
  assign n63996 = decrypt_pad & ~\u0_uk_K_r5_reg[23]/NET0131  ;
  assign n63997 = ~decrypt_pad & ~\u0_uk_K_r5_reg[43]/NET0131  ;
  assign n63998 = ~n63996 & ~n63997 ;
  assign n63999 = \u0_R5_reg[18]/NET0131  & ~n63998 ;
  assign n64000 = ~\u0_R5_reg[18]/NET0131  & n63998 ;
  assign n64001 = ~n63999 & ~n64000 ;
  assign n63990 = decrypt_pad & ~\u0_uk_K_r5_reg[38]/NET0131  ;
  assign n63991 = ~decrypt_pad & ~\u0_uk_K_r5_reg[30]/NET0131  ;
  assign n63992 = ~n63990 & ~n63991 ;
  assign n63993 = \u0_R5_reg[19]/NET0131  & ~n63992 ;
  assign n63994 = ~\u0_R5_reg[19]/NET0131  & n63992 ;
  assign n63995 = ~n63993 & ~n63994 ;
  assign n64009 = decrypt_pad & ~\u0_uk_K_r5_reg[50]/NET0131  ;
  assign n64010 = ~decrypt_pad & ~\u0_uk_K_r5_reg[15]/NET0131  ;
  assign n64011 = ~n64009 & ~n64010 ;
  assign n64012 = \u0_R5_reg[21]/NET0131  & ~n64011 ;
  assign n64013 = ~\u0_R5_reg[21]/NET0131  & n64011 ;
  assign n64014 = ~n64012 & ~n64013 ;
  assign n64002 = decrypt_pad & ~\u0_uk_K_r5_reg[29]/NET0131  ;
  assign n64003 = ~decrypt_pad & ~\u0_uk_K_r5_reg[49]/NET0131  ;
  assign n64004 = ~n64002 & ~n64003 ;
  assign n64005 = \u0_R5_reg[17]/NET0131  & ~n64004 ;
  assign n64006 = ~\u0_R5_reg[17]/NET0131  & n64004 ;
  assign n64007 = ~n64005 & ~n64006 ;
  assign n64016 = decrypt_pad & ~\u0_uk_K_r5_reg[7]/NET0131  ;
  assign n64017 = ~decrypt_pad & ~\u0_uk_K_r5_reg[31]/NET0131  ;
  assign n64018 = ~n64016 & ~n64017 ;
  assign n64019 = \u0_R5_reg[16]/NET0131  & ~n64018 ;
  assign n64020 = ~\u0_R5_reg[16]/NET0131  & n64018 ;
  assign n64021 = ~n64019 & ~n64020 ;
  assign n64036 = ~n64007 & ~n64021 ;
  assign n64059 = ~n64014 & n64036 ;
  assign n64060 = ~n63995 & n64059 ;
  assign n64022 = n64014 & ~n64021 ;
  assign n64062 = ~n63995 & n64007 ;
  assign n64063 = n64022 & n64062 ;
  assign n64027 = n64007 & n64021 ;
  assign n64052 = ~n64014 & n64027 ;
  assign n64024 = ~n64007 & n64021 ;
  assign n64061 = n64014 & n64024 ;
  assign n64064 = ~n64052 & ~n64061 ;
  assign n64065 = ~n64063 & n64064 ;
  assign n64066 = ~n64060 & n64065 ;
  assign n64067 = ~n64001 & ~n64066 ;
  assign n64041 = ~n64001 & n64007 ;
  assign n64042 = ~n64021 & n64041 ;
  assign n64040 = n64001 & n64021 ;
  assign n64043 = n64014 & ~n64040 ;
  assign n64044 = ~n64042 & n64043 ;
  assign n64053 = ~n64044 & ~n64052 ;
  assign n64054 = n63995 & ~n64053 ;
  assign n64028 = n64014 & n64027 ;
  assign n64055 = ~n63995 & n64001 ;
  assign n64056 = n64028 & n64055 ;
  assign n64034 = ~n64014 & n64021 ;
  assign n64057 = n64001 & ~n64007 ;
  assign n64058 = n64034 & n64057 ;
  assign n64068 = ~n64056 & ~n64058 ;
  assign n64069 = ~n64054 & n64068 ;
  assign n64070 = ~n64067 & n64069 ;
  assign n64071 = n63989 & ~n64070 ;
  assign n64029 = ~n64001 & n64028 ;
  assign n64025 = ~n64001 & ~n64014 ;
  assign n64026 = n64024 & n64025 ;
  assign n64008 = n64001 & n64007 ;
  assign n64015 = n64008 & ~n64014 ;
  assign n64023 = ~n64007 & n64022 ;
  assign n64030 = ~n64015 & ~n64023 ;
  assign n64031 = ~n64026 & n64030 ;
  assign n64032 = ~n64029 & n64031 ;
  assign n64033 = ~n63995 & ~n64032 ;
  assign n64035 = ~n64008 & ~n64034 ;
  assign n64037 = ~n64001 & n64014 ;
  assign n64038 = ~n64036 & ~n64037 ;
  assign n64039 = n64035 & n64038 ;
  assign n64045 = ~n64014 & ~n64036 ;
  assign n64046 = ~n64042 & n64045 ;
  assign n64047 = n63995 & ~n64044 ;
  assign n64048 = ~n64046 & n64047 ;
  assign n64049 = ~n64039 & ~n64048 ;
  assign n64050 = ~n64033 & n64049 ;
  assign n64051 = ~n63989 & ~n64050 ;
  assign n64072 = ~n64027 & ~n64057 ;
  assign n64073 = ~n64014 & ~n64040 ;
  assign n64074 = ~n64072 & n64073 ;
  assign n64075 = n63995 & ~n64074 ;
  assign n64076 = n64001 & n64023 ;
  assign n64077 = ~n64015 & ~n64076 ;
  assign n64078 = ~n64021 & ~n64077 ;
  assign n64079 = ~n63995 & ~n64078 ;
  assign n64080 = ~n64075 & ~n64079 ;
  assign n64081 = ~n64051 & ~n64080 ;
  assign n64082 = ~n64071 & n64081 ;
  assign n64083 = ~\u0_L5_reg[14]/NET0131  & ~n64082 ;
  assign n64084 = \u0_L5_reg[14]/NET0131  & n64082 ;
  assign n64085 = ~n64083 & ~n64084 ;
  assign n64086 = ~n63713 & ~n63739 ;
  assign n64087 = ~n63695 & n64086 ;
  assign n64088 = n63702 & ~n64087 ;
  assign n64089 = n63726 & n63732 ;
  assign n64090 = ~n64088 & ~n64089 ;
  assign n64091 = ~n63724 & ~n64090 ;
  assign n64095 = n63706 & n63742 ;
  assign n64092 = n63672 & n63731 ;
  assign n64094 = n63704 & n63712 ;
  assign n64097 = ~n64092 & ~n64094 ;
  assign n64098 = ~n64095 & n64097 ;
  assign n64093 = n63702 & n63727 ;
  assign n64096 = n63686 & n63692 ;
  assign n64099 = ~n64093 & ~n64096 ;
  assign n64100 = n64098 & n64099 ;
  assign n64101 = n63724 & ~n64100 ;
  assign n64103 = n63679 & ~n63724 ;
  assign n64102 = n63694 & n63731 ;
  assign n64105 = ~n64094 & ~n64102 ;
  assign n64106 = ~n64103 & n64105 ;
  assign n64104 = ~n63686 & ~n63702 ;
  assign n64107 = ~n63728 & n64104 ;
  assign n64108 = n64106 & n64107 ;
  assign n64109 = ~n63685 & n63695 ;
  assign n64110 = n63702 & ~n63748 ;
  assign n64111 = ~n64109 & n64110 ;
  assign n64112 = ~n64108 & ~n64111 ;
  assign n64113 = ~n64101 & ~n64112 ;
  assign n64114 = ~n64091 & n64113 ;
  assign n64115 = \u0_L5_reg[15]/P0001  & n64114 ;
  assign n64116 = ~\u0_L5_reg[15]/P0001  & ~n64114 ;
  assign n64117 = ~n64115 & ~n64116 ;
  assign n64118 = ~n64041 & n64073 ;
  assign n64119 = ~n64028 & ~n64036 ;
  assign n64120 = ~n64118 & n64119 ;
  assign n64121 = n63995 & ~n64120 ;
  assign n64122 = ~n64042 & ~n64061 ;
  assign n64123 = ~n63995 & ~n64122 ;
  assign n64124 = ~n64034 & ~n64037 ;
  assign n64125 = n64007 & ~n64025 ;
  assign n64126 = ~n64124 & n64125 ;
  assign n64127 = ~n64123 & ~n64126 ;
  assign n64128 = ~n64121 & n64127 ;
  assign n64129 = n63989 & ~n64128 ;
  assign n64142 = ~n64052 & ~n64059 ;
  assign n64143 = n64001 & ~n64142 ;
  assign n64144 = ~n64001 & n64022 ;
  assign n64145 = ~n64007 & n64144 ;
  assign n64146 = ~n64143 & ~n64145 ;
  assign n64147 = n63995 & ~n64146 ;
  assign n64135 = ~n63995 & ~n64027 ;
  assign n64136 = ~n64035 & n64135 ;
  assign n64133 = n63995 & ~n64014 ;
  assign n64134 = n64041 & n64133 ;
  assign n64130 = n64008 & n64022 ;
  assign n64131 = ~n63995 & ~n64001 ;
  assign n64132 = n64036 & n64131 ;
  assign n64137 = ~n64130 & ~n64132 ;
  assign n64138 = ~n64134 & n64137 ;
  assign n64139 = ~n64136 & n64138 ;
  assign n64140 = ~n63989 & ~n64139 ;
  assign n64141 = n64024 & n64055 ;
  assign n64148 = ~n64029 & ~n64141 ;
  assign n64149 = ~n64140 & n64148 ;
  assign n64150 = ~n64147 & n64149 ;
  assign n64151 = ~n64129 & n64150 ;
  assign n64152 = ~\u0_L5_reg[25]/NET0131  & ~n64151 ;
  assign n64153 = \u0_L5_reg[25]/NET0131  & n64151 ;
  assign n64154 = ~n64152 & ~n64153 ;
  assign n64157 = ~n63706 & n63732 ;
  assign n64158 = ~n63702 & ~n64157 ;
  assign n64159 = ~n64096 & n64158 ;
  assign n64161 = ~n63739 & ~n63749 ;
  assign n64162 = ~n64157 & ~n64161 ;
  assign n64160 = n63678 & n63694 ;
  assign n64163 = n63702 & ~n64160 ;
  assign n64164 = ~n64162 & n64163 ;
  assign n64165 = ~n64159 & ~n64164 ;
  assign n64155 = ~n63727 & ~n63740 ;
  assign n64156 = n63685 & ~n64155 ;
  assign n64166 = n63724 & ~n64109 ;
  assign n64167 = ~n64156 & n64166 ;
  assign n64168 = ~n64165 & n64167 ;
  assign n64169 = ~n63740 & ~n63750 ;
  assign n64170 = ~n63686 & n64169 ;
  assign n64171 = n63702 & ~n64170 ;
  assign n64175 = n63678 & n63704 ;
  assign n64179 = ~n63724 & ~n64175 ;
  assign n64180 = ~n63693 & n64179 ;
  assign n64176 = n63672 & n63692 ;
  assign n64177 = ~n63709 & ~n63731 ;
  assign n64178 = n64176 & ~n64177 ;
  assign n64172 = ~n63672 & ~n63702 ;
  assign n64173 = ~n63710 & ~n63712 ;
  assign n64174 = n64172 & ~n64173 ;
  assign n64181 = ~n63728 & ~n64174 ;
  assign n64182 = ~n64178 & n64181 ;
  assign n64183 = n64180 & n64182 ;
  assign n64184 = ~n64171 & n64183 ;
  assign n64185 = ~n64168 & ~n64184 ;
  assign n64186 = ~\u0_L5_reg[21]/NET0131  & n64185 ;
  assign n64187 = \u0_L5_reg[21]/NET0131  & ~n64185 ;
  assign n64188 = ~n64186 & ~n64187 ;
  assign n64204 = ~n63606 & n63634 ;
  assign n64205 = n63658 & ~n64204 ;
  assign n64207 = n63598 & n63606 ;
  assign n64206 = ~n63583 & n63621 ;
  assign n64208 = ~n63577 & ~n64206 ;
  assign n64209 = ~n64207 & n64208 ;
  assign n64210 = ~n64205 & ~n64209 ;
  assign n64211 = n63621 & n63623 ;
  assign n64212 = ~n63624 & ~n64211 ;
  assign n64213 = ~n63628 & n64212 ;
  assign n64214 = ~n64210 & n64213 ;
  assign n64215 = ~n63615 & ~n64214 ;
  assign n64196 = ~n63621 & n63623 ;
  assign n64197 = n63590 & n63607 ;
  assign n64198 = ~n64196 & ~n64197 ;
  assign n64199 = ~n63577 & ~n64198 ;
  assign n64194 = n63590 & n63639 ;
  assign n64200 = ~n63596 & n63656 ;
  assign n64201 = ~n64194 & ~n64200 ;
  assign n64202 = ~n64199 & n64201 ;
  assign n64203 = n63615 & ~n64202 ;
  assign n64189 = ~n63648 & n63933 ;
  assign n64190 = n63577 & ~n64189 ;
  assign n64195 = ~n63577 & n64194 ;
  assign n64191 = ~n63638 & ~n63643 ;
  assign n64192 = n63577 & n63615 ;
  assign n64193 = ~n64191 & n64192 ;
  assign n64216 = ~n63619 & ~n64193 ;
  assign n64217 = ~n64195 & n64216 ;
  assign n64218 = ~n64190 & n64217 ;
  assign n64219 = ~n64203 & n64218 ;
  assign n64220 = ~n64215 & n64219 ;
  assign n64221 = ~\u0_L5_reg[1]/NET0131  & ~n64220 ;
  assign n64222 = \u0_L5_reg[1]/NET0131  & n64220 ;
  assign n64223 = ~n64221 & ~n64222 ;
  assign n64246 = n63863 & n63894 ;
  assign n64247 = n63870 & n64246 ;
  assign n64248 = ~n63899 & ~n63901 ;
  assign n64249 = ~n64247 & n64248 ;
  assign n64250 = n63844 & ~n64249 ;
  assign n64228 = n63863 & n63873 ;
  assign n64229 = ~n63870 & n63894 ;
  assign n64230 = ~n64228 & ~n64229 ;
  assign n64245 = ~n63844 & ~n64230 ;
  assign n64242 = n63844 & n63850 ;
  assign n64243 = ~n63864 & ~n64242 ;
  assign n64244 = ~n63870 & ~n64243 ;
  assign n64251 = n63873 & n63916 ;
  assign n64252 = ~n64244 & ~n64251 ;
  assign n64253 = ~n64245 & n64252 ;
  assign n64254 = ~n64250 & n64253 ;
  assign n64255 = n63838 & ~n64254 ;
  assign n64224 = n63876 & n63887 ;
  assign n64225 = ~n63863 & n63896 ;
  assign n64226 = ~n64224 & ~n64225 ;
  assign n64227 = ~n63844 & ~n64226 ;
  assign n64231 = n63844 & n64230 ;
  assign n64232 = ~n63870 & n63876 ;
  assign n64233 = ~n63844 & ~n63875 ;
  assign n64234 = ~n63874 & n64233 ;
  assign n64235 = ~n64232 & n64234 ;
  assign n64236 = ~n64231 & ~n64235 ;
  assign n64237 = ~n63873 & ~n63876 ;
  assign n64238 = n63916 & n64237 ;
  assign n64239 = ~n64224 & ~n64238 ;
  assign n64240 = ~n64236 & n64239 ;
  assign n64241 = ~n63838 & ~n64240 ;
  assign n64256 = ~n64227 & ~n64241 ;
  assign n64257 = ~n64255 & n64256 ;
  assign n64258 = ~\u0_L5_reg[28]/NET0131  & ~n64257 ;
  assign n64259 = \u0_L5_reg[28]/NET0131  & n64257 ;
  assign n64260 = ~n64258 & ~n64259 ;
  assign n64279 = ~n63484 & n63805 ;
  assign n64280 = ~n63517 & ~n64279 ;
  assign n64281 = ~n63532 & n64280 ;
  assign n64282 = n63508 & ~n64281 ;
  assign n64277 = ~n63500 & ~n63823 ;
  assign n64278 = ~n63508 & ~n64277 ;
  assign n64283 = ~n63548 & ~n63553 ;
  assign n64284 = ~n64278 & n64283 ;
  assign n64285 = ~n64282 & n64284 ;
  assign n64286 = ~n63526 & ~n64285 ;
  assign n64270 = n63491 & ~n63818 ;
  assign n64271 = ~n63478 & n63538 ;
  assign n64272 = ~n64270 & ~n64271 ;
  assign n64273 = ~n63508 & ~n64272 ;
  assign n64262 = ~n63478 & n63528 ;
  assign n64263 = ~n63538 & ~n64262 ;
  assign n64264 = ~n63508 & ~n64263 ;
  assign n64261 = n63485 & n63813 ;
  assign n64265 = n63491 & n63555 ;
  assign n64266 = ~n64261 & ~n64265 ;
  assign n64267 = ~n63501 & n64266 ;
  assign n64268 = ~n64264 & n64267 ;
  assign n64269 = n63526 & ~n64268 ;
  assign n64274 = ~n63512 & ~n63556 ;
  assign n64275 = ~n63517 & n64274 ;
  assign n64276 = n63534 & ~n64275 ;
  assign n64287 = ~n64269 & ~n64276 ;
  assign n64288 = ~n64273 & n64287 ;
  assign n64289 = ~n64286 & n64288 ;
  assign n64290 = ~\u0_L5_reg[4]/NET0131  & ~n64289 ;
  assign n64291 = \u0_L5_reg[4]/NET0131  & n64289 ;
  assign n64292 = ~n64290 & ~n64291 ;
  assign n64297 = ~n63902 & ~n64224 ;
  assign n64298 = ~n64246 & ~n64251 ;
  assign n64299 = ~n63900 & n64298 ;
  assign n64300 = n64297 & n64299 ;
  assign n64301 = ~n63844 & ~n64300 ;
  assign n64302 = n63863 & ~n64232 ;
  assign n64303 = n63844 & ~n63874 ;
  assign n64304 = ~n63899 & n64303 ;
  assign n64305 = ~n64302 & n64304 ;
  assign n64295 = n63870 & ~n63881 ;
  assign n64296 = n64242 & n64295 ;
  assign n64293 = ~n63850 & ~n63884 ;
  assign n64294 = n63885 & n64293 ;
  assign n64306 = ~n63838 & ~n64294 ;
  assign n64307 = ~n64296 & n64306 ;
  assign n64308 = ~n64305 & n64307 ;
  assign n64309 = ~n64301 & n64308 ;
  assign n64312 = ~n63856 & n63911 ;
  assign n64311 = n63856 & n63896 ;
  assign n64313 = n63844 & ~n64311 ;
  assign n64314 = ~n64312 & n64313 ;
  assign n64315 = ~n63844 & ~n63864 ;
  assign n64316 = ~n63917 & n64315 ;
  assign n64317 = ~n64314 & ~n64316 ;
  assign n64310 = n63863 & n64229 ;
  assign n64318 = n63838 & n63889 ;
  assign n64319 = ~n64310 & n64318 ;
  assign n64320 = n64297 & n64319 ;
  assign n64321 = ~n64317 & n64320 ;
  assign n64322 = ~n64309 & ~n64321 ;
  assign n64323 = ~\u0_L5_reg[13]/NET0131  & ~n64322 ;
  assign n64324 = \u0_L5_reg[13]/NET0131  & n64322 ;
  assign n64325 = ~n64323 & ~n64324 ;
  assign n64329 = ~n64160 & n64169 ;
  assign n64330 = ~n63702 & ~n64329 ;
  assign n64327 = n63702 & ~n63730 ;
  assign n64328 = ~n64086 & n64327 ;
  assign n64326 = ~n63685 & n63706 ;
  assign n64331 = ~n63693 & ~n64326 ;
  assign n64332 = ~n63748 & n64331 ;
  assign n64333 = ~n64328 & n64332 ;
  assign n64334 = ~n64330 & n64333 ;
  assign n64335 = n63724 & ~n64334 ;
  assign n64339 = n63702 & ~n63713 ;
  assign n64338 = n63692 & ~n63731 ;
  assign n64340 = ~n64175 & ~n64338 ;
  assign n64341 = n64339 & n64340 ;
  assign n64337 = n63742 & n64176 ;
  assign n64336 = n63712 & n64172 ;
  assign n64342 = ~n63729 & ~n64336 ;
  assign n64343 = ~n64337 & n64342 ;
  assign n64344 = ~n64341 & n64343 ;
  assign n64345 = ~n63724 & ~n64344 ;
  assign n64348 = ~n63702 & n63735 ;
  assign n64346 = n63685 & n63702 ;
  assign n64347 = n63726 & n64346 ;
  assign n64349 = ~n63741 & ~n64347 ;
  assign n64350 = ~n64348 & n64349 ;
  assign n64351 = ~n64345 & n64350 ;
  assign n64352 = ~n64335 & n64351 ;
  assign n64353 = ~\u0_L5_reg[27]/NET0131  & ~n64352 ;
  assign n64354 = \u0_L5_reg[27]/NET0131  & n64352 ;
  assign n64355 = ~n64353 & ~n64354 ;
  assign n64375 = ~n63427 & ~n63435 ;
  assign n64376 = ~n63410 & ~n64375 ;
  assign n64377 = ~n63426 & ~n64376 ;
  assign n64378 = ~n63391 & ~n64377 ;
  assign n64379 = n63391 & ~n63775 ;
  assign n64380 = n63422 & n64379 ;
  assign n64381 = ~n63413 & ~n63780 ;
  assign n64382 = ~n64380 & n64381 ;
  assign n64383 = ~n64378 & n64382 ;
  assign n64384 = n63419 & ~n64383 ;
  assign n64357 = n63404 & ~n63410 ;
  assign n64358 = n63398 & n64357 ;
  assign n64362 = ~n63451 & ~n63779 ;
  assign n64363 = ~n64358 & n64362 ;
  assign n64356 = n63391 & n63435 ;
  assign n64359 = ~n63385 & ~n63778 ;
  assign n64360 = ~n63391 & n63410 ;
  assign n64361 = ~n64359 & n64360 ;
  assign n64364 = ~n64356 & ~n64361 ;
  assign n64365 = n64363 & n64364 ;
  assign n64366 = ~n63419 & ~n64365 ;
  assign n64369 = n63427 & n63428 ;
  assign n64370 = ~n63783 & ~n64369 ;
  assign n64371 = ~n63391 & ~n64370 ;
  assign n64367 = ~n63424 & ~n63435 ;
  assign n64368 = n63391 & ~n64367 ;
  assign n64372 = ~n63460 & ~n64368 ;
  assign n64373 = ~n64371 & n64372 ;
  assign n64374 = ~n63398 & ~n64373 ;
  assign n64385 = ~n64366 & ~n64374 ;
  assign n64386 = ~n64384 & n64385 ;
  assign n64387 = \u0_L5_reg[23]/NET0131  & ~n64386 ;
  assign n64388 = ~\u0_L5_reg[23]/NET0131  & n64386 ;
  assign n64389 = ~n64387 & ~n64388 ;
  assign n64390 = n63300 & n63356 ;
  assign n64392 = n63326 & ~n63962 ;
  assign n64391 = n63316 & n63325 ;
  assign n64393 = ~n63324 & ~n63350 ;
  assign n64394 = ~n64391 & n64393 ;
  assign n64395 = ~n64392 & n64394 ;
  assign n64396 = n63300 & n63307 ;
  assign n64397 = ~n63959 & ~n64396 ;
  assign n64398 = ~n63313 & n63349 ;
  assign n64399 = n63324 & ~n64398 ;
  assign n64400 = ~n64397 & n64399 ;
  assign n64401 = ~n64395 & ~n64400 ;
  assign n64402 = ~n64390 & ~n64401 ;
  assign n64403 = n63288 & ~n64402 ;
  assign n64406 = ~n63328 & ~n63357 ;
  assign n64407 = ~n64398 & n64406 ;
  assign n64408 = ~n63324 & ~n64407 ;
  assign n64411 = ~n63335 & ~n63962 ;
  assign n64409 = n63294 & ~n63328 ;
  assign n64410 = ~n63300 & ~n64409 ;
  assign n64412 = ~n63313 & ~n63332 ;
  assign n64413 = ~n64410 & ~n64412 ;
  assign n64414 = ~n64411 & n64413 ;
  assign n64415 = ~n64408 & ~n64414 ;
  assign n64416 = ~n63288 & ~n64415 ;
  assign n64404 = n63288 & ~n63324 ;
  assign n64405 = n63318 & ~n64404 ;
  assign n64417 = n63346 & ~n63366 ;
  assign n64418 = n63345 & n64417 ;
  assign n64419 = ~n64405 & ~n64418 ;
  assign n64420 = ~n64416 & n64419 ;
  assign n64421 = ~n64403 & n64420 ;
  assign n64422 = \u0_L5_reg[32]/NET0131  & n64421 ;
  assign n64423 = ~\u0_L5_reg[32]/NET0131  & ~n64421 ;
  assign n64424 = ~n64422 & ~n64423 ;
  assign n64428 = ~n63333 & ~n63962 ;
  assign n64425 = n63300 & ~n63317 ;
  assign n64426 = ~n64409 & n64425 ;
  assign n64427 = ~n63288 & n63324 ;
  assign n64429 = ~n64426 & n64427 ;
  assign n64430 = ~n64428 & n64429 ;
  assign n64431 = n63333 & n63962 ;
  assign n64432 = ~n63314 & ~n64428 ;
  assign n64433 = ~n64431 & n64432 ;
  assign n64434 = ~n64404 & ~n64427 ;
  assign n64435 = ~n64433 & n64434 ;
  assign n64436 = ~n64430 & ~n64435 ;
  assign n64437 = ~n63358 & ~n64436 ;
  assign n64440 = n63313 & ~n63962 ;
  assign n64439 = ~n63294 & ~n63334 ;
  assign n64438 = ~n63328 & n63344 ;
  assign n64441 = n64404 & ~n64438 ;
  assign n64442 = ~n64439 & n64441 ;
  assign n64443 = ~n64440 & n64442 ;
  assign n64444 = ~n64437 & ~n64443 ;
  assign n64445 = ~\u0_L5_reg[7]/NET0131  & n64444 ;
  assign n64446 = \u0_L5_reg[7]/NET0131  & ~n64444 ;
  assign n64447 = ~n64445 & ~n64446 ;
  assign n64461 = n64025 & n64036 ;
  assign n64462 = ~n64061 & ~n64461 ;
  assign n64463 = n63995 & ~n64462 ;
  assign n64464 = n64021 & n64131 ;
  assign n64465 = ~n64463 & ~n64464 ;
  assign n64466 = ~n64078 & n64465 ;
  assign n64467 = n63989 & ~n64466 ;
  assign n64452 = n63995 & ~n64026 ;
  assign n64453 = ~n64028 & n64452 ;
  assign n64454 = n64022 & ~n64057 ;
  assign n64455 = ~n63995 & ~n64061 ;
  assign n64456 = ~n64454 & n64455 ;
  assign n64457 = ~n64453 & ~n64456 ;
  assign n64458 = ~n64042 & ~n64143 ;
  assign n64459 = ~n64457 & n64458 ;
  assign n64460 = ~n63989 & ~n64459 ;
  assign n64448 = ~n64014 & n64141 ;
  assign n64449 = n64007 & n64144 ;
  assign n64450 = n64077 & ~n64449 ;
  assign n64451 = n63995 & ~n64450 ;
  assign n64468 = ~n64448 & ~n64451 ;
  assign n64469 = ~n64460 & n64468 ;
  assign n64470 = ~n64467 & n64469 ;
  assign n64471 = ~\u0_L5_reg[8]/NET0131  & ~n64470 ;
  assign n64472 = \u0_L5_reg[8]/NET0131  & n64470 ;
  assign n64473 = ~n64471 & ~n64472 ;
  assign n64476 = ~n63514 & ~n63529 ;
  assign n64477 = n63508 & ~n64476 ;
  assign n64475 = ~n63508 & n63533 ;
  assign n64478 = n63526 & ~n64262 ;
  assign n64479 = ~n64475 & n64478 ;
  assign n64474 = n63491 & n63556 ;
  assign n64480 = ~n63807 & ~n64474 ;
  assign n64481 = n64479 & n64480 ;
  assign n64482 = ~n64477 & n64481 ;
  assign n64485 = n63484 & ~n63528 ;
  assign n64486 = ~n63500 & ~n64485 ;
  assign n64487 = n63508 & ~n64486 ;
  assign n64484 = ~n63508 & ~n64274 ;
  assign n64483 = n63491 & n63549 ;
  assign n64488 = ~n63526 & ~n64483 ;
  assign n64489 = ~n64484 & n64488 ;
  assign n64490 = ~n64487 & n64489 ;
  assign n64491 = ~n64482 & ~n64490 ;
  assign n64492 = ~n63520 & ~n63554 ;
  assign n64493 = ~n64491 & n64492 ;
  assign n64494 = ~\u0_L5_reg[19]/P0001  & ~n64493 ;
  assign n64495 = \u0_L5_reg[19]/P0001  & n64493 ;
  assign n64496 = ~n64494 & ~n64495 ;
  assign n64533 = decrypt_pad & ~\u0_uk_K_r5_reg[32]/NET0131  ;
  assign n64534 = ~decrypt_pad & ~\u0_uk_K_r5_reg[54]/NET0131  ;
  assign n64535 = ~n64533 & ~n64534 ;
  assign n64536 = \u0_R5_reg[11]/P0001  & ~n64535 ;
  assign n64537 = ~\u0_R5_reg[11]/P0001  & n64535 ;
  assign n64538 = ~n64536 & ~n64537 ;
  assign n64503 = decrypt_pad & ~\u0_uk_K_r5_reg[55]/NET0131  ;
  assign n64504 = ~decrypt_pad & ~\u0_uk_K_r5_reg[20]/NET0131  ;
  assign n64505 = ~n64503 & ~n64504 ;
  assign n64506 = \u0_R5_reg[9]/NET0131  & ~n64505 ;
  assign n64507 = ~\u0_R5_reg[9]/NET0131  & n64505 ;
  assign n64508 = ~n64506 & ~n64507 ;
  assign n64509 = decrypt_pad & ~\u0_uk_K_r5_reg[3]/NET0131  ;
  assign n64510 = ~decrypt_pad & ~\u0_uk_K_r5_reg[25]/NET0131  ;
  assign n64511 = ~n64509 & ~n64510 ;
  assign n64512 = \u0_R5_reg[13]/NET0131  & ~n64511 ;
  assign n64513 = ~\u0_R5_reg[13]/NET0131  & n64511 ;
  assign n64514 = ~n64512 & ~n64513 ;
  assign n64515 = n64508 & ~n64514 ;
  assign n64516 = decrypt_pad & ~\u0_uk_K_r5_reg[6]/NET0131  ;
  assign n64517 = ~decrypt_pad & ~\u0_uk_K_r5_reg[53]/NET0131  ;
  assign n64518 = ~n64516 & ~n64517 ;
  assign n64519 = \u0_R5_reg[10]/NET0131  & ~n64518 ;
  assign n64520 = ~\u0_R5_reg[10]/NET0131  & n64518 ;
  assign n64521 = ~n64519 & ~n64520 ;
  assign n64522 = decrypt_pad & ~\u0_uk_K_r5_reg[26]/NET0131  ;
  assign n64523 = ~decrypt_pad & ~\u0_uk_K_r5_reg[48]/NET0131  ;
  assign n64524 = ~n64522 & ~n64523 ;
  assign n64525 = \u0_R5_reg[8]/NET0131  & ~n64524 ;
  assign n64526 = ~\u0_R5_reg[8]/NET0131  & n64524 ;
  assign n64527 = ~n64525 & ~n64526 ;
  assign n64528 = n64521 & ~n64527 ;
  assign n64529 = ~n64508 & n64514 ;
  assign n64530 = ~n64528 & ~n64529 ;
  assign n64531 = ~n64515 & n64530 ;
  assign n64497 = decrypt_pad & ~\u0_uk_K_r5_reg[47]/NET0131  ;
  assign n64498 = ~decrypt_pad & ~\u0_uk_K_r5_reg[12]/NET0131  ;
  assign n64499 = ~n64497 & ~n64498 ;
  assign n64500 = \u0_R5_reg[12]/NET0131  & ~n64499 ;
  assign n64501 = ~\u0_R5_reg[12]/NET0131  & n64499 ;
  assign n64502 = ~n64500 & ~n64501 ;
  assign n64562 = ~n64514 & ~n64527 ;
  assign n64563 = n64502 & ~n64562 ;
  assign n64564 = ~n64531 & n64563 ;
  assign n64532 = ~n64508 & ~n64527 ;
  assign n64559 = ~n64514 & n64532 ;
  assign n64560 = ~n64521 & n64559 ;
  assign n64561 = n64521 & n64529 ;
  assign n64565 = ~n64560 & ~n64561 ;
  assign n64566 = ~n64564 & n64565 ;
  assign n64567 = n64538 & ~n64566 ;
  assign n64539 = ~n64532 & ~n64538 ;
  assign n64540 = n64531 & n64539 ;
  assign n64541 = n64508 & n64521 ;
  assign n64542 = ~n64514 & n64541 ;
  assign n64543 = ~n64527 & n64542 ;
  assign n64544 = ~n64540 & ~n64543 ;
  assign n64545 = n64502 & ~n64544 ;
  assign n64548 = n64514 & n64538 ;
  assign n64554 = n64508 & n64548 ;
  assign n64546 = ~n64508 & ~n64521 ;
  assign n64547 = ~n64541 & ~n64546 ;
  assign n64549 = n64514 & ~n64527 ;
  assign n64550 = ~n64514 & n64527 ;
  assign n64551 = ~n64549 & ~n64550 ;
  assign n64555 = n64547 & ~n64551 ;
  assign n64556 = ~n64554 & n64555 ;
  assign n64552 = ~n64548 & ~n64551 ;
  assign n64553 = ~n64547 & ~n64552 ;
  assign n64557 = ~n64502 & ~n64553 ;
  assign n64558 = ~n64556 & n64557 ;
  assign n64568 = ~n64545 & ~n64558 ;
  assign n64569 = ~n64567 & n64568 ;
  assign n64570 = ~\u0_L5_reg[6]/NET0131  & ~n64569 ;
  assign n64571 = \u0_L5_reg[6]/NET0131  & n64569 ;
  assign n64572 = ~n64570 & ~n64571 ;
  assign n64575 = n64538 & ~n64549 ;
  assign n64576 = ~n64552 & ~n64575 ;
  assign n64577 = n64546 & ~n64576 ;
  assign n64573 = ~n64538 & ~n64546 ;
  assign n64574 = n64551 & n64573 ;
  assign n64578 = n64502 & ~n64574 ;
  assign n64579 = ~n64577 & n64578 ;
  assign n64583 = ~n64521 & n64549 ;
  assign n64584 = n64521 & n64562 ;
  assign n64585 = ~n64583 & ~n64584 ;
  assign n64580 = n64521 & n64527 ;
  assign n64581 = ~n64508 & n64580 ;
  assign n64586 = n64508 & n64562 ;
  assign n64587 = ~n64581 & ~n64586 ;
  assign n64588 = n64585 & n64587 ;
  assign n64589 = n64538 & ~n64588 ;
  assign n64582 = ~n64514 & n64581 ;
  assign n64590 = ~n64502 & ~n64582 ;
  assign n64591 = ~n64589 & n64590 ;
  assign n64592 = ~n64579 & ~n64591 ;
  assign n64597 = ~n64532 & ~n64551 ;
  assign n64598 = ~n64515 & ~n64521 ;
  assign n64599 = n64597 & n64598 ;
  assign n64593 = n64521 & n64549 ;
  assign n64594 = n64508 & n64580 ;
  assign n64595 = ~n64593 & ~n64594 ;
  assign n64596 = n64502 & ~n64595 ;
  assign n64600 = n64538 & ~n64596 ;
  assign n64601 = ~n64599 & n64600 ;
  assign n64603 = n64546 & n64551 ;
  assign n64602 = n64508 & n64550 ;
  assign n64604 = ~n64593 & ~n64602 ;
  assign n64605 = ~n64603 & n64604 ;
  assign n64606 = ~n64502 & ~n64605 ;
  assign n64607 = n64514 & n64527 ;
  assign n64608 = n64508 & n64607 ;
  assign n64609 = n64521 & n64608 ;
  assign n64610 = ~n64538 & ~n64609 ;
  assign n64611 = ~n64606 & n64610 ;
  assign n64612 = ~n64601 & ~n64611 ;
  assign n64613 = ~n64592 & ~n64612 ;
  assign n64614 = ~\u0_L5_reg[24]/NET0131  & ~n64613 ;
  assign n64615 = \u0_L5_reg[24]/NET0131  & n64613 ;
  assign n64616 = ~n64614 & ~n64615 ;
  assign n64618 = ~n64508 & ~n64607 ;
  assign n64619 = ~n64608 & ~n64618 ;
  assign n64620 = ~n64562 & ~n64619 ;
  assign n64621 = n64538 & n64586 ;
  assign n64622 = ~n64620 & ~n64621 ;
  assign n64623 = ~n64521 & ~n64622 ;
  assign n64617 = n64541 & n64549 ;
  assign n64624 = ~n64538 & ~n64580 ;
  assign n64625 = ~n64521 & ~n64527 ;
  assign n64626 = ~n64514 & ~n64625 ;
  assign n64627 = n64624 & n64626 ;
  assign n64628 = ~n64617 & ~n64627 ;
  assign n64629 = ~n64623 & n64628 ;
  assign n64630 = n64502 & ~n64629 ;
  assign n64631 = ~n64530 & ~n64549 ;
  assign n64632 = ~n64502 & ~n64597 ;
  assign n64633 = ~n64631 & n64632 ;
  assign n64634 = ~n64581 & ~n64633 ;
  assign n64635 = ~n64538 & ~n64634 ;
  assign n64636 = n64538 & ~n64562 ;
  assign n64637 = n64619 & n64636 ;
  assign n64638 = ~n64560 & ~n64637 ;
  assign n64639 = ~n64502 & ~n64638 ;
  assign n64640 = ~n64559 & ~n64602 ;
  assign n64641 = n64521 & n64538 ;
  assign n64642 = ~n64640 & n64641 ;
  assign n64643 = ~n64639 & ~n64642 ;
  assign n64644 = ~n64635 & n64643 ;
  assign n64645 = ~n64630 & n64644 ;
  assign n64646 = ~\u0_L5_reg[16]/NET0131  & ~n64645 ;
  assign n64647 = \u0_L5_reg[16]/NET0131  & n64645 ;
  assign n64648 = ~n64646 & ~n64647 ;
  assign n64649 = ~n64076 & n64452 ;
  assign n64650 = ~n64001 & ~n64142 ;
  assign n64651 = ~n64131 & ~n64455 ;
  assign n64652 = ~n64650 & ~n64651 ;
  assign n64653 = ~n64649 & ~n64652 ;
  assign n64656 = ~n64052 & ~n64144 ;
  assign n64657 = n63995 & ~n64656 ;
  assign n64654 = ~n64061 & ~n64124 ;
  assign n64655 = ~n63995 & ~n64654 ;
  assign n64658 = ~n64034 & n64057 ;
  assign n64659 = ~n63989 & ~n64658 ;
  assign n64660 = ~n64655 & n64659 ;
  assign n64661 = ~n64657 & n64660 ;
  assign n64662 = ~n64001 & n64021 ;
  assign n64663 = ~n64045 & ~n64662 ;
  assign n64664 = n63995 & ~n64034 ;
  assign n64665 = ~n64663 & n64664 ;
  assign n64666 = n63989 & ~n64058 ;
  assign n64667 = ~n64063 & n64666 ;
  assign n64668 = ~n64029 & n64667 ;
  assign n64669 = ~n64665 & n64668 ;
  assign n64670 = ~n64661 & ~n64669 ;
  assign n64671 = ~n64653 & ~n64670 ;
  assign n64672 = ~\u0_L5_reg[3]/NET0131  & ~n64671 ;
  assign n64673 = \u0_L5_reg[3]/NET0131  & n64671 ;
  assign n64674 = ~n64672 & ~n64673 ;
  assign n64687 = ~n64515 & ~n64580 ;
  assign n64689 = n64538 & ~n64542 ;
  assign n64690 = ~n64687 & n64689 ;
  assign n64688 = n64539 & n64687 ;
  assign n64686 = n64528 & n64529 ;
  assign n64691 = ~n64603 & ~n64686 ;
  assign n64692 = ~n64688 & n64691 ;
  assign n64693 = ~n64690 & n64692 ;
  assign n64694 = ~n64502 & ~n64693 ;
  assign n64675 = n64548 & n64581 ;
  assign n64676 = ~n64538 & n64542 ;
  assign n64677 = ~n64502 & ~n64676 ;
  assign n64678 = n64541 & ~n64607 ;
  assign n64679 = ~n64586 & n64624 ;
  assign n64680 = n64546 & n64550 ;
  assign n64681 = n64538 & ~n64680 ;
  assign n64682 = n64585 & n64681 ;
  assign n64683 = ~n64679 & ~n64682 ;
  assign n64684 = ~n64678 & ~n64683 ;
  assign n64685 = ~n64677 & ~n64684 ;
  assign n64695 = ~n64675 & ~n64685 ;
  assign n64696 = ~n64694 & n64695 ;
  assign n64697 = \u0_L5_reg[30]/NET0131  & ~n64696 ;
  assign n64698 = ~\u0_L5_reg[30]/NET0131  & n64696 ;
  assign n64699 = ~n64697 & ~n64698 ;
  assign n64704 = n63404 & ~n63445 ;
  assign n64705 = ~n63434 & ~n64704 ;
  assign n64712 = ~n63391 & ~n64705 ;
  assign n64713 = n63391 & ~n63769 ;
  assign n64714 = n64375 & n64713 ;
  assign n64715 = ~n64712 & ~n64714 ;
  assign n64700 = ~n63397 & n63459 ;
  assign n64716 = n63397 & n63764 ;
  assign n64717 = ~n64700 & ~n64716 ;
  assign n64718 = ~n64715 & n64717 ;
  assign n64719 = ~n63419 & ~n64718 ;
  assign n64701 = ~n63410 & n63779 ;
  assign n64702 = ~n64700 & ~n64701 ;
  assign n64703 = ~n63391 & ~n64702 ;
  assign n64707 = n63397 & ~n63422 ;
  assign n64708 = ~n63764 & n64707 ;
  assign n64706 = n63448 & n64705 ;
  assign n64709 = ~n63783 & ~n64706 ;
  assign n64710 = ~n64708 & n64709 ;
  assign n64711 = n63419 & ~n64710 ;
  assign n64720 = ~n64703 & ~n64711 ;
  assign n64721 = ~n64719 & n64720 ;
  assign n64722 = ~\u0_L5_reg[9]/NET0131  & ~n64721 ;
  assign n64723 = \u0_L5_reg[9]/NET0131  & n64721 ;
  assign n64724 = ~n64722 & ~n64723 ;
  assign n64729 = n63844 & ~n63882 ;
  assign n64726 = n63850 & n63885 ;
  assign n64727 = ~n63899 & ~n64726 ;
  assign n64728 = ~n63844 & ~n64727 ;
  assign n64730 = ~n63918 & ~n64728 ;
  assign n64731 = ~n64729 & n64730 ;
  assign n64732 = n63838 & ~n64731 ;
  assign n64733 = n63857 & n63897 ;
  assign n64736 = ~n64224 & ~n64312 ;
  assign n64737 = ~n64733 & n64736 ;
  assign n64734 = ~n63850 & ~n63897 ;
  assign n64735 = ~n63912 & n64734 ;
  assign n64738 = ~n63871 & ~n64735 ;
  assign n64739 = n64737 & n64738 ;
  assign n64740 = ~n63838 & ~n64739 ;
  assign n64725 = ~n63844 & n64228 ;
  assign n64741 = n63857 & n63870 ;
  assign n64742 = ~n64310 & ~n64741 ;
  assign n64743 = n63844 & ~n64742 ;
  assign n64744 = ~n64725 & ~n64743 ;
  assign n64745 = ~n64740 & n64744 ;
  assign n64746 = ~n64732 & n64745 ;
  assign n64747 = \u0_L5_reg[18]/NET0131  & n64746 ;
  assign n64748 = ~\u0_L5_reg[18]/NET0131  & ~n64746 ;
  assign n64749 = ~n64747 & ~n64748 ;
  assign n64801 = decrypt_pad & ~\u0_uk_K_r4_reg[25]/NET0131  ;
  assign n64802 = ~decrypt_pad & ~\u0_uk_K_r4_reg[19]/NET0131  ;
  assign n64803 = ~n64801 & ~n64802 ;
  assign n64804 = \u0_R4_reg[4]/NET0131  & ~n64803 ;
  assign n64805 = ~\u0_R4_reg[4]/NET0131  & n64803 ;
  assign n64806 = ~n64804 & ~n64805 ;
  assign n64756 = decrypt_pad & ~\u0_uk_K_r4_reg[13]/NET0131  ;
  assign n64757 = ~decrypt_pad & ~\u0_uk_K_r4_reg[32]/NET0131  ;
  assign n64758 = ~n64756 & ~n64757 ;
  assign n64759 = \u0_R4_reg[2]/NET0131  & ~n64758 ;
  assign n64760 = ~\u0_R4_reg[2]/NET0131  & n64758 ;
  assign n64761 = ~n64759 & ~n64760 ;
  assign n64750 = decrypt_pad & ~\u0_uk_K_r4_reg[47]/NET0131  ;
  assign n64751 = ~decrypt_pad & ~\u0_uk_K_r4_reg[41]/NET0131  ;
  assign n64752 = ~n64750 & ~n64751 ;
  assign n64753 = \u0_R4_reg[3]/NET0131  & ~n64752 ;
  assign n64754 = ~\u0_R4_reg[3]/NET0131  & n64752 ;
  assign n64755 = ~n64753 & ~n64754 ;
  assign n64769 = decrypt_pad & ~\u0_uk_K_r4_reg[55]/NET0131  ;
  assign n64770 = ~decrypt_pad & ~\u0_uk_K_r4_reg[17]/NET0131  ;
  assign n64771 = ~n64769 & ~n64770 ;
  assign n64772 = \u0_R4_reg[1]/NET0131  & ~n64771 ;
  assign n64773 = ~\u0_R4_reg[1]/NET0131  & n64771 ;
  assign n64774 = ~n64772 & ~n64773 ;
  assign n64777 = ~n64755 & n64774 ;
  assign n64763 = decrypt_pad & ~\u0_uk_K_r4_reg[34]/NET0131  ;
  assign n64764 = ~decrypt_pad & ~\u0_uk_K_r4_reg[53]/NET0131  ;
  assign n64765 = ~n64763 & ~n64764 ;
  assign n64766 = \u0_R4_reg[32]/NET0131  & ~n64765 ;
  assign n64767 = ~\u0_R4_reg[32]/NET0131  & n64765 ;
  assign n64768 = ~n64766 & ~n64767 ;
  assign n64778 = decrypt_pad & ~\u0_uk_K_r4_reg[53]/NET0131  ;
  assign n64779 = ~decrypt_pad & ~\u0_uk_K_r4_reg[47]/NET0131  ;
  assign n64780 = ~n64778 & ~n64779 ;
  assign n64781 = \u0_R4_reg[5]/NET0131  & ~n64780 ;
  assign n64782 = ~\u0_R4_reg[5]/NET0131  & n64780 ;
  assign n64783 = ~n64781 & ~n64782 ;
  assign n64818 = n64768 & n64783 ;
  assign n64819 = ~n64777 & n64818 ;
  assign n64820 = n64774 & ~n64783 ;
  assign n64821 = ~n64768 & n64820 ;
  assign n64822 = ~n64819 & ~n64821 ;
  assign n64823 = ~n64761 & ~n64822 ;
  assign n64808 = n64755 & n64761 ;
  assign n64789 = n64768 & ~n64783 ;
  assign n64793 = ~n64768 & n64783 ;
  assign n64809 = ~n64789 & ~n64793 ;
  assign n64810 = n64774 & ~n64809 ;
  assign n64811 = n64808 & n64810 ;
  assign n64812 = ~n64774 & n64783 ;
  assign n64813 = ~n64761 & ~n64768 ;
  assign n64814 = ~n64812 & n64813 ;
  assign n64796 = n64761 & ~n64774 ;
  assign n64815 = n64789 & n64796 ;
  assign n64816 = ~n64814 & ~n64815 ;
  assign n64817 = ~n64755 & ~n64816 ;
  assign n64824 = ~n64811 & ~n64817 ;
  assign n64825 = ~n64823 & n64824 ;
  assign n64826 = ~n64806 & ~n64825 ;
  assign n64784 = ~n64761 & ~n64783 ;
  assign n64785 = ~n64774 & n64784 ;
  assign n64786 = ~n64777 & ~n64785 ;
  assign n64787 = n64768 & ~n64786 ;
  assign n64762 = n64755 & ~n64761 ;
  assign n64794 = ~n64762 & n64774 ;
  assign n64795 = n64793 & ~n64794 ;
  assign n64788 = n64755 & ~n64784 ;
  assign n64790 = n64774 & n64783 ;
  assign n64791 = ~n64789 & ~n64790 ;
  assign n64792 = n64788 & n64791 ;
  assign n64797 = ~n64768 & n64796 ;
  assign n64798 = ~n64792 & ~n64797 ;
  assign n64799 = ~n64795 & n64798 ;
  assign n64800 = ~n64787 & n64799 ;
  assign n64807 = ~n64800 & n64806 ;
  assign n64827 = n64761 & n64818 ;
  assign n64828 = ~n64784 & ~n64827 ;
  assign n64829 = n64774 & ~n64828 ;
  assign n64830 = n64783 & n64797 ;
  assign n64831 = ~n64829 & ~n64830 ;
  assign n64832 = ~n64755 & ~n64831 ;
  assign n64775 = n64768 & ~n64774 ;
  assign n64776 = n64762 & n64775 ;
  assign n64833 = n64755 & ~n64783 ;
  assign n64834 = n64797 & n64833 ;
  assign n64835 = ~n64776 & ~n64834 ;
  assign n64836 = ~n64832 & n64835 ;
  assign n64837 = ~n64807 & n64836 ;
  assign n64838 = ~n64826 & n64837 ;
  assign n64839 = ~\u0_L4_reg[31]/NET0131  & ~n64838 ;
  assign n64840 = \u0_L4_reg[31]/NET0131  & n64838 ;
  assign n64841 = ~n64839 & ~n64840 ;
  assign n64891 = decrypt_pad & ~\u0_uk_K_r4_reg[51]/NET0131  ;
  assign n64892 = ~decrypt_pad & ~\u0_uk_K_r4_reg[43]/NET0131  ;
  assign n64893 = ~n64891 & ~n64892 ;
  assign n64894 = \u0_R4_reg[24]/NET0131  & ~n64893 ;
  assign n64895 = ~\u0_R4_reg[24]/NET0131  & n64893 ;
  assign n64896 = ~n64894 & ~n64895 ;
  assign n64855 = decrypt_pad & ~\u0_uk_K_r4_reg[36]/NET0131  ;
  assign n64856 = ~decrypt_pad & ~\u0_uk_K_r4_reg[28]/NET0131  ;
  assign n64857 = ~n64855 & ~n64856 ;
  assign n64858 = \u0_R4_reg[22]/NET0131  & ~n64857 ;
  assign n64859 = ~\u0_R4_reg[22]/NET0131  & n64857 ;
  assign n64860 = ~n64858 & ~n64859 ;
  assign n64862 = decrypt_pad & ~\u0_uk_K_r4_reg[14]/NET0131  ;
  assign n64863 = ~decrypt_pad & ~\u0_uk_K_r4_reg[37]/NET0131  ;
  assign n64864 = ~n64862 & ~n64863 ;
  assign n64865 = \u0_R4_reg[21]/NET0131  & ~n64864 ;
  assign n64866 = ~\u0_R4_reg[21]/NET0131  & n64864 ;
  assign n64867 = ~n64865 & ~n64866 ;
  assign n64842 = decrypt_pad & ~\u0_uk_K_r4_reg[30]/NET0131  ;
  assign n64843 = ~decrypt_pad & ~\u0_uk_K_r4_reg[22]/NET0131  ;
  assign n64844 = ~n64842 & ~n64843 ;
  assign n64845 = \u0_R4_reg[20]/NET0131  & ~n64844 ;
  assign n64846 = ~\u0_R4_reg[20]/NET0131  & n64844 ;
  assign n64847 = ~n64845 & ~n64846 ;
  assign n64848 = decrypt_pad & ~\u0_uk_K_r4_reg[15]/NET0131  ;
  assign n64849 = ~decrypt_pad & ~\u0_uk_K_r4_reg[7]/NET0131  ;
  assign n64850 = ~n64848 & ~n64849 ;
  assign n64851 = \u0_R4_reg[25]/NET0131  & ~n64850 ;
  assign n64852 = ~\u0_R4_reg[25]/NET0131  & n64850 ;
  assign n64853 = ~n64851 & ~n64852 ;
  assign n64883 = ~n64847 & n64853 ;
  assign n64926 = n64867 & n64883 ;
  assign n64927 = ~n64860 & ~n64926 ;
  assign n64897 = n64860 & n64867 ;
  assign n64898 = ~n64847 & n64897 ;
  assign n64854 = n64847 & n64853 ;
  assign n64861 = n64854 & n64860 ;
  assign n64872 = decrypt_pad & ~\u0_uk_K_r4_reg[49]/NET0131  ;
  assign n64873 = ~decrypt_pad & ~\u0_uk_K_r4_reg[45]/NET0131  ;
  assign n64874 = ~n64872 & ~n64873 ;
  assign n64875 = \u0_R4_reg[23]/NET0131  & ~n64874 ;
  assign n64876 = ~\u0_R4_reg[23]/NET0131  & n64874 ;
  assign n64877 = ~n64875 & ~n64876 ;
  assign n64928 = ~n64861 & ~n64877 ;
  assign n64929 = ~n64898 & n64928 ;
  assign n64930 = ~n64927 & n64929 ;
  assign n64886 = n64847 & ~n64853 ;
  assign n64919 = ~n64867 & n64886 ;
  assign n64920 = ~n64860 & n64919 ;
  assign n64918 = n64854 & n64867 ;
  assign n64921 = ~n64898 & ~n64918 ;
  assign n64922 = ~n64920 & n64921 ;
  assign n64923 = n64877 & ~n64922 ;
  assign n64879 = ~n64860 & ~n64877 ;
  assign n64924 = n64854 & n64879 ;
  assign n64925 = ~n64867 & n64924 ;
  assign n64931 = ~n64923 & ~n64925 ;
  assign n64932 = ~n64930 & n64931 ;
  assign n64933 = n64896 & ~n64932 ;
  assign n64899 = n64847 & ~n64860 ;
  assign n64900 = n64867 & n64899 ;
  assign n64901 = ~n64898 & ~n64900 ;
  assign n64902 = ~n64877 & ~n64901 ;
  assign n64868 = ~n64853 & n64867 ;
  assign n64904 = n64868 & n64899 ;
  assign n64905 = n64847 & ~n64867 ;
  assign n64906 = n64860 & n64877 ;
  assign n64907 = n64905 & n64906 ;
  assign n64911 = ~n64904 & ~n64907 ;
  assign n64908 = ~n64860 & n64877 ;
  assign n64909 = ~n64847 & n64908 ;
  assign n64910 = n64879 & n64886 ;
  assign n64912 = ~n64909 & ~n64910 ;
  assign n64913 = n64911 & n64912 ;
  assign n64884 = ~n64867 & n64883 ;
  assign n64885 = n64877 & n64884 ;
  assign n64903 = n64861 & ~n64867 ;
  assign n64914 = ~n64885 & ~n64903 ;
  assign n64915 = n64913 & n64914 ;
  assign n64916 = ~n64902 & n64915 ;
  assign n64917 = ~n64896 & ~n64916 ;
  assign n64887 = n64867 & n64886 ;
  assign n64888 = ~n64877 & n64887 ;
  assign n64889 = ~n64885 & ~n64888 ;
  assign n64890 = ~n64860 & ~n64889 ;
  assign n64869 = ~n64860 & n64868 ;
  assign n64870 = ~n64847 & n64869 ;
  assign n64871 = ~n64861 & ~n64870 ;
  assign n64878 = ~n64871 & n64877 ;
  assign n64880 = ~n64847 & ~n64853 ;
  assign n64881 = ~n64867 & n64880 ;
  assign n64882 = n64879 & n64881 ;
  assign n64934 = ~n64878 & ~n64882 ;
  assign n64935 = ~n64890 & n64934 ;
  assign n64936 = ~n64917 & n64935 ;
  assign n64937 = ~n64933 & n64936 ;
  assign n64938 = ~\u0_L4_reg[11]/NET0131  & n64937 ;
  assign n64939 = \u0_L4_reg[11]/NET0131  & ~n64937 ;
  assign n64940 = ~n64938 & ~n64939 ;
  assign n64947 = decrypt_pad & ~\u0_uk_K_r4_reg[42]/NET0131  ;
  assign n64948 = ~decrypt_pad & ~\u0_uk_K_r4_reg[38]/NET0131  ;
  assign n64949 = ~n64947 & ~n64948 ;
  assign n64950 = \u0_R4_reg[24]/NET0131  & ~n64949 ;
  assign n64951 = ~\u0_R4_reg[24]/NET0131  & n64949 ;
  assign n64952 = ~n64950 & ~n64951 ;
  assign n64956 = decrypt_pad & ~\u0_uk_K_r4_reg[22]/NET0131  ;
  assign n64957 = ~decrypt_pad & ~\u0_uk_K_r4_reg[14]/NET0131  ;
  assign n64958 = ~n64956 & ~n64957 ;
  assign n64959 = \u0_R4_reg[25]/NET0131  & ~n64958 ;
  assign n64960 = ~\u0_R4_reg[25]/NET0131  & n64958 ;
  assign n64961 = ~n64959 & ~n64960 ;
  assign n64978 = ~n64952 & ~n64961 ;
  assign n64941 = decrypt_pad & ~\u0_uk_K_r4_reg[7]/NET0131  ;
  assign n64942 = ~decrypt_pad & ~\u0_uk_K_r4_reg[30]/NET0131  ;
  assign n64943 = ~n64941 & ~n64942 ;
  assign n64944 = \u0_R4_reg[26]/NET0131  & ~n64943 ;
  assign n64945 = ~\u0_R4_reg[26]/NET0131  & n64943 ;
  assign n64946 = ~n64944 & ~n64945 ;
  assign n64970 = decrypt_pad & ~\u0_uk_K_r4_reg[50]/NET0131  ;
  assign n64971 = ~decrypt_pad & ~\u0_uk_K_r4_reg[42]/NET0131  ;
  assign n64972 = ~n64970 & ~n64971 ;
  assign n64973 = \u0_R4_reg[29]/NET0131  & ~n64972 ;
  assign n64974 = ~\u0_R4_reg[29]/NET0131  & n64972 ;
  assign n64975 = ~n64973 & ~n64974 ;
  assign n64979 = n64946 & n64975 ;
  assign n64988 = ~n64946 & ~n64975 ;
  assign n64991 = ~n64979 & ~n64988 ;
  assign n64992 = n64978 & ~n64991 ;
  assign n64993 = decrypt_pad & ~\u0_uk_K_r4_reg[31]/P0001  ;
  assign n64994 = ~decrypt_pad & ~\u0_uk_K_r4_reg[50]/NET0131  ;
  assign n64995 = ~n64993 & ~n64994 ;
  assign n64996 = \u0_R4_reg[28]/NET0131  & ~n64995 ;
  assign n64997 = ~\u0_R4_reg[28]/NET0131  & n64995 ;
  assign n64998 = ~n64996 & ~n64997 ;
  assign n65009 = ~n64992 & n64998 ;
  assign n64981 = n64946 & n64961 ;
  assign n65000 = ~n64981 & ~n64988 ;
  assign n64999 = ~n64946 & ~n64961 ;
  assign n64963 = decrypt_pad & ~\u0_uk_K_r4_reg[16]/NET0131  ;
  assign n64964 = ~decrypt_pad & ~\u0_uk_K_r4_reg[8]/NET0131  ;
  assign n64965 = ~n64963 & ~n64964 ;
  assign n64966 = \u0_R4_reg[27]/NET0131  & ~n64965 ;
  assign n64967 = ~\u0_R4_reg[27]/NET0131  & n64965 ;
  assign n64968 = ~n64966 & ~n64967 ;
  assign n65001 = n64952 & n64968 ;
  assign n65002 = ~n64999 & n65001 ;
  assign n65003 = n65000 & n65002 ;
  assign n65004 = n64952 & n64961 ;
  assign n65005 = ~n64978 & ~n65004 ;
  assign n64953 = n64946 & n64952 ;
  assign n65006 = ~n64968 & n64975 ;
  assign n65007 = ~n64953 & n65006 ;
  assign n65008 = n65005 & n65007 ;
  assign n65010 = ~n65003 & ~n65008 ;
  assign n65011 = n65009 & n65010 ;
  assign n65014 = n64946 & ~n64968 ;
  assign n65015 = ~n65001 & ~n65014 ;
  assign n65016 = ~n64952 & n64975 ;
  assign n65017 = ~n64953 & ~n64961 ;
  assign n65018 = ~n65016 & n65017 ;
  assign n65019 = ~n65015 & n65018 ;
  assign n64954 = ~n64946 & ~n64952 ;
  assign n64955 = ~n64953 & ~n64954 ;
  assign n64989 = ~n64961 & n64968 ;
  assign n65020 = n64975 & ~n64989 ;
  assign n65021 = ~n64955 & n65020 ;
  assign n65012 = n64952 & ~n64968 ;
  assign n65013 = ~n65000 & n65012 ;
  assign n65022 = ~n64998 & ~n65013 ;
  assign n65023 = ~n65021 & n65022 ;
  assign n65024 = ~n65019 & n65023 ;
  assign n65025 = ~n65011 & ~n65024 ;
  assign n64962 = ~n64955 & n64961 ;
  assign n64969 = ~n64962 & ~n64968 ;
  assign n64980 = n64978 & n64979 ;
  assign n64982 = ~n64952 & ~n64975 ;
  assign n64983 = n64981 & n64982 ;
  assign n64984 = ~n64980 & ~n64983 ;
  assign n64976 = ~n64961 & ~n64975 ;
  assign n64977 = n64952 & n64976 ;
  assign n64985 = n64968 & ~n64977 ;
  assign n64986 = n64984 & n64985 ;
  assign n64987 = ~n64969 & ~n64986 ;
  assign n64990 = n64988 & n64989 ;
  assign n65026 = ~n64987 & ~n64990 ;
  assign n65027 = ~n65025 & n65026 ;
  assign n65028 = ~\u0_L4_reg[22]/NET0131  & ~n65027 ;
  assign n65029 = \u0_L4_reg[22]/NET0131  & n65027 ;
  assign n65030 = ~n65028 & ~n65029 ;
  assign n65034 = ~n64761 & ~n64774 ;
  assign n65035 = ~n64768 & ~n65034 ;
  assign n65039 = n64818 & n65034 ;
  assign n65040 = ~n65035 & ~n65039 ;
  assign n65041 = n64755 & ~n65040 ;
  assign n65036 = ~n64761 & n64768 ;
  assign n65037 = ~n64755 & ~n65036 ;
  assign n65038 = ~n65035 & n65037 ;
  assign n65031 = n64768 & n64774 ;
  assign n65032 = n64784 & n65031 ;
  assign n65033 = n64806 & ~n65032 ;
  assign n65042 = n64761 & n64790 ;
  assign n65043 = n65033 & ~n65042 ;
  assign n65044 = ~n65038 & n65043 ;
  assign n65045 = ~n65041 & n65044 ;
  assign n65046 = n64774 & ~n64784 ;
  assign n65047 = n64809 & ~n65046 ;
  assign n65048 = ~n64755 & ~n65047 ;
  assign n65052 = n64761 & n64821 ;
  assign n65050 = ~n64812 & ~n64820 ;
  assign n65051 = n64768 & n65050 ;
  assign n65049 = n64790 & n64813 ;
  assign n65053 = n64755 & ~n65049 ;
  assign n65054 = ~n65051 & n65053 ;
  assign n65055 = ~n65052 & n65054 ;
  assign n65056 = ~n65048 & ~n65055 ;
  assign n65057 = n64761 & n64768 ;
  assign n65058 = n64820 & n65057 ;
  assign n65059 = ~n64806 & ~n65058 ;
  assign n65060 = ~n64830 & n65059 ;
  assign n65061 = ~n65056 & n65060 ;
  assign n65062 = ~n65045 & ~n65061 ;
  assign n65063 = ~\u0_L4_reg[17]/NET0131  & n65062 ;
  assign n65064 = \u0_L4_reg[17]/NET0131  & ~n65062 ;
  assign n65065 = ~n65063 & ~n65064 ;
  assign n65066 = decrypt_pad & ~\u0_uk_K_r4_reg[26]/NET0131  ;
  assign n65067 = ~decrypt_pad & ~\u0_uk_K_r4_reg[20]/NET0131  ;
  assign n65068 = ~n65066 & ~n65067 ;
  assign n65069 = \u0_R4_reg[8]/NET0131  & ~n65068 ;
  assign n65070 = ~\u0_R4_reg[8]/NET0131  & n65068 ;
  assign n65071 = ~n65069 & ~n65070 ;
  assign n65072 = decrypt_pad & ~\u0_uk_K_r4_reg[3]/NET0131  ;
  assign n65073 = ~decrypt_pad & ~\u0_uk_K_r4_reg[54]/NET0131  ;
  assign n65074 = ~n65072 & ~n65073 ;
  assign n65075 = \u0_R4_reg[7]/NET0131  & ~n65074 ;
  assign n65076 = ~\u0_R4_reg[7]/NET0131  & n65074 ;
  assign n65077 = ~n65075 & ~n65076 ;
  assign n65091 = decrypt_pad & ~\u0_uk_K_r4_reg[18]/NET0131  ;
  assign n65092 = ~decrypt_pad & ~\u0_uk_K_r4_reg[12]/NET0131  ;
  assign n65093 = ~n65091 & ~n65092 ;
  assign n65094 = \u0_R4_reg[5]/NET0131  & ~n65093 ;
  assign n65095 = ~\u0_R4_reg[5]/NET0131  & n65093 ;
  assign n65096 = ~n65094 & ~n65095 ;
  assign n65078 = decrypt_pad & ~\u0_uk_K_r4_reg[39]/NET0131  ;
  assign n65079 = ~decrypt_pad & ~\u0_uk_K_r4_reg[33]/NET0131  ;
  assign n65080 = ~n65078 & ~n65079 ;
  assign n65081 = \u0_R4_reg[4]/NET0131  & ~n65080 ;
  assign n65082 = ~\u0_R4_reg[4]/NET0131  & n65080 ;
  assign n65083 = ~n65081 & ~n65082 ;
  assign n65084 = decrypt_pad & ~\u0_uk_K_r4_reg[6]/NET0131  ;
  assign n65085 = ~decrypt_pad & ~\u0_uk_K_r4_reg[25]/NET0131  ;
  assign n65086 = ~n65084 & ~n65085 ;
  assign n65087 = \u0_R4_reg[9]/NET0131  & ~n65086 ;
  assign n65088 = ~\u0_R4_reg[9]/NET0131  & n65086 ;
  assign n65089 = ~n65087 & ~n65088 ;
  assign n65106 = ~n65083 & n65089 ;
  assign n65107 = ~n65096 & n65106 ;
  assign n65098 = decrypt_pad & ~\u0_uk_K_r4_reg[41]/NET0131  ;
  assign n65099 = ~decrypt_pad & ~\u0_uk_K_r4_reg[3]/NET0131  ;
  assign n65100 = ~n65098 & ~n65099 ;
  assign n65101 = \u0_R4_reg[6]/NET0131  & ~n65100 ;
  assign n65102 = ~\u0_R4_reg[6]/NET0131  & n65100 ;
  assign n65103 = ~n65101 & ~n65102 ;
  assign n65108 = n65083 & n65096 ;
  assign n65109 = n65083 & ~n65089 ;
  assign n65110 = ~n65108 & ~n65109 ;
  assign n65111 = n65103 & ~n65110 ;
  assign n65112 = ~n65107 & ~n65111 ;
  assign n65113 = ~n65077 & ~n65112 ;
  assign n65114 = ~n65089 & n65096 ;
  assign n65115 = ~n65107 & ~n65114 ;
  assign n65116 = ~n65103 & ~n65115 ;
  assign n65090 = n65083 & n65089 ;
  assign n65097 = n65090 & ~n65096 ;
  assign n65104 = n65097 & n65103 ;
  assign n65105 = n65077 & n65104 ;
  assign n65117 = ~n65077 & ~n65096 ;
  assign n65118 = n65089 & ~n65103 ;
  assign n65119 = n65117 & n65118 ;
  assign n65120 = n65096 & n65103 ;
  assign n65121 = n65106 & n65120 ;
  assign n65122 = ~n65119 & ~n65121 ;
  assign n65123 = ~n65105 & n65122 ;
  assign n65124 = ~n65116 & n65123 ;
  assign n65125 = ~n65113 & n65124 ;
  assign n65126 = ~n65071 & ~n65125 ;
  assign n65143 = ~n65083 & ~n65089 ;
  assign n65144 = ~n65104 & ~n65143 ;
  assign n65145 = n65071 & ~n65144 ;
  assign n65127 = ~n65096 & n65103 ;
  assign n65146 = n65106 & ~n65127 ;
  assign n65147 = ~n65145 & ~n65146 ;
  assign n65130 = n65096 & ~n65103 ;
  assign n65148 = ~n65077 & ~n65130 ;
  assign n65149 = ~n65147 & n65148 ;
  assign n65128 = ~n65089 & n65127 ;
  assign n65129 = ~n65083 & n65128 ;
  assign n65131 = n65083 & n65130 ;
  assign n65132 = ~n65129 & ~n65131 ;
  assign n65133 = n65077 & ~n65132 ;
  assign n65134 = ~n65096 & n65109 ;
  assign n65135 = ~n65103 & n65134 ;
  assign n65136 = n65108 & n65118 ;
  assign n65137 = ~n65083 & n65103 ;
  assign n65138 = n65077 & n65096 ;
  assign n65139 = ~n65137 & n65138 ;
  assign n65140 = ~n65136 & ~n65139 ;
  assign n65141 = ~n65135 & n65140 ;
  assign n65142 = n65071 & ~n65141 ;
  assign n65150 = ~n65133 & ~n65142 ;
  assign n65151 = ~n65149 & n65150 ;
  assign n65152 = ~n65126 & n65151 ;
  assign n65153 = \u0_L4_reg[2]/NET0131  & n65152 ;
  assign n65154 = ~\u0_L4_reg[2]/NET0131  & ~n65152 ;
  assign n65155 = ~n65153 & ~n65154 ;
  assign n65177 = ~n64860 & n64883 ;
  assign n65178 = ~n64887 & ~n65177 ;
  assign n65179 = ~n64903 & n65178 ;
  assign n65180 = n64877 & ~n65179 ;
  assign n65173 = n64860 & n64884 ;
  assign n65174 = ~n64847 & n64868 ;
  assign n65175 = ~n65173 & ~n65174 ;
  assign n65176 = ~n64877 & ~n65175 ;
  assign n65181 = ~n64920 & ~n64924 ;
  assign n65182 = ~n65176 & n65181 ;
  assign n65183 = ~n65180 & n65182 ;
  assign n65184 = ~n64896 & ~n65183 ;
  assign n65158 = n64847 & ~n64868 ;
  assign n65159 = n64879 & ~n65158 ;
  assign n65156 = n64853 & n64867 ;
  assign n65157 = n64860 & n65156 ;
  assign n65160 = n64854 & n64908 ;
  assign n65161 = ~n65157 & ~n65160 ;
  assign n65162 = ~n64870 & n65161 ;
  assign n65163 = ~n65159 & n65162 ;
  assign n65164 = n64896 & ~n65163 ;
  assign n65165 = ~n64881 & ~n64926 ;
  assign n65166 = ~n64887 & n65165 ;
  assign n65167 = n64906 & ~n65166 ;
  assign n65168 = ~n64918 & ~n64919 ;
  assign n65169 = n64860 & n65168 ;
  assign n65170 = ~n64860 & ~n64880 ;
  assign n65171 = ~n64877 & ~n65170 ;
  assign n65172 = ~n65169 & n65171 ;
  assign n65185 = ~n65167 & ~n65172 ;
  assign n65186 = ~n65164 & n65185 ;
  assign n65187 = ~n65184 & n65186 ;
  assign n65188 = ~\u0_L4_reg[4]/NET0131  & ~n65187 ;
  assign n65189 = \u0_L4_reg[4]/NET0131  & n65187 ;
  assign n65190 = ~n65188 & ~n65189 ;
  assign n65191 = decrypt_pad & ~\u0_uk_K_r4_reg[45]/NET0131  ;
  assign n65192 = ~decrypt_pad & ~\u0_uk_K_r4_reg[9]/NET0131  ;
  assign n65193 = ~n65191 & ~n65192 ;
  assign n65194 = \u0_R4_reg[31]/P0001  & ~n65193 ;
  assign n65195 = ~\u0_R4_reg[31]/P0001  & n65193 ;
  assign n65196 = ~n65194 & ~n65195 ;
  assign n65197 = decrypt_pad & ~\u0_uk_K_r4_reg[28]/NET0131  ;
  assign n65198 = ~decrypt_pad & ~\u0_uk_K_r4_reg[51]/NET0131  ;
  assign n65199 = ~n65197 & ~n65198 ;
  assign n65200 = \u0_R4_reg[29]/NET0131  & ~n65199 ;
  assign n65201 = ~\u0_R4_reg[29]/NET0131  & n65199 ;
  assign n65202 = ~n65200 & ~n65201 ;
  assign n65210 = decrypt_pad & ~\u0_uk_K_r4_reg[29]/NET0131  ;
  assign n65211 = ~decrypt_pad & ~\u0_uk_K_r4_reg[21]/NET0131  ;
  assign n65212 = ~n65210 & ~n65211 ;
  assign n65213 = \u0_R4_reg[30]/NET0131  & ~n65212 ;
  assign n65214 = ~\u0_R4_reg[30]/NET0131  & n65212 ;
  assign n65215 = ~n65213 & ~n65214 ;
  assign n65203 = decrypt_pad & ~\u0_uk_K_r4_reg[44]/NET0131  ;
  assign n65204 = ~decrypt_pad & ~\u0_uk_K_r4_reg[36]/NET0131  ;
  assign n65205 = ~n65203 & ~n65204 ;
  assign n65206 = \u0_R4_reg[1]/NET0131  & ~n65205 ;
  assign n65207 = ~\u0_R4_reg[1]/NET0131  & n65205 ;
  assign n65208 = ~n65206 & ~n65207 ;
  assign n65216 = decrypt_pad & ~\u0_uk_K_r4_reg[1]/NET0131  ;
  assign n65217 = ~decrypt_pad & ~\u0_uk_K_r4_reg[52]/NET0131  ;
  assign n65218 = ~n65216 & ~n65217 ;
  assign n65219 = \u0_R4_reg[28]/NET0131  & ~n65218 ;
  assign n65220 = ~\u0_R4_reg[28]/NET0131  & n65218 ;
  assign n65221 = ~n65219 & ~n65220 ;
  assign n65240 = ~n65208 & n65221 ;
  assign n65241 = ~n65215 & n65240 ;
  assign n65242 = n65202 & n65241 ;
  assign n65233 = decrypt_pad & ~\u0_uk_K_r4_reg[23]/P0001  ;
  assign n65234 = ~decrypt_pad & ~\u0_uk_K_r4_reg[15]/NET0131  ;
  assign n65235 = ~n65233 & ~n65234 ;
  assign n65236 = \u0_R4_reg[32]/NET0131  & ~n65235 ;
  assign n65237 = ~\u0_R4_reg[32]/NET0131  & n65235 ;
  assign n65238 = ~n65236 & ~n65237 ;
  assign n65209 = n65202 & ~n65208 ;
  assign n65224 = ~n65215 & n65221 ;
  assign n65239 = ~n65209 & ~n65224 ;
  assign n65243 = n65238 & ~n65239 ;
  assign n65244 = ~n65242 & n65243 ;
  assign n65228 = ~n65202 & ~n65221 ;
  assign n65231 = n65208 & n65228 ;
  assign n65232 = n65215 & n65231 ;
  assign n65222 = n65215 & ~n65221 ;
  assign n65223 = n65209 & n65222 ;
  assign n65225 = ~n65202 & n65208 ;
  assign n65226 = n65224 & n65225 ;
  assign n65227 = ~n65223 & ~n65226 ;
  assign n65229 = ~n65215 & n65228 ;
  assign n65230 = ~n65208 & n65229 ;
  assign n65245 = n65227 & ~n65230 ;
  assign n65246 = ~n65232 & n65245 ;
  assign n65247 = ~n65244 & n65246 ;
  assign n65248 = n65196 & ~n65247 ;
  assign n65262 = n65209 & ~n65215 ;
  assign n65263 = n65196 & ~n65262 ;
  assign n65264 = ~n65215 & n65263 ;
  assign n65249 = n65202 & n65208 ;
  assign n65261 = n65215 & ~n65249 ;
  assign n65265 = n65221 & ~n65261 ;
  assign n65266 = ~n65264 & n65265 ;
  assign n65250 = ~n65208 & ~n65221 ;
  assign n65251 = n65215 & n65250 ;
  assign n65252 = ~n65196 & ~n65249 ;
  assign n65253 = ~n65251 & n65252 ;
  assign n65254 = ~n65242 & n65253 ;
  assign n65255 = n65215 & n65221 ;
  assign n65256 = ~n65202 & n65255 ;
  assign n65257 = ~n65208 & n65256 ;
  assign n65258 = n65196 & ~n65231 ;
  assign n65259 = ~n65257 & n65258 ;
  assign n65260 = ~n65254 & ~n65259 ;
  assign n65267 = ~n65238 & ~n65260 ;
  assign n65268 = ~n65266 & n65267 ;
  assign n65269 = ~n65229 & ~n65256 ;
  assign n65270 = ~n65242 & n65269 ;
  assign n65271 = ~n65196 & ~n65270 ;
  assign n65272 = ~n65221 & n65249 ;
  assign n65273 = n65215 & n65272 ;
  assign n65274 = n65238 & ~n65273 ;
  assign n65275 = ~n65271 & n65274 ;
  assign n65276 = ~n65268 & ~n65275 ;
  assign n65277 = ~n65248 & ~n65276 ;
  assign n65278 = \u0_L4_reg[5]/NET0131  & ~n65277 ;
  assign n65279 = ~\u0_L4_reg[5]/NET0131  & n65277 ;
  assign n65280 = ~n65278 & ~n65279 ;
  assign n65290 = ~n64860 & ~n64867 ;
  assign n65299 = ~n64898 & ~n65290 ;
  assign n65300 = ~n64853 & ~n65299 ;
  assign n65301 = n65168 & ~n65300 ;
  assign n65302 = n64877 & ~n65301 ;
  assign n65281 = n64860 & ~n64886 ;
  assign n65282 = n64867 & ~n64899 ;
  assign n65283 = ~n65281 & n65282 ;
  assign n65303 = ~n64877 & n65283 ;
  assign n65304 = ~n64924 & ~n65173 ;
  assign n65305 = ~n65303 & n65304 ;
  assign n65306 = ~n65302 & n65305 ;
  assign n65307 = ~n64896 & ~n65306 ;
  assign n65286 = ~n64883 & n65281 ;
  assign n65287 = ~n64881 & ~n65286 ;
  assign n65288 = ~n64877 & ~n65287 ;
  assign n65284 = ~n64926 & ~n65283 ;
  assign n65285 = n64877 & ~n65284 ;
  assign n65289 = n64860 & n64881 ;
  assign n65291 = n64883 & n65290 ;
  assign n65292 = ~n65289 & ~n65291 ;
  assign n65293 = ~n64903 & ~n64910 ;
  assign n65294 = n65292 & n65293 ;
  assign n65295 = ~n65285 & n65294 ;
  assign n65296 = ~n65288 & n65295 ;
  assign n65297 = n64896 & ~n65296 ;
  assign n65298 = n64908 & n65156 ;
  assign n65308 = ~n64920 & ~n65298 ;
  assign n65309 = ~n65297 & n65308 ;
  assign n65310 = ~n65307 & n65309 ;
  assign n65311 = \u0_L4_reg[29]/NET0131  & ~n65310 ;
  assign n65312 = ~\u0_L4_reg[29]/NET0131  & n65310 ;
  assign n65313 = ~n65311 & ~n65312 ;
  assign n65314 = decrypt_pad & ~\u0_uk_K_r4_reg[10]/NET0131  ;
  assign n65315 = ~decrypt_pad & ~\u0_uk_K_r4_reg[4]/NET0131  ;
  assign n65316 = ~n65314 & ~n65315 ;
  assign n65317 = \u0_R4_reg[13]/NET0131  & ~n65316 ;
  assign n65318 = ~\u0_R4_reg[13]/NET0131  & n65316 ;
  assign n65319 = ~n65317 & ~n65318 ;
  assign n65320 = decrypt_pad & ~\u0_uk_K_r4_reg[19]/NET0131  ;
  assign n65321 = ~decrypt_pad & ~\u0_uk_K_r4_reg[13]/NET0131  ;
  assign n65322 = ~n65320 & ~n65321 ;
  assign n65323 = \u0_R4_reg[15]/NET0131  & ~n65322 ;
  assign n65324 = ~\u0_R4_reg[15]/NET0131  & n65322 ;
  assign n65325 = ~n65323 & ~n65324 ;
  assign n65326 = n65319 & n65325 ;
  assign n65327 = decrypt_pad & ~\u0_uk_K_r4_reg[11]/NET0131  ;
  assign n65328 = ~decrypt_pad & ~\u0_uk_K_r4_reg[5]/NET0131  ;
  assign n65329 = ~n65327 & ~n65328 ;
  assign n65330 = \u0_R4_reg[14]/NET0131  & ~n65329 ;
  assign n65331 = ~\u0_R4_reg[14]/NET0131  & n65329 ;
  assign n65332 = ~n65330 & ~n65331 ;
  assign n65333 = n65326 & n65332 ;
  assign n65334 = decrypt_pad & ~\u0_uk_K_r4_reg[48]/NET0131  ;
  assign n65335 = ~decrypt_pad & ~\u0_uk_K_r4_reg[10]/NET0131  ;
  assign n65336 = ~n65334 & ~n65335 ;
  assign n65337 = \u0_R4_reg[12]/NET0131  & ~n65336 ;
  assign n65338 = ~\u0_R4_reg[12]/NET0131  & n65336 ;
  assign n65339 = ~n65337 & ~n65338 ;
  assign n65340 = n65333 & ~n65339 ;
  assign n65341 = decrypt_pad & ~\u0_uk_K_r4_reg[32]/NET0131  ;
  assign n65342 = ~decrypt_pad & ~\u0_uk_K_r4_reg[26]/NET0131  ;
  assign n65343 = ~n65341 & ~n65342 ;
  assign n65344 = \u0_R4_reg[17]/NET0131  & ~n65343 ;
  assign n65345 = ~\u0_R4_reg[17]/NET0131  & n65343 ;
  assign n65346 = ~n65344 & ~n65345 ;
  assign n65347 = n65339 & n65346 ;
  assign n65348 = n65326 & n65347 ;
  assign n65352 = decrypt_pad & ~\u0_uk_K_r4_reg[27]/P0001  ;
  assign n65353 = ~decrypt_pad & ~\u0_uk_K_r4_reg[46]/NET0131  ;
  assign n65354 = ~n65352 & ~n65353 ;
  assign n65355 = \u0_R4_reg[16]/NET0131  & ~n65354 ;
  assign n65356 = ~\u0_R4_reg[16]/NET0131  & n65354 ;
  assign n65357 = ~n65355 & ~n65356 ;
  assign n65371 = ~n65348 & ~n65357 ;
  assign n65349 = ~n65319 & n65325 ;
  assign n65350 = ~n65339 & ~n65346 ;
  assign n65351 = n65349 & n65350 ;
  assign n65366 = ~n65319 & n65346 ;
  assign n65369 = ~n65332 & n65339 ;
  assign n65370 = n65366 & n65369 ;
  assign n65372 = ~n65351 & ~n65370 ;
  assign n65373 = n65371 & n65372 ;
  assign n65374 = ~n65340 & n65373 ;
  assign n65358 = n65319 & n65350 ;
  assign n65359 = n65332 & n65358 ;
  assign n65360 = ~n65319 & ~n65339 ;
  assign n65361 = ~n65332 & ~n65346 ;
  assign n65362 = n65360 & n65361 ;
  assign n65363 = ~n65359 & ~n65362 ;
  assign n65364 = n65339 & ~n65346 ;
  assign n65365 = n65332 & n65364 ;
  assign n65367 = ~n65365 & ~n65366 ;
  assign n65368 = ~n65325 & ~n65367 ;
  assign n65375 = n65363 & ~n65368 ;
  assign n65376 = n65374 & n65375 ;
  assign n65392 = n65325 & n65366 ;
  assign n65393 = ~n65339 & n65392 ;
  assign n65381 = ~n65325 & ~n65332 ;
  assign n65382 = n65319 & n65339 ;
  assign n65383 = ~n65360 & ~n65382 ;
  assign n65384 = n65381 & n65383 ;
  assign n65385 = n65332 & n65346 ;
  assign n65386 = n65382 & n65385 ;
  assign n65394 = n65357 & ~n65386 ;
  assign n65395 = ~n65384 & n65394 ;
  assign n65396 = ~n65393 & n65395 ;
  assign n65377 = ~n65319 & ~n65346 ;
  assign n65378 = ~n65325 & n65377 ;
  assign n65379 = ~n65339 & n65378 ;
  assign n65380 = n65332 & n65379 ;
  assign n65387 = n65326 & n65364 ;
  assign n65388 = ~n65339 & n65346 ;
  assign n65389 = n65319 & n65388 ;
  assign n65390 = ~n65332 & n65389 ;
  assign n65391 = ~n65387 & ~n65390 ;
  assign n65397 = ~n65380 & n65391 ;
  assign n65398 = n65396 & n65397 ;
  assign n65399 = ~n65376 & ~n65398 ;
  assign n65400 = ~n65339 & n65361 ;
  assign n65401 = ~n65365 & ~n65400 ;
  assign n65402 = n65349 & ~n65401 ;
  assign n65403 = ~n65332 & n65387 ;
  assign n65404 = n65381 & n65389 ;
  assign n65405 = ~n65403 & ~n65404 ;
  assign n65406 = ~n65402 & n65405 ;
  assign n65407 = ~n65399 & n65406 ;
  assign n65408 = ~\u0_L4_reg[20]/NET0131  & ~n65407 ;
  assign n65409 = \u0_L4_reg[20]/NET0131  & n65407 ;
  assign n65410 = ~n65408 & ~n65409 ;
  assign n65412 = n65103 & n65107 ;
  assign n65411 = ~n65083 & n65114 ;
  assign n65413 = ~n65135 & ~n65411 ;
  assign n65414 = ~n65412 & n65413 ;
  assign n65415 = ~n65077 & ~n65414 ;
  assign n65423 = n65077 & ~n65134 ;
  assign n65421 = ~n65103 & n65109 ;
  assign n65422 = n65096 & ~n65421 ;
  assign n65424 = ~n65107 & ~n65422 ;
  assign n65425 = n65423 & n65424 ;
  assign n65416 = n65077 & n65083 ;
  assign n65417 = n65103 & ~n65114 ;
  assign n65418 = n65416 & n65417 ;
  assign n65419 = ~n65083 & ~n65117 ;
  assign n65420 = n65118 & n65419 ;
  assign n65426 = ~n65418 & ~n65420 ;
  assign n65427 = ~n65425 & n65426 ;
  assign n65428 = ~n65415 & n65427 ;
  assign n65429 = ~n65071 & ~n65428 ;
  assign n65430 = n65109 & n65120 ;
  assign n65431 = ~n65136 & ~n65430 ;
  assign n65432 = ~n65077 & ~n65431 ;
  assign n65433 = ~n65077 & ~n65097 ;
  assign n65434 = ~n65128 & n65433 ;
  assign n65437 = n65089 & n65137 ;
  assign n65435 = ~n65096 & ~n65103 ;
  assign n65436 = ~n65089 & n65435 ;
  assign n65438 = n65077 & ~n65436 ;
  assign n65439 = ~n65437 & n65438 ;
  assign n65440 = ~n65434 & ~n65439 ;
  assign n65441 = ~n65103 & n65143 ;
  assign n65442 = n65096 & n65441 ;
  assign n65443 = n65122 & n65431 ;
  assign n65444 = ~n65442 & n65443 ;
  assign n65445 = ~n65440 & n65444 ;
  assign n65446 = n65071 & ~n65445 ;
  assign n65447 = ~n65432 & ~n65446 ;
  assign n65448 = ~n65429 & n65447 ;
  assign n65449 = ~\u0_L4_reg[13]/NET0131  & n65448 ;
  assign n65450 = \u0_L4_reg[13]/NET0131  & ~n65448 ;
  assign n65451 = ~n65449 & ~n65450 ;
  assign n65452 = n65319 & ~n65332 ;
  assign n65454 = n65339 & n65452 ;
  assign n65464 = n65347 & n65381 ;
  assign n65470 = ~n65454 & ~n65464 ;
  assign n65471 = ~n65379 & n65470 ;
  assign n65465 = ~n65332 & n65346 ;
  assign n65466 = n65339 & n65349 ;
  assign n65467 = ~n65465 & n65466 ;
  assign n65468 = n65325 & n65388 ;
  assign n65469 = ~n65332 & n65468 ;
  assign n65472 = ~n65467 & ~n65469 ;
  assign n65473 = n65471 & n65472 ;
  assign n65474 = n65363 & n65473 ;
  assign n65475 = ~n65357 & ~n65474 ;
  assign n65458 = ~n65358 & ~n65370 ;
  assign n65459 = n65325 & ~n65458 ;
  assign n65453 = n65346 & ~n65452 ;
  assign n65455 = ~n65325 & ~n65350 ;
  assign n65456 = ~n65453 & n65455 ;
  assign n65457 = ~n65454 & n65456 ;
  assign n65460 = ~n65383 & n65385 ;
  assign n65461 = ~n65457 & ~n65460 ;
  assign n65462 = ~n65459 & n65461 ;
  assign n65463 = n65357 & ~n65462 ;
  assign n65476 = ~n65362 & ~n65460 ;
  assign n65477 = ~n65325 & ~n65476 ;
  assign n65478 = ~n65340 & ~n65403 ;
  assign n65479 = ~n65477 & n65478 ;
  assign n65480 = ~n65463 & n65479 ;
  assign n65481 = ~n65475 & n65480 ;
  assign n65482 = ~\u0_L4_reg[10]/NET0131  & ~n65481 ;
  assign n65483 = \u0_L4_reg[10]/NET0131  & n65481 ;
  assign n65484 = ~n65482 & ~n65483 ;
  assign n65487 = n64978 & n64988 ;
  assign n65488 = ~n65004 & ~n65487 ;
  assign n65489 = n64968 & ~n65488 ;
  assign n65486 = n64991 & n65005 ;
  assign n65485 = ~n64968 & n64980 ;
  assign n65490 = n64998 & ~n65485 ;
  assign n65491 = ~n65486 & n65490 ;
  assign n65492 = ~n65489 & n65491 ;
  assign n65498 = ~n64981 & ~n64999 ;
  assign n65499 = n64952 & n64975 ;
  assign n65500 = ~n64982 & ~n65499 ;
  assign n65502 = n65498 & n65500 ;
  assign n65497 = ~n64976 & n64991 ;
  assign n65501 = ~n65498 & ~n65500 ;
  assign n65503 = ~n65497 & ~n65501 ;
  assign n65504 = ~n65502 & n65503 ;
  assign n65494 = n64961 & n64975 ;
  assign n65495 = ~n64976 & ~n65494 ;
  assign n65496 = ~n64968 & ~n65495 ;
  assign n65505 = n64952 & n65014 ;
  assign n65493 = n64989 & n65016 ;
  assign n65506 = ~n64998 & ~n65493 ;
  assign n65507 = ~n65505 & n65506 ;
  assign n65508 = ~n65496 & n65507 ;
  assign n65509 = ~n65504 & n65508 ;
  assign n65510 = ~n65492 & ~n65509 ;
  assign n65511 = \u0_L4_reg[12]/NET0131  & n65510 ;
  assign n65512 = ~\u0_L4_reg[12]/NET0131  & ~n65510 ;
  assign n65513 = ~n65511 & ~n65512 ;
  assign n65526 = ~n64827 & ~n65031 ;
  assign n65527 = ~n64755 & ~n65526 ;
  assign n65528 = n64755 & n64821 ;
  assign n65529 = ~n64785 & ~n64806 ;
  assign n65525 = n64793 & n64808 ;
  assign n65530 = ~n65042 & ~n65525 ;
  assign n65531 = n65529 & n65530 ;
  assign n65532 = ~n65528 & n65531 ;
  assign n65533 = ~n65527 & n65532 ;
  assign n65534 = n64788 & n64810 ;
  assign n65535 = n64806 & ~n65039 ;
  assign n65536 = ~n64834 & n65535 ;
  assign n65537 = ~n65534 & n65536 ;
  assign n65538 = ~n65533 & ~n65537 ;
  assign n65514 = ~n64768 & ~n65050 ;
  assign n65515 = ~n64815 & ~n65514 ;
  assign n65516 = n64806 & ~n65515 ;
  assign n65517 = ~n64761 & ~n64809 ;
  assign n65518 = ~n65050 & n65517 ;
  assign n65519 = ~n65516 & ~n65518 ;
  assign n65520 = ~n64755 & ~n65519 ;
  assign n65521 = ~n64755 & n64790 ;
  assign n65522 = n65057 & n65521 ;
  assign n65523 = ~n64775 & ~n64821 ;
  assign n65524 = n64762 & ~n65523 ;
  assign n65539 = ~n65522 & ~n65524 ;
  assign n65540 = ~n65520 & n65539 ;
  assign n65541 = ~n65538 & n65540 ;
  assign n65542 = \u0_L4_reg[23]/NET0131  & ~n65541 ;
  assign n65543 = ~\u0_L4_reg[23]/NET0131  & n65541 ;
  assign n65544 = ~n65542 & ~n65543 ;
  assign n65545 = n65202 & n65221 ;
  assign n65546 = ~n65262 & ~n65545 ;
  assign n65547 = ~n65231 & n65546 ;
  assign n65548 = n65196 & ~n65547 ;
  assign n65549 = ~n65202 & ~n65208 ;
  assign n65550 = n65224 & n65549 ;
  assign n65551 = ~n65548 & ~n65550 ;
  assign n65552 = ~n65238 & ~n65551 ;
  assign n65571 = ~n65215 & n65272 ;
  assign n65568 = ~n65202 & n65221 ;
  assign n65569 = ~n65215 & n65238 ;
  assign n65570 = n65568 & ~n65569 ;
  assign n65572 = ~n65223 & ~n65570 ;
  assign n65573 = ~n65230 & n65572 ;
  assign n65574 = ~n65571 & n65573 ;
  assign n65575 = ~n65196 & ~n65574 ;
  assign n65553 = n65208 & n65229 ;
  assign n65554 = ~n65273 & ~n65553 ;
  assign n65555 = n65196 & ~n65554 ;
  assign n65556 = n65196 & ~n65202 ;
  assign n65557 = n65250 & n65556 ;
  assign n65563 = ~n65223 & ~n65557 ;
  assign n65562 = n65225 & n65255 ;
  assign n65558 = ~n65215 & n65545 ;
  assign n65559 = ~n65202 & n65215 ;
  assign n65560 = ~n65196 & n65208 ;
  assign n65561 = n65559 & n65560 ;
  assign n65564 = ~n65558 & ~n65561 ;
  assign n65565 = ~n65562 & n65564 ;
  assign n65566 = n65563 & n65565 ;
  assign n65567 = n65238 & ~n65566 ;
  assign n65576 = ~n65555 & ~n65567 ;
  assign n65577 = ~n65575 & n65576 ;
  assign n65578 = ~n65552 & n65577 ;
  assign n65579 = \u0_L4_reg[15]/P0001  & n65578 ;
  assign n65580 = ~\u0_L4_reg[15]/P0001  & ~n65578 ;
  assign n65581 = ~n65579 & ~n65580 ;
  assign n65585 = n65096 & n65106 ;
  assign n65586 = ~n65441 & ~n65585 ;
  assign n65587 = n65077 & n65586 ;
  assign n65588 = ~n65096 & n65137 ;
  assign n65589 = ~n65077 & ~n65430 ;
  assign n65590 = ~n65588 & n65589 ;
  assign n65591 = ~n65107 & ~n65108 ;
  assign n65592 = ~n65421 & n65591 ;
  assign n65593 = n65590 & n65592 ;
  assign n65594 = ~n65587 & ~n65593 ;
  assign n65582 = ~n65106 & ~n65109 ;
  assign n65583 = n65127 & n65582 ;
  assign n65584 = ~n65071 & ~n65430 ;
  assign n65595 = ~n65583 & n65584 ;
  assign n65596 = ~n65594 & n65595 ;
  assign n65597 = n65586 & n65590 ;
  assign n65599 = n65103 & n65411 ;
  assign n65598 = n65090 & n65096 ;
  assign n65600 = n65423 & ~n65598 ;
  assign n65601 = ~n65599 & n65600 ;
  assign n65602 = ~n65597 & ~n65601 ;
  assign n65603 = ~n65097 & ~n65416 ;
  assign n65604 = ~n65103 & ~n65603 ;
  assign n65605 = n65071 & ~n65412 ;
  assign n65606 = ~n65604 & n65605 ;
  assign n65607 = ~n65602 & n65606 ;
  assign n65608 = ~n65596 & ~n65607 ;
  assign n65609 = ~\u0_L4_reg[28]/NET0131  & n65608 ;
  assign n65610 = \u0_L4_reg[28]/NET0131  & ~n65608 ;
  assign n65611 = ~n65609 & ~n65610 ;
  assign n65612 = decrypt_pad & ~\u0_uk_K_r4_reg[9]/NET0131  ;
  assign n65613 = ~decrypt_pad & ~\u0_uk_K_r4_reg[1]/NET0131  ;
  assign n65614 = ~n65612 & ~n65613 ;
  assign n65615 = \u0_R4_reg[21]/NET0131  & ~n65614 ;
  assign n65616 = ~\u0_R4_reg[21]/NET0131  & n65614 ;
  assign n65617 = ~n65615 & ~n65616 ;
  assign n65618 = decrypt_pad & ~\u0_uk_K_r4_reg[21]/NET0131  ;
  assign n65619 = ~decrypt_pad & ~\u0_uk_K_r4_reg[44]/NET0131  ;
  assign n65620 = ~n65618 & ~n65619 ;
  assign n65621 = \u0_R4_reg[16]/NET0131  & ~n65620 ;
  assign n65622 = ~\u0_R4_reg[16]/NET0131  & n65620 ;
  assign n65623 = ~n65621 & ~n65622 ;
  assign n65624 = ~n65617 & n65623 ;
  assign n65625 = decrypt_pad & ~\u0_uk_K_r4_reg[43]/NET0131  ;
  assign n65626 = ~decrypt_pad & ~\u0_uk_K_r4_reg[35]/NET0131  ;
  assign n65627 = ~n65625 & ~n65626 ;
  assign n65628 = \u0_R4_reg[17]/NET0131  & ~n65627 ;
  assign n65629 = ~\u0_R4_reg[17]/NET0131  & n65627 ;
  assign n65630 = ~n65628 & ~n65629 ;
  assign n65631 = decrypt_pad & ~\u0_uk_K_r4_reg[37]/NET0131  ;
  assign n65632 = ~decrypt_pad & ~\u0_uk_K_r4_reg[29]/NET0131  ;
  assign n65633 = ~n65631 & ~n65632 ;
  assign n65634 = \u0_R4_reg[18]/NET0131  & ~n65633 ;
  assign n65635 = ~\u0_R4_reg[18]/NET0131  & n65633 ;
  assign n65636 = ~n65634 & ~n65635 ;
  assign n65637 = ~n65630 & n65636 ;
  assign n65638 = n65624 & n65637 ;
  assign n65639 = decrypt_pad & ~\u0_uk_K_r4_reg[52]/NET0131  ;
  assign n65640 = ~decrypt_pad & ~\u0_uk_K_r4_reg[16]/NET0131  ;
  assign n65641 = ~n65639 & ~n65640 ;
  assign n65642 = \u0_R4_reg[19]/NET0131  & ~n65641 ;
  assign n65643 = ~\u0_R4_reg[19]/NET0131  & n65641 ;
  assign n65644 = ~n65642 & ~n65643 ;
  assign n65645 = ~n65638 & ~n65644 ;
  assign n65646 = n65617 & ~n65623 ;
  assign n65647 = ~n65630 & n65646 ;
  assign n65648 = n65636 & n65647 ;
  assign n65649 = n65644 & ~n65648 ;
  assign n65650 = ~n65617 & n65630 ;
  assign n65651 = n65636 & n65650 ;
  assign n65652 = n65630 & ~n65636 ;
  assign n65653 = ~n65623 & n65652 ;
  assign n65654 = n65617 & n65653 ;
  assign n65655 = ~n65651 & ~n65654 ;
  assign n65656 = n65649 & n65655 ;
  assign n65657 = ~n65645 & ~n65656 ;
  assign n65666 = ~n65623 & ~n65630 ;
  assign n65667 = ~n65617 & n65666 ;
  assign n65668 = ~n65636 & n65667 ;
  assign n65669 = n65617 & n65623 ;
  assign n65670 = ~n65630 & n65669 ;
  assign n65671 = ~n65668 & ~n65670 ;
  assign n65672 = n65644 & ~n65671 ;
  assign n65673 = ~n65623 & n65650 ;
  assign n65674 = ~n65647 & ~n65673 ;
  assign n65675 = n65636 & ~n65674 ;
  assign n65658 = decrypt_pad & ~\u0_uk_K_r4_reg[8]/NET0131  ;
  assign n65659 = ~decrypt_pad & ~\u0_uk_K_r4_reg[0]/P0001  ;
  assign n65660 = ~n65658 & ~n65659 ;
  assign n65661 = \u0_R4_reg[20]/NET0131  & ~n65660 ;
  assign n65662 = ~\u0_R4_reg[20]/NET0131  & n65660 ;
  assign n65663 = ~n65661 & ~n65662 ;
  assign n65664 = n65623 & ~n65636 ;
  assign n65665 = ~n65644 & n65664 ;
  assign n65676 = n65663 & ~n65665 ;
  assign n65677 = ~n65675 & n65676 ;
  assign n65678 = ~n65672 & n65677 ;
  assign n65684 = ~n65630 & ~n65636 ;
  assign n65685 = n65624 & n65684 ;
  assign n65683 = n65630 & n65669 ;
  assign n65686 = n65644 & ~n65683 ;
  assign n65687 = ~n65685 & n65686 ;
  assign n65688 = ~n65637 & n65646 ;
  assign n65689 = ~n65644 & ~n65670 ;
  assign n65690 = ~n65688 & n65689 ;
  assign n65691 = ~n65687 & ~n65690 ;
  assign n65679 = n65636 & n65667 ;
  assign n65680 = n65623 & n65650 ;
  assign n65681 = n65636 & n65680 ;
  assign n65682 = ~n65679 & ~n65681 ;
  assign n65692 = ~n65653 & ~n65663 ;
  assign n65693 = n65682 & n65692 ;
  assign n65694 = ~n65691 & n65693 ;
  assign n65695 = ~n65678 & ~n65694 ;
  assign n65696 = ~n65657 & ~n65695 ;
  assign n65697 = ~\u0_L4_reg[8]/NET0131  & ~n65696 ;
  assign n65698 = \u0_L4_reg[8]/NET0131  & n65696 ;
  assign n65699 = ~n65697 & ~n65698 ;
  assign n65715 = ~n65361 & ~n65366 ;
  assign n65716 = n65339 & ~n65715 ;
  assign n65717 = ~n65325 & ~n65716 ;
  assign n65718 = ~n65319 & n65365 ;
  assign n65719 = n65325 & ~n65400 ;
  assign n65720 = ~n65718 & n65719 ;
  assign n65721 = ~n65717 & ~n65720 ;
  assign n65722 = ~n65364 & ~n65388 ;
  assign n65723 = n65452 & ~n65722 ;
  assign n65724 = ~n65386 & ~n65723 ;
  assign n65725 = ~n65721 & n65724 ;
  assign n65726 = ~n65357 & ~n65725 ;
  assign n65709 = ~n65319 & n65369 ;
  assign n65710 = ~n65366 & ~n65709 ;
  assign n65711 = n65357 & ~n65710 ;
  assign n65712 = ~n65359 & ~n65460 ;
  assign n65713 = ~n65711 & n65712 ;
  assign n65714 = n65325 & ~n65713 ;
  assign n65700 = n65319 & n65365 ;
  assign n65701 = ~n65364 & n65452 ;
  assign n65702 = ~n65389 & ~n65701 ;
  assign n65703 = n65357 & ~n65702 ;
  assign n65704 = ~n65700 & ~n65703 ;
  assign n65705 = ~n65325 & ~n65704 ;
  assign n65706 = n65332 & n65360 ;
  assign n65707 = ~n65700 & ~n65706 ;
  assign n65708 = n65357 & ~n65707 ;
  assign n65727 = ~n65380 & ~n65708 ;
  assign n65728 = ~n65705 & n65727 ;
  assign n65729 = ~n65714 & n65728 ;
  assign n65730 = ~n65726 & n65729 ;
  assign n65731 = ~\u0_L4_reg[1]/NET0131  & ~n65730 ;
  assign n65732 = \u0_L4_reg[1]/NET0131  & n65730 ;
  assign n65733 = ~n65731 & ~n65732 ;
  assign n65744 = n65636 & n65669 ;
  assign n65734 = n65617 & ~n65636 ;
  assign n65751 = ~n65623 & n65734 ;
  assign n65752 = ~n65744 & ~n65751 ;
  assign n65753 = n65630 & ~n65752 ;
  assign n65754 = ~n65668 & ~n65753 ;
  assign n65755 = ~n65644 & ~n65754 ;
  assign n65761 = n65636 & ~n65644 ;
  assign n65762 = n65630 & n65761 ;
  assign n65763 = n65624 & ~n65684 ;
  assign n65764 = ~n65762 & n65763 ;
  assign n65756 = n65630 & ~n65644 ;
  assign n65757 = ~n65636 & n65669 ;
  assign n65758 = ~n65756 & n65757 ;
  assign n65759 = n65644 & n65646 ;
  assign n65760 = ~n65652 & n65759 ;
  assign n65765 = ~n65758 & ~n65760 ;
  assign n65766 = ~n65764 & n65765 ;
  assign n65767 = ~n65755 & n65766 ;
  assign n65768 = n65663 & ~n65767 ;
  assign n65735 = ~n65624 & ~n65734 ;
  assign n65736 = n65623 & ~n65630 ;
  assign n65737 = ~n65652 & ~n65736 ;
  assign n65738 = n65735 & ~n65737 ;
  assign n65739 = ~n65636 & n65683 ;
  assign n65740 = ~n65644 & ~n65647 ;
  assign n65741 = ~n65651 & ~n65685 ;
  assign n65742 = n65740 & n65741 ;
  assign n65743 = ~n65739 & n65742 ;
  assign n65745 = n65644 & ~n65653 ;
  assign n65746 = ~n65667 & ~n65744 ;
  assign n65747 = n65745 & n65746 ;
  assign n65748 = ~n65743 & ~n65747 ;
  assign n65749 = ~n65738 & ~n65748 ;
  assign n65750 = ~n65663 & ~n65749 ;
  assign n65769 = ~n65644 & ~n65675 ;
  assign n65770 = ~n65636 & n65680 ;
  assign n65771 = n65644 & ~n65679 ;
  assign n65772 = ~n65770 & n65771 ;
  assign n65773 = ~n65769 & ~n65772 ;
  assign n65774 = ~n65750 & ~n65773 ;
  assign n65775 = ~n65768 & n65774 ;
  assign n65776 = ~\u0_L4_reg[14]/NET0131  & ~n65775 ;
  assign n65777 = \u0_L4_reg[14]/NET0131  & n65775 ;
  assign n65778 = ~n65776 & ~n65777 ;
  assign n65780 = ~n64884 & ~n64900 ;
  assign n65781 = n64877 & ~n65780 ;
  assign n65783 = ~n64869 & n64896 ;
  assign n65779 = n64883 & n64897 ;
  assign n65782 = ~n64877 & n64905 ;
  assign n65784 = ~n65779 & ~n65782 ;
  assign n65785 = n65783 & n65784 ;
  assign n65786 = n65292 & n65785 ;
  assign n65787 = ~n65781 & n65786 ;
  assign n65790 = ~n64847 & ~n64868 ;
  assign n65791 = n64877 & ~n64900 ;
  assign n65792 = ~n65790 & n65791 ;
  assign n65788 = ~n64877 & ~n65165 ;
  assign n65789 = n64861 & n64867 ;
  assign n65793 = ~n64896 & ~n65789 ;
  assign n65794 = ~n65788 & n65793 ;
  assign n65795 = ~n65792 & n65794 ;
  assign n65796 = ~n65787 & ~n65795 ;
  assign n65797 = ~n64890 & ~n64925 ;
  assign n65798 = ~n65796 & n65797 ;
  assign n65799 = ~\u0_L4_reg[19]/NET0131  & ~n65798 ;
  assign n65800 = \u0_L4_reg[19]/NET0131  & n65798 ;
  assign n65801 = ~n65799 & ~n65800 ;
  assign n65803 = ~n65623 & n65636 ;
  assign n65804 = ~n65684 & ~n65803 ;
  assign n65805 = ~n65617 & ~n65804 ;
  assign n65806 = ~n65666 & ~n65683 ;
  assign n65807 = ~n65805 & n65806 ;
  assign n65808 = n65644 & ~n65807 ;
  assign n65809 = ~n65653 & ~n65670 ;
  assign n65810 = ~n65644 & ~n65809 ;
  assign n65802 = n65630 & n65734 ;
  assign n65811 = ~n65681 & ~n65802 ;
  assign n65812 = ~n65810 & n65811 ;
  assign n65813 = ~n65808 & n65812 ;
  assign n65814 = n65663 & ~n65813 ;
  assign n65826 = ~n65636 & n65647 ;
  assign n65827 = n65682 & ~n65826 ;
  assign n65828 = n65644 & ~n65827 ;
  assign n65816 = ~n65624 & ~n65630 ;
  assign n65815 = n65630 & ~n65803 ;
  assign n65817 = ~n65617 & n65644 ;
  assign n65818 = ~n65815 & ~n65817 ;
  assign n65819 = ~n65816 & n65818 ;
  assign n65821 = n65644 & ~n65650 ;
  assign n65820 = ~n65644 & ~n65666 ;
  assign n65822 = ~n65636 & ~n65820 ;
  assign n65823 = ~n65821 & n65822 ;
  assign n65824 = ~n65819 & ~n65823 ;
  assign n65825 = ~n65663 & ~n65824 ;
  assign n65829 = n65736 & n65761 ;
  assign n65830 = ~n65739 & ~n65829 ;
  assign n65831 = ~n65825 & n65830 ;
  assign n65832 = ~n65828 & n65831 ;
  assign n65833 = ~n65814 & n65832 ;
  assign n65834 = ~\u0_L4_reg[25]/NET0131  & ~n65833 ;
  assign n65835 = \u0_L4_reg[25]/NET0131  & n65833 ;
  assign n65836 = ~n65834 & ~n65835 ;
  assign n65838 = ~n65389 & ~n65468 ;
  assign n65839 = n65332 & ~n65838 ;
  assign n65845 = ~n65351 & ~n65839 ;
  assign n65840 = ~n65319 & n65465 ;
  assign n65841 = ~n65347 & ~n65840 ;
  assign n65842 = ~n65325 & ~n65369 ;
  assign n65843 = ~n65841 & n65842 ;
  assign n65844 = n65319 & ~n65401 ;
  assign n65846 = ~n65843 & ~n65844 ;
  assign n65847 = n65845 & n65846 ;
  assign n65848 = n65357 & ~n65847 ;
  assign n65856 = n65333 & ~n65388 ;
  assign n65857 = ~n65709 & ~n65856 ;
  assign n65858 = n65391 & n65857 ;
  assign n65859 = ~n65357 & ~n65858 ;
  assign n65849 = ~n65377 & ~n65706 ;
  assign n65850 = ~n65357 & ~n65849 ;
  assign n65851 = n65452 & n65722 ;
  assign n65852 = ~n65850 & ~n65851 ;
  assign n65853 = ~n65325 & ~n65852 ;
  assign n65837 = n65319 & n65469 ;
  assign n65854 = ~n65378 & ~n65392 ;
  assign n65855 = n65369 & ~n65854 ;
  assign n65860 = ~n65837 & ~n65855 ;
  assign n65861 = ~n65853 & n65860 ;
  assign n65862 = ~n65859 & n65861 ;
  assign n65863 = ~n65848 & n65862 ;
  assign n65864 = ~\u0_L4_reg[26]/NET0131  & ~n65863 ;
  assign n65865 = \u0_L4_reg[26]/NET0131  & n65863 ;
  assign n65866 = ~n65864 & ~n65865 ;
  assign n65871 = n65196 & ~n65272 ;
  assign n65869 = n65215 & n65545 ;
  assign n65870 = ~n65215 & n65225 ;
  assign n65872 = ~n65869 & ~n65870 ;
  assign n65873 = n65871 & n65872 ;
  assign n65874 = ~n65196 & ~n65241 ;
  assign n65875 = ~n65562 & n65874 ;
  assign n65876 = ~n65873 & ~n65875 ;
  assign n65877 = ~n65240 & ~n65549 ;
  assign n65878 = n65215 & ~n65568 ;
  assign n65879 = ~n65877 & n65878 ;
  assign n65880 = n65238 & ~n65553 ;
  assign n65881 = ~n65879 & n65880 ;
  assign n65882 = ~n65876 & n65881 ;
  assign n65883 = ~n65208 & ~n65269 ;
  assign n65884 = ~n65196 & n65202 ;
  assign n65885 = n65250 & n65884 ;
  assign n65893 = ~n65238 & ~n65885 ;
  assign n65894 = ~n65883 & n65893 ;
  assign n65886 = ~n65208 & n65545 ;
  assign n65887 = ~n65256 & ~n65886 ;
  assign n65888 = n65196 & ~n65887 ;
  assign n65889 = n65208 & n65224 ;
  assign n65890 = n65222 & ~n65549 ;
  assign n65891 = ~n65889 & ~n65890 ;
  assign n65892 = ~n65556 & ~n65891 ;
  assign n65895 = ~n65888 & ~n65892 ;
  assign n65896 = n65894 & n65895 ;
  assign n65897 = ~n65882 & ~n65896 ;
  assign n65867 = n65196 & n65229 ;
  assign n65868 = n65558 & n65560 ;
  assign n65898 = ~n65867 & ~n65868 ;
  assign n65899 = ~n65897 & n65898 ;
  assign n65900 = ~\u0_L4_reg[21]/NET0131  & ~n65899 ;
  assign n65901 = \u0_L4_reg[21]/NET0131  & n65899 ;
  assign n65902 = ~n65900 & ~n65901 ;
  assign n65915 = ~n65240 & ~n65546 ;
  assign n65916 = n65196 & ~n65915 ;
  assign n65917 = ~n65196 & ~n65229 ;
  assign n65918 = ~n65272 & ~n65886 ;
  assign n65919 = n65917 & n65918 ;
  assign n65920 = ~n65916 & ~n65919 ;
  assign n65921 = ~n65257 & ~n65870 ;
  assign n65922 = ~n65273 & n65921 ;
  assign n65923 = ~n65920 & n65922 ;
  assign n65924 = n65238 & ~n65923 ;
  assign n65903 = n65202 & ~n65215 ;
  assign n65904 = n65877 & ~n65903 ;
  assign n65905 = n65263 & ~n65904 ;
  assign n65906 = n65255 & n65560 ;
  assign n65907 = ~n65885 & ~n65906 ;
  assign n65908 = ~n65232 & n65907 ;
  assign n65909 = ~n65905 & n65908 ;
  assign n65910 = ~n65238 & ~n65909 ;
  assign n65911 = n65227 & ~n65242 ;
  assign n65912 = ~n65196 & ~n65911 ;
  assign n65913 = n65196 & ~n65208 ;
  assign n65914 = n65559 & n65913 ;
  assign n65925 = ~n65912 & ~n65914 ;
  assign n65926 = ~n65910 & n65925 ;
  assign n65927 = ~n65924 & n65926 ;
  assign n65928 = ~\u0_L4_reg[27]/NET0131  & ~n65927 ;
  assign n65929 = \u0_L4_reg[27]/NET0131  & n65927 ;
  assign n65930 = ~n65928 & ~n65929 ;
  assign n65931 = ~n64952 & n64976 ;
  assign n65932 = n64946 & n65931 ;
  assign n65933 = n64968 & ~n64998 ;
  assign n65935 = n64981 & n65500 ;
  assign n65934 = ~n64946 & ~n65500 ;
  assign n65936 = ~n64961 & n65499 ;
  assign n65937 = ~n65934 & ~n65936 ;
  assign n65938 = ~n65935 & n65937 ;
  assign n65939 = n65933 & ~n65938 ;
  assign n65943 = ~n64978 & n65934 ;
  assign n65940 = n64946 & n65936 ;
  assign n65941 = ~n65935 & ~n65940 ;
  assign n65942 = ~n64968 & n64998 ;
  assign n65944 = ~n65933 & ~n65942 ;
  assign n65945 = n65941 & n65944 ;
  assign n65946 = ~n65943 & n65945 ;
  assign n65947 = ~n65939 & ~n65946 ;
  assign n65948 = ~n65932 & ~n65947 ;
  assign n65949 = ~n64975 & ~n64999 ;
  assign n65950 = n64952 & ~n65949 ;
  assign n65951 = ~n64952 & ~n65494 ;
  assign n65952 = n65498 & n65951 ;
  assign n65953 = ~n65950 & ~n65952 ;
  assign n65954 = n65941 & n65942 ;
  assign n65955 = ~n65953 & n65954 ;
  assign n65956 = ~n65948 & ~n65955 ;
  assign n65957 = ~\u0_L4_reg[7]/NET0131  & n65956 ;
  assign n65958 = \u0_L4_reg[7]/NET0131  & ~n65956 ;
  assign n65959 = ~n65957 & ~n65958 ;
  assign n65961 = ~n65644 & ~n65668 ;
  assign n65960 = n65636 & n65670 ;
  assign n65962 = ~n65770 & ~n65960 ;
  assign n65963 = n65961 & n65962 ;
  assign n65964 = n65649 & ~n65685 ;
  assign n65965 = ~n65963 & ~n65964 ;
  assign n65969 = ~n65680 & ~n65751 ;
  assign n65970 = n65644 & ~n65969 ;
  assign n65966 = ~n65637 & n65644 ;
  assign n65967 = ~n65670 & ~n65735 ;
  assign n65968 = ~n65966 & ~n65967 ;
  assign n65971 = ~n65663 & ~n65968 ;
  assign n65972 = ~n65970 & n65971 ;
  assign n65973 = ~n65673 & ~n65757 ;
  assign n65974 = n65644 & ~n65973 ;
  assign n65975 = n65646 & n65756 ;
  assign n65976 = ~n65638 & n65663 ;
  assign n65977 = ~n65975 & n65976 ;
  assign n65978 = ~n65739 & n65977 ;
  assign n65979 = ~n65974 & n65978 ;
  assign n65980 = ~n65972 & ~n65979 ;
  assign n65981 = ~n65965 & ~n65980 ;
  assign n65982 = ~\u0_L4_reg[3]/NET0131  & ~n65981 ;
  assign n65983 = \u0_L4_reg[3]/NET0131  & n65981 ;
  assign n65984 = ~n65982 & ~n65983 ;
  assign n65991 = decrypt_pad & ~\u0_uk_K_r4_reg[17]/NET0131  ;
  assign n65992 = ~decrypt_pad & ~\u0_uk_K_r4_reg[11]/NET0131  ;
  assign n65993 = ~n65991 & ~n65992 ;
  assign n65994 = \u0_R4_reg[13]/NET0131  & ~n65993 ;
  assign n65995 = ~\u0_R4_reg[13]/NET0131  & n65993 ;
  assign n65996 = ~n65994 & ~n65995 ;
  assign n65998 = decrypt_pad & ~\u0_uk_K_r4_reg[12]/NET0131  ;
  assign n65999 = ~decrypt_pad & ~\u0_uk_K_r4_reg[6]/NET0131  ;
  assign n66000 = ~n65998 & ~n65999 ;
  assign n66001 = \u0_R4_reg[9]/NET0131  & ~n66000 ;
  assign n66002 = ~\u0_R4_reg[9]/NET0131  & n66000 ;
  assign n66003 = ~n66001 & ~n66002 ;
  assign n66020 = n65996 & ~n66003 ;
  assign n66021 = ~n65996 & n66003 ;
  assign n66022 = ~n66020 & ~n66021 ;
  assign n66012 = decrypt_pad & ~\u0_uk_K_r4_reg[46]/NET0131  ;
  assign n66013 = ~decrypt_pad & ~\u0_uk_K_r4_reg[40]/NET0131  ;
  assign n66014 = ~n66012 & ~n66013 ;
  assign n66015 = \u0_R4_reg[11]/NET0131  & ~n66014 ;
  assign n66016 = ~\u0_R4_reg[11]/NET0131  & n66014 ;
  assign n66017 = ~n66015 & ~n66016 ;
  assign n65985 = decrypt_pad & ~\u0_uk_K_r4_reg[40]/NET0131  ;
  assign n65986 = ~decrypt_pad & ~\u0_uk_K_r4_reg[34]/NET0131  ;
  assign n65987 = ~n65985 & ~n65986 ;
  assign n65988 = \u0_R4_reg[8]/NET0131  & ~n65987 ;
  assign n65989 = ~\u0_R4_reg[8]/NET0131  & n65987 ;
  assign n65990 = ~n65988 & ~n65989 ;
  assign n66004 = decrypt_pad & ~\u0_uk_K_r4_reg[20]/NET0131  ;
  assign n66005 = ~decrypt_pad & ~\u0_uk_K_r4_reg[39]/NET0131  ;
  assign n66006 = ~n66004 & ~n66005 ;
  assign n66007 = \u0_R4_reg[10]/NET0131  & ~n66006 ;
  assign n66008 = ~\u0_R4_reg[10]/NET0131  & n66006 ;
  assign n66009 = ~n66007 & ~n66008 ;
  assign n66018 = n66003 & ~n66009 ;
  assign n66019 = ~n65990 & ~n66018 ;
  assign n66023 = ~n66017 & ~n66019 ;
  assign n66024 = n66022 & n66023 ;
  assign n65997 = ~n65990 & ~n65996 ;
  assign n66010 = n66003 & n66009 ;
  assign n66011 = n65997 & n66010 ;
  assign n66025 = decrypt_pad & ~\u0_uk_K_r4_reg[4]/NET0131  ;
  assign n66026 = ~decrypt_pad & ~\u0_uk_K_r4_reg[55]/NET0131  ;
  assign n66027 = ~n66025 & ~n66026 ;
  assign n66028 = \u0_R4_reg[12]/NET0131  & ~n66027 ;
  assign n66029 = ~\u0_R4_reg[12]/NET0131  & n66027 ;
  assign n66030 = ~n66028 & ~n66029 ;
  assign n66031 = ~n66011 & n66030 ;
  assign n66032 = ~n66024 & n66031 ;
  assign n66036 = ~n66003 & ~n66009 ;
  assign n66037 = n65990 & n65996 ;
  assign n66038 = ~n65997 & ~n66037 ;
  assign n66039 = ~n66036 & ~n66038 ;
  assign n66040 = ~n66010 & n66039 ;
  assign n66033 = ~n65990 & n65996 ;
  assign n66034 = n66010 & ~n66017 ;
  assign n66035 = n66033 & n66034 ;
  assign n66041 = ~n65990 & n66017 ;
  assign n66042 = n66018 & n66041 ;
  assign n66047 = ~n66030 & ~n66042 ;
  assign n66048 = ~n66035 & n66047 ;
  assign n66043 = ~n65996 & n66010 ;
  assign n66044 = n65990 & n66043 ;
  assign n66045 = n66036 & ~n66041 ;
  assign n66046 = n66038 & n66045 ;
  assign n66049 = ~n66044 & ~n66046 ;
  assign n66050 = n66048 & n66049 ;
  assign n66051 = ~n66040 & n66050 ;
  assign n66052 = ~n66032 & ~n66051 ;
  assign n66054 = n66009 & n66033 ;
  assign n66055 = n65990 & ~n65996 ;
  assign n66056 = n66003 & n66055 ;
  assign n66057 = ~n66054 & ~n66056 ;
  assign n66058 = ~n66020 & n66057 ;
  assign n66059 = n66030 & ~n66058 ;
  assign n66053 = n66009 & n66020 ;
  assign n66060 = n65997 & n66036 ;
  assign n66061 = ~n66053 & ~n66060 ;
  assign n66062 = ~n66059 & n66061 ;
  assign n66063 = n66017 & ~n66062 ;
  assign n66064 = ~n66052 & ~n66063 ;
  assign n66065 = ~\u0_L4_reg[6]/NET0131  & ~n66064 ;
  assign n66066 = \u0_L4_reg[6]/NET0131  & n66064 ;
  assign n66067 = ~n66065 & ~n66066 ;
  assign n66069 = n64953 & ~n64975 ;
  assign n66070 = n64961 & n66069 ;
  assign n66072 = n64999 & n65500 ;
  assign n66071 = n64961 & n64982 ;
  assign n66073 = ~n64968 & ~n66071 ;
  assign n66074 = ~n65940 & n66073 ;
  assign n66075 = ~n66072 & n66074 ;
  assign n66077 = n64968 & ~n65931 ;
  assign n66076 = ~n64946 & n65494 ;
  assign n66078 = ~n66069 & ~n66076 ;
  assign n66079 = n66077 & n66078 ;
  assign n66080 = ~n66075 & ~n66079 ;
  assign n66081 = ~n66070 & ~n66080 ;
  assign n66082 = n64998 & ~n66081 ;
  assign n66083 = n64952 & n64988 ;
  assign n66085 = ~n65936 & ~n66083 ;
  assign n66086 = n64968 & ~n66085 ;
  assign n66084 = n65496 & ~n66083 ;
  assign n66087 = ~n64991 & n65004 ;
  assign n66088 = n64984 & ~n66087 ;
  assign n66089 = ~n66084 & n66088 ;
  assign n66090 = ~n66086 & n66089 ;
  assign n66091 = ~n64998 & ~n66090 ;
  assign n66068 = n64946 & n65493 ;
  assign n66092 = ~n64952 & n64961 ;
  assign n66093 = ~n66076 & ~n66092 ;
  assign n66094 = ~n64954 & ~n64968 ;
  assign n66095 = ~n66093 & n66094 ;
  assign n66096 = ~n66068 & ~n66095 ;
  assign n66097 = ~n66091 & n66096 ;
  assign n66098 = ~n66082 & n66097 ;
  assign n66099 = \u0_L4_reg[32]/NET0131  & n66098 ;
  assign n66100 = ~\u0_L4_reg[32]/NET0131  & ~n66098 ;
  assign n66101 = ~n66099 & ~n66100 ;
  assign n66102 = ~n65031 & n65050 ;
  assign n66103 = ~n64755 & n66102 ;
  assign n66109 = ~n64806 & ~n66103 ;
  assign n66104 = ~n64761 & n65031 ;
  assign n66105 = ~n64796 & ~n66104 ;
  assign n66106 = n64809 & ~n66105 ;
  assign n66107 = n64755 & ~n65050 ;
  assign n66108 = ~n66104 & n66107 ;
  assign n66110 = ~n66106 & ~n66108 ;
  assign n66111 = n66109 & n66110 ;
  assign n66113 = ~n65051 & ~n65514 ;
  assign n66114 = n64761 & ~n66113 ;
  assign n66112 = n64762 & n66102 ;
  assign n66115 = n65033 & ~n66112 ;
  assign n66116 = ~n66114 & n66115 ;
  assign n66117 = ~n66111 & ~n66116 ;
  assign n66118 = ~n64813 & ~n65057 ;
  assign n66119 = n65521 & n66118 ;
  assign n66120 = ~n66117 & ~n66119 ;
  assign n66121 = ~\u0_L4_reg[9]/NET0131  & ~n66120 ;
  assign n66122 = \u0_L4_reg[9]/NET0131  & n66120 ;
  assign n66123 = ~n66121 & ~n66122 ;
  assign n66126 = n65990 & n66009 ;
  assign n66127 = ~n66021 & ~n66126 ;
  assign n66131 = n66017 & ~n66043 ;
  assign n66132 = ~n66127 & n66131 ;
  assign n66128 = ~n65990 & ~n66003 ;
  assign n66129 = ~n66017 & ~n66128 ;
  assign n66130 = n66127 & n66129 ;
  assign n66124 = n66036 & ~n66038 ;
  assign n66125 = ~n66003 & n66054 ;
  assign n66133 = ~n66124 & ~n66125 ;
  assign n66134 = ~n66130 & n66133 ;
  assign n66135 = ~n66132 & n66134 ;
  assign n66136 = ~n66030 & ~n66135 ;
  assign n66137 = n65997 & n66009 ;
  assign n66138 = ~n66009 & n66033 ;
  assign n66139 = ~n66137 & ~n66138 ;
  assign n66140 = n66036 & n66055 ;
  assign n66141 = n66017 & ~n66140 ;
  assign n66142 = n66139 & n66141 ;
  assign n66143 = n65997 & n66003 ;
  assign n66144 = ~n66017 & ~n66126 ;
  assign n66145 = ~n66143 & n66144 ;
  assign n66146 = n66030 & ~n66145 ;
  assign n66147 = ~n66142 & n66146 ;
  assign n66148 = ~n66003 & n66126 ;
  assign n66149 = n65996 & n66017 ;
  assign n66150 = n66148 & n66149 ;
  assign n66151 = ~n65996 & ~n66017 ;
  assign n66152 = ~n66030 & ~n66151 ;
  assign n66153 = n66010 & ~n66037 ;
  assign n66154 = ~n66152 & n66153 ;
  assign n66155 = ~n66150 & ~n66154 ;
  assign n66156 = ~n66147 & n66155 ;
  assign n66157 = ~n66136 & n66156 ;
  assign n66158 = \u0_L4_reg[30]/NET0131  & ~n66157 ;
  assign n66159 = ~\u0_L4_reg[30]/NET0131  & n66157 ;
  assign n66160 = ~n66158 & ~n66159 ;
  assign n66162 = n66003 & n66037 ;
  assign n66163 = ~n66003 & ~n66037 ;
  assign n66164 = ~n66162 & ~n66163 ;
  assign n66165 = ~n65997 & ~n66164 ;
  assign n66166 = n66017 & n66143 ;
  assign n66167 = ~n66165 & ~n66166 ;
  assign n66168 = ~n66009 & ~n66167 ;
  assign n66161 = n66010 & n66033 ;
  assign n66169 = ~n66009 & n66055 ;
  assign n66170 = ~n66137 & ~n66169 ;
  assign n66171 = ~n66017 & ~n66170 ;
  assign n66172 = ~n66161 & ~n66171 ;
  assign n66173 = ~n66168 & n66172 ;
  assign n66174 = n66030 & ~n66173 ;
  assign n66176 = n65996 & n66128 ;
  assign n66175 = n65997 & ~n66009 ;
  assign n66177 = ~n66162 & ~n66175 ;
  assign n66178 = ~n66176 & n66177 ;
  assign n66179 = ~n66017 & ~n66178 ;
  assign n66180 = ~n65997 & n66017 ;
  assign n66181 = n66164 & n66180 ;
  assign n66182 = ~n66060 & ~n66181 ;
  assign n66183 = ~n66179 & n66182 ;
  assign n66184 = ~n66030 & ~n66183 ;
  assign n66185 = ~n66003 & n66137 ;
  assign n66186 = ~n66044 & ~n66185 ;
  assign n66187 = n66017 & ~n66186 ;
  assign n66188 = ~n66017 & n66148 ;
  assign n66189 = ~n66187 & ~n66188 ;
  assign n66190 = ~n66184 & n66189 ;
  assign n66191 = ~n66174 & n66190 ;
  assign n66192 = ~\u0_L4_reg[16]/NET0131  & ~n66191 ;
  assign n66193 = \u0_L4_reg[16]/NET0131  & n66191 ;
  assign n66194 = ~n66192 & ~n66193 ;
  assign n66195 = ~n65077 & n65120 ;
  assign n66196 = ~n65435 & ~n66195 ;
  assign n66197 = ~n65083 & ~n66196 ;
  assign n66199 = ~n65104 & ~n65436 ;
  assign n66198 = n65077 & n65598 ;
  assign n66200 = n65584 & ~n66198 ;
  assign n66201 = n66199 & n66200 ;
  assign n66202 = ~n66197 & n66201 ;
  assign n66204 = n65083 & n65118 ;
  assign n66205 = ~n65134 & ~n66204 ;
  assign n66206 = ~n65077 & ~n66205 ;
  assign n66203 = n65077 & ~n65115 ;
  assign n66207 = n65071 & ~n65129 ;
  assign n66208 = ~n66203 & n66207 ;
  assign n66209 = ~n66206 & n66208 ;
  assign n66210 = ~n66202 & ~n66209 ;
  assign n66211 = n65090 & n65103 ;
  assign n66212 = ~n65442 & ~n66211 ;
  assign n66213 = n65077 & ~n66212 ;
  assign n66214 = ~n65077 & n65585 ;
  assign n66215 = ~n66213 & ~n66214 ;
  assign n66216 = ~n66210 & n66215 ;
  assign n66217 = \u0_L4_reg[18]/NET0131  & n66216 ;
  assign n66218 = ~\u0_L4_reg[18]/NET0131  & ~n66216 ;
  assign n66219 = ~n66217 & ~n66218 ;
  assign n66232 = ~n65996 & n66148 ;
  assign n66233 = ~n66143 & ~n66148 ;
  assign n66234 = n66139 & n66233 ;
  assign n66235 = n66017 & ~n66234 ;
  assign n66236 = ~n66232 & ~n66235 ;
  assign n66237 = ~n66030 & ~n66236 ;
  assign n66227 = ~n66017 & n66039 ;
  assign n66221 = n66003 & n66126 ;
  assign n66222 = ~n66054 & ~n66221 ;
  assign n66223 = n66017 & ~n66222 ;
  assign n66224 = ~n66009 & n66017 ;
  assign n66225 = ~n66003 & ~n66033 ;
  assign n66226 = n66224 & n66225 ;
  assign n66228 = ~n66046 & ~n66226 ;
  assign n66229 = ~n66223 & n66228 ;
  assign n66230 = ~n66227 & n66229 ;
  assign n66231 = n66030 & ~n66230 ;
  assign n66238 = n66057 & ~n66124 ;
  assign n66239 = ~n66017 & ~n66030 ;
  assign n66240 = ~n66238 & n66239 ;
  assign n66220 = n66034 & n66037 ;
  assign n66241 = n66022 & n66224 ;
  assign n66242 = n66038 & n66241 ;
  assign n66243 = ~n66220 & ~n66242 ;
  assign n66244 = ~n66240 & n66243 ;
  assign n66245 = ~n66231 & n66244 ;
  assign n66246 = ~n66237 & n66245 ;
  assign n66247 = ~\u0_L4_reg[24]/NET0131  & ~n66246 ;
  assign n66248 = \u0_L4_reg[24]/NET0131  & n66246 ;
  assign n66249 = ~n66247 & ~n66248 ;
  assign n66250 = decrypt_pad & ~\u0_uk_K_r3_reg[45]/P0001  ;
  assign n66251 = ~decrypt_pad & ~\u0_uk_K_r3_reg[36]/NET0131  ;
  assign n66252 = ~n66250 & ~n66251 ;
  assign n66253 = \u0_R3_reg[28]/NET0131  & ~n66252 ;
  assign n66254 = ~\u0_R3_reg[28]/NET0131  & n66252 ;
  assign n66255 = ~n66253 & ~n66254 ;
  assign n66283 = decrypt_pad & ~\u0_uk_K_r3_reg[30]/NET0131  ;
  assign n66284 = ~decrypt_pad & ~\u0_uk_K_r3_reg[49]/NET0131  ;
  assign n66285 = ~n66283 & ~n66284 ;
  assign n66286 = \u0_R3_reg[27]/NET0131  & ~n66285 ;
  assign n66287 = ~\u0_R3_reg[27]/NET0131  & n66285 ;
  assign n66288 = ~n66286 & ~n66287 ;
  assign n66269 = decrypt_pad & ~\u0_uk_K_r3_reg[21]/NET0131  ;
  assign n66270 = ~decrypt_pad & ~\u0_uk_K_r3_reg[16]/NET0131  ;
  assign n66271 = ~n66269 & ~n66270 ;
  assign n66272 = \u0_R3_reg[26]/NET0131  & ~n66271 ;
  assign n66273 = ~\u0_R3_reg[26]/NET0131  & n66271 ;
  assign n66274 = ~n66272 & ~n66273 ;
  assign n66256 = decrypt_pad & ~\u0_uk_K_r3_reg[1]/NET0131  ;
  assign n66257 = ~decrypt_pad & ~\u0_uk_K_r3_reg[51]/NET0131  ;
  assign n66258 = ~n66256 & ~n66257 ;
  assign n66259 = \u0_R3_reg[24]/NET0131  & ~n66258 ;
  assign n66260 = ~\u0_R3_reg[24]/NET0131  & n66258 ;
  assign n66261 = ~n66259 & ~n66260 ;
  assign n66275 = decrypt_pad & ~\u0_uk_K_r3_reg[9]/NET0131  ;
  assign n66276 = ~decrypt_pad & ~\u0_uk_K_r3_reg[28]/NET0131  ;
  assign n66277 = ~n66275 & ~n66276 ;
  assign n66278 = \u0_R3_reg[29]/NET0131  & ~n66277 ;
  assign n66279 = ~\u0_R3_reg[29]/NET0131  & n66277 ;
  assign n66280 = ~n66278 & ~n66279 ;
  assign n66289 = n66261 & ~n66280 ;
  assign n66290 = ~n66261 & n66280 ;
  assign n66291 = ~n66289 & ~n66290 ;
  assign n66262 = decrypt_pad & ~\u0_uk_K_r3_reg[36]/NET0131  ;
  assign n66263 = ~decrypt_pad & ~\u0_uk_K_r3_reg[0]/NET0131  ;
  assign n66264 = ~n66262 & ~n66263 ;
  assign n66265 = \u0_R3_reg[25]/NET0131  & ~n66264 ;
  assign n66266 = ~\u0_R3_reg[25]/NET0131  & n66264 ;
  assign n66267 = ~n66265 & ~n66266 ;
  assign n66292 = ~n66261 & n66267 ;
  assign n66293 = n66291 & ~n66292 ;
  assign n66294 = n66274 & n66293 ;
  assign n66295 = n66267 & n66289 ;
  assign n66296 = ~n66294 & ~n66295 ;
  assign n66297 = ~n66288 & ~n66296 ;
  assign n66298 = ~n66267 & n66288 ;
  assign n66299 = n66290 & ~n66298 ;
  assign n66300 = ~n66267 & n66289 ;
  assign n66301 = ~n66299 & ~n66300 ;
  assign n66302 = ~n66274 & ~n66301 ;
  assign n66268 = n66261 & n66267 ;
  assign n66281 = n66274 & n66280 ;
  assign n66282 = n66268 & n66281 ;
  assign n66303 = n66261 & n66288 ;
  assign n66304 = ~n66267 & ~n66274 ;
  assign n66305 = n66303 & n66304 ;
  assign n66306 = ~n66282 & ~n66305 ;
  assign n66307 = ~n66302 & n66306 ;
  assign n66308 = ~n66297 & n66307 ;
  assign n66309 = ~n66255 & ~n66308 ;
  assign n66321 = n66267 & n66274 ;
  assign n66322 = ~n66304 & ~n66321 ;
  assign n66310 = ~n66274 & ~n66280 ;
  assign n66323 = n66303 & ~n66310 ;
  assign n66324 = n66322 & n66323 ;
  assign n66312 = ~n66261 & ~n66267 ;
  assign n66313 = ~n66281 & ~n66310 ;
  assign n66314 = n66312 & ~n66313 ;
  assign n66315 = n66261 & ~n66267 ;
  assign n66316 = ~n66292 & ~n66315 ;
  assign n66317 = n66261 & n66274 ;
  assign n66318 = n66280 & ~n66288 ;
  assign n66319 = ~n66317 & n66318 ;
  assign n66320 = ~n66316 & n66319 ;
  assign n66325 = ~n66314 & ~n66320 ;
  assign n66326 = ~n66324 & n66325 ;
  assign n66327 = n66255 & ~n66326 ;
  assign n66328 = n66281 & n66312 ;
  assign n66329 = n66274 & ~n66280 ;
  assign n66330 = n66292 & n66329 ;
  assign n66331 = ~n66328 & ~n66330 ;
  assign n66332 = ~n66300 & n66331 ;
  assign n66333 = n66288 & ~n66332 ;
  assign n66311 = n66298 & n66310 ;
  assign n66334 = ~n66261 & ~n66274 ;
  assign n66335 = ~n66317 & ~n66334 ;
  assign n66336 = n66267 & ~n66288 ;
  assign n66337 = ~n66335 & n66336 ;
  assign n66338 = ~n66311 & ~n66337 ;
  assign n66339 = ~n66333 & n66338 ;
  assign n66340 = ~n66327 & n66339 ;
  assign n66341 = ~n66309 & n66340 ;
  assign n66342 = ~\u0_L3_reg[22]/NET0131  & ~n66341 ;
  assign n66343 = \u0_L3_reg[22]/NET0131  & n66341 ;
  assign n66344 = ~n66342 & ~n66343 ;
  assign n66395 = decrypt_pad & ~\u0_uk_K_r3_reg[39]/NET0131  ;
  assign n66396 = ~decrypt_pad & ~\u0_uk_K_r3_reg[5]/NET0131  ;
  assign n66397 = ~n66395 & ~n66396 ;
  assign n66398 = \u0_R3_reg[4]/NET0131  & ~n66397 ;
  assign n66399 = ~\u0_R3_reg[4]/NET0131  & n66397 ;
  assign n66400 = ~n66398 & ~n66399 ;
  assign n66372 = decrypt_pad & ~\u0_uk_K_r3_reg[4]/NET0131  ;
  assign n66373 = ~decrypt_pad & ~\u0_uk_K_r3_reg[27]/NET0131  ;
  assign n66374 = ~n66372 & ~n66373 ;
  assign n66375 = \u0_R3_reg[3]/NET0131  & ~n66374 ;
  assign n66376 = ~\u0_R3_reg[3]/NET0131  & n66374 ;
  assign n66377 = ~n66375 & ~n66376 ;
  assign n66345 = decrypt_pad & ~\u0_uk_K_r3_reg[48]/NET0131  ;
  assign n66346 = ~decrypt_pad & ~\u0_uk_K_r3_reg[39]/NET0131  ;
  assign n66347 = ~n66345 & ~n66346 ;
  assign n66348 = \u0_R3_reg[32]/NET0131  & ~n66347 ;
  assign n66349 = ~\u0_R3_reg[32]/NET0131  & n66347 ;
  assign n66350 = ~n66348 & ~n66349 ;
  assign n66358 = decrypt_pad & ~\u0_uk_K_r3_reg[12]/NET0131  ;
  assign n66359 = ~decrypt_pad & ~\u0_uk_K_r3_reg[3]/NET0131  ;
  assign n66360 = ~n66358 & ~n66359 ;
  assign n66361 = \u0_R3_reg[1]/NET0131  & ~n66360 ;
  assign n66362 = ~\u0_R3_reg[1]/NET0131  & n66360 ;
  assign n66363 = ~n66361 & ~n66362 ;
  assign n66351 = decrypt_pad & ~\u0_uk_K_r3_reg[10]/NET0131  ;
  assign n66352 = ~decrypt_pad & ~\u0_uk_K_r3_reg[33]/NET0131  ;
  assign n66353 = ~n66351 & ~n66352 ;
  assign n66354 = \u0_R3_reg[5]/NET0131  & ~n66353 ;
  assign n66355 = ~\u0_R3_reg[5]/NET0131  & n66353 ;
  assign n66356 = ~n66354 & ~n66355 ;
  assign n66364 = decrypt_pad & ~\u0_uk_K_r3_reg[27]/NET0131  ;
  assign n66365 = ~decrypt_pad & ~\u0_uk_K_r3_reg[18]/NET0131  ;
  assign n66366 = ~n66364 & ~n66365 ;
  assign n66367 = \u0_R3_reg[2]/NET0131  & ~n66366 ;
  assign n66368 = ~\u0_R3_reg[2]/NET0131  & n66366 ;
  assign n66369 = ~n66367 & ~n66368 ;
  assign n66405 = n66356 & n66369 ;
  assign n66406 = n66363 & n66405 ;
  assign n66407 = ~n66350 & n66406 ;
  assign n66384 = ~n66356 & n66369 ;
  assign n66408 = n66350 & n66363 ;
  assign n66409 = n66384 & n66408 ;
  assign n66410 = ~n66407 & ~n66409 ;
  assign n66411 = n66377 & ~n66410 ;
  assign n66402 = ~n66356 & n66363 ;
  assign n66403 = ~n66369 & n66402 ;
  assign n66404 = ~n66350 & n66403 ;
  assign n66412 = n66350 & n66356 ;
  assign n66370 = ~n66363 & ~n66369 ;
  assign n66378 = ~n66369 & n66377 ;
  assign n66413 = ~n66370 & ~n66378 ;
  assign n66414 = n66412 & ~n66413 ;
  assign n66415 = ~n66404 & ~n66414 ;
  assign n66416 = ~n66411 & n66415 ;
  assign n66417 = ~n66400 & ~n66416 ;
  assign n66357 = ~n66350 & ~n66356 ;
  assign n66371 = ~n66356 & n66370 ;
  assign n66379 = n66363 & ~n66378 ;
  assign n66380 = ~n66350 & ~n66379 ;
  assign n66381 = ~n66371 & ~n66380 ;
  assign n66382 = ~n66357 & ~n66381 ;
  assign n66383 = n66356 & ~n66363 ;
  assign n66385 = ~n66350 & n66384 ;
  assign n66386 = ~n66383 & ~n66385 ;
  assign n66387 = n66377 & ~n66386 ;
  assign n66388 = n66350 & ~n66363 ;
  assign n66389 = ~n66363 & n66369 ;
  assign n66390 = n66350 & ~n66377 ;
  assign n66391 = ~n66389 & ~n66390 ;
  assign n66392 = ~n66388 & ~n66391 ;
  assign n66393 = ~n66387 & ~n66392 ;
  assign n66394 = ~n66382 & n66393 ;
  assign n66401 = ~n66394 & n66400 ;
  assign n66425 = n66350 & n66406 ;
  assign n66426 = ~n66350 & n66356 ;
  assign n66427 = n66389 & n66426 ;
  assign n66428 = ~n66403 & ~n66427 ;
  assign n66429 = ~n66425 & n66428 ;
  assign n66430 = ~n66377 & ~n66429 ;
  assign n66421 = n66369 & ~n66388 ;
  assign n66419 = n66350 & ~n66369 ;
  assign n66420 = ~n66377 & ~n66419 ;
  assign n66422 = ~n66383 & ~n66400 ;
  assign n66423 = n66420 & n66422 ;
  assign n66424 = ~n66421 & n66423 ;
  assign n66418 = n66378 & n66388 ;
  assign n66431 = ~n66350 & n66377 ;
  assign n66432 = ~n66356 & n66389 ;
  assign n66433 = n66431 & n66432 ;
  assign n66434 = ~n66418 & ~n66433 ;
  assign n66435 = ~n66424 & n66434 ;
  assign n66436 = ~n66430 & n66435 ;
  assign n66437 = ~n66401 & n66436 ;
  assign n66438 = ~n66417 & n66437 ;
  assign n66439 = ~\u0_L3_reg[31]/NET0131  & ~n66438 ;
  assign n66440 = \u0_L3_reg[31]/NET0131  & n66438 ;
  assign n66441 = ~n66439 & ~n66440 ;
  assign n66442 = decrypt_pad & ~\u0_uk_K_r3_reg[33]/NET0131  ;
  assign n66443 = ~decrypt_pad & ~\u0_uk_K_r3_reg[24]/NET0131  ;
  assign n66444 = ~n66442 & ~n66443 ;
  assign n66445 = \u0_R3_reg[15]/NET0131  & ~n66444 ;
  assign n66446 = ~\u0_R3_reg[15]/NET0131  & n66444 ;
  assign n66447 = ~n66445 & ~n66446 ;
  assign n66448 = decrypt_pad & ~\u0_uk_K_r3_reg[24]/NET0131  ;
  assign n66449 = ~decrypt_pad & ~\u0_uk_K_r3_reg[47]/NET0131  ;
  assign n66450 = ~n66448 & ~n66449 ;
  assign n66451 = \u0_R3_reg[13]/NET0131  & ~n66450 ;
  assign n66452 = ~\u0_R3_reg[13]/NET0131  & n66450 ;
  assign n66453 = ~n66451 & ~n66452 ;
  assign n66454 = decrypt_pad & ~\u0_uk_K_r3_reg[5]/NET0131  ;
  assign n66455 = ~decrypt_pad & ~\u0_uk_K_r3_reg[53]/NET0131  ;
  assign n66456 = ~n66454 & ~n66455 ;
  assign n66457 = \u0_R3_reg[12]/NET0131  & ~n66456 ;
  assign n66458 = ~\u0_R3_reg[12]/NET0131  & n66456 ;
  assign n66459 = ~n66457 & ~n66458 ;
  assign n66460 = n66453 & ~n66459 ;
  assign n66461 = decrypt_pad & ~\u0_uk_K_r3_reg[25]/NET0131  ;
  assign n66462 = ~decrypt_pad & ~\u0_uk_K_r3_reg[48]/NET0131  ;
  assign n66463 = ~n66461 & ~n66462 ;
  assign n66464 = \u0_R3_reg[14]/NET0131  & ~n66463 ;
  assign n66465 = ~\u0_R3_reg[14]/NET0131  & n66463 ;
  assign n66466 = ~n66464 & ~n66465 ;
  assign n66467 = decrypt_pad & ~\u0_uk_K_r3_reg[46]/NET0131  ;
  assign n66468 = ~decrypt_pad & ~\u0_uk_K_r3_reg[12]/NET0131  ;
  assign n66469 = ~n66467 & ~n66468 ;
  assign n66470 = \u0_R3_reg[17]/NET0131  & ~n66469 ;
  assign n66471 = ~\u0_R3_reg[17]/NET0131  & n66469 ;
  assign n66472 = ~n66470 & ~n66471 ;
  assign n66473 = ~n66466 & n66472 ;
  assign n66474 = n66460 & n66473 ;
  assign n66475 = ~n66447 & ~n66474 ;
  assign n66482 = ~n66453 & ~n66472 ;
  assign n66483 = ~n66459 & n66482 ;
  assign n66484 = ~n66466 & n66483 ;
  assign n66476 = n66459 & ~n66472 ;
  assign n66477 = ~n66453 & n66466 ;
  assign n66478 = n66476 & n66477 ;
  assign n66479 = n66447 & ~n66478 ;
  assign n66480 = n66453 & ~n66466 ;
  assign n66481 = n66476 & n66480 ;
  assign n66485 = n66479 & ~n66481 ;
  assign n66486 = ~n66484 & n66485 ;
  assign n66487 = ~n66475 & ~n66486 ;
  assign n66488 = ~n66459 & n66472 ;
  assign n66489 = n66447 & n66488 ;
  assign n66490 = ~n66453 & n66489 ;
  assign n66491 = decrypt_pad & ~\u0_uk_K_r3_reg[41]/NET0131  ;
  assign n66492 = ~decrypt_pad & ~\u0_uk_K_r3_reg[32]/NET0131  ;
  assign n66493 = ~n66491 & ~n66492 ;
  assign n66494 = \u0_R3_reg[16]/NET0131  & ~n66493 ;
  assign n66495 = ~\u0_R3_reg[16]/NET0131  & n66493 ;
  assign n66496 = ~n66494 & ~n66495 ;
  assign n66509 = ~n66490 & n66496 ;
  assign n66497 = n66453 & n66476 ;
  assign n66498 = n66447 & n66497 ;
  assign n66505 = ~n66447 & ~n66466 ;
  assign n66506 = ~n66453 & n66459 ;
  assign n66507 = ~n66460 & ~n66506 ;
  assign n66508 = n66505 & ~n66507 ;
  assign n66510 = ~n66498 & ~n66508 ;
  assign n66511 = n66509 & n66510 ;
  assign n66499 = n66459 & n66472 ;
  assign n66500 = n66453 & n66499 ;
  assign n66501 = n66466 & n66500 ;
  assign n66502 = ~n66474 & ~n66501 ;
  assign n66503 = ~n66447 & n66483 ;
  assign n66504 = n66466 & n66503 ;
  assign n66512 = n66502 & ~n66504 ;
  assign n66513 = n66511 & n66512 ;
  assign n66520 = n66447 & ~n66483 ;
  assign n66521 = ~n66500 & n66520 ;
  assign n66522 = n66466 & n66476 ;
  assign n66517 = ~n66453 & n66472 ;
  assign n66523 = ~n66447 & ~n66517 ;
  assign n66524 = ~n66522 & n66523 ;
  assign n66525 = ~n66521 & ~n66524 ;
  assign n66514 = n66460 & ~n66472 ;
  assign n66515 = n66466 & n66514 ;
  assign n66516 = ~n66484 & ~n66515 ;
  assign n66526 = n66447 & n66466 ;
  assign n66527 = n66460 & n66526 ;
  assign n66518 = n66459 & ~n66466 ;
  assign n66519 = n66517 & n66518 ;
  assign n66528 = ~n66496 & ~n66519 ;
  assign n66529 = ~n66527 & n66528 ;
  assign n66530 = n66516 & n66529 ;
  assign n66531 = ~n66525 & n66530 ;
  assign n66532 = ~n66513 & ~n66531 ;
  assign n66533 = ~n66487 & ~n66532 ;
  assign n66534 = ~\u0_L3_reg[20]/NET0131  & ~n66533 ;
  assign n66535 = \u0_L3_reg[20]/NET0131  & n66533 ;
  assign n66536 = ~n66534 & ~n66535 ;
  assign n66586 = decrypt_pad & ~\u0_uk_K_r3_reg[37]/NET0131  ;
  assign n66587 = ~decrypt_pad & ~\u0_uk_K_r3_reg[1]/NET0131  ;
  assign n66588 = ~n66586 & ~n66587 ;
  assign n66589 = \u0_R3_reg[32]/NET0131  & ~n66588 ;
  assign n66590 = ~\u0_R3_reg[32]/NET0131  & n66588 ;
  assign n66591 = ~n66589 & ~n66590 ;
  assign n66537 = decrypt_pad & ~\u0_uk_K_r3_reg[15]/NET0131  ;
  assign n66538 = ~decrypt_pad & ~\u0_uk_K_r3_reg[38]/NET0131  ;
  assign n66539 = ~n66537 & ~n66538 ;
  assign n66540 = \u0_R3_reg[28]/NET0131  & ~n66539 ;
  assign n66541 = ~\u0_R3_reg[28]/NET0131  & n66539 ;
  assign n66542 = ~n66540 & ~n66541 ;
  assign n66567 = decrypt_pad & ~\u0_uk_K_r3_reg[31]/NET0131  ;
  assign n66568 = ~decrypt_pad & ~\u0_uk_K_r3_reg[22]/NET0131  ;
  assign n66569 = ~n66567 & ~n66568 ;
  assign n66570 = \u0_R3_reg[1]/NET0131  & ~n66569 ;
  assign n66571 = ~\u0_R3_reg[1]/NET0131  & n66569 ;
  assign n66572 = ~n66570 & ~n66571 ;
  assign n66543 = decrypt_pad & ~\u0_uk_K_r3_reg[43]/NET0131  ;
  assign n66544 = ~decrypt_pad & ~\u0_uk_K_r3_reg[7]/NET0131  ;
  assign n66545 = ~n66543 & ~n66544 ;
  assign n66546 = \u0_R3_reg[30]/NET0131  & ~n66545 ;
  assign n66547 = ~\u0_R3_reg[30]/NET0131  & n66545 ;
  assign n66548 = ~n66546 & ~n66547 ;
  assign n66550 = decrypt_pad & ~\u0_uk_K_r3_reg[42]/NET0131  ;
  assign n66551 = ~decrypt_pad & ~\u0_uk_K_r3_reg[37]/NET0131  ;
  assign n66552 = ~n66550 & ~n66551 ;
  assign n66553 = \u0_R3_reg[29]/NET0131  & ~n66552 ;
  assign n66554 = ~\u0_R3_reg[29]/NET0131  & n66552 ;
  assign n66555 = ~n66553 & ~n66554 ;
  assign n66593 = ~n66548 & n66555 ;
  assign n66594 = ~n66572 & n66593 ;
  assign n66577 = n66555 & n66572 ;
  assign n66578 = n66548 & n66577 ;
  assign n66560 = decrypt_pad & ~\u0_uk_K_r3_reg[0]/NET0131  ;
  assign n66561 = ~decrypt_pad & ~\u0_uk_K_r3_reg[50]/NET0131  ;
  assign n66562 = ~n66560 & ~n66561 ;
  assign n66563 = \u0_R3_reg[31]/P0001  & ~n66562 ;
  assign n66564 = ~\u0_R3_reg[31]/P0001  & n66562 ;
  assign n66565 = ~n66563 & ~n66564 ;
  assign n66595 = ~n66548 & ~n66565 ;
  assign n66596 = ~n66578 & ~n66595 ;
  assign n66597 = ~n66594 & n66596 ;
  assign n66598 = n66542 & ~n66597 ;
  assign n66557 = n66542 & ~n66555 ;
  assign n66558 = n66548 & n66557 ;
  assign n66601 = n66558 & ~n66572 ;
  assign n66599 = ~n66555 & n66572 ;
  assign n66600 = ~n66542 & n66599 ;
  assign n66602 = n66565 & ~n66600 ;
  assign n66603 = ~n66601 & n66602 ;
  assign n66604 = ~n66542 & ~n66572 ;
  assign n66605 = n66548 & n66604 ;
  assign n66606 = ~n66565 & ~n66577 ;
  assign n66607 = ~n66605 & n66606 ;
  assign n66608 = ~n66603 & ~n66607 ;
  assign n66609 = ~n66598 & ~n66608 ;
  assign n66610 = ~n66591 & ~n66609 ;
  assign n66549 = ~n66542 & ~n66548 ;
  assign n66556 = n66549 & ~n66555 ;
  assign n66559 = ~n66556 & ~n66558 ;
  assign n66566 = ~n66559 & ~n66565 ;
  assign n66573 = n66555 & ~n66572 ;
  assign n66574 = n66542 & ~n66548 ;
  assign n66575 = ~n66573 & ~n66574 ;
  assign n66576 = n66565 & ~n66575 ;
  assign n66579 = ~n66542 & n66578 ;
  assign n66580 = ~n66576 & ~n66579 ;
  assign n66581 = n66542 & n66555 ;
  assign n66582 = ~n66548 & n66581 ;
  assign n66583 = ~n66572 & n66582 ;
  assign n66584 = ~n66580 & ~n66583 ;
  assign n66585 = ~n66566 & ~n66584 ;
  assign n66592 = ~n66585 & n66591 ;
  assign n66611 = n66548 & ~n66572 ;
  assign n66612 = ~n66542 & n66555 ;
  assign n66613 = n66611 & n66612 ;
  assign n66614 = ~n66548 & n66599 ;
  assign n66615 = n66542 & n66614 ;
  assign n66616 = ~n66613 & ~n66615 ;
  assign n66617 = n66556 & ~n66572 ;
  assign n66618 = ~n66542 & n66548 ;
  assign n66619 = n66599 & n66618 ;
  assign n66620 = ~n66617 & ~n66619 ;
  assign n66621 = n66616 & n66620 ;
  assign n66622 = n66565 & ~n66621 ;
  assign n66623 = ~n66565 & ~n66572 ;
  assign n66624 = n66582 & n66623 ;
  assign n66625 = ~n66622 & ~n66624 ;
  assign n66626 = ~n66592 & n66625 ;
  assign n66627 = ~n66610 & n66626 ;
  assign n66628 = \u0_L3_reg[5]/NET0131  & ~n66627 ;
  assign n66629 = ~\u0_L3_reg[5]/NET0131  & n66627 ;
  assign n66630 = ~n66628 & ~n66629 ;
  assign n66631 = decrypt_pad & ~\u0_uk_K_r3_reg[38]/NET0131  ;
  assign n66632 = ~decrypt_pad & ~\u0_uk_K_r3_reg[29]/NET0131  ;
  assign n66633 = ~n66631 & ~n66632 ;
  assign n66634 = \u0_R3_reg[24]/NET0131  & ~n66633 ;
  assign n66635 = ~\u0_R3_reg[24]/NET0131  & n66633 ;
  assign n66636 = ~n66634 & ~n66635 ;
  assign n66637 = decrypt_pad & ~\u0_uk_K_r3_reg[50]/NET0131  ;
  assign n66638 = ~decrypt_pad & ~\u0_uk_K_r3_reg[14]/NET0131  ;
  assign n66639 = ~n66637 & ~n66638 ;
  assign n66640 = \u0_R3_reg[22]/NET0131  & ~n66639 ;
  assign n66641 = ~\u0_R3_reg[22]/NET0131  & n66639 ;
  assign n66642 = ~n66640 & ~n66641 ;
  assign n66643 = decrypt_pad & ~\u0_uk_K_r3_reg[44]/NET0131  ;
  assign n66644 = ~decrypt_pad & ~\u0_uk_K_r3_reg[8]/NET0131  ;
  assign n66645 = ~n66643 & ~n66644 ;
  assign n66646 = \u0_R3_reg[20]/NET0131  & ~n66645 ;
  assign n66647 = ~\u0_R3_reg[20]/NET0131  & n66645 ;
  assign n66648 = ~n66646 & ~n66647 ;
  assign n66650 = decrypt_pad & ~\u0_uk_K_r3_reg[28]/NET0131  ;
  assign n66651 = ~decrypt_pad & ~\u0_uk_K_r3_reg[23]/NET0131  ;
  assign n66652 = ~n66650 & ~n66651 ;
  assign n66653 = \u0_R3_reg[21]/NET0131  & ~n66652 ;
  assign n66654 = ~\u0_R3_reg[21]/NET0131  & n66652 ;
  assign n66655 = ~n66653 & ~n66654 ;
  assign n66675 = ~n66648 & n66655 ;
  assign n66656 = decrypt_pad & ~\u0_uk_K_r3_reg[29]/NET0131  ;
  assign n66657 = ~decrypt_pad & ~\u0_uk_K_r3_reg[52]/NET0131  ;
  assign n66658 = ~n66656 & ~n66657 ;
  assign n66659 = \u0_R3_reg[25]/NET0131  & ~n66658 ;
  assign n66660 = ~\u0_R3_reg[25]/NET0131  & n66658 ;
  assign n66661 = ~n66659 & ~n66660 ;
  assign n66681 = n66648 & n66661 ;
  assign n66704 = ~n66675 & ~n66681 ;
  assign n66705 = n66642 & ~n66704 ;
  assign n66664 = decrypt_pad & ~\u0_uk_K_r3_reg[8]/NET0131  ;
  assign n66665 = ~decrypt_pad & ~\u0_uk_K_r3_reg[31]/NET0131  ;
  assign n66666 = ~n66664 & ~n66665 ;
  assign n66667 = \u0_R3_reg[23]/NET0131  & ~n66666 ;
  assign n66668 = ~\u0_R3_reg[23]/NET0131  & n66666 ;
  assign n66669 = ~n66667 & ~n66668 ;
  assign n66701 = ~n66648 & n66661 ;
  assign n66702 = n66655 & n66701 ;
  assign n66703 = ~n66642 & ~n66702 ;
  assign n66706 = ~n66669 & ~n66703 ;
  assign n66707 = ~n66705 & n66706 ;
  assign n66687 = ~n66642 & ~n66669 ;
  assign n66708 = n66681 & n66687 ;
  assign n66709 = ~n66655 & n66708 ;
  assign n66692 = n66655 & ~n66661 ;
  assign n66693 = n66648 & n66692 ;
  assign n66710 = n66669 & ~n66693 ;
  assign n66649 = ~n66642 & ~n66648 ;
  assign n66671 = ~n66642 & ~n66661 ;
  assign n66711 = ~n66655 & ~n66671 ;
  assign n66712 = ~n66649 & ~n66711 ;
  assign n66713 = n66710 & n66712 ;
  assign n66714 = ~n66709 & ~n66713 ;
  assign n66715 = ~n66707 & n66714 ;
  assign n66716 = n66636 & ~n66715 ;
  assign n66672 = n66655 & n66671 ;
  assign n66673 = ~n66649 & ~n66672 ;
  assign n66674 = n66669 & n66673 ;
  assign n66662 = ~n66655 & n66661 ;
  assign n66663 = ~n66649 & ~n66662 ;
  assign n66670 = ~n66663 & ~n66669 ;
  assign n66676 = n66642 & ~n66675 ;
  assign n66677 = ~n66670 & ~n66676 ;
  assign n66678 = ~n66674 & n66677 ;
  assign n66682 = ~n66669 & ~n66681 ;
  assign n66679 = ~n66648 & ~n66661 ;
  assign n66680 = n66642 & ~n66679 ;
  assign n66683 = ~n66655 & n66680 ;
  assign n66684 = ~n66682 & n66683 ;
  assign n66685 = ~n66678 & ~n66684 ;
  assign n66686 = ~n66636 & ~n66685 ;
  assign n66690 = ~n66648 & n66662 ;
  assign n66691 = n66669 & n66690 ;
  assign n66694 = ~n66669 & n66693 ;
  assign n66695 = ~n66691 & ~n66694 ;
  assign n66696 = ~n66642 & ~n66695 ;
  assign n66688 = n66679 & n66687 ;
  assign n66689 = ~n66655 & n66688 ;
  assign n66697 = n66642 & n66681 ;
  assign n66698 = n66649 & n66692 ;
  assign n66699 = ~n66697 & ~n66698 ;
  assign n66700 = n66669 & ~n66699 ;
  assign n66717 = ~n66689 & ~n66700 ;
  assign n66718 = ~n66696 & n66717 ;
  assign n66719 = ~n66686 & n66718 ;
  assign n66720 = ~n66716 & n66719 ;
  assign n66721 = \u0_L3_reg[11]/NET0131  & ~n66720 ;
  assign n66722 = ~\u0_L3_reg[11]/NET0131  & n66720 ;
  assign n66723 = ~n66721 & ~n66722 ;
  assign n66724 = n66556 & n66565 ;
  assign n66725 = ~n66591 & ~n66724 ;
  assign n66729 = n66555 & ~n66604 ;
  assign n66730 = ~n66574 & n66729 ;
  assign n66731 = ~n66556 & n66565 ;
  assign n66732 = ~n66614 & n66731 ;
  assign n66733 = ~n66730 & n66732 ;
  assign n66735 = n66558 & n66572 ;
  assign n66734 = ~n66572 & n66574 ;
  assign n66736 = ~n66565 & ~n66734 ;
  assign n66737 = ~n66735 & n66736 ;
  assign n66738 = ~n66733 & ~n66737 ;
  assign n66726 = ~n66572 & ~n66612 ;
  assign n66727 = n66548 & ~n66557 ;
  assign n66728 = n66726 & n66727 ;
  assign n66739 = n66556 & n66572 ;
  assign n66740 = ~n66728 & ~n66739 ;
  assign n66741 = ~n66738 & n66740 ;
  assign n66742 = ~n66725 & ~n66741 ;
  assign n66743 = n66542 & n66577 ;
  assign n66744 = n66595 & n66743 ;
  assign n66745 = ~n66555 & n66565 ;
  assign n66747 = n66618 & ~n66726 ;
  assign n66746 = n66612 & n66623 ;
  assign n66748 = n66542 & n66572 ;
  assign n66749 = ~n66548 & n66748 ;
  assign n66750 = ~n66746 & ~n66749 ;
  assign n66751 = ~n66747 & n66750 ;
  assign n66752 = ~n66745 & ~n66751 ;
  assign n66753 = ~n66572 & n66581 ;
  assign n66754 = ~n66558 & ~n66753 ;
  assign n66755 = n66565 & ~n66754 ;
  assign n66756 = ~n66601 & ~n66617 ;
  assign n66757 = ~n66755 & n66756 ;
  assign n66758 = ~n66752 & n66757 ;
  assign n66759 = ~n66591 & ~n66758 ;
  assign n66760 = ~n66744 & ~n66759 ;
  assign n66761 = ~n66742 & n66760 ;
  assign n66762 = ~\u0_L3_reg[21]/NET0131  & ~n66761 ;
  assign n66763 = \u0_L3_reg[21]/NET0131  & n66761 ;
  assign n66764 = ~n66762 & ~n66763 ;
  assign n66765 = decrypt_pad & ~\u0_uk_K_r3_reg[22]/NET0131  ;
  assign n66766 = ~decrypt_pad & ~\u0_uk_K_r3_reg[45]/P0001  ;
  assign n66767 = ~n66765 & ~n66766 ;
  assign n66768 = \u0_R3_reg[20]/NET0131  & ~n66767 ;
  assign n66769 = ~\u0_R3_reg[20]/NET0131  & n66767 ;
  assign n66770 = ~n66768 & ~n66769 ;
  assign n66798 = decrypt_pad & ~\u0_uk_K_r3_reg[7]/NET0131  ;
  assign n66799 = ~decrypt_pad & ~\u0_uk_K_r3_reg[2]/NET0131  ;
  assign n66800 = ~n66798 & ~n66799 ;
  assign n66801 = \u0_R3_reg[19]/NET0131  & ~n66800 ;
  assign n66802 = ~\u0_R3_reg[19]/NET0131  & n66800 ;
  assign n66803 = ~n66801 & ~n66802 ;
  assign n66771 = decrypt_pad & ~\u0_uk_K_r3_reg[2]/NET0131  ;
  assign n66772 = ~decrypt_pad & ~\u0_uk_K_r3_reg[21]/NET0131  ;
  assign n66773 = ~n66771 & ~n66772 ;
  assign n66774 = \u0_R3_reg[17]/NET0131  & ~n66773 ;
  assign n66775 = ~\u0_R3_reg[17]/NET0131  & n66773 ;
  assign n66776 = ~n66774 & ~n66775 ;
  assign n66784 = decrypt_pad & ~\u0_uk_K_r3_reg[35]/NET0131  ;
  assign n66785 = ~decrypt_pad & ~\u0_uk_K_r3_reg[30]/NET0131  ;
  assign n66786 = ~n66784 & ~n66785 ;
  assign n66787 = \u0_R3_reg[16]/NET0131  & ~n66786 ;
  assign n66788 = ~\u0_R3_reg[16]/NET0131  & n66786 ;
  assign n66789 = ~n66787 & ~n66788 ;
  assign n66791 = decrypt_pad & ~\u0_uk_K_r3_reg[23]/NET0131  ;
  assign n66792 = ~decrypt_pad & ~\u0_uk_K_r3_reg[42]/NET0131  ;
  assign n66793 = ~n66791 & ~n66792 ;
  assign n66794 = \u0_R3_reg[21]/NET0131  & ~n66793 ;
  assign n66795 = ~\u0_R3_reg[21]/NET0131  & n66793 ;
  assign n66796 = ~n66794 & ~n66795 ;
  assign n66804 = n66789 & ~n66796 ;
  assign n66831 = n66776 & n66804 ;
  assign n66777 = decrypt_pad & ~\u0_uk_K_r3_reg[51]/NET0131  ;
  assign n66778 = ~decrypt_pad & ~\u0_uk_K_r3_reg[15]/NET0131  ;
  assign n66779 = ~n66777 & ~n66778 ;
  assign n66780 = \u0_R3_reg[18]/NET0131  & ~n66779 ;
  assign n66781 = ~\u0_R3_reg[18]/NET0131  & n66779 ;
  assign n66782 = ~n66780 & ~n66781 ;
  assign n66783 = n66776 & ~n66782 ;
  assign n66790 = n66783 & ~n66789 ;
  assign n66822 = n66782 & n66789 ;
  assign n66832 = n66796 & ~n66822 ;
  assign n66833 = ~n66790 & n66832 ;
  assign n66834 = ~n66831 & ~n66833 ;
  assign n66835 = n66803 & ~n66834 ;
  assign n66820 = ~n66789 & ~n66796 ;
  assign n66821 = ~n66776 & n66820 ;
  assign n66811 = ~n66789 & n66796 ;
  assign n66840 = n66776 & n66811 ;
  assign n66841 = ~n66821 & ~n66840 ;
  assign n66842 = ~n66782 & ~n66803 ;
  assign n66843 = ~n66841 & n66842 ;
  assign n66817 = n66789 & n66796 ;
  assign n66805 = ~n66776 & ~n66782 ;
  assign n66809 = n66776 & n66782 ;
  assign n66836 = ~n66803 & n66809 ;
  assign n66837 = ~n66805 & ~n66836 ;
  assign n66838 = n66817 & ~n66837 ;
  assign n66839 = ~n66782 & n66831 ;
  assign n66844 = ~n66776 & n66782 ;
  assign n66845 = n66804 & n66844 ;
  assign n66846 = ~n66839 & ~n66845 ;
  assign n66847 = ~n66838 & n66846 ;
  assign n66848 = ~n66843 & n66847 ;
  assign n66849 = ~n66835 & n66848 ;
  assign n66850 = n66770 & ~n66849 ;
  assign n66807 = n66783 & n66796 ;
  assign n66808 = n66789 & n66807 ;
  assign n66812 = ~n66776 & n66811 ;
  assign n66806 = n66804 & n66805 ;
  assign n66810 = ~n66796 & n66809 ;
  assign n66813 = ~n66806 & ~n66810 ;
  assign n66814 = ~n66812 & n66813 ;
  assign n66815 = ~n66808 & n66814 ;
  assign n66816 = ~n66803 & ~n66815 ;
  assign n66823 = n66796 & n66822 ;
  assign n66824 = ~n66790 & ~n66821 ;
  assign n66825 = ~n66823 & n66824 ;
  assign n66826 = n66803 & ~n66825 ;
  assign n66797 = n66790 & ~n66796 ;
  assign n66818 = ~n66776 & n66817 ;
  assign n66819 = n66782 & n66818 ;
  assign n66827 = ~n66797 & ~n66819 ;
  assign n66828 = ~n66826 & n66827 ;
  assign n66829 = ~n66816 & n66828 ;
  assign n66830 = ~n66770 & ~n66829 ;
  assign n66851 = n66782 & n66821 ;
  assign n66852 = ~n66839 & ~n66851 ;
  assign n66853 = n66803 & ~n66852 ;
  assign n66854 = n66811 & n66844 ;
  assign n66855 = ~n66789 & n66810 ;
  assign n66856 = ~n66854 & ~n66855 ;
  assign n66857 = ~n66803 & ~n66856 ;
  assign n66858 = ~n66853 & ~n66857 ;
  assign n66859 = ~n66830 & n66858 ;
  assign n66860 = ~n66850 & n66859 ;
  assign n66861 = ~\u0_L3_reg[14]/NET0131  & ~n66860 ;
  assign n66862 = \u0_L3_reg[14]/NET0131  & n66860 ;
  assign n66863 = ~n66861 & ~n66862 ;
  assign n66864 = decrypt_pad & ~\u0_uk_K_r3_reg[40]/NET0131  ;
  assign n66865 = ~decrypt_pad & ~\u0_uk_K_r3_reg[6]/NET0131  ;
  assign n66866 = ~n66864 & ~n66865 ;
  assign n66867 = \u0_R3_reg[8]/NET0131  & ~n66866 ;
  assign n66868 = ~\u0_R3_reg[8]/NET0131  & n66866 ;
  assign n66869 = ~n66867 & ~n66868 ;
  assign n66870 = decrypt_pad & ~\u0_uk_K_r3_reg[55]/NET0131  ;
  assign n66871 = ~decrypt_pad & ~\u0_uk_K_r3_reg[46]/NET0131  ;
  assign n66872 = ~n66870 & ~n66871 ;
  assign n66873 = \u0_R3_reg[6]/NET0131  & ~n66872 ;
  assign n66874 = ~\u0_R3_reg[6]/NET0131  & n66872 ;
  assign n66875 = ~n66873 & ~n66874 ;
  assign n66876 = decrypt_pad & ~\u0_uk_K_r3_reg[20]/NET0131  ;
  assign n66877 = ~decrypt_pad & ~\u0_uk_K_r3_reg[11]/NET0131  ;
  assign n66878 = ~n66876 & ~n66877 ;
  assign n66879 = \u0_R3_reg[9]/NET0131  & ~n66878 ;
  assign n66880 = ~\u0_R3_reg[9]/NET0131  & n66878 ;
  assign n66881 = ~n66879 & ~n66880 ;
  assign n66882 = ~n66875 & n66881 ;
  assign n66883 = decrypt_pad & ~\u0_uk_K_r3_reg[32]/NET0131  ;
  assign n66884 = ~decrypt_pad & ~\u0_uk_K_r3_reg[55]/NET0131  ;
  assign n66885 = ~n66883 & ~n66884 ;
  assign n66886 = \u0_R3_reg[5]/NET0131  & ~n66885 ;
  assign n66887 = ~\u0_R3_reg[5]/NET0131  & n66885 ;
  assign n66888 = ~n66886 & ~n66887 ;
  assign n66889 = decrypt_pad & ~\u0_uk_K_r3_reg[17]/NET0131  ;
  assign n66890 = ~decrypt_pad & ~\u0_uk_K_r3_reg[40]/NET0131  ;
  assign n66891 = ~n66889 & ~n66890 ;
  assign n66892 = \u0_R3_reg[7]/NET0131  & ~n66891 ;
  assign n66893 = ~\u0_R3_reg[7]/NET0131  & n66891 ;
  assign n66894 = ~n66892 & ~n66893 ;
  assign n66895 = ~n66888 & ~n66894 ;
  assign n66896 = n66882 & n66895 ;
  assign n66897 = decrypt_pad & ~\u0_uk_K_r3_reg[53]/NET0131  ;
  assign n66898 = ~decrypt_pad & ~\u0_uk_K_r3_reg[19]/NET0131  ;
  assign n66899 = ~n66897 & ~n66898 ;
  assign n66900 = \u0_R3_reg[4]/NET0131  & ~n66899 ;
  assign n66901 = ~\u0_R3_reg[4]/NET0131  & n66899 ;
  assign n66902 = ~n66900 & ~n66901 ;
  assign n66903 = n66881 & ~n66902 ;
  assign n66904 = n66888 & n66903 ;
  assign n66905 = n66875 & n66904 ;
  assign n66906 = ~n66896 & ~n66905 ;
  assign n66908 = n66881 & ~n66888 ;
  assign n66913 = n66875 & n66902 ;
  assign n66914 = n66908 & n66913 ;
  assign n66915 = n66894 & n66914 ;
  assign n66920 = n66906 & ~n66915 ;
  assign n66907 = n66881 & n66902 ;
  assign n66909 = ~n66881 & n66888 ;
  assign n66910 = ~n66908 & ~n66909 ;
  assign n66911 = ~n66907 & ~n66910 ;
  assign n66912 = ~n66875 & n66911 ;
  assign n66916 = ~n66888 & n66907 ;
  assign n66917 = ~n66894 & ~n66916 ;
  assign n66918 = ~n66908 & ~n66913 ;
  assign n66919 = n66917 & ~n66918 ;
  assign n66921 = ~n66912 & ~n66919 ;
  assign n66922 = n66920 & n66921 ;
  assign n66923 = ~n66869 & ~n66922 ;
  assign n66925 = ~n66881 & ~n66902 ;
  assign n66942 = ~n66914 & ~n66925 ;
  assign n66943 = n66869 & ~n66942 ;
  assign n66924 = n66875 & ~n66888 ;
  assign n66944 = n66903 & ~n66924 ;
  assign n66945 = ~n66943 & ~n66944 ;
  assign n66941 = ~n66875 & n66888 ;
  assign n66946 = ~n66894 & ~n66941 ;
  assign n66947 = ~n66945 & n66946 ;
  assign n66926 = n66924 & n66925 ;
  assign n66927 = n66888 & n66902 ;
  assign n66928 = ~n66875 & n66927 ;
  assign n66929 = ~n66926 & ~n66928 ;
  assign n66930 = n66894 & ~n66929 ;
  assign n66931 = ~n66881 & ~n66888 ;
  assign n66932 = ~n66875 & n66931 ;
  assign n66933 = n66902 & n66932 ;
  assign n66934 = n66875 & ~n66902 ;
  assign n66935 = n66888 & n66894 ;
  assign n66936 = ~n66934 & n66935 ;
  assign n66937 = n66882 & n66927 ;
  assign n66938 = ~n66936 & ~n66937 ;
  assign n66939 = ~n66933 & n66938 ;
  assign n66940 = n66869 & ~n66939 ;
  assign n66948 = ~n66930 & ~n66940 ;
  assign n66949 = ~n66947 & n66948 ;
  assign n66950 = ~n66923 & n66949 ;
  assign n66951 = \u0_L3_reg[2]/NET0131  & n66950 ;
  assign n66952 = ~\u0_L3_reg[2]/NET0131  & ~n66950 ;
  assign n66953 = ~n66951 & ~n66952 ;
  assign n66959 = n66642 & n66690 ;
  assign n66960 = n66655 & n66679 ;
  assign n66961 = ~n66959 & ~n66960 ;
  assign n66962 = ~n66669 & ~n66961 ;
  assign n66954 = ~n66655 & n66697 ;
  assign n66955 = ~n66642 & n66701 ;
  assign n66956 = ~n66693 & ~n66955 ;
  assign n66957 = ~n66954 & n66956 ;
  assign n66958 = n66669 & ~n66957 ;
  assign n66963 = n66648 & ~n66655 ;
  assign n66964 = n66671 & n66963 ;
  assign n66965 = ~n66708 & ~n66964 ;
  assign n66966 = ~n66958 & n66965 ;
  assign n66967 = ~n66962 & n66966 ;
  assign n66968 = ~n66636 & ~n66967 ;
  assign n66976 = ~n66669 & ~n66673 ;
  assign n66979 = n66655 & n66661 ;
  assign n66980 = n66642 & n66979 ;
  assign n66977 = ~n66642 & n66669 ;
  assign n66978 = n66681 & n66977 ;
  assign n66981 = ~n66698 & ~n66978 ;
  assign n66982 = ~n66980 & n66981 ;
  assign n66983 = ~n66976 & n66982 ;
  assign n66984 = n66636 & ~n66983 ;
  assign n66969 = ~n66662 & ~n66692 ;
  assign n66972 = n66648 & n66969 ;
  assign n66973 = ~n66669 & ~n66972 ;
  assign n66970 = ~n66648 & n66969 ;
  assign n66971 = n66710 & ~n66970 ;
  assign n66974 = n66642 & ~n66971 ;
  assign n66975 = ~n66973 & n66974 ;
  assign n66985 = ~n66688 & ~n66975 ;
  assign n66986 = ~n66984 & n66985 ;
  assign n66987 = ~n66968 & n66986 ;
  assign n66988 = ~\u0_L3_reg[4]/NET0131  & ~n66987 ;
  assign n66989 = \u0_L3_reg[4]/NET0131  & n66987 ;
  assign n66990 = ~n66988 & ~n66989 ;
  assign n67015 = ~n66459 & n66477 ;
  assign n67016 = ~n66482 & ~n67015 ;
  assign n67017 = ~n66447 & ~n67016 ;
  assign n67019 = n66453 & ~n66488 ;
  assign n67020 = n66526 & n67019 ;
  assign n67018 = ~n66466 & n66506 ;
  assign n67021 = ~n66474 & ~n67018 ;
  assign n67022 = ~n66498 & n67021 ;
  assign n67023 = ~n67020 & n67022 ;
  assign n67024 = ~n67017 & n67023 ;
  assign n67025 = ~n66496 & ~n67024 ;
  assign n66991 = n66466 & n66488 ;
  assign n66992 = ~n66483 & ~n66991 ;
  assign n66993 = n66447 & ~n66992 ;
  assign n66994 = ~n66466 & ~n66472 ;
  assign n66995 = ~n66459 & n66994 ;
  assign n66996 = n66453 & n66995 ;
  assign n67004 = ~n66993 & ~n66996 ;
  assign n66997 = n66453 & n66488 ;
  assign n66998 = ~n66497 & ~n66997 ;
  assign n66999 = n66466 & ~n66998 ;
  assign n67000 = ~n66453 & n66473 ;
  assign n67001 = ~n66499 & ~n67000 ;
  assign n67002 = ~n66447 & ~n66518 ;
  assign n67003 = ~n67001 & n67002 ;
  assign n67005 = ~n66999 & ~n67003 ;
  assign n67006 = n67004 & n67005 ;
  assign n67007 = n66496 & ~n67006 ;
  assign n67010 = ~n66472 & ~n66507 ;
  assign n67011 = ~n66447 & ~n66500 ;
  assign n67012 = ~n67010 & n67011 ;
  assign n67008 = n66472 & ~n66507 ;
  assign n67009 = n66447 & ~n67008 ;
  assign n67013 = ~n66466 & ~n67009 ;
  assign n67014 = ~n67012 & n67013 ;
  assign n67026 = ~n67007 & ~n67014 ;
  assign n67027 = ~n67025 & n67026 ;
  assign n67028 = ~\u0_L3_reg[26]/NET0131  & ~n67027 ;
  assign n67029 = \u0_L3_reg[26]/NET0131  & n67027 ;
  assign n67030 = ~n67028 & ~n67029 ;
  assign n67031 = ~n66555 & n66734 ;
  assign n67032 = ~n66581 & ~n66594 ;
  assign n67033 = ~n66600 & n67032 ;
  assign n67034 = n66565 & ~n67033 ;
  assign n67035 = ~n67031 & ~n67034 ;
  assign n67036 = ~n66591 & ~n67035 ;
  assign n67042 = ~n66582 & ~n66613 ;
  assign n67039 = n66548 & ~n66565 ;
  assign n67040 = n66599 & n67039 ;
  assign n67041 = n66604 & n66745 ;
  assign n67043 = ~n67040 & ~n67041 ;
  assign n67044 = n67042 & n67043 ;
  assign n67045 = ~n66735 & n67044 ;
  assign n67046 = n66591 & ~n67045 ;
  assign n67037 = ~n66579 & ~n66739 ;
  assign n67038 = n66565 & ~n67037 ;
  assign n67049 = n66549 & ~n66573 ;
  assign n67050 = ~n66599 & n67049 ;
  assign n67047 = ~n66548 & n66591 ;
  assign n67048 = n66557 & ~n67047 ;
  assign n67051 = ~n66613 & ~n67048 ;
  assign n67052 = ~n67050 & n67051 ;
  assign n67053 = ~n66565 & ~n67052 ;
  assign n67054 = ~n67038 & ~n67053 ;
  assign n67055 = ~n67046 & n67054 ;
  assign n67056 = ~n67036 & n67055 ;
  assign n67057 = \u0_L3_reg[15]/P0001  & n67056 ;
  assign n67058 = ~\u0_L3_reg[15]/P0001  & ~n67056 ;
  assign n67059 = ~n67057 & ~n67058 ;
  assign n67075 = ~n66517 & ~n66994 ;
  assign n67076 = n66459 & ~n67075 ;
  assign n67077 = ~n66447 & ~n67076 ;
  assign n67078 = n66479 & ~n66995 ;
  assign n67079 = ~n67077 & ~n67078 ;
  assign n67080 = ~n66481 & n66502 ;
  assign n67081 = ~n67079 & n67080 ;
  assign n67082 = ~n66496 & ~n67081 ;
  assign n67069 = ~n66476 & n66480 ;
  assign n67070 = ~n66997 & ~n67069 ;
  assign n67071 = ~n66447 & ~n67070 ;
  assign n67067 = n66466 & n66497 ;
  assign n67072 = ~n67015 & ~n67067 ;
  assign n67073 = ~n67071 & n67072 ;
  assign n67074 = n66496 & ~n67073 ;
  assign n67060 = n66477 & n66488 ;
  assign n67061 = ~n66501 & ~n67060 ;
  assign n67062 = ~n66515 & n67061 ;
  assign n67063 = n66447 & ~n67062 ;
  assign n67068 = ~n66447 & n67067 ;
  assign n67064 = ~n66517 & ~n67018 ;
  assign n67065 = n66447 & n66496 ;
  assign n67066 = ~n67064 & n67065 ;
  assign n67083 = ~n66504 & ~n67066 ;
  assign n67084 = ~n67068 & n67083 ;
  assign n67085 = ~n67063 & n67084 ;
  assign n67086 = ~n67074 & n67085 ;
  assign n67087 = ~n67082 & n67086 ;
  assign n67088 = ~\u0_L3_reg[1]/NET0131  & ~n67087 ;
  assign n67089 = \u0_L3_reg[1]/NET0131  & n67087 ;
  assign n67090 = ~n67088 & ~n67089 ;
  assign n67094 = ~n66875 & n66925 ;
  assign n67095 = ~n66904 & ~n67094 ;
  assign n67096 = n66894 & n67095 ;
  assign n67100 = ~n66888 & n66934 ;
  assign n67101 = ~n66894 & ~n67100 ;
  assign n67098 = ~n66881 & n66902 ;
  assign n67099 = ~n66875 & n67098 ;
  assign n67097 = ~n66888 & n66903 ;
  assign n67102 = ~n66927 & ~n67097 ;
  assign n67103 = ~n67099 & n67102 ;
  assign n67104 = n67101 & n67103 ;
  assign n67105 = ~n67096 & ~n67104 ;
  assign n67092 = ~n66907 & ~n66925 ;
  assign n67093 = n66924 & ~n67092 ;
  assign n67091 = n66909 & n66913 ;
  assign n67106 = ~n66869 & ~n67091 ;
  assign n67107 = ~n67093 & n67106 ;
  assign n67108 = ~n67105 & n67107 ;
  assign n67114 = n66902 & n66910 ;
  assign n67113 = n66909 & n66934 ;
  assign n67115 = n66894 & ~n67113 ;
  assign n67116 = ~n67114 & n67115 ;
  assign n67117 = ~n67091 & n67095 ;
  assign n67118 = n67101 & n67117 ;
  assign n67119 = ~n67116 & ~n67118 ;
  assign n67109 = n66894 & n66902 ;
  assign n67110 = ~n66916 & ~n67109 ;
  assign n67111 = ~n66875 & ~n67110 ;
  assign n67112 = n66903 & n66924 ;
  assign n67120 = n66869 & ~n67112 ;
  assign n67121 = ~n67111 & n67120 ;
  assign n67122 = ~n67119 & n67121 ;
  assign n67123 = ~n67108 & ~n67122 ;
  assign n67124 = ~\u0_L3_reg[28]/NET0131  & n67123 ;
  assign n67125 = \u0_L3_reg[28]/NET0131  & ~n67123 ;
  assign n67126 = ~n67124 & ~n67125 ;
  assign n67136 = n66499 & n66505 ;
  assign n67140 = n66453 & n66518 ;
  assign n67141 = ~n67136 & ~n67140 ;
  assign n67142 = ~n66503 & n67141 ;
  assign n67137 = ~n66466 & n66489 ;
  assign n67138 = n66447 & ~n66473 ;
  assign n67139 = n66506 & n67138 ;
  assign n67143 = ~n67137 & ~n67139 ;
  assign n67144 = n67142 & n67143 ;
  assign n67145 = n66516 & n67144 ;
  assign n67146 = ~n66496 & ~n67145 ;
  assign n67130 = n66476 & ~n66480 ;
  assign n67131 = ~n66474 & ~n67130 ;
  assign n67132 = ~n66447 & ~n67131 ;
  assign n67128 = ~n66514 & ~n66519 ;
  assign n67129 = n66447 & ~n67128 ;
  assign n67133 = n67061 & ~n67129 ;
  assign n67134 = ~n67132 & n67133 ;
  assign n67135 = n66496 & ~n67134 ;
  assign n67147 = ~n66484 & n67061 ;
  assign n67148 = ~n66447 & ~n67147 ;
  assign n67127 = n66447 & n66481 ;
  assign n67149 = ~n66527 & ~n67127 ;
  assign n67150 = ~n67148 & n67149 ;
  assign n67151 = ~n67135 & n67150 ;
  assign n67152 = ~n67146 & n67151 ;
  assign n67153 = ~\u0_L3_reg[10]/NET0131  & ~n67152 ;
  assign n67154 = \u0_L3_reg[10]/NET0131  & n67152 ;
  assign n67155 = ~n67153 & ~n67154 ;
  assign n67162 = ~n66642 & ~n66704 ;
  assign n67163 = n66642 & n66693 ;
  assign n67164 = ~n67162 & ~n67163 ;
  assign n67165 = ~n66669 & ~n67164 ;
  assign n67157 = ~n66642 & n66655 ;
  assign n67158 = ~n66661 & ~n67157 ;
  assign n67159 = ~n66676 & n67158 ;
  assign n67160 = ~n66972 & ~n67159 ;
  assign n67161 = n66669 & ~n67160 ;
  assign n67166 = ~n66636 & ~n66959 ;
  assign n67167 = ~n67161 & n67166 ;
  assign n67168 = ~n67165 & n67167 ;
  assign n67174 = n66680 & ~n66681 ;
  assign n67173 = n66669 & ~n66711 ;
  assign n67175 = ~n67162 & ~n67173 ;
  assign n67176 = ~n67174 & n67175 ;
  assign n67169 = n66642 & ~n66661 ;
  assign n67170 = n66675 & ~n67169 ;
  assign n67171 = ~n67163 & ~n67170 ;
  assign n67172 = n66669 & ~n67171 ;
  assign n67177 = n66636 & ~n67172 ;
  assign n67178 = ~n67176 & n67177 ;
  assign n67179 = ~n67168 & ~n67178 ;
  assign n67156 = n66977 & n66979 ;
  assign n67180 = ~n66964 & ~n67156 ;
  assign n67181 = ~n67179 & n67180 ;
  assign n67182 = \u0_L3_reg[29]/NET0131  & ~n67181 ;
  assign n67183 = ~\u0_L3_reg[29]/NET0131  & n67181 ;
  assign n67184 = ~n67182 & ~n67183 ;
  assign n67202 = ~n66383 & ~n66402 ;
  assign n67203 = n66350 & n67202 ;
  assign n67204 = ~n66350 & ~n67202 ;
  assign n67205 = ~n67203 & ~n67204 ;
  assign n67194 = n66350 & ~n66384 ;
  assign n67206 = n66400 & ~n67194 ;
  assign n67207 = ~n67205 & n67206 ;
  assign n67208 = n66350 & n66403 ;
  assign n67209 = n66370 & n66426 ;
  assign n67210 = ~n66425 & ~n67209 ;
  assign n67211 = ~n67208 & n67210 ;
  assign n67212 = ~n67207 & n67211 ;
  assign n67213 = ~n66377 & ~n67212 ;
  assign n67189 = ~n66371 & ~n66400 ;
  assign n67190 = ~n66406 & n67189 ;
  assign n67185 = ~n66363 & ~n66405 ;
  assign n67186 = n66390 & ~n67185 ;
  assign n67187 = ~n66402 & ~n66405 ;
  assign n67188 = n66431 & ~n67187 ;
  assign n67191 = ~n67186 & ~n67188 ;
  assign n67192 = n67190 & n67191 ;
  assign n67195 = n66363 & n66377 ;
  assign n67196 = ~n66385 & n67195 ;
  assign n67197 = ~n67194 & n67196 ;
  assign n67193 = n66370 & n66412 ;
  assign n67198 = n66400 & ~n67193 ;
  assign n67199 = ~n66433 & n67198 ;
  assign n67200 = ~n67197 & n67199 ;
  assign n67201 = ~n67192 & ~n67200 ;
  assign n67214 = ~n66418 & ~n67201 ;
  assign n67215 = ~n67213 & n67214 ;
  assign n67216 = \u0_L3_reg[23]/NET0131  & ~n67215 ;
  assign n67217 = ~\u0_L3_reg[23]/NET0131  & n67215 ;
  assign n67218 = ~n67216 & ~n67217 ;
  assign n67220 = n66805 & n66820 ;
  assign n67221 = ~n66818 & ~n67220 ;
  assign n67222 = n66803 & ~n67221 ;
  assign n67219 = n66789 & n66842 ;
  assign n67223 = n66770 & ~n67219 ;
  assign n67224 = n66856 & n67223 ;
  assign n67225 = ~n67222 & n67224 ;
  assign n67226 = n66776 & n66817 ;
  assign n67227 = ~n66806 & ~n67226 ;
  assign n67228 = n66803 & ~n67227 ;
  assign n67234 = ~n66770 & ~n66790 ;
  assign n67235 = ~n67228 & n67234 ;
  assign n67229 = n66811 & ~n66844 ;
  assign n67230 = ~n66818 & ~n67229 ;
  assign n67231 = ~n66803 & ~n67230 ;
  assign n67232 = n66782 & n66831 ;
  assign n67233 = ~n66851 & ~n67232 ;
  assign n67236 = ~n67231 & n67233 ;
  assign n67237 = n67235 & n67236 ;
  assign n67238 = ~n67225 & ~n67237 ;
  assign n67239 = ~n66803 & ~n66845 ;
  assign n67241 = n66790 & n66796 ;
  assign n67240 = n66803 & ~n66854 ;
  assign n67242 = ~n66810 & n67240 ;
  assign n67243 = ~n67241 & n67242 ;
  assign n67244 = ~n67239 & ~n67243 ;
  assign n67245 = ~n67238 & ~n67244 ;
  assign n67246 = ~\u0_L3_reg[8]/NET0131  & ~n67245 ;
  assign n67247 = \u0_L3_reg[8]/NET0131  & n67245 ;
  assign n67248 = ~n67246 & ~n67247 ;
  assign n67249 = ~n66291 & ~n66304 ;
  assign n67250 = ~n66267 & n66317 ;
  assign n67251 = n66293 & ~n67250 ;
  assign n67252 = ~n67249 & ~n67251 ;
  assign n67253 = ~n66288 & ~n67252 ;
  assign n67254 = ~n66280 & n66312 ;
  assign n67258 = n66288 & ~n67254 ;
  assign n67255 = n66267 & n66280 ;
  assign n67256 = ~n66274 & n67255 ;
  assign n67257 = ~n66280 & n66317 ;
  assign n67259 = ~n67256 & ~n67257 ;
  assign n67260 = n67258 & n67259 ;
  assign n67261 = ~n67253 & ~n67260 ;
  assign n67262 = n66289 & n66321 ;
  assign n67263 = ~n67261 & ~n67262 ;
  assign n67264 = n66255 & ~n67263 ;
  assign n67268 = ~n66274 & n66289 ;
  assign n67271 = n66280 & n66315 ;
  assign n67272 = ~n67268 & ~n67271 ;
  assign n67273 = n66288 & ~n67272 ;
  assign n67266 = ~n66267 & ~n66280 ;
  assign n67267 = ~n67255 & ~n67266 ;
  assign n67269 = ~n66288 & ~n67267 ;
  assign n67270 = ~n67268 & n67269 ;
  assign n67265 = n66268 & ~n66313 ;
  assign n67274 = n66331 & ~n67265 ;
  assign n67275 = ~n67270 & n67274 ;
  assign n67276 = ~n67273 & n67275 ;
  assign n67277 = ~n66255 & ~n67276 ;
  assign n67278 = n66288 & n66328 ;
  assign n67279 = ~n66292 & ~n67256 ;
  assign n67280 = ~n66288 & ~n66334 ;
  assign n67281 = ~n67279 & n67280 ;
  assign n67282 = ~n67278 & ~n67281 ;
  assign n67283 = ~n67277 & n67282 ;
  assign n67284 = ~n67264 & n67283 ;
  assign n67285 = \u0_L3_reg[32]/NET0131  & n67284 ;
  assign n67286 = ~\u0_L3_reg[32]/NET0131  & ~n67284 ;
  assign n67287 = ~n67285 & ~n67286 ;
  assign n67289 = n66648 & n67157 ;
  assign n67290 = n66669 & ~n67289 ;
  assign n67300 = ~n66980 & ~n67290 ;
  assign n67301 = n66648 & ~n67300 ;
  assign n67299 = ~n66669 & n66970 ;
  assign n67302 = n66692 & n67290 ;
  assign n67303 = ~n67299 & ~n67302 ;
  assign n67304 = ~n67301 & n67303 ;
  assign n67305 = ~n66636 & ~n67304 ;
  assign n67291 = ~n66669 & ~n66963 ;
  assign n67292 = ~n67290 & ~n67291 ;
  assign n67288 = n66642 & n66970 ;
  assign n67293 = ~n66642 & ~n66963 ;
  assign n67294 = ~n66969 & n67293 ;
  assign n67295 = ~n66691 & ~n67294 ;
  assign n67296 = ~n67288 & n67295 ;
  assign n67297 = ~n67292 & n67296 ;
  assign n67298 = n66636 & ~n67297 ;
  assign n67306 = ~n66696 & ~n66709 ;
  assign n67307 = ~n67298 & n67306 ;
  assign n67308 = ~n67305 & n67307 ;
  assign n67309 = ~\u0_L3_reg[19]/P0001  & ~n67308 ;
  assign n67310 = \u0_L3_reg[19]/P0001  & n67308 ;
  assign n67311 = ~n67309 & ~n67310 ;
  assign n67312 = n66549 & n66573 ;
  assign n67313 = n66565 & ~n66743 ;
  assign n67314 = ~n67312 & n67313 ;
  assign n67315 = n66729 & ~n66748 ;
  assign n67316 = ~n66556 & ~n66565 ;
  assign n67317 = ~n67315 & n67316 ;
  assign n67318 = ~n67314 & ~n67317 ;
  assign n67319 = ~n66579 & ~n66614 ;
  assign n67320 = ~n66601 & n67319 ;
  assign n67321 = ~n67318 & n67320 ;
  assign n67322 = n66591 & ~n67321 ;
  assign n67324 = ~n66593 & ~n66726 ;
  assign n67325 = n66565 & ~n66594 ;
  assign n67326 = ~n67324 & n67325 ;
  assign n67323 = n66748 & n67039 ;
  assign n67327 = ~n66619 & ~n66746 ;
  assign n67328 = ~n67323 & n67327 ;
  assign n67329 = ~n67326 & n67328 ;
  assign n67330 = ~n66591 & ~n67329 ;
  assign n67331 = ~n66565 & ~n66616 ;
  assign n67332 = n66611 & n66745 ;
  assign n67333 = ~n66624 & ~n67332 ;
  assign n67334 = ~n67331 & n67333 ;
  assign n67335 = ~n67330 & n67334 ;
  assign n67336 = ~n67322 & n67335 ;
  assign n67337 = ~\u0_L3_reg[27]/NET0131  & ~n67336 ;
  assign n67338 = \u0_L3_reg[27]/NET0131  & n67336 ;
  assign n67339 = ~n67337 & ~n67338 ;
  assign n67374 = decrypt_pad & ~\u0_uk_K_r3_reg[3]/NET0131  ;
  assign n67375 = ~decrypt_pad & ~\u0_uk_K_r3_reg[26]/NET0131  ;
  assign n67376 = ~n67374 & ~n67375 ;
  assign n67377 = \u0_R3_reg[11]/NET0131  & ~n67376 ;
  assign n67378 = ~\u0_R3_reg[11]/NET0131  & n67376 ;
  assign n67379 = ~n67377 & ~n67378 ;
  assign n67366 = decrypt_pad & ~\u0_uk_K_r3_reg[18]/NET0131  ;
  assign n67367 = ~decrypt_pad & ~\u0_uk_K_r3_reg[41]/NET0131  ;
  assign n67368 = ~n67366 & ~n67367 ;
  assign n67369 = \u0_R3_reg[12]/NET0131  & ~n67368 ;
  assign n67370 = ~\u0_R3_reg[12]/NET0131  & n67368 ;
  assign n67371 = ~n67369 & ~n67370 ;
  assign n67340 = decrypt_pad & ~\u0_uk_K_r3_reg[6]/NET0131  ;
  assign n67341 = ~decrypt_pad & ~\u0_uk_K_r3_reg[54]/NET0131  ;
  assign n67342 = ~n67340 & ~n67341 ;
  assign n67343 = \u0_R3_reg[13]/NET0131  & ~n67342 ;
  assign n67344 = ~\u0_R3_reg[13]/NET0131  & n67342 ;
  assign n67345 = ~n67343 & ~n67344 ;
  assign n67353 = decrypt_pad & ~\u0_uk_K_r3_reg[26]/NET0131  ;
  assign n67354 = ~decrypt_pad & ~\u0_uk_K_r3_reg[17]/NET0131  ;
  assign n67355 = ~n67353 & ~n67354 ;
  assign n67356 = \u0_R3_reg[9]/NET0131  & ~n67355 ;
  assign n67357 = ~\u0_R3_reg[9]/NET0131  & n67355 ;
  assign n67358 = ~n67356 & ~n67357 ;
  assign n67380 = n67345 & ~n67358 ;
  assign n67359 = decrypt_pad & ~\u0_uk_K_r3_reg[34]/NET0131  ;
  assign n67360 = ~decrypt_pad & ~\u0_uk_K_r3_reg[25]/NET0131  ;
  assign n67361 = ~n67359 & ~n67360 ;
  assign n67362 = \u0_R3_reg[10]/NET0131  & ~n67361 ;
  assign n67363 = ~\u0_R3_reg[10]/NET0131  & n67361 ;
  assign n67364 = ~n67362 & ~n67363 ;
  assign n67346 = decrypt_pad & ~\u0_uk_K_r3_reg[54]/NET0131  ;
  assign n67347 = ~decrypt_pad & ~\u0_uk_K_r3_reg[20]/NET0131  ;
  assign n67348 = ~n67346 & ~n67347 ;
  assign n67349 = \u0_R3_reg[8]/NET0131  & ~n67348 ;
  assign n67350 = ~\u0_R3_reg[8]/NET0131  & n67348 ;
  assign n67351 = ~n67349 & ~n67350 ;
  assign n67382 = n67345 & ~n67351 ;
  assign n67383 = n67364 & n67382 ;
  assign n67384 = ~n67345 & n67358 ;
  assign n67385 = n67351 & n67384 ;
  assign n67386 = ~n67383 & ~n67385 ;
  assign n67387 = ~n67380 & n67386 ;
  assign n67388 = n67371 & ~n67387 ;
  assign n67381 = n67364 & n67380 ;
  assign n67389 = ~n67351 & ~n67358 ;
  assign n67390 = ~n67345 & n67389 ;
  assign n67391 = ~n67364 & n67390 ;
  assign n67392 = ~n67381 & ~n67391 ;
  assign n67393 = ~n67388 & n67392 ;
  assign n67394 = n67379 & ~n67393 ;
  assign n67365 = n67358 & n67364 ;
  assign n67401 = ~n67358 & ~n67364 ;
  assign n67402 = ~n67365 & ~n67401 ;
  assign n67403 = ~n67351 & n67379 ;
  assign n67352 = ~n67345 & ~n67351 ;
  assign n67405 = n67345 & n67351 ;
  assign n67406 = ~n67352 & ~n67405 ;
  assign n67409 = ~n67403 & n67406 ;
  assign n67410 = ~n67402 & ~n67409 ;
  assign n67404 = ~n67364 & n67403 ;
  assign n67407 = n67402 & ~n67404 ;
  assign n67408 = n67406 & n67407 ;
  assign n67411 = ~n67371 & ~n67408 ;
  assign n67412 = ~n67410 & n67411 ;
  assign n67372 = n67365 & n67371 ;
  assign n67373 = n67352 & n67372 ;
  assign n67395 = n67358 & ~n67364 ;
  assign n67396 = ~n67351 & ~n67395 ;
  assign n67397 = n67371 & ~n67379 ;
  assign n67398 = ~n67380 & n67397 ;
  assign n67399 = ~n67384 & n67398 ;
  assign n67400 = ~n67396 & n67399 ;
  assign n67413 = ~n67373 & ~n67400 ;
  assign n67414 = ~n67412 & n67413 ;
  assign n67415 = ~n67394 & n67414 ;
  assign n67416 = ~\u0_L3_reg[6]/NET0131  & ~n67415 ;
  assign n67417 = \u0_L3_reg[6]/NET0131  & n67415 ;
  assign n67418 = ~n67416 & ~n67417 ;
  assign n67420 = ~n66261 & ~n66322 ;
  assign n67419 = n66267 & ~n66291 ;
  assign n67421 = ~n67257 & ~n67419 ;
  assign n67422 = ~n67420 & n67421 ;
  assign n67423 = ~n66288 & ~n67422 ;
  assign n67424 = ~n67271 & ~n67419 ;
  assign n67425 = n66274 & ~n67424 ;
  assign n67426 = ~n66274 & ~n67266 ;
  assign n67427 = n66291 & n67426 ;
  assign n67428 = n66288 & n67427 ;
  assign n67429 = n66255 & ~n67428 ;
  assign n67430 = ~n67425 & n67429 ;
  assign n67431 = ~n67423 & n67430 ;
  assign n67434 = n66274 & n67419 ;
  assign n67432 = n66274 & ~n66315 ;
  assign n67433 = n66291 & ~n67432 ;
  assign n67435 = n66288 & ~n67433 ;
  assign n67436 = ~n67434 & n67435 ;
  assign n67437 = ~n66255 & ~n67436 ;
  assign n67438 = ~n67431 & ~n67437 ;
  assign n67439 = ~n66288 & n67425 ;
  assign n67440 = n66255 & ~n66288 ;
  assign n67441 = ~n66288 & n67427 ;
  assign n67442 = n66274 & n67254 ;
  assign n67443 = ~n67441 & ~n67442 ;
  assign n67444 = ~n67440 & ~n67443 ;
  assign n67445 = ~n67439 & ~n67444 ;
  assign n67446 = ~n67438 & n67445 ;
  assign n67447 = ~\u0_L3_reg[7]/NET0131  & ~n67446 ;
  assign n67448 = \u0_L3_reg[7]/NET0131  & n67446 ;
  assign n67449 = ~n67447 & ~n67448 ;
  assign n67450 = ~n66937 & ~n67091 ;
  assign n67451 = ~n66902 & n66909 ;
  assign n67452 = ~n67112 & ~n67451 ;
  assign n67453 = ~n66933 & n67452 ;
  assign n67454 = ~n66869 & ~n67453 ;
  assign n67455 = n67450 & ~n67454 ;
  assign n67456 = ~n66894 & ~n67455 ;
  assign n67462 = ~n66888 & n67092 ;
  assign n67461 = n66888 & ~n67099 ;
  assign n67463 = n66894 & ~n67461 ;
  assign n67464 = ~n67462 & n67463 ;
  assign n67459 = ~n66875 & ~n66895 ;
  assign n67460 = n66903 & n67459 ;
  assign n67457 = n66875 & ~n66909 ;
  assign n67458 = n67109 & n67457 ;
  assign n67465 = ~n66869 & ~n67458 ;
  assign n67466 = ~n67460 & n67465 ;
  assign n67467 = ~n67464 & n67466 ;
  assign n67468 = ~n66881 & n66924 ;
  assign n67469 = n66917 & ~n67468 ;
  assign n67470 = n66875 & n66903 ;
  assign n67471 = n66894 & ~n66932 ;
  assign n67472 = ~n67470 & n67471 ;
  assign n67473 = ~n67469 & ~n67472 ;
  assign n67474 = ~n66875 & n67451 ;
  assign n67475 = n66869 & n67450 ;
  assign n67476 = ~n67474 & n67475 ;
  assign n67477 = n66906 & n67476 ;
  assign n67478 = ~n67473 & n67477 ;
  assign n67479 = ~n67467 & ~n67478 ;
  assign n67480 = ~n67456 & ~n67479 ;
  assign n67481 = ~\u0_L3_reg[13]/NET0131  & n67480 ;
  assign n67482 = \u0_L3_reg[13]/NET0131  & ~n67480 ;
  assign n67483 = ~n67481 & ~n67482 ;
  assign n67484 = n66770 & ~n66845 ;
  assign n67487 = ~n66804 & ~n66811 ;
  assign n67485 = ~n66776 & ~n66789 ;
  assign n67486 = n66782 & n66796 ;
  assign n67488 = ~n67485 & ~n67486 ;
  assign n67489 = n67487 & n67488 ;
  assign n67490 = n67484 & ~n67489 ;
  assign n67491 = ~n66804 & n66844 ;
  assign n67492 = ~n66770 & ~n67491 ;
  assign n67493 = ~n66782 & n66811 ;
  assign n67494 = ~n66831 & ~n67493 ;
  assign n67495 = n67492 & n67494 ;
  assign n67496 = ~n67490 & ~n67495 ;
  assign n67497 = ~n66806 & n67240 ;
  assign n67498 = ~n67496 & n67497 ;
  assign n67499 = ~n66820 & ~n67486 ;
  assign n67500 = ~n66818 & n67499 ;
  assign n67501 = n67492 & n67500 ;
  assign n67502 = ~n66808 & ~n66840 ;
  assign n67503 = n67484 & n67502 ;
  assign n67504 = ~n67501 & ~n67503 ;
  assign n67505 = ~n66803 & ~n67220 ;
  assign n67506 = ~n66819 & n67505 ;
  assign n67507 = ~n66839 & n67506 ;
  assign n67508 = ~n67504 & n67507 ;
  assign n67509 = ~n67498 & ~n67508 ;
  assign n67510 = ~\u0_L3_reg[3]/NET0131  & n67509 ;
  assign n67511 = \u0_L3_reg[3]/NET0131  & ~n67509 ;
  assign n67512 = ~n67510 & ~n67511 ;
  assign n67513 = n67351 & n67364 ;
  assign n67514 = ~n67358 & n67513 ;
  assign n67515 = ~n67345 & n67514 ;
  assign n67516 = n67352 & n67364 ;
  assign n67517 = ~n67364 & n67382 ;
  assign n67518 = ~n67516 & ~n67517 ;
  assign n67519 = n67352 & n67358 ;
  assign n67520 = ~n67514 & ~n67519 ;
  assign n67521 = n67518 & n67520 ;
  assign n67522 = n67379 & ~n67521 ;
  assign n67523 = ~n67515 & ~n67522 ;
  assign n67524 = ~n67371 & ~n67523 ;
  assign n67533 = n67401 & n67409 ;
  assign n67535 = ~n67345 & n67351 ;
  assign n67536 = ~n67401 & ~n67535 ;
  assign n67537 = ~n67379 & ~n67536 ;
  assign n67534 = n67379 & ~n67401 ;
  assign n67538 = ~n67382 & ~n67534 ;
  assign n67539 = ~n67537 & n67538 ;
  assign n67540 = ~n67533 & ~n67539 ;
  assign n67541 = n67371 & ~n67540 ;
  assign n67525 = n67358 & n67513 ;
  assign n67526 = ~n67383 & ~n67525 ;
  assign n67527 = n67371 & ~n67526 ;
  assign n67528 = ~n67384 & ~n67389 ;
  assign n67529 = ~n67364 & ~n67405 ;
  assign n67530 = n67528 & n67529 ;
  assign n67531 = ~n67527 & ~n67530 ;
  assign n67532 = n67379 & ~n67531 ;
  assign n67542 = n67358 & n67405 ;
  assign n67543 = n67364 & ~n67379 ;
  assign n67544 = n67542 & n67543 ;
  assign n67545 = n67401 & ~n67406 ;
  assign n67546 = n67386 & ~n67545 ;
  assign n67547 = ~n67371 & ~n67379 ;
  assign n67548 = ~n67546 & n67547 ;
  assign n67549 = ~n67544 & ~n67548 ;
  assign n67550 = ~n67532 & n67549 ;
  assign n67551 = ~n67541 & n67550 ;
  assign n67552 = ~n67524 & n67551 ;
  assign n67553 = ~\u0_L3_reg[24]/NET0131  & ~n67552 ;
  assign n67554 = \u0_L3_reg[24]/NET0131  & n67552 ;
  assign n67555 = ~n67553 & ~n67554 ;
  assign n67556 = n67401 & n67535 ;
  assign n67557 = n67379 & ~n67556 ;
  assign n67558 = n67518 & n67557 ;
  assign n67559 = ~n67379 & ~n67513 ;
  assign n67560 = ~n67519 & n67559 ;
  assign n67561 = ~n67558 & ~n67560 ;
  assign n67562 = n67371 & ~n67561 ;
  assign n67565 = ~n67513 & n67528 ;
  assign n67566 = ~n67379 & ~n67565 ;
  assign n67568 = ~n67384 & n67513 ;
  assign n67567 = ~n67345 & n67395 ;
  assign n67569 = n67379 & ~n67567 ;
  assign n67570 = ~n67568 & n67569 ;
  assign n67571 = ~n67566 & ~n67570 ;
  assign n67563 = ~n67358 & n67382 ;
  assign n67564 = n67364 & n67563 ;
  assign n67572 = ~n67371 & ~n67545 ;
  assign n67573 = ~n67564 & n67572 ;
  assign n67574 = ~n67571 & n67573 ;
  assign n67575 = ~n67562 & ~n67574 ;
  assign n67578 = n67364 & n67379 ;
  assign n67579 = ~n67358 & n67405 ;
  assign n67580 = n67578 & n67579 ;
  assign n67576 = n67372 & ~n67405 ;
  assign n67577 = n67384 & n67543 ;
  assign n67581 = ~n67576 & ~n67577 ;
  assign n67582 = ~n67580 & n67581 ;
  assign n67583 = ~n67575 & n67582 ;
  assign n67584 = \u0_L3_reg[30]/NET0131  & ~n67583 ;
  assign n67585 = ~\u0_L3_reg[30]/NET0131  & n67583 ;
  assign n67586 = ~n67584 & ~n67585 ;
  assign n67602 = n66369 & ~n67205 ;
  assign n67590 = ~n66412 & n67202 ;
  assign n67601 = n66378 & n67590 ;
  assign n67603 = ~n67208 & ~n67601 ;
  assign n67604 = ~n67602 & n67603 ;
  assign n67605 = n66400 & ~n67604 ;
  assign n67591 = ~n66377 & n67590 ;
  assign n67587 = n66363 & n66419 ;
  assign n67588 = n66377 & ~n67202 ;
  assign n67589 = ~n67587 & n67588 ;
  assign n67592 = ~n66357 & ~n66412 ;
  assign n67593 = n66389 & ~n67592 ;
  assign n67594 = n66356 & n67587 ;
  assign n67595 = ~n67593 & ~n67594 ;
  assign n67596 = ~n67589 & n67595 ;
  assign n67597 = ~n67591 & n67596 ;
  assign n67598 = ~n66400 & ~n67597 ;
  assign n67599 = ~n66407 & ~n67594 ;
  assign n67600 = ~n66377 & ~n67599 ;
  assign n67606 = ~n67598 & ~n67600 ;
  assign n67607 = ~n67605 & n67606 ;
  assign n67608 = ~\u0_L3_reg[9]/NET0131  & ~n67607 ;
  assign n67609 = \u0_L3_reg[9]/NET0131  & n67607 ;
  assign n67610 = ~n67608 & ~n67609 ;
  assign n67611 = ~n67542 & ~n67563 ;
  assign n67627 = n67352 & ~n67364 ;
  assign n67628 = n67611 & ~n67627 ;
  assign n67629 = ~n67379 & ~n67628 ;
  assign n67630 = ~n67358 & ~n67405 ;
  assign n67631 = ~n67352 & n67379 ;
  assign n67632 = ~n67542 & n67631 ;
  assign n67633 = ~n67630 & n67632 ;
  assign n67634 = ~n67391 & ~n67633 ;
  assign n67635 = ~n67629 & n67634 ;
  assign n67636 = ~n67371 & ~n67635 ;
  assign n67612 = n67358 & ~n67403 ;
  assign n67613 = ~n67345 & ~n67389 ;
  assign n67614 = ~n67612 & n67613 ;
  assign n67615 = n67611 & ~n67614 ;
  assign n67616 = ~n67364 & ~n67615 ;
  assign n67617 = n67365 & n67382 ;
  assign n67618 = ~n67616 & ~n67617 ;
  assign n67619 = n67371 & ~n67618 ;
  assign n67620 = ~n67364 & n67535 ;
  assign n67621 = ~n67516 & ~n67620 ;
  assign n67622 = n67371 & ~n67621 ;
  assign n67623 = ~n67514 & ~n67622 ;
  assign n67624 = ~n67379 & ~n67623 ;
  assign n67625 = ~n67385 & ~n67390 ;
  assign n67626 = n67578 & ~n67625 ;
  assign n67637 = ~n67624 & ~n67626 ;
  assign n67638 = ~n67619 & n67637 ;
  assign n67639 = ~n67636 & n67638 ;
  assign n67640 = ~\u0_L3_reg[16]/NET0131  & ~n67639 ;
  assign n67641 = \u0_L3_reg[16]/NET0131  & n67639 ;
  assign n67642 = ~n67640 & ~n67641 ;
  assign n67655 = ~n66924 & ~n66935 ;
  assign n67657 = n66907 & ~n67655 ;
  assign n67651 = ~n66902 & ~n66941 ;
  assign n67656 = n67651 & n67655 ;
  assign n67658 = ~n66932 & ~n67091 ;
  assign n67659 = ~n67656 & n67658 ;
  assign n67660 = ~n67657 & n67659 ;
  assign n67661 = ~n66869 & ~n67660 ;
  assign n67648 = n66894 & n66911 ;
  assign n67649 = ~n66926 & ~n67648 ;
  assign n67650 = n66869 & ~n67649 ;
  assign n67643 = ~n66882 & ~n66931 ;
  assign n67644 = n66869 & n66902 ;
  assign n67645 = ~n67643 & n67644 ;
  assign n67646 = ~n66904 & ~n67645 ;
  assign n67647 = ~n66894 & ~n67646 ;
  assign n67652 = ~n66882 & n66894 ;
  assign n67653 = ~n67098 & n67652 ;
  assign n67654 = ~n67651 & n67653 ;
  assign n67662 = ~n67647 & ~n67654 ;
  assign n67663 = ~n67650 & n67662 ;
  assign n67664 = ~n67661 & n67663 ;
  assign n67665 = \u0_L3_reg[18]/NET0131  & n67664 ;
  assign n67666 = ~\u0_L3_reg[18]/NET0131  & ~n67664 ;
  assign n67667 = ~n67665 & ~n67666 ;
  assign n67695 = decrypt_pad & ~\u0_uk_K_r2_reg[53]/P0001  ;
  assign n67696 = ~decrypt_pad & ~\u0_uk_K_r2_reg[48]/NET0131  ;
  assign n67697 = ~n67695 & ~n67696 ;
  assign n67698 = \u0_R2_reg[4]/NET0131  & ~n67697 ;
  assign n67699 = ~\u0_R2_reg[4]/NET0131  & n67697 ;
  assign n67700 = ~n67698 & ~n67699 ;
  assign n67674 = decrypt_pad & ~\u0_uk_K_r2_reg[18]/NET0131  ;
  assign n67675 = ~decrypt_pad & ~\u0_uk_K_r2_reg[13]/NET0131  ;
  assign n67676 = ~n67674 & ~n67675 ;
  assign n67677 = \u0_R2_reg[3]/NET0131  & ~n67676 ;
  assign n67678 = ~\u0_R2_reg[3]/NET0131  & n67676 ;
  assign n67679 = ~n67677 & ~n67678 ;
  assign n67681 = decrypt_pad & ~\u0_uk_K_r2_reg[26]/NET0131  ;
  assign n67682 = ~decrypt_pad & ~\u0_uk_K_r2_reg[46]/NET0131  ;
  assign n67683 = ~n67681 & ~n67682 ;
  assign n67684 = \u0_R2_reg[1]/NET0131  & ~n67683 ;
  assign n67685 = ~\u0_R2_reg[1]/NET0131  & n67683 ;
  assign n67686 = ~n67684 & ~n67685 ;
  assign n67705 = decrypt_pad & ~\u0_uk_K_r2_reg[24]/NET0131  ;
  assign n67706 = ~decrypt_pad & ~\u0_uk_K_r2_reg[19]/NET0131  ;
  assign n67707 = ~n67705 & ~n67706 ;
  assign n67708 = \u0_R2_reg[5]/NET0131  & ~n67707 ;
  assign n67709 = ~\u0_R2_reg[5]/NET0131  & n67707 ;
  assign n67710 = ~n67708 & ~n67709 ;
  assign n67711 = ~n67686 & n67710 ;
  assign n67668 = decrypt_pad & ~\u0_uk_K_r2_reg[41]/NET0131  ;
  assign n67669 = ~decrypt_pad & ~\u0_uk_K_r2_reg[4]/NET0131  ;
  assign n67670 = ~n67668 & ~n67669 ;
  assign n67671 = \u0_R2_reg[2]/NET0131  & ~n67670 ;
  assign n67672 = ~\u0_R2_reg[2]/NET0131  & n67670 ;
  assign n67673 = ~n67671 & ~n67672 ;
  assign n67687 = decrypt_pad & ~\u0_uk_K_r2_reg[5]/NET0131  ;
  assign n67688 = ~decrypt_pad & ~\u0_uk_K_r2_reg[25]/NET0131  ;
  assign n67689 = ~n67687 & ~n67688 ;
  assign n67690 = \u0_R2_reg[32]/NET0131  & ~n67689 ;
  assign n67691 = ~\u0_R2_reg[32]/NET0131  & n67689 ;
  assign n67692 = ~n67690 & ~n67691 ;
  assign n67701 = n67673 & ~n67692 ;
  assign n67729 = n67701 & ~n67710 ;
  assign n67730 = ~n67711 & ~n67729 ;
  assign n67731 = n67679 & ~n67730 ;
  assign n67702 = ~n67673 & n67692 ;
  assign n67703 = ~n67701 & ~n67702 ;
  assign n67715 = n67692 & n67710 ;
  assign n67736 = ~n67686 & ~n67715 ;
  assign n67737 = ~n67703 & n67736 ;
  assign n67721 = ~n67679 & n67686 ;
  assign n67732 = n67692 & n67721 ;
  assign n67733 = ~n67692 & n67710 ;
  assign n67680 = ~n67673 & n67679 ;
  assign n67734 = ~n67680 & n67686 ;
  assign n67735 = n67733 & ~n67734 ;
  assign n67738 = ~n67732 & ~n67735 ;
  assign n67739 = ~n67737 & n67738 ;
  assign n67740 = ~n67731 & n67739 ;
  assign n67741 = n67700 & ~n67740 ;
  assign n67716 = ~n67692 & ~n67710 ;
  assign n67717 = ~n67715 & ~n67716 ;
  assign n67718 = n67686 & n67717 ;
  assign n67719 = n67679 & n67718 ;
  assign n67720 = n67673 & n67719 ;
  assign n67704 = n67673 & n67686 ;
  assign n67712 = ~n67679 & ~n67704 ;
  assign n67713 = ~n67711 & n67712 ;
  assign n67714 = n67703 & n67713 ;
  assign n67722 = n67715 & ~n67721 ;
  assign n67723 = n67686 & n67716 ;
  assign n67724 = ~n67722 & ~n67723 ;
  assign n67725 = ~n67673 & ~n67724 ;
  assign n67726 = ~n67714 & ~n67725 ;
  assign n67727 = ~n67720 & n67726 ;
  assign n67728 = ~n67700 & ~n67727 ;
  assign n67745 = n67686 & n67715 ;
  assign n67746 = n67673 & n67745 ;
  assign n67747 = ~n67673 & n67686 ;
  assign n67748 = ~n67710 & n67747 ;
  assign n67749 = n67701 & n67711 ;
  assign n67750 = ~n67748 & ~n67749 ;
  assign n67751 = ~n67746 & n67750 ;
  assign n67752 = ~n67679 & ~n67751 ;
  assign n67693 = ~n67686 & n67692 ;
  assign n67694 = n67680 & n67693 ;
  assign n67742 = ~n67686 & ~n67710 ;
  assign n67743 = n67679 & n67701 ;
  assign n67744 = n67742 & n67743 ;
  assign n67753 = ~n67694 & ~n67744 ;
  assign n67754 = ~n67752 & n67753 ;
  assign n67755 = ~n67728 & n67754 ;
  assign n67756 = ~n67741 & n67755 ;
  assign n67757 = ~\u0_L2_reg[31]/NET0131  & ~n67756 ;
  assign n67758 = \u0_L2_reg[31]/NET0131  & n67756 ;
  assign n67759 = ~n67757 & ~n67758 ;
  assign n67760 = decrypt_pad & ~\u0_uk_K_r2_reg[52]/NET0131  ;
  assign n67761 = ~decrypt_pad & ~\u0_uk_K_r2_reg[15]/NET0131  ;
  assign n67762 = ~n67760 & ~n67761 ;
  assign n67763 = \u0_R2_reg[24]/NET0131  & ~n67762 ;
  assign n67764 = ~\u0_R2_reg[24]/NET0131  & n67762 ;
  assign n67765 = ~n67763 & ~n67764 ;
  assign n67797 = decrypt_pad & ~\u0_uk_K_r2_reg[22]/NET0131  ;
  assign n67798 = ~decrypt_pad & ~\u0_uk_K_r2_reg[44]/NET0131  ;
  assign n67799 = ~n67797 & ~n67798 ;
  assign n67800 = \u0_R2_reg[23]/NET0131  & ~n67799 ;
  assign n67801 = ~\u0_R2_reg[23]/NET0131  & n67799 ;
  assign n67802 = ~n67800 & ~n67801 ;
  assign n67772 = decrypt_pad & ~\u0_uk_K_r2_reg[9]/NET0131  ;
  assign n67773 = ~decrypt_pad & ~\u0_uk_K_r2_reg[0]/NET0131  ;
  assign n67774 = ~n67772 & ~n67773 ;
  assign n67775 = \u0_R2_reg[22]/NET0131  & ~n67774 ;
  assign n67776 = ~\u0_R2_reg[22]/NET0131  & n67774 ;
  assign n67777 = ~n67775 & ~n67776 ;
  assign n67766 = decrypt_pad & ~\u0_uk_K_r2_reg[42]/NET0131  ;
  assign n67767 = ~decrypt_pad & ~\u0_uk_K_r2_reg[9]/NET0131  ;
  assign n67768 = ~n67766 & ~n67767 ;
  assign n67769 = \u0_R2_reg[21]/NET0131  & ~n67768 ;
  assign n67770 = ~\u0_R2_reg[21]/NET0131  & n67768 ;
  assign n67771 = ~n67769 & ~n67770 ;
  assign n67779 = decrypt_pad & ~\u0_uk_K_r2_reg[31]/NET0131  ;
  assign n67780 = ~decrypt_pad & ~\u0_uk_K_r2_reg[49]/NET0131  ;
  assign n67781 = ~n67779 & ~n67780 ;
  assign n67782 = \u0_R2_reg[20]/NET0131  & ~n67781 ;
  assign n67783 = ~\u0_R2_reg[20]/NET0131  & n67781 ;
  assign n67784 = ~n67782 & ~n67783 ;
  assign n67785 = decrypt_pad & ~\u0_uk_K_r2_reg[43]/NET0131  ;
  assign n67786 = ~decrypt_pad & ~\u0_uk_K_r2_reg[38]/NET0131  ;
  assign n67787 = ~n67785 & ~n67786 ;
  assign n67788 = \u0_R2_reg[25]/NET0131  & ~n67787 ;
  assign n67789 = ~\u0_R2_reg[25]/NET0131  & n67787 ;
  assign n67790 = ~n67788 & ~n67789 ;
  assign n67791 = n67784 & ~n67790 ;
  assign n67836 = ~n67771 & n67791 ;
  assign n67837 = ~n67777 & n67836 ;
  assign n67793 = n67771 & ~n67784 ;
  assign n67794 = n67777 & n67793 ;
  assign n67804 = n67784 & n67790 ;
  assign n67835 = n67771 & n67804 ;
  assign n67838 = ~n67794 & ~n67835 ;
  assign n67839 = ~n67837 & n67838 ;
  assign n67840 = n67802 & ~n67839 ;
  assign n67813 = ~n67777 & ~n67802 ;
  assign n67841 = n67804 & n67813 ;
  assign n67842 = ~n67771 & n67841 ;
  assign n67843 = n67771 & n67790 ;
  assign n67844 = ~n67777 & ~n67843 ;
  assign n67845 = ~n67802 & ~n67804 ;
  assign n67846 = ~n67794 & n67845 ;
  assign n67847 = ~n67844 & n67846 ;
  assign n67848 = ~n67842 & ~n67847 ;
  assign n67849 = ~n67840 & n67848 ;
  assign n67850 = n67765 & ~n67849 ;
  assign n67778 = n67771 & ~n67777 ;
  assign n67795 = n67778 & n67784 ;
  assign n67796 = ~n67794 & ~n67795 ;
  assign n67803 = ~n67796 & ~n67802 ;
  assign n67792 = n67778 & n67791 ;
  assign n67810 = ~n67771 & n67784 ;
  assign n67811 = n67777 & n67802 ;
  assign n67812 = n67810 & n67811 ;
  assign n67817 = ~n67792 & ~n67812 ;
  assign n67814 = n67791 & n67813 ;
  assign n67815 = ~n67777 & ~n67784 ;
  assign n67816 = n67802 & n67815 ;
  assign n67818 = ~n67814 & ~n67816 ;
  assign n67819 = n67817 & n67818 ;
  assign n67805 = n67777 & n67804 ;
  assign n67806 = ~n67771 & n67805 ;
  assign n67807 = ~n67784 & n67790 ;
  assign n67808 = ~n67771 & n67807 ;
  assign n67809 = n67802 & n67808 ;
  assign n67820 = ~n67806 & ~n67809 ;
  assign n67821 = n67819 & n67820 ;
  assign n67822 = ~n67803 & n67821 ;
  assign n67823 = ~n67765 & ~n67822 ;
  assign n67831 = n67771 & n67791 ;
  assign n67832 = ~n67802 & n67831 ;
  assign n67833 = ~n67809 & ~n67832 ;
  assign n67834 = ~n67777 & ~n67833 ;
  assign n67824 = ~n67771 & ~n67784 ;
  assign n67825 = ~n67790 & n67824 ;
  assign n67826 = n67813 & n67825 ;
  assign n67827 = ~n67790 & n67793 ;
  assign n67828 = ~n67777 & n67827 ;
  assign n67829 = ~n67805 & ~n67828 ;
  assign n67830 = n67802 & ~n67829 ;
  assign n67851 = ~n67826 & ~n67830 ;
  assign n67852 = ~n67834 & n67851 ;
  assign n67853 = ~n67823 & n67852 ;
  assign n67854 = ~n67850 & n67853 ;
  assign n67855 = \u0_L2_reg[11]/NET0131  & ~n67854 ;
  assign n67856 = ~\u0_L2_reg[11]/NET0131  & n67854 ;
  assign n67857 = ~n67855 & ~n67856 ;
  assign n67858 = decrypt_pad & ~\u0_uk_K_r2_reg[35]/NET0131  ;
  assign n67859 = ~decrypt_pad & ~\u0_uk_K_r2_reg[2]/NET0131  ;
  assign n67860 = ~n67858 & ~n67859 ;
  assign n67861 = \u0_R2_reg[26]/NET0131  & ~n67860 ;
  assign n67862 = ~\u0_R2_reg[26]/NET0131  & n67860 ;
  assign n67863 = ~n67861 & ~n67862 ;
  assign n67864 = decrypt_pad & ~\u0_uk_K_r2_reg[50]/NET0131  ;
  assign n67865 = ~decrypt_pad & ~\u0_uk_K_r2_reg[45]/NET0131  ;
  assign n67866 = ~n67864 & ~n67865 ;
  assign n67867 = \u0_R2_reg[25]/NET0131  & ~n67866 ;
  assign n67868 = ~\u0_R2_reg[25]/NET0131  & n67866 ;
  assign n67869 = ~n67867 & ~n67868 ;
  assign n67870 = n67863 & ~n67869 ;
  assign n67871 = decrypt_pad & ~\u0_uk_K_r2_reg[15]/NET0131  ;
  assign n67872 = ~decrypt_pad & ~\u0_uk_K_r2_reg[37]/NET0131  ;
  assign n67873 = ~n67871 & ~n67872 ;
  assign n67874 = \u0_R2_reg[24]/NET0131  & ~n67873 ;
  assign n67875 = ~\u0_R2_reg[24]/NET0131  & n67873 ;
  assign n67876 = ~n67874 & ~n67875 ;
  assign n67877 = decrypt_pad & ~\u0_uk_K_r2_reg[23]/NET0131  ;
  assign n67878 = ~decrypt_pad & ~\u0_uk_K_r2_reg[14]/NET0131  ;
  assign n67879 = ~n67877 & ~n67878 ;
  assign n67880 = \u0_R2_reg[29]/NET0131  & ~n67879 ;
  assign n67881 = ~\u0_R2_reg[29]/NET0131  & n67879 ;
  assign n67882 = ~n67880 & ~n67881 ;
  assign n67883 = ~n67876 & n67882 ;
  assign n67884 = n67870 & n67883 ;
  assign n67885 = ~n67876 & ~n67882 ;
  assign n67886 = n67863 & n67869 ;
  assign n67887 = n67885 & n67886 ;
  assign n67888 = ~n67884 & ~n67887 ;
  assign n67889 = ~n67869 & ~n67882 ;
  assign n67890 = n67869 & n67882 ;
  assign n67891 = ~n67863 & n67890 ;
  assign n67892 = ~n67870 & ~n67891 ;
  assign n67893 = decrypt_pad & ~\u0_uk_K_r2_reg[0]/NET0131  ;
  assign n67894 = ~decrypt_pad & ~\u0_uk_K_r2_reg[22]/NET0131  ;
  assign n67895 = ~n67893 & ~n67894 ;
  assign n67896 = \u0_R2_reg[28]/NET0131  & ~n67895 ;
  assign n67897 = ~\u0_R2_reg[28]/NET0131  & n67895 ;
  assign n67898 = ~n67896 & ~n67897 ;
  assign n67899 = ~n67892 & n67898 ;
  assign n67900 = ~n67889 & ~n67899 ;
  assign n67901 = n67876 & ~n67900 ;
  assign n67902 = n67888 & ~n67901 ;
  assign n67903 = decrypt_pad & ~\u0_uk_K_r2_reg[44]/NET0131  ;
  assign n67904 = ~decrypt_pad & ~\u0_uk_K_r2_reg[35]/NET0131  ;
  assign n67905 = ~n67903 & ~n67904 ;
  assign n67906 = \u0_R2_reg[27]/NET0131  & ~n67905 ;
  assign n67907 = ~\u0_R2_reg[27]/NET0131  & n67905 ;
  assign n67908 = ~n67906 & ~n67907 ;
  assign n67909 = ~n67902 & n67908 ;
  assign n67910 = ~n67869 & n67908 ;
  assign n67911 = ~n67863 & n67910 ;
  assign n67912 = ~n67863 & n67882 ;
  assign n67913 = ~n67870 & ~n67908 ;
  assign n67914 = ~n67912 & n67913 ;
  assign n67915 = ~n67911 & ~n67914 ;
  assign n67916 = n67876 & ~n67915 ;
  assign n67917 = ~n67876 & n67889 ;
  assign n67918 = n67863 & n67917 ;
  assign n67919 = ~n67908 & n67918 ;
  assign n67920 = ~n67863 & ~n67876 ;
  assign n67921 = n67863 & n67876 ;
  assign n67922 = ~n67920 & ~n67921 ;
  assign n67923 = n67882 & ~n67910 ;
  assign n67924 = ~n67922 & n67923 ;
  assign n67925 = ~n67919 & ~n67924 ;
  assign n67926 = ~n67916 & n67925 ;
  assign n67927 = ~n67898 & ~n67926 ;
  assign n67931 = n67876 & n67882 ;
  assign n67932 = ~n67863 & ~n67869 ;
  assign n67933 = n67931 & n67932 ;
  assign n67934 = n67869 & n67883 ;
  assign n67935 = ~n67933 & ~n67934 ;
  assign n67936 = ~n67908 & ~n67935 ;
  assign n67937 = n67889 & n67920 ;
  assign n67938 = ~n67884 & ~n67937 ;
  assign n67939 = ~n67936 & n67938 ;
  assign n67940 = n67898 & ~n67939 ;
  assign n67928 = n67869 & ~n67908 ;
  assign n67929 = ~n67922 & n67928 ;
  assign n67930 = ~n67882 & n67911 ;
  assign n67941 = ~n67929 & ~n67930 ;
  assign n67942 = ~n67940 & n67941 ;
  assign n67943 = ~n67927 & n67942 ;
  assign n67944 = ~n67909 & n67943 ;
  assign n67945 = ~\u0_L2_reg[22]/NET0131  & ~n67944 ;
  assign n67946 = \u0_L2_reg[22]/NET0131  & n67944 ;
  assign n67947 = ~n67945 & ~n67946 ;
  assign n67948 = decrypt_pad & ~\u0_uk_K_r2_reg[54]/NET0131  ;
  assign n67949 = ~decrypt_pad & ~\u0_uk_K_r2_reg[17]/NET0131  ;
  assign n67950 = ~n67948 & ~n67949 ;
  assign n67951 = \u0_R2_reg[8]/NET0131  & ~n67950 ;
  assign n67952 = ~\u0_R2_reg[8]/NET0131  & n67950 ;
  assign n67953 = ~n67951 & ~n67952 ;
  assign n67954 = decrypt_pad & ~\u0_uk_K_r2_reg[10]/NET0131  ;
  assign n67955 = ~decrypt_pad & ~\u0_uk_K_r2_reg[5]/NET0131  ;
  assign n67956 = ~n67954 & ~n67955 ;
  assign n67957 = \u0_R2_reg[4]/NET0131  & ~n67956 ;
  assign n67958 = ~\u0_R2_reg[4]/NET0131  & n67956 ;
  assign n67959 = ~n67957 & ~n67958 ;
  assign n67960 = decrypt_pad & ~\u0_uk_K_r2_reg[34]/NET0131  ;
  assign n67961 = ~decrypt_pad & ~\u0_uk_K_r2_reg[54]/NET0131  ;
  assign n67962 = ~n67960 & ~n67961 ;
  assign n67963 = \u0_R2_reg[9]/NET0131  & ~n67962 ;
  assign n67964 = ~\u0_R2_reg[9]/NET0131  & n67962 ;
  assign n67965 = ~n67963 & ~n67964 ;
  assign n67966 = ~n67959 & n67965 ;
  assign n67967 = decrypt_pad & ~\u0_uk_K_r2_reg[46]/NET0131  ;
  assign n67968 = ~decrypt_pad & ~\u0_uk_K_r2_reg[41]/NET0131  ;
  assign n67969 = ~n67967 & ~n67968 ;
  assign n67970 = \u0_R2_reg[5]/NET0131  & ~n67969 ;
  assign n67971 = ~\u0_R2_reg[5]/NET0131  & n67969 ;
  assign n67972 = ~n67970 & ~n67971 ;
  assign n67973 = n67966 & ~n67972 ;
  assign n67976 = decrypt_pad & ~\u0_uk_K_r2_reg[12]/NET0131  ;
  assign n67977 = ~decrypt_pad & ~\u0_uk_K_r2_reg[32]/NET0131  ;
  assign n67978 = ~n67976 & ~n67977 ;
  assign n67979 = \u0_R2_reg[6]/NET0131  & ~n67978 ;
  assign n67980 = ~\u0_R2_reg[6]/NET0131  & n67978 ;
  assign n67981 = ~n67979 & ~n67980 ;
  assign n67983 = n67959 & n67972 ;
  assign n67984 = n67959 & ~n67965 ;
  assign n67985 = ~n67983 & ~n67984 ;
  assign n67986 = n67981 & ~n67985 ;
  assign n67987 = ~n67973 & ~n67986 ;
  assign n67988 = decrypt_pad & ~\u0_uk_K_r2_reg[6]/NET0131  ;
  assign n67989 = ~decrypt_pad & ~\u0_uk_K_r2_reg[26]/NET0131  ;
  assign n67990 = ~n67988 & ~n67989 ;
  assign n67991 = \u0_R2_reg[7]/NET0131  & ~n67990 ;
  assign n67992 = ~\u0_R2_reg[7]/NET0131  & n67990 ;
  assign n67993 = ~n67991 & ~n67992 ;
  assign n67994 = ~n67987 & ~n67993 ;
  assign n67999 = n67966 & n67972 ;
  assign n68000 = n67981 & ~n67999 ;
  assign n68001 = ~n67972 & ~n67993 ;
  assign n68002 = n67965 & n68001 ;
  assign n68003 = ~n67981 & ~n68002 ;
  assign n68004 = ~n68000 & ~n68003 ;
  assign n67974 = ~n67965 & n67972 ;
  assign n67975 = ~n67973 & ~n67974 ;
  assign n67982 = ~n67975 & ~n67981 ;
  assign n67995 = n67959 & n67965 ;
  assign n67996 = ~n67972 & n67981 ;
  assign n67997 = n67995 & n67996 ;
  assign n67998 = n67993 & n67997 ;
  assign n68005 = ~n67982 & ~n67998 ;
  assign n68006 = ~n68004 & n68005 ;
  assign n68007 = ~n67994 & n68006 ;
  assign n68008 = ~n67953 & ~n68007 ;
  assign n68024 = ~n67959 & ~n67965 ;
  assign n68025 = ~n67997 & ~n68024 ;
  assign n68026 = n67953 & ~n68025 ;
  assign n68027 = n67966 & ~n67996 ;
  assign n68028 = ~n68026 & ~n68027 ;
  assign n68012 = n67972 & ~n67981 ;
  assign n68029 = ~n67993 & ~n68012 ;
  assign n68030 = ~n68028 & n68029 ;
  assign n68009 = ~n67959 & n67981 ;
  assign n68010 = ~n67965 & ~n67972 ;
  assign n68011 = n68009 & n68010 ;
  assign n68013 = n67959 & n68012 ;
  assign n68014 = ~n68011 & ~n68013 ;
  assign n68015 = n67993 & ~n68014 ;
  assign n68020 = n67965 & n68013 ;
  assign n68016 = ~n67972 & n67984 ;
  assign n68017 = ~n67981 & n68016 ;
  assign n68018 = n67972 & n67993 ;
  assign n68019 = ~n68009 & n68018 ;
  assign n68021 = ~n68017 & ~n68019 ;
  assign n68022 = ~n68020 & n68021 ;
  assign n68023 = n67953 & ~n68022 ;
  assign n68031 = ~n68015 & ~n68023 ;
  assign n68032 = ~n68030 & n68031 ;
  assign n68033 = ~n68008 & n68032 ;
  assign n68034 = \u0_L2_reg[2]/NET0131  & n68033 ;
  assign n68035 = ~\u0_L2_reg[2]/NET0131  & ~n68033 ;
  assign n68036 = ~n68034 & ~n68035 ;
  assign n68039 = ~n67686 & ~n67717 ;
  assign n68041 = n67673 & ~n68039 ;
  assign n68040 = ~n67716 & ~n68039 ;
  assign n68042 = ~n67679 & ~n68040 ;
  assign n68043 = ~n68041 & n68042 ;
  assign n68044 = n67692 & n67742 ;
  assign n68045 = ~n67745 & ~n68044 ;
  assign n68046 = n67679 & ~n68045 ;
  assign n68037 = n67704 & ~n67710 ;
  assign n68038 = n67692 & n68037 ;
  assign n68047 = ~n67749 & ~n68038 ;
  assign n68048 = ~n68046 & n68047 ;
  assign n68049 = ~n68043 & n68048 ;
  assign n68050 = ~n67700 & ~n68049 ;
  assign n68051 = ~n67673 & ~n67686 ;
  assign n68052 = ~n67692 & ~n68051 ;
  assign n68053 = n67715 & n68051 ;
  assign n68054 = ~n68052 & ~n68053 ;
  assign n68055 = n67679 & ~n68054 ;
  assign n68058 = n67692 & n67748 ;
  assign n68056 = ~n67679 & ~n67702 ;
  assign n68057 = ~n68052 & n68056 ;
  assign n68059 = n67704 & n67710 ;
  assign n68060 = ~n68057 & ~n68059 ;
  assign n68061 = ~n68058 & n68060 ;
  assign n68062 = ~n68055 & n68061 ;
  assign n68063 = n67700 & ~n68062 ;
  assign n68064 = n67710 & n67747 ;
  assign n68065 = ~n68037 & ~n68064 ;
  assign n68066 = n67679 & ~n67692 ;
  assign n68067 = ~n68065 & n68066 ;
  assign n68068 = ~n68063 & ~n68067 ;
  assign n68069 = ~n68050 & n68068 ;
  assign n68070 = ~\u0_L2_reg[17]/NET0131  & ~n68069 ;
  assign n68071 = \u0_L2_reg[17]/NET0131  & n68069 ;
  assign n68072 = ~n68070 & ~n68071 ;
  assign n68094 = ~n67835 & ~n67836 ;
  assign n68079 = ~n67777 & ~n67790 ;
  assign n68095 = ~n67827 & ~n68079 ;
  assign n68096 = ~n67778 & ~n68095 ;
  assign n68097 = n68094 & ~n68096 ;
  assign n68098 = n67802 & ~n68097 ;
  assign n68074 = n67777 & n67831 ;
  assign n68084 = ~n67777 & ~n67791 ;
  assign n68085 = ~n67824 & n68084 ;
  assign n68092 = ~n68074 & ~n68085 ;
  assign n68093 = ~n67802 & ~n68092 ;
  assign n68099 = n67777 & n67808 ;
  assign n68100 = ~n68093 & ~n68099 ;
  assign n68101 = ~n68098 & n68100 ;
  assign n68102 = ~n67765 & ~n68101 ;
  assign n68073 = n67790 & n67793 ;
  assign n68075 = n67771 & n67815 ;
  assign n68076 = ~n68073 & ~n68075 ;
  assign n68077 = ~n68074 & n68076 ;
  assign n68078 = n67802 & ~n68077 ;
  assign n68080 = ~n67771 & ~n68079 ;
  assign n68081 = n67802 & ~n68080 ;
  assign n68082 = ~n67791 & ~n67807 ;
  assign n68083 = n67777 & ~n68082 ;
  assign n68086 = ~n68081 & ~n68083 ;
  assign n68087 = ~n68085 & n68086 ;
  assign n68088 = ~n68078 & ~n68087 ;
  assign n68089 = n67765 & ~n68088 ;
  assign n68090 = ~n67777 & n67802 ;
  assign n68091 = n67843 & n68090 ;
  assign n68103 = ~n67837 & ~n68091 ;
  assign n68104 = ~n68089 & n68103 ;
  assign n68105 = ~n68102 & n68104 ;
  assign n68106 = \u0_L2_reg[29]/NET0131  & ~n68105 ;
  assign n68107 = ~\u0_L2_reg[29]/NET0131  & n68105 ;
  assign n68108 = ~n68106 & ~n68107 ;
  assign n68129 = ~n67827 & ~n68099 ;
  assign n68130 = ~n67802 & ~n68129 ;
  assign n68125 = ~n67777 & n67807 ;
  assign n68126 = ~n67831 & ~n68125 ;
  assign n68127 = ~n67806 & n68126 ;
  assign n68128 = n67802 & ~n68127 ;
  assign n68131 = ~n67837 & ~n67841 ;
  assign n68132 = ~n68128 & n68131 ;
  assign n68133 = ~n68130 & n68132 ;
  assign n68134 = ~n67765 & ~n68133 ;
  assign n68118 = n67778 & ~n67790 ;
  assign n68119 = ~n67815 & ~n68118 ;
  assign n68120 = ~n67802 & ~n68119 ;
  assign n68116 = n67804 & n68090 ;
  assign n68117 = n67777 & n67843 ;
  assign n68121 = ~n68116 & ~n68117 ;
  assign n68122 = ~n67828 & n68121 ;
  assign n68123 = ~n68120 & n68122 ;
  assign n68124 = n67765 & ~n68123 ;
  assign n68109 = n67777 & ~n68094 ;
  assign n68110 = ~n67784 & n68079 ;
  assign n68111 = ~n68109 & ~n68110 ;
  assign n68112 = ~n67802 & ~n68111 ;
  assign n68113 = ~n67825 & ~n68073 ;
  assign n68114 = ~n67831 & n68113 ;
  assign n68115 = n67811 & ~n68114 ;
  assign n68135 = ~n68112 & ~n68115 ;
  assign n68136 = ~n68124 & n68135 ;
  assign n68137 = ~n68134 & n68136 ;
  assign n68138 = ~\u0_L2_reg[4]/NET0131  & ~n68137 ;
  assign n68139 = \u0_L2_reg[4]/NET0131  & n68137 ;
  assign n68140 = ~n68138 & ~n68139 ;
  assign n68147 = decrypt_pad & ~\u0_uk_K_r2_reg[14]/NET0131  ;
  assign n68148 = ~decrypt_pad & ~\u0_uk_K_r2_reg[36]/NET0131  ;
  assign n68149 = ~n68147 & ~n68148 ;
  assign n68150 = \u0_R2_reg[31]/NET0131  & ~n68149 ;
  assign n68151 = ~\u0_R2_reg[31]/NET0131  & n68149 ;
  assign n68152 = ~n68150 & ~n68151 ;
  assign n68153 = decrypt_pad & ~\u0_uk_K_r2_reg[29]/NET0131  ;
  assign n68154 = ~decrypt_pad & ~\u0_uk_K_r2_reg[51]/NET0131  ;
  assign n68155 = ~n68153 & ~n68154 ;
  assign n68156 = \u0_R2_reg[28]/NET0131  & ~n68155 ;
  assign n68157 = ~\u0_R2_reg[28]/NET0131  & n68155 ;
  assign n68158 = ~n68156 & ~n68157 ;
  assign n68174 = decrypt_pad & ~\u0_uk_K_r2_reg[2]/NET0131  ;
  assign n68175 = ~decrypt_pad & ~\u0_uk_K_r2_reg[52]/NET0131  ;
  assign n68176 = ~n68174 & ~n68175 ;
  assign n68177 = \u0_R2_reg[30]/NET0131  & ~n68176 ;
  assign n68178 = ~\u0_R2_reg[30]/NET0131  & n68176 ;
  assign n68179 = ~n68177 & ~n68178 ;
  assign n68190 = n68158 & ~n68179 ;
  assign n68159 = decrypt_pad & ~\u0_uk_K_r2_reg[45]/NET0131  ;
  assign n68160 = ~decrypt_pad & ~\u0_uk_K_r2_reg[8]/NET0131  ;
  assign n68161 = ~n68159 & ~n68160 ;
  assign n68162 = \u0_R2_reg[1]/NET0131  & ~n68161 ;
  assign n68163 = ~\u0_R2_reg[1]/NET0131  & n68161 ;
  assign n68164 = ~n68162 & ~n68163 ;
  assign n68166 = decrypt_pad & ~\u0_uk_K_r2_reg[1]/NET0131  ;
  assign n68167 = ~decrypt_pad & ~\u0_uk_K_r2_reg[23]/NET0131  ;
  assign n68168 = ~n68166 & ~n68167 ;
  assign n68169 = \u0_R2_reg[29]/NET0131  & ~n68168 ;
  assign n68170 = ~\u0_R2_reg[29]/NET0131  & n68168 ;
  assign n68171 = ~n68169 & ~n68170 ;
  assign n68191 = ~n68164 & n68171 ;
  assign n68216 = ~n68190 & ~n68191 ;
  assign n68141 = decrypt_pad & ~\u0_uk_K_r2_reg[51]/NET0131  ;
  assign n68142 = ~decrypt_pad & ~\u0_uk_K_r2_reg[42]/NET0131  ;
  assign n68143 = ~n68141 & ~n68142 ;
  assign n68144 = \u0_R2_reg[32]/NET0131  & ~n68143 ;
  assign n68145 = ~\u0_R2_reg[32]/NET0131  & n68143 ;
  assign n68146 = ~n68144 & ~n68145 ;
  assign n68192 = n68190 & n68191 ;
  assign n68217 = n68146 & ~n68192 ;
  assign n68218 = ~n68216 & n68217 ;
  assign n68184 = ~n68158 & ~n68164 ;
  assign n68194 = n68171 & n68179 ;
  assign n68210 = n68184 & n68194 ;
  assign n68204 = ~n68171 & ~n68179 ;
  assign n68211 = n68164 & n68204 ;
  assign n68212 = n68158 & n68211 ;
  assign n68213 = ~n68210 & ~n68212 ;
  assign n68165 = ~n68158 & n68164 ;
  assign n68172 = n68165 & ~n68171 ;
  assign n68214 = n68172 & n68179 ;
  assign n68205 = ~n68158 & n68204 ;
  assign n68215 = ~n68164 & n68205 ;
  assign n68219 = ~n68214 & ~n68215 ;
  assign n68220 = n68213 & n68219 ;
  assign n68221 = ~n68218 & n68220 ;
  assign n68222 = n68152 & ~n68221 ;
  assign n68173 = n68158 & ~n68171 ;
  assign n68180 = n68173 & n68179 ;
  assign n68181 = ~n68164 & n68180 ;
  assign n68182 = n68152 & ~n68172 ;
  assign n68183 = ~n68181 & n68182 ;
  assign n68185 = n68179 & n68184 ;
  assign n68186 = n68164 & n68171 ;
  assign n68187 = ~n68152 & ~n68186 ;
  assign n68188 = ~n68185 & n68187 ;
  assign n68189 = ~n68183 & ~n68188 ;
  assign n68195 = n68158 & n68164 ;
  assign n68196 = n68194 & n68195 ;
  assign n68193 = ~n68152 & n68190 ;
  assign n68197 = ~n68192 & ~n68193 ;
  assign n68198 = ~n68196 & n68197 ;
  assign n68199 = ~n68189 & n68198 ;
  assign n68200 = ~n68146 & ~n68199 ;
  assign n68201 = ~n68152 & n68192 ;
  assign n68202 = n68165 & n68194 ;
  assign n68206 = ~n68180 & ~n68202 ;
  assign n68207 = ~n68205 & n68206 ;
  assign n68203 = n68152 & ~n68202 ;
  assign n68208 = n68146 & ~n68203 ;
  assign n68209 = ~n68207 & n68208 ;
  assign n68223 = ~n68201 & ~n68209 ;
  assign n68224 = ~n68200 & n68223 ;
  assign n68225 = ~n68222 & n68224 ;
  assign n68226 = \u0_L2_reg[5]/NET0131  & ~n68225 ;
  assign n68227 = ~\u0_L2_reg[5]/NET0131  & n68225 ;
  assign n68228 = ~n68226 & ~n68227 ;
  assign n68229 = decrypt_pad & ~\u0_uk_K_r2_reg[55]/NET0131  ;
  assign n68230 = ~decrypt_pad & ~\u0_uk_K_r2_reg[18]/NET0131  ;
  assign n68231 = ~n68229 & ~n68230 ;
  assign n68232 = \u0_R2_reg[16]/NET0131  & ~n68231 ;
  assign n68233 = ~\u0_R2_reg[16]/NET0131  & n68231 ;
  assign n68234 = ~n68232 & ~n68233 ;
  assign n68248 = decrypt_pad & ~\u0_uk_K_r2_reg[19]/NET0131  ;
  assign n68249 = ~decrypt_pad & ~\u0_uk_K_r2_reg[39]/NET0131  ;
  assign n68250 = ~n68248 & ~n68249 ;
  assign n68251 = \u0_R2_reg[12]/NET0131  & ~n68250 ;
  assign n68252 = ~\u0_R2_reg[12]/NET0131  & n68250 ;
  assign n68253 = ~n68251 & ~n68252 ;
  assign n68235 = decrypt_pad & ~\u0_uk_K_r2_reg[47]/NET0131  ;
  assign n68236 = ~decrypt_pad & ~\u0_uk_K_r2_reg[10]/NET0131  ;
  assign n68237 = ~n68235 & ~n68236 ;
  assign n68238 = \u0_R2_reg[15]/NET0131  & ~n68237 ;
  assign n68239 = ~\u0_R2_reg[15]/NET0131  & n68237 ;
  assign n68240 = ~n68238 & ~n68239 ;
  assign n68241 = decrypt_pad & ~\u0_uk_K_r2_reg[13]/NET0131  ;
  assign n68242 = ~decrypt_pad & ~\u0_uk_K_r2_reg[33]/NET0131  ;
  assign n68243 = ~n68241 & ~n68242 ;
  assign n68244 = \u0_R2_reg[13]/NET0131  & ~n68243 ;
  assign n68245 = ~\u0_R2_reg[13]/NET0131  & n68243 ;
  assign n68246 = ~n68244 & ~n68245 ;
  assign n68247 = n68240 & n68246 ;
  assign n68262 = decrypt_pad & ~\u0_uk_K_r2_reg[39]/NET0131  ;
  assign n68263 = ~decrypt_pad & ~\u0_uk_K_r2_reg[34]/NET0131  ;
  assign n68264 = ~n68262 & ~n68263 ;
  assign n68265 = \u0_R2_reg[14]/NET0131  & ~n68264 ;
  assign n68266 = ~\u0_R2_reg[14]/NET0131  & n68264 ;
  assign n68267 = ~n68265 & ~n68266 ;
  assign n68304 = n68247 & n68267 ;
  assign n68305 = ~n68253 & n68304 ;
  assign n68254 = decrypt_pad & ~\u0_uk_K_r2_reg[3]/NET0131  ;
  assign n68255 = ~decrypt_pad & ~\u0_uk_K_r2_reg[55]/NET0131  ;
  assign n68256 = ~n68254 & ~n68255 ;
  assign n68257 = \u0_R2_reg[17]/NET0131  & ~n68256 ;
  assign n68258 = ~\u0_R2_reg[17]/NET0131  & n68256 ;
  assign n68259 = ~n68257 & ~n68258 ;
  assign n68291 = ~n68253 & ~n68259 ;
  assign n68294 = ~n68246 & n68291 ;
  assign n68301 = n68240 & n68294 ;
  assign n68272 = n68253 & n68259 ;
  assign n68275 = ~n68246 & ~n68267 ;
  assign n68302 = ~n68247 & ~n68275 ;
  assign n68303 = n68272 & ~n68302 ;
  assign n68306 = ~n68301 & ~n68303 ;
  assign n68307 = ~n68305 & n68306 ;
  assign n68292 = n68246 & n68291 ;
  assign n68293 = n68267 & n68292 ;
  assign n68295 = ~n68267 & n68294 ;
  assign n68296 = ~n68293 & ~n68295 ;
  assign n68260 = n68253 & ~n68259 ;
  assign n68297 = n68260 & n68267 ;
  assign n68298 = ~n68246 & n68259 ;
  assign n68299 = ~n68297 & ~n68298 ;
  assign n68300 = ~n68240 & ~n68299 ;
  assign n68308 = n68296 & ~n68300 ;
  assign n68309 = n68307 & n68308 ;
  assign n68310 = ~n68234 & ~n68309 ;
  assign n68268 = n68246 & ~n68267 ;
  assign n68269 = ~n68253 & n68268 ;
  assign n68276 = n68253 & n68275 ;
  assign n68277 = ~n68269 & ~n68276 ;
  assign n68278 = ~n68246 & n68267 ;
  assign n68279 = ~n68253 & n68278 ;
  assign n68280 = ~n68259 & n68279 ;
  assign n68281 = n68277 & ~n68280 ;
  assign n68282 = ~n68240 & ~n68281 ;
  assign n68261 = n68247 & n68260 ;
  assign n68270 = n68259 & n68269 ;
  assign n68271 = ~n68261 & ~n68270 ;
  assign n68273 = n68267 & n68272 ;
  assign n68274 = n68246 & n68273 ;
  assign n68283 = ~n68253 & n68259 ;
  assign n68284 = n68240 & n68283 ;
  assign n68285 = ~n68246 & n68284 ;
  assign n68286 = ~n68274 & ~n68285 ;
  assign n68287 = n68271 & n68286 ;
  assign n68288 = ~n68282 & n68287 ;
  assign n68289 = n68234 & ~n68288 ;
  assign n68311 = n68260 & n68278 ;
  assign n68312 = ~n68295 & ~n68311 ;
  assign n68313 = n68240 & ~n68312 ;
  assign n68290 = n68261 & ~n68267 ;
  assign n68314 = ~n68240 & n68270 ;
  assign n68315 = ~n68290 & ~n68314 ;
  assign n68316 = ~n68313 & n68315 ;
  assign n68317 = ~n68289 & n68316 ;
  assign n68318 = ~n68310 & n68317 ;
  assign n68319 = ~\u0_L2_reg[20]/NET0131  & ~n68318 ;
  assign n68320 = \u0_L2_reg[20]/NET0131  & n68318 ;
  assign n68321 = ~n68319 & ~n68320 ;
  assign n68327 = ~n67966 & ~n67984 ;
  assign n68333 = ~n67959 & ~n67981 ;
  assign n68345 = n67972 & ~n68333 ;
  assign n68346 = n68327 & n68345 ;
  assign n68347 = ~n68016 & ~n68346 ;
  assign n68348 = n67993 & ~n68347 ;
  assign n68334 = ~n67965 & n68333 ;
  assign n68335 = ~n67999 & ~n68334 ;
  assign n68349 = ~n67993 & ~n68335 ;
  assign n68341 = ~n67972 & n67995 ;
  assign n68342 = n67959 & n67993 ;
  assign n68343 = ~n68341 & ~n68342 ;
  assign n68344 = ~n67981 & ~n68343 ;
  assign n68350 = n67966 & n67996 ;
  assign n68351 = ~n68344 & ~n68350 ;
  assign n68352 = ~n68349 & n68351 ;
  assign n68353 = ~n68348 & n68352 ;
  assign n68354 = n67953 & ~n68353 ;
  assign n68322 = ~n67965 & n67981 ;
  assign n68323 = n67983 & n68322 ;
  assign n68324 = ~n67959 & n67996 ;
  assign n68325 = ~n68323 & ~n68324 ;
  assign n68326 = ~n67993 & ~n68325 ;
  assign n68329 = ~n67981 & n67984 ;
  assign n68330 = ~n67973 & ~n67983 ;
  assign n68331 = ~n68329 & n68330 ;
  assign n68332 = ~n67993 & ~n68331 ;
  assign n68336 = n67993 & ~n68335 ;
  assign n68328 = n67996 & n68327 ;
  assign n68337 = ~n68323 & ~n68328 ;
  assign n68338 = ~n68336 & n68337 ;
  assign n68339 = ~n68332 & n68338 ;
  assign n68340 = ~n67953 & ~n68339 ;
  assign n68355 = ~n68326 & ~n68340 ;
  assign n68356 = ~n68354 & n68355 ;
  assign n68357 = ~\u0_L2_reg[28]/NET0131  & ~n68356 ;
  assign n68358 = \u0_L2_reg[28]/NET0131  & n68356 ;
  assign n68359 = ~n68357 & ~n68358 ;
  assign n68360 = n68246 & n68297 ;
  assign n68361 = ~n68240 & ~n68280 ;
  assign n68362 = ~n68360 & n68361 ;
  assign n68365 = ~n68276 & ~n68298 ;
  assign n68366 = n68234 & ~n68365 ;
  assign n68363 = n68278 & n68283 ;
  assign n68364 = ~n68274 & ~n68363 ;
  assign n68367 = n68240 & ~n68293 ;
  assign n68368 = n68364 & n68367 ;
  assign n68369 = ~n68366 & n68368 ;
  assign n68370 = ~n68362 & ~n68369 ;
  assign n68371 = n68246 & n68283 ;
  assign n68372 = ~n68268 & ~n68371 ;
  assign n68373 = ~n68240 & ~n68260 ;
  assign n68374 = ~n68372 & n68373 ;
  assign n68375 = n68234 & ~n68279 ;
  assign n68376 = ~n68360 & n68375 ;
  assign n68377 = ~n68374 & n68376 ;
  assign n68381 = ~n68267 & n68291 ;
  assign n68382 = n68240 & ~n68311 ;
  assign n68383 = ~n68381 & n68382 ;
  assign n68384 = n68253 & n68298 ;
  assign n68378 = n68260 & ~n68267 ;
  assign n68385 = ~n68240 & ~n68378 ;
  assign n68386 = ~n68384 & n68385 ;
  assign n68387 = ~n68383 & ~n68386 ;
  assign n68379 = ~n68273 & ~n68378 ;
  assign n68380 = n68246 & ~n68379 ;
  assign n68388 = ~n68234 & ~n68270 ;
  assign n68389 = ~n68380 & n68388 ;
  assign n68390 = ~n68387 & n68389 ;
  assign n68391 = ~n68377 & ~n68390 ;
  assign n68392 = ~n68370 & ~n68391 ;
  assign n68393 = ~\u0_L2_reg[1]/NET0131  & ~n68392 ;
  assign n68394 = \u0_L2_reg[1]/NET0131  & n68392 ;
  assign n68395 = ~n68393 & ~n68394 ;
  assign n68412 = n68260 & ~n68268 ;
  assign n68413 = ~n68270 & ~n68412 ;
  assign n68414 = ~n68240 & ~n68413 ;
  assign n68409 = n68259 & n68276 ;
  assign n68410 = ~n68292 & ~n68409 ;
  assign n68411 = n68240 & ~n68410 ;
  assign n68415 = n68364 & ~n68411 ;
  assign n68416 = ~n68414 & n68415 ;
  assign n68417 = n68234 & ~n68416 ;
  assign n68397 = ~n68246 & ~n68259 ;
  assign n68398 = ~n68278 & ~n68397 ;
  assign n68399 = n68240 & ~n68398 ;
  assign n68400 = ~n68268 & ~n68399 ;
  assign n68401 = n68253 & ~n68400 ;
  assign n68402 = ~n68240 & n68272 ;
  assign n68403 = ~n68284 & ~n68402 ;
  assign n68404 = ~n68267 & ~n68403 ;
  assign n68396 = ~n68240 & n68294 ;
  assign n68405 = n68296 & ~n68396 ;
  assign n68406 = ~n68404 & n68405 ;
  assign n68407 = ~n68401 & n68406 ;
  assign n68408 = ~n68234 & ~n68407 ;
  assign n68418 = ~n68295 & n68364 ;
  assign n68419 = ~n68240 & ~n68418 ;
  assign n68420 = ~n68290 & ~n68305 ;
  assign n68421 = ~n68419 & n68420 ;
  assign n68422 = ~n68408 & n68421 ;
  assign n68423 = ~n68417 & n68422 ;
  assign n68424 = ~\u0_L2_reg[10]/NET0131  & ~n68423 ;
  assign n68425 = \u0_L2_reg[10]/NET0131  & n68423 ;
  assign n68426 = ~n68424 & ~n68425 ;
  assign n68486 = decrypt_pad & ~\u0_uk_K_r2_reg[36]/NET0131  ;
  assign n68487 = ~decrypt_pad & ~\u0_uk_K_r2_reg[31]/NET0131  ;
  assign n68488 = ~n68486 & ~n68487 ;
  assign n68489 = \u0_R2_reg[20]/NET0131  & ~n68488 ;
  assign n68490 = ~\u0_R2_reg[20]/NET0131  & n68488 ;
  assign n68491 = ~n68489 & ~n68490 ;
  assign n68427 = decrypt_pad & ~\u0_uk_K_r2_reg[21]/NET0131  ;
  assign n68428 = ~decrypt_pad & ~\u0_uk_K_r2_reg[43]/NET0131  ;
  assign n68429 = ~n68427 & ~n68428 ;
  assign n68430 = \u0_R2_reg[19]/NET0131  & ~n68429 ;
  assign n68431 = ~\u0_R2_reg[19]/NET0131  & n68429 ;
  assign n68432 = ~n68430 & ~n68431 ;
  assign n68446 = decrypt_pad & ~\u0_uk_K_r2_reg[49]/NET0131  ;
  assign n68447 = ~decrypt_pad & ~\u0_uk_K_r2_reg[16]/NET0131  ;
  assign n68448 = ~n68446 & ~n68447 ;
  assign n68449 = \u0_R2_reg[16]/NET0131  & ~n68448 ;
  assign n68450 = ~\u0_R2_reg[16]/NET0131  & n68448 ;
  assign n68451 = ~n68449 & ~n68450 ;
  assign n68439 = decrypt_pad & ~\u0_uk_K_r2_reg[16]/NET0131  ;
  assign n68440 = ~decrypt_pad & ~\u0_uk_K_r2_reg[7]/NET0131  ;
  assign n68441 = ~n68439 & ~n68440 ;
  assign n68442 = \u0_R2_reg[17]/NET0131  & ~n68441 ;
  assign n68443 = ~\u0_R2_reg[17]/NET0131  & n68441 ;
  assign n68444 = ~n68442 & ~n68443 ;
  assign n68453 = decrypt_pad & ~\u0_uk_K_r2_reg[37]/NET0131  ;
  assign n68454 = ~decrypt_pad & ~\u0_uk_K_r2_reg[28]/NET0131  ;
  assign n68455 = ~n68453 & ~n68454 ;
  assign n68456 = \u0_R2_reg[21]/NET0131  & ~n68455 ;
  assign n68457 = ~\u0_R2_reg[21]/NET0131  & n68455 ;
  assign n68458 = ~n68456 & ~n68457 ;
  assign n68462 = n68444 & ~n68458 ;
  assign n68493 = n68451 & n68462 ;
  assign n68433 = decrypt_pad & ~\u0_uk_K_r2_reg[38]/NET0131  ;
  assign n68434 = ~decrypt_pad & ~\u0_uk_K_r2_reg[1]/NET0131  ;
  assign n68435 = ~n68433 & ~n68434 ;
  assign n68436 = \u0_R2_reg[18]/NET0131  & ~n68435 ;
  assign n68437 = ~\u0_R2_reg[18]/NET0131  & n68435 ;
  assign n68438 = ~n68436 & ~n68437 ;
  assign n68445 = ~n68438 & n68444 ;
  assign n68452 = n68445 & ~n68451 ;
  assign n68460 = n68438 & n68451 ;
  assign n68461 = n68458 & ~n68460 ;
  assign n68504 = ~n68452 & n68461 ;
  assign n68505 = ~n68493 & ~n68504 ;
  assign n68506 = n68432 & ~n68505 ;
  assign n68495 = ~n68432 & ~n68438 ;
  assign n68467 = ~n68451 & n68458 ;
  assign n68496 = n68444 & n68467 ;
  assign n68481 = ~n68444 & ~n68451 ;
  assign n68497 = ~n68458 & n68481 ;
  assign n68498 = ~n68496 & ~n68497 ;
  assign n68499 = n68495 & ~n68498 ;
  assign n68459 = n68451 & ~n68458 ;
  assign n68471 = ~n68444 & n68459 ;
  assign n68507 = n68438 & n68471 ;
  assign n68494 = ~n68438 & n68493 ;
  assign n68500 = ~n68432 & n68444 ;
  assign n68501 = n68438 & ~n68500 ;
  assign n68473 = n68451 & n68458 ;
  assign n68502 = ~n68445 & n68473 ;
  assign n68503 = ~n68501 & n68502 ;
  assign n68508 = ~n68494 & ~n68503 ;
  assign n68509 = ~n68507 & n68508 ;
  assign n68510 = ~n68499 & n68509 ;
  assign n68511 = ~n68506 & n68510 ;
  assign n68512 = n68491 & ~n68511 ;
  assign n68472 = ~n68438 & n68471 ;
  assign n68474 = n68445 & n68473 ;
  assign n68468 = ~n68444 & n68467 ;
  assign n68469 = n68438 & n68444 ;
  assign n68470 = ~n68458 & n68469 ;
  assign n68475 = ~n68468 & ~n68470 ;
  assign n68476 = ~n68474 & n68475 ;
  assign n68477 = ~n68472 & n68476 ;
  assign n68478 = ~n68432 & ~n68477 ;
  assign n68463 = ~n68459 & ~n68462 ;
  assign n68464 = ~n68461 & n68463 ;
  assign n68465 = ~n68452 & ~n68464 ;
  assign n68466 = n68432 & ~n68465 ;
  assign n68479 = ~n68438 & n68458 ;
  assign n68480 = ~n68459 & ~n68479 ;
  assign n68482 = ~n68469 & ~n68481 ;
  assign n68483 = n68480 & n68482 ;
  assign n68484 = ~n68466 & ~n68483 ;
  assign n68485 = ~n68478 & n68484 ;
  assign n68492 = ~n68485 & ~n68491 ;
  assign n68513 = ~n68451 & n68462 ;
  assign n68514 = ~n68468 & ~n68513 ;
  assign n68515 = n68438 & ~n68514 ;
  assign n68516 = ~n68432 & n68515 ;
  assign n68517 = n68438 & n68497 ;
  assign n68518 = ~n68494 & ~n68517 ;
  assign n68519 = n68432 & ~n68518 ;
  assign n68520 = ~n68516 & ~n68519 ;
  assign n68521 = ~n68492 & n68520 ;
  assign n68522 = ~n68512 & n68521 ;
  assign n68523 = ~\u0_L2_reg[14]/NET0131  & ~n68522 ;
  assign n68524 = \u0_L2_reg[14]/NET0131  & n68522 ;
  assign n68525 = ~n68523 & ~n68524 ;
  assign n68529 = ~n67981 & n68010 ;
  assign n68530 = n67965 & n68009 ;
  assign n68531 = ~n68529 & ~n68530 ;
  assign n68532 = n67993 & ~n68531 ;
  assign n68527 = ~n67995 & ~n68322 ;
  assign n68528 = n68001 & ~n68527 ;
  assign n68526 = n67974 & n68333 ;
  assign n68533 = n67953 & ~n68526 ;
  assign n68534 = ~n68528 & n68533 ;
  assign n68535 = ~n68004 & n68534 ;
  assign n68536 = ~n68532 & n68535 ;
  assign n68539 = n67965 & ~n68001 ;
  assign n68540 = n68333 & n68539 ;
  assign n68537 = ~n67974 & n67981 ;
  assign n68538 = n68342 & n68537 ;
  assign n68541 = ~n67953 & ~n68538 ;
  assign n68542 = ~n68540 & n68541 ;
  assign n68543 = n67972 & n68024 ;
  assign n68544 = ~n67993 & ~n68350 ;
  assign n68545 = ~n68543 & n68544 ;
  assign n68546 = ~n68017 & n68545 ;
  assign n68547 = n68542 & n68546 ;
  assign n68548 = ~n68536 & ~n68547 ;
  assign n68549 = ~n68020 & ~n68323 ;
  assign n68550 = ~n68548 & n68549 ;
  assign n68551 = n67972 & ~n68329 ;
  assign n68552 = ~n67973 & ~n68016 ;
  assign n68553 = ~n68551 & n68552 ;
  assign n68554 = n67993 & ~n68553 ;
  assign n68555 = n68542 & n68554 ;
  assign n68556 = ~n68550 & ~n68555 ;
  assign n68557 = ~\u0_L2_reg[13]/NET0131  & ~n68556 ;
  assign n68558 = \u0_L2_reg[13]/NET0131  & n68556 ;
  assign n68559 = ~n68557 & ~n68558 ;
  assign n68560 = n68158 & n68171 ;
  assign n68561 = ~n68179 & n68191 ;
  assign n68562 = ~n68560 & ~n68561 ;
  assign n68563 = ~n68172 & n68562 ;
  assign n68564 = n68152 & ~n68563 ;
  assign n68565 = n68158 & ~n68164 ;
  assign n68566 = ~n68179 & n68565 ;
  assign n68567 = ~n68171 & n68566 ;
  assign n68568 = ~n68564 & ~n68567 ;
  assign n68569 = ~n68146 & ~n68568 ;
  assign n68570 = n68164 & n68205 ;
  assign n68571 = n68203 & ~n68570 ;
  assign n68576 = ~n68152 & ~n68210 ;
  assign n68572 = n68171 & ~n68179 ;
  assign n68573 = n68165 & n68572 ;
  assign n68574 = n68146 & ~n68179 ;
  assign n68575 = n68173 & ~n68574 ;
  assign n68577 = ~n68573 & ~n68575 ;
  assign n68578 = n68576 & n68577 ;
  assign n68579 = ~n68215 & n68578 ;
  assign n68580 = ~n68571 & ~n68579 ;
  assign n68584 = ~n68152 & n68179 ;
  assign n68585 = ~n68184 & ~n68584 ;
  assign n68583 = ~n68152 & ~n68164 ;
  assign n68586 = ~n68171 & ~n68583 ;
  assign n68587 = ~n68585 & n68586 ;
  assign n68582 = n68164 & n68180 ;
  assign n68581 = n68158 & n68572 ;
  assign n68588 = ~n68210 & ~n68581 ;
  assign n68589 = ~n68582 & n68588 ;
  assign n68590 = ~n68587 & n68589 ;
  assign n68591 = n68146 & ~n68590 ;
  assign n68592 = ~n68580 & ~n68591 ;
  assign n68593 = ~n68569 & n68592 ;
  assign n68594 = \u0_L2_reg[15]/P0001  & n68593 ;
  assign n68595 = ~\u0_L2_reg[15]/P0001  & ~n68593 ;
  assign n68596 = ~n68594 & ~n68595 ;
  assign n68597 = ~n68152 & ~n68566 ;
  assign n68598 = ~n68582 & n68597 ;
  assign n68599 = n68171 & ~n68184 ;
  assign n68600 = ~n68190 & n68599 ;
  assign n68601 = n68152 & ~n68211 ;
  assign n68602 = ~n68600 & n68601 ;
  assign n68603 = ~n68598 & ~n68602 ;
  assign n68604 = ~n68164 & ~n68171 ;
  assign n68605 = ~n68565 & ~n68604 ;
  assign n68606 = ~n68173 & n68179 ;
  assign n68607 = ~n68605 & n68606 ;
  assign n68608 = n68146 & ~n68570 ;
  assign n68609 = ~n68607 & n68608 ;
  assign n68610 = ~n68603 & n68609 ;
  assign n68623 = ~n68181 & ~n68215 ;
  assign n68611 = n68164 & n68193 ;
  assign n68618 = n68152 & n68158 ;
  assign n68619 = ~n68186 & n68618 ;
  assign n68620 = ~n68204 & n68619 ;
  assign n68624 = ~n68611 & ~n68620 ;
  assign n68625 = n68623 & n68624 ;
  assign n68612 = ~n68158 & n68171 ;
  assign n68614 = ~n68152 & n68165 ;
  assign n68615 = ~n68612 & ~n68614 ;
  assign n68616 = n68179 & ~n68615 ;
  assign n68617 = n68195 & n68572 ;
  assign n68613 = n68583 & n68612 ;
  assign n68621 = ~n68146 & ~n68613 ;
  assign n68622 = ~n68617 & n68621 ;
  assign n68626 = ~n68616 & n68622 ;
  assign n68627 = n68625 & n68626 ;
  assign n68628 = ~n68610 & ~n68627 ;
  assign n68629 = n68152 & n68205 ;
  assign n68630 = ~n68152 & n68617 ;
  assign n68631 = ~n68629 & ~n68630 ;
  assign n68632 = ~n68628 & n68631 ;
  assign n68633 = ~\u0_L2_reg[21]/NET0131  & ~n68632 ;
  assign n68634 = \u0_L2_reg[21]/NET0131  & n68632 ;
  assign n68635 = ~n68633 & ~n68634 ;
  assign n68636 = n67673 & n68044 ;
  assign n68637 = ~n67711 & ~n67723 ;
  assign n68638 = ~n67692 & ~n68637 ;
  assign n68639 = ~n68636 & ~n68638 ;
  assign n68640 = ~n67679 & ~n68639 ;
  assign n68641 = ~n67702 & n67719 ;
  assign n68642 = ~n67744 & ~n68053 ;
  assign n68643 = ~n68641 & n68642 ;
  assign n68644 = ~n68640 & n68643 ;
  assign n68645 = n67700 & ~n68644 ;
  assign n68647 = ~n67704 & ~n67743 ;
  assign n68648 = n67710 & ~n68647 ;
  assign n68650 = ~n67679 & n67692 ;
  assign n68651 = ~n67742 & n68650 ;
  assign n68652 = ~n68051 & n68651 ;
  assign n68646 = ~n67710 & n68051 ;
  assign n68649 = n67679 & n67723 ;
  assign n68653 = ~n68646 & ~n68649 ;
  assign n68654 = ~n68652 & n68653 ;
  assign n68655 = ~n68648 & n68654 ;
  assign n68656 = ~n67700 & ~n68655 ;
  assign n68657 = ~n67693 & ~n67723 ;
  assign n68658 = n67680 & ~n68657 ;
  assign n68659 = n67733 & n68051 ;
  assign n68660 = ~n67746 & ~n68659 ;
  assign n68661 = ~n68058 & n68660 ;
  assign n68662 = ~n67679 & ~n68661 ;
  assign n68663 = ~n68658 & ~n68662 ;
  assign n68664 = ~n68656 & n68663 ;
  assign n68665 = ~n68645 & n68664 ;
  assign n68666 = \u0_L2_reg[23]/NET0131  & ~n68665 ;
  assign n68667 = ~\u0_L2_reg[23]/NET0131  & n68665 ;
  assign n68668 = ~n68666 & ~n68667 ;
  assign n68683 = n67802 & ~n67807 ;
  assign n68684 = ~n67824 & n68683 ;
  assign n68685 = ~n67795 & n68684 ;
  assign n68681 = ~n67802 & ~n68113 ;
  assign n68682 = n67777 & n67835 ;
  assign n68686 = ~n68681 & ~n68682 ;
  assign n68687 = ~n68685 & n68686 ;
  assign n68688 = ~n67765 & ~n68687 ;
  assign n68672 = n67777 & ~n67825 ;
  assign n68673 = ~n67777 & ~n67808 ;
  assign n68674 = ~n68672 & ~n68673 ;
  assign n68669 = ~n67802 & n67810 ;
  assign n68675 = ~n68118 & ~n68669 ;
  assign n68676 = ~n67809 & n68675 ;
  assign n68670 = n67795 & n67802 ;
  assign n68671 = n67777 & n68073 ;
  assign n68677 = ~n68670 & ~n68671 ;
  assign n68678 = n68676 & n68677 ;
  assign n68679 = ~n68674 & n68678 ;
  assign n68680 = n67765 & ~n68679 ;
  assign n68689 = ~n67834 & ~n67842 ;
  assign n68690 = ~n68680 & n68689 ;
  assign n68691 = ~n68688 & n68690 ;
  assign n68692 = ~\u0_L2_reg[19]/P0001  & ~n68691 ;
  assign n68693 = \u0_L2_reg[19]/P0001  & n68691 ;
  assign n68694 = ~n68692 & ~n68693 ;
  assign n68716 = ~n68444 & n68473 ;
  assign n68717 = ~n68432 & ~n68716 ;
  assign n68718 = ~n68452 & n68717 ;
  assign n68721 = ~n68445 & ~n68458 ;
  assign n68722 = ~n68460 & n68721 ;
  assign n68719 = n68444 & n68473 ;
  assign n68720 = n68432 & ~n68719 ;
  assign n68723 = ~n68481 & n68720 ;
  assign n68724 = ~n68722 & n68723 ;
  assign n68725 = ~n68718 & ~n68724 ;
  assign n68695 = n68460 & n68462 ;
  assign n68713 = n68444 & n68479 ;
  assign n68726 = ~n68695 & ~n68713 ;
  assign n68727 = ~n68725 & n68726 ;
  assign n68728 = n68491 & ~n68727 ;
  assign n68705 = n68432 & ~n68462 ;
  assign n68704 = ~n68432 & ~n68481 ;
  assign n68706 = ~n68438 & ~n68704 ;
  assign n68707 = ~n68705 & n68706 ;
  assign n68700 = n68467 & n68469 ;
  assign n68701 = ~n68451 & n68469 ;
  assign n68702 = ~n68471 & ~n68701 ;
  assign n68703 = ~n68432 & ~n68702 ;
  assign n68708 = ~n68700 & ~n68703 ;
  assign n68709 = ~n68707 & n68708 ;
  assign n68710 = ~n68491 & ~n68709 ;
  assign n68696 = ~n68517 & ~n68695 ;
  assign n68697 = ~n68438 & n68468 ;
  assign n68698 = n68696 & ~n68697 ;
  assign n68699 = n68432 & ~n68698 ;
  assign n68711 = n68438 & ~n68444 ;
  assign n68712 = ~n68432 & n68711 ;
  assign n68714 = ~n68712 & ~n68713 ;
  assign n68715 = n68451 & ~n68714 ;
  assign n68729 = ~n68699 & ~n68715 ;
  assign n68730 = ~n68710 & n68729 ;
  assign n68731 = ~n68728 & n68730 ;
  assign n68732 = ~\u0_L2_reg[25]/NET0131  & ~n68731 ;
  assign n68733 = \u0_L2_reg[25]/NET0131  & n68731 ;
  assign n68734 = ~n68732 & ~n68733 ;
  assign n68735 = n68246 & n68381 ;
  assign n68741 = ~n68301 & ~n68360 ;
  assign n68742 = ~n68735 & n68741 ;
  assign n68736 = n68275 & n68283 ;
  assign n68737 = ~n68273 & ~n68736 ;
  assign n68738 = ~n68240 & ~n68737 ;
  assign n68739 = ~n68284 & ~n68371 ;
  assign n68740 = n68267 & ~n68739 ;
  assign n68743 = ~n68738 & ~n68740 ;
  assign n68744 = n68742 & n68743 ;
  assign n68745 = n68234 & ~n68744 ;
  assign n68750 = ~n68279 & ~n68397 ;
  assign n68751 = ~n68234 & ~n68750 ;
  assign n68752 = ~n68268 & ~n68378 ;
  assign n68753 = n68246 & ~n68272 ;
  assign n68754 = ~n68291 & n68753 ;
  assign n68755 = ~n68752 & ~n68754 ;
  assign n68756 = ~n68751 & ~n68755 ;
  assign n68757 = ~n68240 & ~n68756 ;
  assign n68746 = ~n68283 & n68304 ;
  assign n68747 = ~n68276 & ~n68746 ;
  assign n68748 = n68271 & n68747 ;
  assign n68749 = ~n68234 & ~n68748 ;
  assign n68758 = n68240 & n68259 ;
  assign n68759 = ~n68277 & n68758 ;
  assign n68760 = ~n68749 & ~n68759 ;
  assign n68761 = ~n68757 & n68760 ;
  assign n68762 = ~n68745 & n68761 ;
  assign n68763 = ~\u0_L2_reg[26]/NET0131  & ~n68762 ;
  assign n68764 = \u0_L2_reg[26]/NET0131  & n68762 ;
  assign n68765 = ~n68763 & ~n68764 ;
  assign n68766 = ~n68432 & ~n68507 ;
  assign n68767 = n68438 & n68468 ;
  assign n68768 = n68432 & ~n68767 ;
  assign n68769 = n68452 & n68458 ;
  assign n68770 = ~n68470 & ~n68769 ;
  assign n68771 = n68768 & n68770 ;
  assign n68772 = ~n68766 & ~n68771 ;
  assign n68774 = ~n68438 & n68497 ;
  assign n68775 = ~n68716 & ~n68774 ;
  assign n68776 = n68432 & ~n68775 ;
  assign n68773 = n68451 & n68495 ;
  assign n68777 = n68491 & ~n68773 ;
  assign n68778 = ~n68515 & n68777 ;
  assign n68779 = ~n68776 & n68778 ;
  assign n68780 = n68467 & ~n68711 ;
  assign n68781 = n68717 & ~n68780 ;
  assign n68782 = ~n68472 & n68720 ;
  assign n68783 = ~n68781 & ~n68782 ;
  assign n68784 = ~n68452 & ~n68491 ;
  assign n68785 = n68696 & n68784 ;
  assign n68786 = ~n68783 & n68785 ;
  assign n68787 = ~n68779 & ~n68786 ;
  assign n68788 = ~n68772 & ~n68787 ;
  assign n68789 = ~\u0_L2_reg[8]/NET0131  & ~n68788 ;
  assign n68790 = \u0_L2_reg[8]/NET0131  & n68788 ;
  assign n68791 = ~n68789 & ~n68790 ;
  assign n68797 = n67869 & n67876 ;
  assign n68798 = ~n67937 & ~n68797 ;
  assign n68799 = n67908 & ~n68798 ;
  assign n68800 = ~n67887 & n67898 ;
  assign n68801 = ~n67933 & n68800 ;
  assign n68792 = ~n67876 & n67891 ;
  assign n68794 = ~n67885 & ~n67931 ;
  assign n68793 = ~n67876 & n67908 ;
  assign n68795 = n67870 & ~n68793 ;
  assign n68796 = n68794 & n68795 ;
  assign n68802 = ~n68792 & ~n68796 ;
  assign n68803 = n68801 & n68802 ;
  assign n68804 = ~n68799 & n68803 ;
  assign n68807 = ~n67886 & ~n67910 ;
  assign n68808 = n67883 & ~n68807 ;
  assign n68805 = ~n67886 & ~n67932 ;
  assign n68806 = n67885 & n68805 ;
  assign n68817 = ~n67898 & ~n68806 ;
  assign n68818 = ~n68808 & n68817 ;
  assign n68809 = ~n67889 & ~n67890 ;
  assign n68810 = ~n67921 & n68809 ;
  assign n68811 = ~n67908 & ~n68810 ;
  assign n68812 = n67876 & ~n67882 ;
  assign n68813 = ~n67863 & n68812 ;
  assign n68814 = n67882 & n67921 ;
  assign n68815 = ~n68813 & ~n68814 ;
  assign n68816 = ~n67869 & ~n68815 ;
  assign n68819 = ~n68811 & ~n68816 ;
  assign n68820 = n68818 & n68819 ;
  assign n68821 = ~n68804 & ~n68820 ;
  assign n68822 = \u0_L2_reg[12]/NET0131  & n68821 ;
  assign n68823 = ~\u0_L2_reg[12]/NET0131  & ~n68821 ;
  assign n68824 = ~n68822 & ~n68823 ;
  assign n68825 = decrypt_pad & ~\u0_uk_K_r2_reg[20]/NET0131  ;
  assign n68826 = ~decrypt_pad & ~\u0_uk_K_r2_reg[40]/NET0131  ;
  assign n68827 = ~n68825 & ~n68826 ;
  assign n68828 = \u0_R2_reg[13]/NET0131  & ~n68827 ;
  assign n68829 = ~\u0_R2_reg[13]/NET0131  & n68827 ;
  assign n68830 = ~n68828 & ~n68829 ;
  assign n68831 = decrypt_pad & ~\u0_uk_K_r2_reg[48]/NET0131  ;
  assign n68832 = ~decrypt_pad & ~\u0_uk_K_r2_reg[11]/NET0131  ;
  assign n68833 = ~n68831 & ~n68832 ;
  assign n68834 = \u0_R2_reg[10]/NET0131  & ~n68833 ;
  assign n68835 = ~\u0_R2_reg[10]/NET0131  & n68833 ;
  assign n68836 = ~n68834 & ~n68835 ;
  assign n68837 = ~n68830 & ~n68836 ;
  assign n68838 = decrypt_pad & ~\u0_uk_K_r2_reg[11]/NET0131  ;
  assign n68839 = ~decrypt_pad & ~\u0_uk_K_r2_reg[6]/NET0131  ;
  assign n68840 = ~n68838 & ~n68839 ;
  assign n68841 = \u0_R2_reg[8]/NET0131  & ~n68840 ;
  assign n68842 = ~\u0_R2_reg[8]/NET0131  & n68840 ;
  assign n68843 = ~n68841 & ~n68842 ;
  assign n68844 = n68837 & n68843 ;
  assign n68845 = decrypt_pad & ~\u0_uk_K_r2_reg[40]/NET0131  ;
  assign n68846 = ~decrypt_pad & ~\u0_uk_K_r2_reg[3]/NET0131  ;
  assign n68847 = ~n68845 & ~n68846 ;
  assign n68848 = \u0_R2_reg[9]/NET0131  & ~n68847 ;
  assign n68849 = ~\u0_R2_reg[9]/NET0131  & n68847 ;
  assign n68850 = ~n68848 & ~n68849 ;
  assign n68851 = n68844 & ~n68850 ;
  assign n68853 = n68830 & ~n68843 ;
  assign n68852 = ~n68836 & ~n68850 ;
  assign n68854 = decrypt_pad & ~\u0_uk_K_r2_reg[17]/NET0131  ;
  assign n68855 = ~decrypt_pad & ~\u0_uk_K_r2_reg[12]/NET0131  ;
  assign n68856 = ~n68854 & ~n68855 ;
  assign n68857 = \u0_R2_reg[11]/NET0131  & ~n68856 ;
  assign n68858 = ~\u0_R2_reg[11]/NET0131  & n68856 ;
  assign n68859 = ~n68857 & ~n68858 ;
  assign n68860 = n68852 & ~n68859 ;
  assign n68861 = n68853 & n68860 ;
  assign n68862 = ~n68851 & ~n68861 ;
  assign n68875 = ~n68830 & n68850 ;
  assign n68876 = n68836 & n68843 ;
  assign n68877 = n68875 & n68876 ;
  assign n68878 = decrypt_pad & ~\u0_uk_K_r2_reg[32]/NET0131  ;
  assign n68879 = ~decrypt_pad & ~\u0_uk_K_r2_reg[27]/P0001  ;
  assign n68880 = ~n68878 & ~n68879 ;
  assign n68881 = \u0_R2_reg[12]/NET0131  & ~n68880 ;
  assign n68882 = ~\u0_R2_reg[12]/NET0131  & n68880 ;
  assign n68883 = ~n68881 & ~n68882 ;
  assign n68884 = ~n68877 & ~n68883 ;
  assign n68885 = n68862 & n68884 ;
  assign n68863 = ~n68836 & n68859 ;
  assign n68864 = n68836 & ~n68859 ;
  assign n68865 = n68830 & n68864 ;
  assign n68866 = ~n68863 & ~n68865 ;
  assign n68867 = ~n68843 & n68850 ;
  assign n68868 = ~n68866 & n68867 ;
  assign n68869 = n68836 & n68850 ;
  assign n68870 = ~n68830 & ~n68843 ;
  assign n68871 = n68830 & n68843 ;
  assign n68872 = ~n68870 & ~n68871 ;
  assign n68873 = ~n68852 & ~n68872 ;
  assign n68874 = ~n68869 & n68873 ;
  assign n68886 = ~n68868 & ~n68874 ;
  assign n68887 = n68885 & n68886 ;
  assign n68888 = n68836 & ~n68843 ;
  assign n68891 = ~n68875 & ~n68888 ;
  assign n68892 = n68830 & ~n68850 ;
  assign n68893 = n68891 & ~n68892 ;
  assign n68894 = ~n68843 & ~n68850 ;
  assign n68895 = ~n68859 & ~n68894 ;
  assign n68896 = n68893 & n68895 ;
  assign n68889 = ~n68830 & n68888 ;
  assign n68890 = n68850 & n68889 ;
  assign n68897 = n68883 & ~n68890 ;
  assign n68898 = ~n68896 & n68897 ;
  assign n68899 = ~n68887 & ~n68898 ;
  assign n68902 = ~n68870 & n68883 ;
  assign n68903 = ~n68893 & n68902 ;
  assign n68900 = n68852 & n68870 ;
  assign n68901 = n68836 & n68892 ;
  assign n68904 = ~n68900 & ~n68901 ;
  assign n68905 = ~n68903 & n68904 ;
  assign n68906 = n68859 & ~n68905 ;
  assign n68907 = ~n68899 & ~n68906 ;
  assign n68908 = ~\u0_L2_reg[6]/NET0131  & ~n68907 ;
  assign n68909 = \u0_L2_reg[6]/NET0131  & n68907 ;
  assign n68910 = ~n68908 & ~n68909 ;
  assign n68922 = ~n68562 & ~n68565 ;
  assign n68923 = n68152 & ~n68922 ;
  assign n68924 = ~n68195 & n68599 ;
  assign n68925 = ~n68152 & ~n68205 ;
  assign n68926 = ~n68924 & n68925 ;
  assign n68927 = ~n68923 & ~n68926 ;
  assign n68928 = ~n68202 & ~n68211 ;
  assign n68929 = ~n68181 & n68928 ;
  assign n68930 = ~n68927 & n68929 ;
  assign n68931 = n68146 & ~n68930 ;
  assign n68911 = ~n68572 & n68605 ;
  assign n68912 = n68152 & ~n68561 ;
  assign n68913 = ~n68911 & n68912 ;
  assign n68914 = ~n68214 & ~n68913 ;
  assign n68915 = ~n68146 & ~n68914 ;
  assign n68918 = ~n68152 & ~n68213 ;
  assign n68919 = n68195 & n68584 ;
  assign n68920 = ~n68613 & ~n68919 ;
  assign n68921 = ~n68146 & ~n68920 ;
  assign n68916 = n68152 & n68179 ;
  assign n68917 = n68604 & n68916 ;
  assign n68932 = ~n68201 & ~n68917 ;
  assign n68933 = ~n68921 & n68932 ;
  assign n68934 = ~n68918 & n68933 ;
  assign n68935 = ~n68915 & n68934 ;
  assign n68936 = ~n68931 & n68935 ;
  assign n68937 = ~\u0_L2_reg[27]/NET0131  & ~n68936 ;
  assign n68938 = \u0_L2_reg[27]/NET0131  & n68936 ;
  assign n68939 = ~n68937 & ~n68938 ;
  assign n68941 = n68451 & n68479 ;
  assign n68942 = ~n68513 & ~n68941 ;
  assign n68943 = n68432 & ~n68942 ;
  assign n68940 = n68461 & n68500 ;
  assign n68944 = ~n68507 & ~n68940 ;
  assign n68945 = ~n68943 & n68944 ;
  assign n68946 = n68491 & ~n68945 ;
  assign n68948 = ~n68480 & ~n68716 ;
  assign n68949 = ~n68491 & ~n68948 ;
  assign n68947 = ~n68495 & ~n68717 ;
  assign n68950 = ~n68494 & ~n68774 ;
  assign n68951 = ~n68947 & n68950 ;
  assign n68952 = ~n68949 & n68951 ;
  assign n68953 = ~n68459 & ~n68711 ;
  assign n68954 = ~n68471 & ~n68953 ;
  assign n68955 = ~n68438 & n68467 ;
  assign n68956 = ~n68954 & ~n68955 ;
  assign n68957 = ~n68491 & ~n68956 ;
  assign n68958 = ~n68472 & n68768 ;
  assign n68959 = ~n68957 & n68958 ;
  assign n68960 = ~n68952 & ~n68959 ;
  assign n68961 = ~n68946 & ~n68960 ;
  assign n68962 = ~\u0_L2_reg[3]/NET0131  & ~n68961 ;
  assign n68963 = \u0_L2_reg[3]/NET0131  & n68961 ;
  assign n68964 = ~n68962 & ~n68963 ;
  assign n68976 = ~n67718 & n68041 ;
  assign n68967 = n67686 & n67733 ;
  assign n68968 = ~n67742 & ~n68967 ;
  assign n68975 = n67680 & ~n68968 ;
  assign n68977 = ~n68058 & ~n68975 ;
  assign n68978 = ~n68976 & n68977 ;
  assign n68979 = n67700 & ~n68978 ;
  assign n68965 = ~n67673 & ~n67745 ;
  assign n68966 = ~n68041 & ~n68965 ;
  assign n68969 = ~n67679 & n68968 ;
  assign n68970 = n67679 & ~n68037 ;
  assign n68971 = n68637 & n68970 ;
  assign n68972 = ~n68969 & ~n68971 ;
  assign n68973 = ~n68966 & ~n68972 ;
  assign n68974 = ~n67700 & ~n68973 ;
  assign n68980 = n67673 & ~n68967 ;
  assign n68981 = ~n67679 & ~n68965 ;
  assign n68982 = ~n68980 & n68981 ;
  assign n68983 = ~n68974 & ~n68982 ;
  assign n68984 = ~n68979 & n68983 ;
  assign n68985 = ~\u0_L2_reg[9]/NET0131  & ~n68984 ;
  assign n68986 = \u0_L2_reg[9]/NET0131  & n68984 ;
  assign n68987 = ~n68985 & ~n68986 ;
  assign n68992 = ~n67863 & ~n68794 ;
  assign n68993 = ~n67889 & n68992 ;
  assign n68994 = n67908 & ~n68993 ;
  assign n68995 = ~n67876 & ~n68805 ;
  assign n68989 = n67869 & n68794 ;
  assign n68996 = n67863 & n68812 ;
  assign n68997 = ~n67908 & ~n68996 ;
  assign n68998 = ~n68989 & n68997 ;
  assign n68999 = ~n68995 & n68998 ;
  assign n69000 = ~n68994 & ~n68999 ;
  assign n68988 = ~n67869 & n67931 ;
  assign n68990 = ~n68988 & ~n68989 ;
  assign n68991 = n67863 & ~n68990 ;
  assign n69001 = n67898 & ~n68991 ;
  assign n69002 = ~n69000 & n69001 ;
  assign n69004 = n67886 & n68794 ;
  assign n69003 = n67908 & ~n68988 ;
  assign n69005 = ~n68992 & n69003 ;
  assign n69006 = ~n69004 & n69005 ;
  assign n69007 = ~n67898 & ~n69006 ;
  assign n69008 = ~n69002 & ~n69007 ;
  assign n69009 = ~n67908 & n68991 ;
  assign n69010 = ~n67908 & n68993 ;
  assign n69011 = ~n67918 & ~n69010 ;
  assign n69012 = n67898 & ~n67908 ;
  assign n69013 = ~n69011 & ~n69012 ;
  assign n69014 = ~n69009 & ~n69013 ;
  assign n69015 = ~n69008 & n69014 ;
  assign n69016 = ~\u0_L2_reg[7]/NET0131  & ~n69015 ;
  assign n69017 = \u0_L2_reg[7]/NET0131  & n69015 ;
  assign n69018 = ~n69016 & ~n69017 ;
  assign n69020 = ~n67932 & ~n68988 ;
  assign n69021 = ~n68992 & ~n69020 ;
  assign n69019 = n67869 & n67885 ;
  assign n69022 = ~n67908 & ~n69019 ;
  assign n69023 = ~n69021 & n69022 ;
  assign n69024 = ~n67891 & n67908 ;
  assign n69025 = ~n67917 & ~n68996 ;
  assign n69026 = n69024 & n69025 ;
  assign n69027 = ~n69023 & ~n69026 ;
  assign n69028 = n67886 & n68812 ;
  assign n69029 = ~n69027 & ~n69028 ;
  assign n69030 = n67898 & ~n69029 ;
  assign n69031 = ~n68809 & ~n68813 ;
  assign n69032 = ~n67908 & ~n69031 ;
  assign n69033 = ~n68813 & n69003 ;
  assign n69034 = ~n69032 & ~n69033 ;
  assign n69035 = n67869 & ~n68815 ;
  assign n69036 = n67888 & ~n69035 ;
  assign n69037 = ~n69034 & n69036 ;
  assign n69038 = ~n67898 & ~n69037 ;
  assign n69039 = n67884 & n67908 ;
  assign n69040 = n67928 & ~n68812 ;
  assign n69041 = n67922 & n69040 ;
  assign n69042 = ~n69039 & ~n69041 ;
  assign n69043 = ~n69038 & n69042 ;
  assign n69044 = ~n69030 & n69043 ;
  assign n69045 = \u0_L2_reg[32]/NET0131  & n69044 ;
  assign n69046 = ~\u0_L2_reg[32]/NET0131  & ~n69044 ;
  assign n69047 = ~n69045 & ~n69046 ;
  assign n69048 = n68852 & ~n68872 ;
  assign n69052 = ~n68859 & ~n69048 ;
  assign n69049 = ~n68870 & ~n68891 ;
  assign n69050 = ~n68850 & n68876 ;
  assign n69051 = ~n68830 & n69050 ;
  assign n69053 = ~n69049 & ~n69051 ;
  assign n69054 = n69052 & n69053 ;
  assign n69055 = ~n68836 & n68853 ;
  assign n69056 = ~n68889 & ~n69055 ;
  assign n69057 = ~n68843 & n68875 ;
  assign n69058 = n68859 & ~n69050 ;
  assign n69059 = ~n69057 & n69058 ;
  assign n69060 = n69056 & n69059 ;
  assign n69061 = ~n69054 & ~n69060 ;
  assign n69062 = ~n68883 & ~n69061 ;
  assign n69063 = ~n68850 & ~n68853 ;
  assign n69064 = n68863 & n69063 ;
  assign n69070 = n68883 & ~n69064 ;
  assign n69071 = n68862 & n69070 ;
  assign n69065 = ~n68859 & n68873 ;
  assign n69066 = n68836 & n68853 ;
  assign n69067 = n68850 & n68876 ;
  assign n69068 = ~n69066 & ~n69067 ;
  assign n69069 = n68859 & ~n69068 ;
  assign n69072 = ~n69065 & ~n69069 ;
  assign n69073 = n69071 & n69072 ;
  assign n69074 = ~n69062 & ~n69073 ;
  assign n69075 = n68850 & n68871 ;
  assign n69076 = n68864 & n69075 ;
  assign n69077 = ~n68875 & ~n68894 ;
  assign n69078 = n68863 & ~n68871 ;
  assign n69079 = n69077 & n69078 ;
  assign n69080 = ~n69076 & ~n69079 ;
  assign n69081 = ~n69074 & n69080 ;
  assign n69082 = ~\u0_L2_reg[24]/NET0131  & ~n69081 ;
  assign n69083 = \u0_L2_reg[24]/NET0131  & n69081 ;
  assign n69084 = ~n69082 & ~n69083 ;
  assign n69086 = n68859 & n69057 ;
  assign n69087 = ~n68850 & ~n68871 ;
  assign n69088 = ~n69075 & ~n69087 ;
  assign n69089 = ~n68870 & ~n69088 ;
  assign n69090 = ~n69086 & ~n69089 ;
  assign n69091 = ~n68836 & ~n69090 ;
  assign n69092 = ~n68844 & ~n68889 ;
  assign n69093 = ~n68859 & ~n69092 ;
  assign n69085 = n68850 & n69066 ;
  assign n69094 = n68883 & ~n69085 ;
  assign n69095 = ~n69093 & n69094 ;
  assign n69096 = ~n69091 & n69095 ;
  assign n69097 = ~n68837 & ~n68892 ;
  assign n69098 = ~n68843 & ~n69097 ;
  assign n69099 = ~n69075 & ~n69098 ;
  assign n69100 = ~n68859 & ~n69099 ;
  assign n69101 = n68859 & ~n68870 ;
  assign n69102 = n69088 & n69101 ;
  assign n69103 = ~n68883 & ~n68900 ;
  assign n69104 = ~n69102 & n69103 ;
  assign n69105 = ~n69100 & n69104 ;
  assign n69106 = ~n69096 & ~n69105 ;
  assign n69107 = ~n68859 & n69050 ;
  assign n69108 = ~n68850 & n68889 ;
  assign n69109 = ~n68877 & ~n69108 ;
  assign n69110 = n68859 & ~n69109 ;
  assign n69111 = ~n69107 & ~n69110 ;
  assign n69112 = ~n69106 & n69111 ;
  assign n69113 = ~\u0_L2_reg[16]/NET0131  & ~n69112 ;
  assign n69114 = \u0_L2_reg[16]/NET0131  & n69112 ;
  assign n69115 = ~n69113 & ~n69114 ;
  assign n69116 = ~n68859 & ~n68876 ;
  assign n69117 = ~n69057 & n69116 ;
  assign n69118 = ~n68851 & n68859 ;
  assign n69119 = n69056 & n69118 ;
  assign n69120 = ~n69117 & ~n69119 ;
  assign n69121 = n68883 & ~n69120 ;
  assign n69124 = ~n68875 & n68876 ;
  assign n69125 = n68837 & n68850 ;
  assign n69126 = ~n69124 & ~n69125 ;
  assign n69127 = n68859 & ~n69126 ;
  assign n69122 = n69077 & n69116 ;
  assign n69123 = n68888 & n68892 ;
  assign n69128 = ~n68883 & ~n69123 ;
  assign n69129 = ~n69048 & n69128 ;
  assign n69130 = ~n69122 & n69129 ;
  assign n69131 = ~n69127 & n69130 ;
  assign n69132 = ~n69121 & ~n69131 ;
  assign n69136 = n68830 & n68859 ;
  assign n69137 = n69050 & n69136 ;
  assign n69133 = n68864 & n68875 ;
  assign n69134 = n68869 & n68883 ;
  assign n69135 = ~n68871 & n69134 ;
  assign n69138 = ~n69133 & ~n69135 ;
  assign n69139 = ~n69137 & n69138 ;
  assign n69140 = ~n69132 & n69139 ;
  assign n69141 = \u0_L2_reg[30]/NET0131  & ~n69140 ;
  assign n69142 = ~\u0_L2_reg[30]/NET0131  & n69140 ;
  assign n69143 = ~n69141 & ~n69142 ;
  assign n69152 = ~n67996 & ~n68018 ;
  assign n69155 = n67995 & ~n69152 ;
  assign n69153 = ~n67959 & ~n68012 ;
  assign n69154 = n69152 & n69153 ;
  assign n69156 = ~n68323 & ~n68529 ;
  assign n69157 = ~n69154 & n69156 ;
  assign n69158 = ~n69155 & n69157 ;
  assign n69159 = ~n67953 & ~n69158 ;
  assign n69145 = ~n67975 & n67993 ;
  assign n69147 = ~n67974 & ~n68333 ;
  assign n69146 = n67965 & n67981 ;
  assign n69148 = ~n68342 & ~n69146 ;
  assign n69149 = n69147 & n69148 ;
  assign n69150 = ~n69145 & ~n69149 ;
  assign n69151 = n67953 & ~n69150 ;
  assign n69144 = ~n67993 & n67999 ;
  assign n69160 = n67959 & n69146 ;
  assign n69161 = ~n68526 & ~n69160 ;
  assign n69162 = n67993 & ~n69161 ;
  assign n69163 = ~n69144 & ~n69162 ;
  assign n69164 = ~n69151 & n69163 ;
  assign n69165 = ~n69159 & n69164 ;
  assign n69166 = \u0_L2_reg[18]/NET0131  & n69165 ;
  assign n69167 = ~\u0_L2_reg[18]/NET0131  & ~n69165 ;
  assign n69168 = ~n69166 & ~n69167 ;
  assign n69169 = decrypt_pad & ~\u0_uk_K_r1_reg[14]/NET0131  ;
  assign n69170 = ~decrypt_pad & ~\u0_uk_K_r1_reg[8]/NET0131  ;
  assign n69171 = ~n69169 & ~n69170 ;
  assign n69172 = \u0_R1_reg[28]/NET0131  & ~n69171 ;
  assign n69173 = ~\u0_R1_reg[28]/NET0131  & n69171 ;
  assign n69174 = ~n69172 & ~n69173 ;
  assign n69175 = decrypt_pad & ~\u0_uk_K_r1_reg[31]/NET0131  ;
  assign n69176 = ~decrypt_pad & ~\u0_uk_K_r1_reg[21]/NET0131  ;
  assign n69177 = ~n69175 & ~n69176 ;
  assign n69178 = \u0_R1_reg[27]/NET0131  & ~n69177 ;
  assign n69179 = ~\u0_R1_reg[27]/NET0131  & n69177 ;
  assign n69180 = ~n69178 & ~n69179 ;
  assign n69188 = decrypt_pad & ~\u0_uk_K_r1_reg[49]/NET0131  ;
  assign n69189 = ~decrypt_pad & ~\u0_uk_K_r1_reg[43]/NET0131  ;
  assign n69190 = ~n69188 & ~n69189 ;
  assign n69191 = \u0_R1_reg[26]/NET0131  & ~n69190 ;
  assign n69192 = ~\u0_R1_reg[26]/NET0131  & n69190 ;
  assign n69193 = ~n69191 & ~n69192 ;
  assign n69181 = decrypt_pad & ~\u0_uk_K_r1_reg[29]/NET0131  ;
  assign n69182 = ~decrypt_pad & ~\u0_uk_K_r1_reg[23]/NET0131  ;
  assign n69183 = ~n69181 & ~n69182 ;
  assign n69184 = \u0_R1_reg[24]/NET0131  & ~n69183 ;
  assign n69185 = ~\u0_R1_reg[24]/NET0131  & n69183 ;
  assign n69186 = ~n69184 & ~n69185 ;
  assign n69194 = decrypt_pad & ~\u0_uk_K_r1_reg[9]/NET0131  ;
  assign n69195 = ~decrypt_pad & ~\u0_uk_K_r1_reg[31]/NET0131  ;
  assign n69196 = ~n69194 & ~n69195 ;
  assign n69197 = \u0_R1_reg[25]/NET0131  & ~n69196 ;
  assign n69198 = ~\u0_R1_reg[25]/NET0131  & n69196 ;
  assign n69199 = ~n69197 & ~n69198 ;
  assign n69202 = decrypt_pad & ~\u0_uk_K_r1_reg[37]/NET0131  ;
  assign n69203 = ~decrypt_pad & ~\u0_uk_K_r1_reg[0]/NET0131  ;
  assign n69204 = ~n69202 & ~n69203 ;
  assign n69205 = \u0_R1_reg[29]/NET0131  & ~n69204 ;
  assign n69206 = ~\u0_R1_reg[29]/NET0131  & n69204 ;
  assign n69207 = ~n69205 & ~n69206 ;
  assign n69217 = ~n69199 & ~n69207 ;
  assign n69218 = ~n69186 & n69217 ;
  assign n69219 = n69193 & n69218 ;
  assign n69213 = ~n69186 & n69207 ;
  assign n69214 = n69186 & ~n69207 ;
  assign n69215 = ~n69213 & ~n69214 ;
  assign n69216 = ~n69193 & ~n69215 ;
  assign n69209 = n69186 & n69193 ;
  assign n69220 = n69209 & ~n69217 ;
  assign n69221 = ~n69216 & ~n69220 ;
  assign n69222 = ~n69219 & n69221 ;
  assign n69223 = ~n69180 & ~n69222 ;
  assign n69187 = n69180 & n69186 ;
  assign n69200 = ~n69193 & ~n69199 ;
  assign n69201 = n69187 & n69200 ;
  assign n69208 = n69199 & n69207 ;
  assign n69210 = ~n69186 & ~n69193 ;
  assign n69211 = ~n69209 & ~n69210 ;
  assign n69212 = n69208 & ~n69211 ;
  assign n69224 = ~n69201 & ~n69212 ;
  assign n69225 = ~n69223 & n69224 ;
  assign n69226 = ~n69174 & ~n69225 ;
  assign n69228 = n69186 & ~n69199 ;
  assign n69229 = n69207 & n69228 ;
  assign n69230 = ~n69193 & n69229 ;
  assign n69231 = n69199 & n69213 ;
  assign n69232 = ~n69230 & ~n69231 ;
  assign n69233 = ~n69180 & ~n69232 ;
  assign n69237 = ~n69193 & ~n69208 ;
  assign n69236 = n69193 & n69199 ;
  assign n69238 = n69187 & ~n69236 ;
  assign n69239 = ~n69237 & n69238 ;
  assign n69227 = n69210 & n69217 ;
  assign n69234 = ~n69199 & n69213 ;
  assign n69235 = n69193 & n69234 ;
  assign n69240 = ~n69227 & ~n69235 ;
  assign n69241 = ~n69239 & n69240 ;
  assign n69242 = ~n69233 & n69241 ;
  assign n69243 = n69174 & ~n69242 ;
  assign n69244 = ~n69180 & n69199 ;
  assign n69245 = ~n69211 & n69244 ;
  assign n69247 = ~n69186 & n69199 ;
  assign n69248 = ~n69207 & n69247 ;
  assign n69249 = n69193 & n69248 ;
  assign n69246 = n69200 & ~n69207 ;
  assign n69250 = ~n69199 & n69214 ;
  assign n69251 = ~n69246 & ~n69250 ;
  assign n69252 = ~n69235 & n69251 ;
  assign n69253 = ~n69249 & n69252 ;
  assign n69254 = n69180 & ~n69253 ;
  assign n69255 = ~n69245 & ~n69254 ;
  assign n69256 = ~n69243 & n69255 ;
  assign n69257 = ~n69226 & n69256 ;
  assign n69258 = ~\u0_L1_reg[22]/NET0131  & ~n69257 ;
  assign n69259 = \u0_L1_reg[22]/NET0131  & n69257 ;
  assign n69260 = ~n69258 & ~n69259 ;
  assign n69261 = decrypt_pad & ~\u0_uk_K_r1_reg[32]/NET0131  ;
  assign n69262 = ~decrypt_pad & ~\u0_uk_K_r1_reg[24]/NET0131  ;
  assign n69263 = ~n69261 & ~n69262 ;
  assign n69264 = \u0_R1_reg[3]/NET0131  & ~n69263 ;
  assign n69265 = ~\u0_R1_reg[3]/NET0131  & n69263 ;
  assign n69266 = ~n69264 & ~n69265 ;
  assign n69280 = decrypt_pad & ~\u0_uk_K_r1_reg[55]/NET0131  ;
  assign n69281 = ~decrypt_pad & ~\u0_uk_K_r1_reg[47]/NET0131  ;
  assign n69282 = ~n69280 & ~n69281 ;
  assign n69283 = \u0_R1_reg[2]/NET0131  & ~n69282 ;
  assign n69284 = ~\u0_R1_reg[2]/NET0131  & n69282 ;
  assign n69285 = ~n69283 & ~n69284 ;
  assign n69288 = decrypt_pad & ~\u0_uk_K_r1_reg[13]/NET0131  ;
  assign n69289 = ~decrypt_pad & ~\u0_uk_K_r1_reg[5]/NET0131  ;
  assign n69290 = ~n69288 & ~n69289 ;
  assign n69291 = \u0_R1_reg[5]/NET0131  & ~n69290 ;
  assign n69292 = ~\u0_R1_reg[5]/NET0131  & n69290 ;
  assign n69293 = ~n69291 & ~n69292 ;
  assign n69343 = ~n69285 & n69293 ;
  assign n69344 = n69285 & ~n69293 ;
  assign n69345 = ~n69343 & ~n69344 ;
  assign n69267 = decrypt_pad & ~\u0_uk_K_r1_reg[19]/NET0131  ;
  assign n69268 = ~decrypt_pad & ~\u0_uk_K_r1_reg[11]/NET0131  ;
  assign n69269 = ~n69267 & ~n69268 ;
  assign n69270 = \u0_R1_reg[32]/NET0131  & ~n69269 ;
  assign n69271 = ~\u0_R1_reg[32]/NET0131  & n69269 ;
  assign n69272 = ~n69270 & ~n69271 ;
  assign n69320 = n69272 & n69293 ;
  assign n69274 = decrypt_pad & ~\u0_uk_K_r1_reg[40]/NET0131  ;
  assign n69275 = ~decrypt_pad & ~\u0_uk_K_r1_reg[32]/NET0131  ;
  assign n69276 = ~n69274 & ~n69275 ;
  assign n69277 = \u0_R1_reg[1]/NET0131  & ~n69276 ;
  assign n69278 = ~\u0_R1_reg[1]/NET0131  & n69276 ;
  assign n69279 = ~n69277 & ~n69278 ;
  assign n69294 = ~n69279 & ~n69293 ;
  assign n69308 = n69279 & n69293 ;
  assign n69346 = ~n69294 & ~n69308 ;
  assign n69347 = ~n69320 & n69346 ;
  assign n69348 = n69345 & n69347 ;
  assign n69297 = ~n69272 & n69279 ;
  assign n69338 = ~n69294 & ~n69297 ;
  assign n69302 = decrypt_pad & ~\u0_uk_K_r1_reg[10]/P0001  ;
  assign n69303 = ~decrypt_pad & ~\u0_uk_K_r1_reg[34]/NET0131  ;
  assign n69304 = ~n69302 & ~n69303 ;
  assign n69305 = \u0_R1_reg[4]/NET0131  & ~n69304 ;
  assign n69306 = ~\u0_R1_reg[4]/NET0131  & n69304 ;
  assign n69307 = ~n69305 & ~n69306 ;
  assign n69295 = n69272 & ~n69285 ;
  assign n69298 = ~n69272 & n69285 ;
  assign n69337 = ~n69295 & ~n69298 ;
  assign n69339 = ~n69307 & n69337 ;
  assign n69340 = ~n69338 & n69339 ;
  assign n69341 = n69285 & n69308 ;
  assign n69342 = n69272 & n69341 ;
  assign n69349 = ~n69340 & ~n69342 ;
  assign n69350 = ~n69348 & n69349 ;
  assign n69351 = ~n69266 & ~n69350 ;
  assign n69299 = ~n69266 & n69279 ;
  assign n69300 = ~n69298 & ~n69299 ;
  assign n69301 = ~n69297 & ~n69300 ;
  assign n69296 = n69294 & n69295 ;
  assign n69316 = ~n69296 & n69307 ;
  assign n69317 = ~n69301 & n69316 ;
  assign n69309 = ~n69293 & ~n69298 ;
  assign n69310 = n69266 & ~n69308 ;
  assign n69311 = ~n69309 & n69310 ;
  assign n69312 = n69266 & ~n69285 ;
  assign n69313 = n69279 & ~n69312 ;
  assign n69314 = ~n69272 & n69293 ;
  assign n69315 = ~n69313 & n69314 ;
  assign n69318 = ~n69311 & ~n69315 ;
  assign n69319 = n69317 & n69318 ;
  assign n69321 = ~n69285 & n69320 ;
  assign n69322 = ~n69299 & n69321 ;
  assign n69331 = ~n69307 & ~n69322 ;
  assign n69328 = n69279 & ~n69293 ;
  assign n69273 = n69266 & n69272 ;
  assign n69329 = n69273 & n69285 ;
  assign n69330 = n69328 & n69329 ;
  assign n69323 = ~n69272 & ~n69293 ;
  assign n69324 = ~n69285 & n69323 ;
  assign n69325 = n69279 & n69324 ;
  assign n69326 = n69266 & n69298 ;
  assign n69327 = n69308 & n69326 ;
  assign n69332 = ~n69325 & ~n69327 ;
  assign n69333 = ~n69330 & n69332 ;
  assign n69334 = n69331 & n69333 ;
  assign n69335 = ~n69319 & ~n69334 ;
  assign n69286 = ~n69279 & ~n69285 ;
  assign n69287 = n69273 & n69286 ;
  assign n69336 = n69294 & n69326 ;
  assign n69352 = ~n69287 & ~n69336 ;
  assign n69353 = ~n69335 & n69352 ;
  assign n69354 = ~n69351 & n69353 ;
  assign n69355 = ~\u0_L1_reg[31]/NET0131  & ~n69354 ;
  assign n69356 = \u0_L1_reg[31]/NET0131  & n69354 ;
  assign n69357 = ~n69355 & ~n69356 ;
  assign n69358 = decrypt_pad & ~\u0_uk_K_r1_reg[38]/NET0131  ;
  assign n69359 = ~decrypt_pad & ~\u0_uk_K_r1_reg[28]/NET0131  ;
  assign n69360 = ~n69358 & ~n69359 ;
  assign n69361 = \u0_R1_reg[32]/NET0131  & ~n69360 ;
  assign n69362 = ~\u0_R1_reg[32]/NET0131  & n69360 ;
  assign n69363 = ~n69361 & ~n69362 ;
  assign n69397 = decrypt_pad & ~\u0_uk_K_r1_reg[28]/NET0131  ;
  assign n69398 = ~decrypt_pad & ~\u0_uk_K_r1_reg[22]/NET0131  ;
  assign n69399 = ~n69397 & ~n69398 ;
  assign n69400 = \u0_R1_reg[31]/NET0131  & ~n69399 ;
  assign n69401 = ~\u0_R1_reg[31]/NET0131  & n69399 ;
  assign n69402 = ~n69400 & ~n69401 ;
  assign n69383 = decrypt_pad & ~\u0_uk_K_r1_reg[43]/NET0131  ;
  assign n69384 = ~decrypt_pad & ~\u0_uk_K_r1_reg[37]/NET0131  ;
  assign n69385 = ~n69383 & ~n69384 ;
  assign n69386 = \u0_R1_reg[28]/NET0131  & ~n69385 ;
  assign n69387 = ~\u0_R1_reg[28]/NET0131  & n69385 ;
  assign n69388 = ~n69386 & ~n69387 ;
  assign n69364 = decrypt_pad & ~\u0_uk_K_r1_reg[16]/NET0131  ;
  assign n69365 = ~decrypt_pad & ~\u0_uk_K_r1_reg[38]/NET0131  ;
  assign n69366 = ~n69364 & ~n69365 ;
  assign n69367 = \u0_R1_reg[30]/NET0131  & ~n69366 ;
  assign n69368 = ~\u0_R1_reg[30]/NET0131  & n69366 ;
  assign n69369 = ~n69367 & ~n69368 ;
  assign n69370 = decrypt_pad & ~\u0_uk_K_r1_reg[15]/NET0131  ;
  assign n69371 = ~decrypt_pad & ~\u0_uk_K_r1_reg[9]/NET0131  ;
  assign n69372 = ~n69370 & ~n69371 ;
  assign n69373 = \u0_R1_reg[29]/NET0131  & ~n69372 ;
  assign n69374 = ~\u0_R1_reg[29]/NET0131  & n69372 ;
  assign n69375 = ~n69373 & ~n69374 ;
  assign n69418 = ~n69369 & ~n69375 ;
  assign n69419 = ~n69388 & n69418 ;
  assign n69420 = ~n69402 & ~n69419 ;
  assign n69377 = decrypt_pad & ~\u0_uk_K_r1_reg[0]/NET0131  ;
  assign n69378 = ~decrypt_pad & ~\u0_uk_K_r1_reg[49]/NET0131  ;
  assign n69379 = ~n69377 & ~n69378 ;
  assign n69380 = \u0_R1_reg[1]/NET0131  & ~n69379 ;
  assign n69381 = ~\u0_R1_reg[1]/NET0131  & n69379 ;
  assign n69382 = ~n69380 & ~n69381 ;
  assign n69411 = n69375 & ~n69382 ;
  assign n69412 = n69388 & n69411 ;
  assign n69413 = ~n69369 & n69412 ;
  assign n69404 = ~n69369 & n69388 ;
  assign n69421 = ~n69404 & ~n69411 ;
  assign n69422 = ~n69413 & ~n69421 ;
  assign n69423 = n69402 & ~n69422 ;
  assign n69424 = ~n69420 & ~n69423 ;
  assign n69425 = n69382 & ~n69388 ;
  assign n69426 = n69375 & n69425 ;
  assign n69427 = n69369 & n69426 ;
  assign n69428 = ~n69424 & ~n69427 ;
  assign n69429 = n69363 & ~n69428 ;
  assign n69406 = ~n69369 & ~n69382 ;
  assign n69394 = ~n69375 & n69382 ;
  assign n69405 = ~n69382 & n69388 ;
  assign n69407 = ~n69394 & ~n69405 ;
  assign n69408 = ~n69406 & n69407 ;
  assign n69409 = ~n69404 & ~n69408 ;
  assign n69410 = ~n69402 & ~n69409 ;
  assign n69391 = ~n69375 & n69388 ;
  assign n69392 = n69369 & n69391 ;
  assign n69393 = ~n69382 & n69392 ;
  assign n69395 = ~n69388 & n69394 ;
  assign n69396 = ~n69393 & ~n69395 ;
  assign n69403 = ~n69396 & n69402 ;
  assign n69376 = n69369 & n69375 ;
  assign n69389 = n69382 & n69388 ;
  assign n69390 = n69376 & n69389 ;
  assign n69414 = ~n69390 & ~n69413 ;
  assign n69415 = ~n69403 & n69414 ;
  assign n69416 = ~n69410 & n69415 ;
  assign n69417 = ~n69363 & ~n69416 ;
  assign n69430 = ~n69369 & n69375 ;
  assign n69431 = ~n69405 & ~n69430 ;
  assign n69432 = ~n69421 & n69431 ;
  assign n69435 = n69402 & ~n69432 ;
  assign n69433 = ~n69382 & n69419 ;
  assign n69434 = n69369 & n69395 ;
  assign n69436 = ~n69433 & ~n69434 ;
  assign n69437 = n69435 & n69436 ;
  assign n69438 = n69363 & n69392 ;
  assign n69439 = ~n69402 & ~n69413 ;
  assign n69440 = ~n69438 & n69439 ;
  assign n69441 = ~n69437 & ~n69440 ;
  assign n69442 = ~n69417 & ~n69441 ;
  assign n69443 = ~n69429 & n69442 ;
  assign n69444 = \u0_L1_reg[5]/NET0131  & ~n69443 ;
  assign n69445 = ~\u0_L1_reg[5]/NET0131  & n69443 ;
  assign n69446 = ~n69444 & ~n69445 ;
  assign n69502 = decrypt_pad & ~\u0_uk_K_r1_reg[7]/P0001  ;
  assign n69503 = ~decrypt_pad & ~\u0_uk_K_r1_reg[1]/NET0131  ;
  assign n69504 = ~n69502 & ~n69503 ;
  assign n69505 = \u0_R1_reg[24]/NET0131  & ~n69504 ;
  assign n69506 = ~\u0_R1_reg[24]/NET0131  & n69504 ;
  assign n69507 = ~n69505 & ~n69506 ;
  assign n69460 = decrypt_pad & ~\u0_uk_K_r1_reg[23]/NET0131  ;
  assign n69461 = ~decrypt_pad & ~\u0_uk_K_r1_reg[45]/NET0131  ;
  assign n69462 = ~n69460 & ~n69461 ;
  assign n69463 = \u0_R1_reg[22]/NET0131  & ~n69462 ;
  assign n69464 = ~\u0_R1_reg[22]/NET0131  & n69462 ;
  assign n69465 = ~n69463 & ~n69464 ;
  assign n69447 = decrypt_pad & ~\u0_uk_K_r1_reg[1]/NET0131  ;
  assign n69448 = ~decrypt_pad & ~\u0_uk_K_r1_reg[50]/NET0131  ;
  assign n69449 = ~n69447 & ~n69448 ;
  assign n69450 = \u0_R1_reg[21]/NET0131  & ~n69449 ;
  assign n69451 = ~\u0_R1_reg[21]/NET0131  & n69449 ;
  assign n69452 = ~n69450 & ~n69451 ;
  assign n69453 = decrypt_pad & ~\u0_uk_K_r1_reg[45]/NET0131  ;
  assign n69454 = ~decrypt_pad & ~\u0_uk_K_r1_reg[35]/NET0131  ;
  assign n69455 = ~n69453 & ~n69454 ;
  assign n69456 = \u0_R1_reg[20]/NET0131  & ~n69455 ;
  assign n69457 = ~\u0_R1_reg[20]/NET0131  & n69455 ;
  assign n69458 = ~n69456 & ~n69457 ;
  assign n69459 = n69452 & ~n69458 ;
  assign n69477 = decrypt_pad & ~\u0_uk_K_r1_reg[2]/NET0131  ;
  assign n69478 = ~decrypt_pad & ~\u0_uk_K_r1_reg[51]/NET0131  ;
  assign n69479 = ~n69477 & ~n69478 ;
  assign n69480 = \u0_R1_reg[25]/NET0131  & ~n69479 ;
  assign n69481 = ~\u0_R1_reg[25]/NET0131  & n69479 ;
  assign n69482 = ~n69480 & ~n69481 ;
  assign n69491 = n69458 & n69482 ;
  assign n69532 = ~n69459 & ~n69491 ;
  assign n69533 = n69465 & ~n69532 ;
  assign n69470 = decrypt_pad & ~\u0_uk_K_r1_reg[36]/NET0131  ;
  assign n69471 = ~decrypt_pad & ~\u0_uk_K_r1_reg[30]/NET0131  ;
  assign n69472 = ~n69470 & ~n69471 ;
  assign n69473 = \u0_R1_reg[23]/NET0131  & ~n69472 ;
  assign n69474 = ~\u0_R1_reg[23]/NET0131  & n69472 ;
  assign n69475 = ~n69473 & ~n69474 ;
  assign n69529 = n69452 & n69482 ;
  assign n69530 = ~n69458 & n69529 ;
  assign n69531 = ~n69465 & ~n69530 ;
  assign n69534 = ~n69475 & ~n69531 ;
  assign n69535 = ~n69533 & n69534 ;
  assign n69489 = n69458 & ~n69482 ;
  assign n69522 = ~n69452 & n69489 ;
  assign n69523 = ~n69465 & n69522 ;
  assign n69466 = n69459 & n69465 ;
  assign n69521 = n69452 & n69491 ;
  assign n69524 = ~n69466 & ~n69521 ;
  assign n69525 = ~n69523 & n69524 ;
  assign n69526 = n69475 & ~n69525 ;
  assign n69488 = ~n69465 & ~n69475 ;
  assign n69527 = n69488 & n69491 ;
  assign n69528 = ~n69452 & n69527 ;
  assign n69536 = ~n69526 & ~n69528 ;
  assign n69537 = ~n69535 & n69536 ;
  assign n69538 = n69507 & ~n69537 ;
  assign n69467 = n69458 & ~n69465 ;
  assign n69468 = n69452 & n69467 ;
  assign n69469 = ~n69466 & ~n69468 ;
  assign n69476 = ~n69469 & ~n69475 ;
  assign n69496 = ~n69467 & n69475 ;
  assign n69495 = ~n69458 & ~n69482 ;
  assign n69497 = ~n69452 & ~n69495 ;
  assign n69498 = n69496 & n69497 ;
  assign n69483 = n69452 & ~n69482 ;
  assign n69484 = n69458 & ~n69483 ;
  assign n69485 = ~n69458 & ~n69475 ;
  assign n69486 = ~n69465 & ~n69485 ;
  assign n69487 = ~n69484 & n69486 ;
  assign n69490 = n69488 & n69489 ;
  assign n69492 = ~n69452 & n69465 ;
  assign n69493 = n69491 & n69492 ;
  assign n69494 = ~n69490 & ~n69493 ;
  assign n69499 = ~n69487 & n69494 ;
  assign n69500 = ~n69498 & n69499 ;
  assign n69501 = ~n69476 & n69500 ;
  assign n69508 = ~n69501 & ~n69507 ;
  assign n69518 = ~n69465 & n69483 ;
  assign n69519 = ~n69491 & ~n69518 ;
  assign n69520 = n69496 & ~n69519 ;
  assign n69509 = ~n69452 & n69495 ;
  assign n69510 = n69488 & n69509 ;
  assign n69511 = ~n69452 & ~n69465 ;
  assign n69512 = ~n69458 & n69482 ;
  assign n69513 = n69511 & n69512 ;
  assign n69514 = n69475 & n69513 ;
  assign n69515 = n69452 & n69489 ;
  assign n69516 = n69488 & n69515 ;
  assign n69517 = ~n69514 & ~n69516 ;
  assign n69539 = ~n69510 & n69517 ;
  assign n69540 = ~n69520 & n69539 ;
  assign n69541 = ~n69508 & n69540 ;
  assign n69542 = ~n69538 & n69541 ;
  assign n69543 = \u0_L1_reg[11]/NET0131  & ~n69542 ;
  assign n69544 = ~\u0_L1_reg[11]/NET0131  & n69542 ;
  assign n69545 = ~n69543 & ~n69544 ;
  assign n69546 = decrypt_pad & ~\u0_uk_K_r1_reg[12]/NET0131  ;
  assign n69547 = ~decrypt_pad & ~\u0_uk_K_r1_reg[4]/NET0131  ;
  assign n69548 = ~n69546 & ~n69547 ;
  assign n69549 = \u0_R1_reg[16]/NET0131  & ~n69548 ;
  assign n69550 = ~\u0_R1_reg[16]/NET0131  & n69548 ;
  assign n69551 = ~n69549 & ~n69550 ;
  assign n69574 = decrypt_pad & ~\u0_uk_K_r1_reg[4]/NET0131  ;
  assign n69575 = ~decrypt_pad & ~\u0_uk_K_r1_reg[53]/NET0131  ;
  assign n69576 = ~n69574 & ~n69575 ;
  assign n69577 = \u0_R1_reg[15]/NET0131  & ~n69576 ;
  assign n69578 = ~\u0_R1_reg[15]/NET0131  & n69576 ;
  assign n69579 = ~n69577 & ~n69578 ;
  assign n69565 = decrypt_pad & ~\u0_uk_K_r1_reg[27]/NET0131  ;
  assign n69566 = ~decrypt_pad & ~\u0_uk_K_r1_reg[19]/NET0131  ;
  assign n69567 = ~n69565 & ~n69566 ;
  assign n69568 = \u0_R1_reg[13]/NET0131  & ~n69567 ;
  assign n69569 = ~\u0_R1_reg[13]/NET0131  & n69567 ;
  assign n69570 = ~n69568 & ~n69569 ;
  assign n69552 = decrypt_pad & ~\u0_uk_K_r1_reg[17]/NET0131  ;
  assign n69553 = ~decrypt_pad & ~\u0_uk_K_r1_reg[41]/NET0131  ;
  assign n69554 = ~n69552 & ~n69553 ;
  assign n69555 = \u0_R1_reg[17]/NET0131  & ~n69554 ;
  assign n69556 = ~\u0_R1_reg[17]/NET0131  & n69554 ;
  assign n69557 = ~n69555 & ~n69556 ;
  assign n69558 = decrypt_pad & ~\u0_uk_K_r1_reg[33]/NET0131  ;
  assign n69559 = ~decrypt_pad & ~\u0_uk_K_r1_reg[25]/NET0131  ;
  assign n69560 = ~n69558 & ~n69559 ;
  assign n69561 = \u0_R1_reg[12]/NET0131  & ~n69560 ;
  assign n69562 = ~\u0_R1_reg[12]/NET0131  & n69560 ;
  assign n69563 = ~n69561 & ~n69562 ;
  assign n69582 = ~n69557 & n69563 ;
  assign n69617 = n69570 & n69582 ;
  assign n69618 = n69579 & n69617 ;
  assign n69583 = decrypt_pad & ~\u0_uk_K_r1_reg[53]/NET0131  ;
  assign n69584 = ~decrypt_pad & ~\u0_uk_K_r1_reg[20]/NET0131  ;
  assign n69585 = ~n69583 & ~n69584 ;
  assign n69586 = \u0_R1_reg[14]/NET0131  & ~n69585 ;
  assign n69587 = ~\u0_R1_reg[14]/NET0131  & n69585 ;
  assign n69588 = ~n69586 & ~n69587 ;
  assign n69611 = n69557 & ~n69563 ;
  assign n69612 = n69570 & n69611 ;
  assign n69620 = ~n69588 & n69612 ;
  assign n69621 = ~n69618 & ~n69620 ;
  assign n69625 = n69557 & n69579 ;
  assign n69626 = ~n69557 & ~n69579 ;
  assign n69627 = ~n69625 & ~n69626 ;
  assign n69572 = ~n69563 & ~n69570 ;
  assign n69610 = ~n69579 & ~n69588 ;
  assign n69628 = n69572 & ~n69610 ;
  assign n69629 = ~n69627 & n69628 ;
  assign n69594 = ~n69563 & n69570 ;
  assign n69600 = n69563 & ~n69570 ;
  assign n69622 = ~n69594 & ~n69600 ;
  assign n69623 = n69610 & ~n69622 ;
  assign n69564 = n69557 & n69563 ;
  assign n69571 = n69564 & n69570 ;
  assign n69624 = n69571 & n69588 ;
  assign n69630 = ~n69623 & ~n69624 ;
  assign n69631 = ~n69629 & n69630 ;
  assign n69632 = n69621 & n69631 ;
  assign n69633 = n69551 & ~n69632 ;
  assign n69573 = ~n69557 & n69572 ;
  assign n69580 = ~n69573 & n69579 ;
  assign n69581 = ~n69571 & n69580 ;
  assign n69589 = n69582 & n69588 ;
  assign n69590 = n69557 & ~n69570 ;
  assign n69591 = ~n69579 & ~n69590 ;
  assign n69592 = ~n69589 & n69591 ;
  assign n69593 = ~n69581 & ~n69592 ;
  assign n69595 = ~n69557 & n69594 ;
  assign n69596 = n69588 & n69595 ;
  assign n69603 = ~n69557 & ~n69588 ;
  assign n69604 = n69572 & n69603 ;
  assign n69605 = ~n69596 & ~n69604 ;
  assign n69597 = n69579 & n69588 ;
  assign n69598 = n69570 & n69597 ;
  assign n69599 = ~n69563 & n69598 ;
  assign n69601 = ~n69588 & n69600 ;
  assign n69602 = n69557 & n69601 ;
  assign n69606 = ~n69599 & ~n69602 ;
  assign n69607 = n69605 & n69606 ;
  assign n69608 = ~n69593 & n69607 ;
  assign n69609 = ~n69551 & ~n69608 ;
  assign n69614 = ~n69570 & n69589 ;
  assign n69615 = ~n69604 & ~n69614 ;
  assign n69616 = n69579 & ~n69615 ;
  assign n69613 = n69610 & n69612 ;
  assign n69619 = ~n69588 & n69618 ;
  assign n69634 = ~n69613 & ~n69619 ;
  assign n69635 = ~n69616 & n69634 ;
  assign n69636 = ~n69609 & n69635 ;
  assign n69637 = ~n69633 & n69636 ;
  assign n69638 = ~\u0_L1_reg[20]/NET0131  & ~n69637 ;
  assign n69639 = \u0_L1_reg[20]/NET0131  & n69637 ;
  assign n69640 = ~n69638 & ~n69639 ;
  assign n69641 = decrypt_pad & ~\u0_uk_K_r1_reg[35]/NET0131  ;
  assign n69642 = ~decrypt_pad & ~\u0_uk_K_r1_reg[29]/NET0131  ;
  assign n69643 = ~n69641 & ~n69642 ;
  assign n69644 = \u0_R1_reg[19]/NET0131  & ~n69643 ;
  assign n69645 = ~\u0_R1_reg[19]/NET0131  & n69643 ;
  assign n69646 = ~n69644 & ~n69645 ;
  assign n69647 = decrypt_pad & ~\u0_uk_K_r1_reg[8]/NET0131  ;
  assign n69648 = ~decrypt_pad & ~\u0_uk_K_r1_reg[2]/NET0131  ;
  assign n69649 = ~n69647 & ~n69648 ;
  assign n69650 = \u0_R1_reg[16]/NET0131  & ~n69649 ;
  assign n69651 = ~\u0_R1_reg[16]/NET0131  & n69649 ;
  assign n69652 = ~n69650 & ~n69651 ;
  assign n69653 = decrypt_pad & ~\u0_uk_K_r1_reg[51]/NET0131  ;
  assign n69654 = ~decrypt_pad & ~\u0_uk_K_r1_reg[14]/NET0131  ;
  assign n69655 = ~n69653 & ~n69654 ;
  assign n69656 = \u0_R1_reg[21]/NET0131  & ~n69655 ;
  assign n69657 = ~\u0_R1_reg[21]/NET0131  & n69655 ;
  assign n69658 = ~n69656 & ~n69657 ;
  assign n69660 = decrypt_pad & ~\u0_uk_K_r1_reg[52]/NET0131  ;
  assign n69661 = ~decrypt_pad & ~\u0_uk_K_r1_reg[42]/NET0131  ;
  assign n69662 = ~n69660 & ~n69661 ;
  assign n69663 = \u0_R1_reg[18]/NET0131  & ~n69662 ;
  assign n69664 = ~\u0_R1_reg[18]/NET0131  & n69662 ;
  assign n69665 = ~n69663 & ~n69664 ;
  assign n69666 = decrypt_pad & ~\u0_uk_K_r1_reg[30]/NET0131  ;
  assign n69667 = ~decrypt_pad & ~\u0_uk_K_r1_reg[52]/NET0131  ;
  assign n69668 = ~n69666 & ~n69667 ;
  assign n69669 = \u0_R1_reg[17]/NET0131  & ~n69668 ;
  assign n69670 = ~\u0_R1_reg[17]/NET0131  & n69668 ;
  assign n69671 = ~n69669 & ~n69670 ;
  assign n69678 = ~n69665 & n69671 ;
  assign n69679 = n69658 & n69678 ;
  assign n69680 = n69652 & n69679 ;
  assign n69676 = ~n69652 & n69658 ;
  assign n69677 = ~n69671 & n69676 ;
  assign n69659 = n69652 & ~n69658 ;
  assign n69672 = ~n69665 & ~n69671 ;
  assign n69673 = n69659 & n69672 ;
  assign n69674 = n69665 & n69671 ;
  assign n69675 = ~n69658 & n69674 ;
  assign n69681 = ~n69673 & ~n69675 ;
  assign n69682 = ~n69677 & n69681 ;
  assign n69683 = ~n69680 & n69682 ;
  assign n69684 = ~n69646 & ~n69683 ;
  assign n69689 = n69658 & n69665 ;
  assign n69690 = n69652 & n69689 ;
  assign n69685 = ~n69652 & n69678 ;
  assign n69687 = ~n69652 & ~n69658 ;
  assign n69688 = ~n69671 & n69687 ;
  assign n69691 = ~n69685 & ~n69688 ;
  assign n69692 = ~n69690 & n69691 ;
  assign n69693 = n69646 & ~n69692 ;
  assign n69686 = ~n69658 & n69685 ;
  assign n69694 = n69652 & n69658 ;
  assign n69695 = n69665 & ~n69671 ;
  assign n69696 = n69694 & n69695 ;
  assign n69697 = ~n69686 & ~n69696 ;
  assign n69698 = ~n69693 & n69697 ;
  assign n69699 = ~n69684 & n69698 ;
  assign n69700 = decrypt_pad & ~\u0_uk_K_r1_reg[50]/NET0131  ;
  assign n69701 = ~decrypt_pad & ~\u0_uk_K_r1_reg[44]/P0001  ;
  assign n69702 = ~n69700 & ~n69701 ;
  assign n69703 = \u0_R1_reg[20]/NET0131  & ~n69702 ;
  assign n69704 = ~\u0_R1_reg[20]/NET0131  & n69702 ;
  assign n69705 = ~n69703 & ~n69704 ;
  assign n69706 = ~n69699 & ~n69705 ;
  assign n69711 = ~n69658 & n69671 ;
  assign n69712 = n69652 & n69711 ;
  assign n69709 = ~n69665 & n69694 ;
  assign n69710 = n69676 & ~n69678 ;
  assign n69713 = ~n69709 & ~n69710 ;
  assign n69714 = ~n69712 & n69713 ;
  assign n69715 = n69646 & ~n69714 ;
  assign n69707 = ~n69672 & ~n69674 ;
  assign n69708 = n69659 & n69707 ;
  assign n69716 = ~n69646 & n69652 ;
  assign n69717 = n69658 & n69716 ;
  assign n69718 = ~n69707 & n69717 ;
  assign n69719 = ~n69708 & ~n69718 ;
  assign n69720 = ~n69715 & n69719 ;
  assign n69721 = n69705 & ~n69720 ;
  assign n69726 = ~n69652 & n69711 ;
  assign n69727 = ~n69677 & ~n69726 ;
  assign n69728 = n69665 & ~n69727 ;
  assign n69722 = n69671 & n69676 ;
  assign n69723 = ~n69688 & ~n69722 ;
  assign n69724 = ~n69665 & n69705 ;
  assign n69725 = ~n69723 & n69724 ;
  assign n69729 = ~n69646 & ~n69725 ;
  assign n69730 = ~n69728 & n69729 ;
  assign n69733 = ~n69665 & n69712 ;
  assign n69731 = n69665 & n69687 ;
  assign n69732 = ~n69671 & n69731 ;
  assign n69734 = n69646 & ~n69732 ;
  assign n69735 = ~n69733 & n69734 ;
  assign n69736 = ~n69730 & ~n69735 ;
  assign n69737 = ~n69721 & ~n69736 ;
  assign n69738 = ~n69706 & n69737 ;
  assign n69739 = ~\u0_L1_reg[14]/NET0131  & ~n69738 ;
  assign n69740 = \u0_L1_reg[14]/NET0131  & n69738 ;
  assign n69741 = ~n69739 & ~n69740 ;
  assign n69759 = ~n69595 & ~n69602 ;
  assign n69760 = n69579 & ~n69759 ;
  assign n69756 = ~n69563 & n69588 ;
  assign n69757 = n69590 & n69756 ;
  assign n69758 = ~n69624 & ~n69757 ;
  assign n69748 = n69557 & ~n69588 ;
  assign n69761 = n69570 & n69748 ;
  assign n69762 = ~n69582 & ~n69761 ;
  assign n69746 = n69570 & ~n69588 ;
  assign n69747 = n69563 & n69746 ;
  assign n69763 = ~n69579 & ~n69747 ;
  assign n69764 = ~n69762 & n69763 ;
  assign n69765 = n69758 & ~n69764 ;
  assign n69766 = ~n69760 & n69765 ;
  assign n69767 = n69551 & ~n69766 ;
  assign n69742 = n69579 & n69611 ;
  assign n69743 = ~n69573 & ~n69742 ;
  assign n69744 = ~n69597 & ~n69743 ;
  assign n69749 = n69579 & n69600 ;
  assign n69750 = ~n69748 & n69749 ;
  assign n69745 = n69564 & n69610 ;
  assign n69751 = ~n69745 & ~n69747 ;
  assign n69752 = ~n69596 & n69751 ;
  assign n69753 = ~n69750 & n69752 ;
  assign n69754 = ~n69744 & n69753 ;
  assign n69755 = ~n69551 & ~n69754 ;
  assign n69768 = ~n69604 & n69758 ;
  assign n69769 = ~n69579 & ~n69768 ;
  assign n69770 = ~n69599 & ~n69619 ;
  assign n69771 = ~n69769 & n69770 ;
  assign n69772 = ~n69755 & n69771 ;
  assign n69773 = ~n69767 & n69772 ;
  assign n69774 = ~\u0_L1_reg[10]/NET0131  & ~n69773 ;
  assign n69775 = \u0_L1_reg[10]/NET0131  & n69773 ;
  assign n69776 = ~n69774 & ~n69775 ;
  assign n69796 = ~n69671 & n69694 ;
  assign n69797 = ~n69646 & ~n69796 ;
  assign n69798 = ~n69685 & n69797 ;
  assign n69788 = ~n69652 & ~n69671 ;
  assign n69801 = n69646 & ~n69788 ;
  assign n69802 = ~n69731 & n69801 ;
  assign n69799 = ~n69658 & n69672 ;
  assign n69800 = n69671 & n69694 ;
  assign n69803 = ~n69799 & ~n69800 ;
  assign n69804 = n69802 & n69803 ;
  assign n69805 = ~n69798 & ~n69804 ;
  assign n69777 = n69659 & n69674 ;
  assign n69806 = ~n69679 & ~n69777 ;
  assign n69807 = ~n69805 & n69806 ;
  assign n69808 = n69705 & ~n69807 ;
  assign n69790 = n69646 & ~n69711 ;
  assign n69789 = ~n69646 & ~n69788 ;
  assign n69791 = ~n69665 & ~n69789 ;
  assign n69792 = ~n69790 & n69791 ;
  assign n69783 = n69674 & n69676 ;
  assign n69784 = n69659 & ~n69671 ;
  assign n69785 = ~n69652 & n69674 ;
  assign n69786 = ~n69784 & ~n69785 ;
  assign n69787 = ~n69646 & ~n69786 ;
  assign n69793 = ~n69783 & ~n69787 ;
  assign n69794 = ~n69792 & n69793 ;
  assign n69795 = ~n69705 & ~n69794 ;
  assign n69778 = ~n69732 & ~n69777 ;
  assign n69779 = n69672 & n69676 ;
  assign n69780 = n69778 & ~n69779 ;
  assign n69781 = n69646 & ~n69780 ;
  assign n69782 = n69695 & n69716 ;
  assign n69809 = ~n69680 & ~n69782 ;
  assign n69810 = ~n69781 & n69809 ;
  assign n69811 = ~n69795 & n69810 ;
  assign n69812 = ~n69808 & n69811 ;
  assign n69813 = ~\u0_L1_reg[25]/NET0131  & ~n69812 ;
  assign n69814 = \u0_L1_reg[25]/NET0131  & n69812 ;
  assign n69815 = ~n69813 & ~n69814 ;
  assign n69820 = n69193 & n69229 ;
  assign n69817 = ~n69193 & n69248 ;
  assign n69818 = ~n69208 & ~n69217 ;
  assign n69819 = ~n69180 & ~n69818 ;
  assign n69827 = ~n69817 & ~n69819 ;
  assign n69828 = ~n69820 & n69827 ;
  assign n69822 = ~n69186 & n69818 ;
  assign n69823 = ~n69187 & n69193 ;
  assign n69824 = ~n69822 & n69823 ;
  assign n69816 = n69180 & n69234 ;
  assign n69821 = n69200 & n69214 ;
  assign n69825 = ~n69174 & ~n69821 ;
  assign n69826 = ~n69816 & n69825 ;
  assign n69829 = ~n69824 & n69826 ;
  assign n69830 = n69828 & n69829 ;
  assign n69837 = n69174 & ~n69230 ;
  assign n69838 = ~n69249 & n69837 ;
  assign n69834 = ~n69186 & ~n69246 ;
  assign n69835 = n69180 & ~n69228 ;
  assign n69836 = ~n69834 & n69835 ;
  assign n69831 = ~n69180 & n69235 ;
  assign n69832 = ~n69210 & ~n69250 ;
  assign n69833 = ~n69237 & ~n69832 ;
  assign n69839 = ~n69831 & ~n69833 ;
  assign n69840 = ~n69836 & n69839 ;
  assign n69841 = n69838 & n69840 ;
  assign n69842 = ~n69830 & ~n69841 ;
  assign n69843 = \u0_L1_reg[12]/NET0131  & n69842 ;
  assign n69844 = ~\u0_L1_reg[12]/NET0131  & ~n69842 ;
  assign n69845 = ~n69843 & ~n69844 ;
  assign n69846 = n69266 & n69297 ;
  assign n69847 = ~n69345 & n69846 ;
  assign n69853 = ~n69323 & n69347 ;
  assign n69854 = n69285 & n69853 ;
  assign n69848 = ~n69320 & ~n69323 ;
  assign n69849 = ~n69279 & ~n69848 ;
  assign n69850 = ~n69324 & ~n69849 ;
  assign n69851 = ~n69266 & ~n69850 ;
  assign n69852 = n69273 & ~n69346 ;
  assign n69855 = ~n69307 & ~n69852 ;
  assign n69856 = ~n69851 & n69855 ;
  assign n69857 = ~n69854 & n69856 ;
  assign n69858 = n69286 & n69320 ;
  assign n69859 = ~n69297 & ~n69298 ;
  assign n69860 = ~n69858 & n69859 ;
  assign n69861 = n69266 & ~n69860 ;
  assign n69864 = ~n69266 & ~n69297 ;
  assign n69865 = n69337 & n69864 ;
  assign n69862 = n69295 & n69328 ;
  assign n69863 = n69307 & ~n69862 ;
  assign n69866 = ~n69341 & n69863 ;
  assign n69867 = ~n69865 & n69866 ;
  assign n69868 = ~n69861 & n69867 ;
  assign n69869 = ~n69857 & ~n69868 ;
  assign n69870 = ~n69847 & ~n69869 ;
  assign n69871 = ~\u0_L1_reg[17]/NET0131  & ~n69870 ;
  assign n69872 = \u0_L1_reg[17]/NET0131  & n69870 ;
  assign n69873 = ~n69871 & ~n69872 ;
  assign n69874 = n69571 & ~n69579 ;
  assign n69875 = ~n69622 & ~n69627 ;
  assign n69876 = ~n69874 & ~n69875 ;
  assign n69877 = ~n69588 & ~n69876 ;
  assign n69880 = n69557 & n69756 ;
  assign n69881 = n69580 & ~n69880 ;
  assign n69883 = n69564 & n69588 ;
  assign n69882 = n69572 & n69748 ;
  assign n69884 = ~n69579 & ~n69882 ;
  assign n69885 = ~n69883 & n69884 ;
  assign n69886 = ~n69881 & ~n69885 ;
  assign n69878 = ~n69612 & ~n69617 ;
  assign n69879 = n69588 & ~n69878 ;
  assign n69887 = ~n69588 & n69595 ;
  assign n69888 = n69551 & ~n69887 ;
  assign n69889 = ~n69879 & n69888 ;
  assign n69890 = ~n69886 & n69889 ;
  assign n69894 = n69598 & ~n69611 ;
  assign n69891 = n69557 & ~n69756 ;
  assign n69892 = ~n69570 & ~n69579 ;
  assign n69893 = ~n69891 & n69892 ;
  assign n69895 = ~n69551 & ~n69601 ;
  assign n69896 = ~n69893 & n69895 ;
  assign n69897 = ~n69894 & n69896 ;
  assign n69898 = n69621 & n69897 ;
  assign n69899 = ~n69890 & ~n69898 ;
  assign n69900 = ~n69877 & ~n69899 ;
  assign n69901 = ~\u0_L1_reg[26]/NET0131  & ~n69900 ;
  assign n69902 = \u0_L1_reg[26]/NET0131  & n69900 ;
  assign n69903 = ~n69901 & ~n69902 ;
  assign n69941 = decrypt_pad & ~\u0_uk_K_r1_reg[11]/NET0131  ;
  assign n69942 = ~decrypt_pad & ~\u0_uk_K_r1_reg[3]/NET0131  ;
  assign n69943 = ~n69941 & ~n69942 ;
  assign n69944 = \u0_R1_reg[8]/NET0131  & ~n69943 ;
  assign n69945 = ~\u0_R1_reg[8]/NET0131  & n69943 ;
  assign n69946 = ~n69944 & ~n69945 ;
  assign n69934 = decrypt_pad & ~\u0_uk_K_r1_reg[20]/NET0131  ;
  assign n69935 = ~decrypt_pad & ~\u0_uk_K_r1_reg[12]/NET0131  ;
  assign n69936 = ~n69934 & ~n69935 ;
  assign n69937 = \u0_R1_reg[7]/NET0131  & ~n69936 ;
  assign n69938 = ~\u0_R1_reg[7]/NET0131  & n69936 ;
  assign n69939 = ~n69937 & ~n69938 ;
  assign n69904 = decrypt_pad & ~\u0_uk_K_r1_reg[26]/NET0131  ;
  assign n69905 = ~decrypt_pad & ~\u0_uk_K_r1_reg[18]/NET0131  ;
  assign n69906 = ~n69904 & ~n69905 ;
  assign n69907 = \u0_R1_reg[6]/NET0131  & ~n69906 ;
  assign n69908 = ~\u0_R1_reg[6]/NET0131  & n69906 ;
  assign n69909 = ~n69907 & ~n69908 ;
  assign n69910 = decrypt_pad & ~\u0_uk_K_r1_reg[3]/NET0131  ;
  assign n69911 = ~decrypt_pad & ~\u0_uk_K_r1_reg[27]/NET0131  ;
  assign n69912 = ~n69910 & ~n69911 ;
  assign n69913 = \u0_R1_reg[5]/NET0131  & ~n69912 ;
  assign n69914 = ~\u0_R1_reg[5]/NET0131  & n69912 ;
  assign n69915 = ~n69913 & ~n69914 ;
  assign n69917 = decrypt_pad & ~\u0_uk_K_r1_reg[24]/NET0131  ;
  assign n69918 = ~decrypt_pad & ~\u0_uk_K_r1_reg[48]/NET0131  ;
  assign n69919 = ~n69917 & ~n69918 ;
  assign n69920 = \u0_R1_reg[4]/NET0131  & ~n69919 ;
  assign n69921 = ~\u0_R1_reg[4]/NET0131  & n69919 ;
  assign n69922 = ~n69920 & ~n69921 ;
  assign n69924 = decrypt_pad & ~\u0_uk_K_r1_reg[48]/NET0131  ;
  assign n69925 = ~decrypt_pad & ~\u0_uk_K_r1_reg[40]/NET0131  ;
  assign n69926 = ~n69924 & ~n69925 ;
  assign n69927 = \u0_R1_reg[9]/NET0131  & ~n69926 ;
  assign n69928 = ~\u0_R1_reg[9]/NET0131  & n69926 ;
  assign n69929 = ~n69927 & ~n69928 ;
  assign n69947 = ~n69922 & ~n69929 ;
  assign n69971 = n69915 & n69947 ;
  assign n69972 = n69909 & n69971 ;
  assign n69930 = n69915 & ~n69929 ;
  assign n69968 = ~n69915 & n69929 ;
  assign n69973 = ~n69930 & ~n69968 ;
  assign n69974 = n69922 & n69973 ;
  assign n69975 = ~n69972 & ~n69974 ;
  assign n69976 = n69939 & ~n69975 ;
  assign n69948 = ~n69909 & n69947 ;
  assign n69949 = ~n69922 & n69929 ;
  assign n69950 = n69915 & n69949 ;
  assign n69951 = ~n69948 & ~n69950 ;
  assign n69967 = ~n69939 & ~n69951 ;
  assign n69955 = ~n69909 & n69922 ;
  assign n69969 = ~n69939 & ~n69968 ;
  assign n69970 = n69955 & ~n69969 ;
  assign n69977 = n69909 & n69949 ;
  assign n69978 = ~n69915 & n69977 ;
  assign n69979 = ~n69970 & ~n69978 ;
  assign n69980 = ~n69967 & n69979 ;
  assign n69981 = ~n69976 & n69980 ;
  assign n69982 = n69946 & ~n69981 ;
  assign n69916 = n69909 & ~n69915 ;
  assign n69923 = n69916 & ~n69922 ;
  assign n69931 = n69909 & n69922 ;
  assign n69932 = n69930 & n69931 ;
  assign n69933 = ~n69923 & ~n69932 ;
  assign n69940 = ~n69933 & ~n69939 ;
  assign n69952 = n69939 & n69951 ;
  assign n69957 = ~n69915 & n69949 ;
  assign n69953 = n69915 & n69922 ;
  assign n69954 = ~n69939 & ~n69953 ;
  assign n69956 = ~n69929 & n69955 ;
  assign n69958 = n69954 & ~n69956 ;
  assign n69959 = ~n69957 & n69958 ;
  assign n69960 = ~n69952 & ~n69959 ;
  assign n69961 = n69922 & n69929 ;
  assign n69962 = ~n69947 & ~n69961 ;
  assign n69963 = n69916 & ~n69962 ;
  assign n69964 = ~n69932 & ~n69963 ;
  assign n69965 = ~n69960 & n69964 ;
  assign n69966 = ~n69946 & ~n69965 ;
  assign n69983 = ~n69940 & ~n69966 ;
  assign n69984 = ~n69982 & n69983 ;
  assign n69985 = ~\u0_L1_reg[28]/NET0131  & ~n69984 ;
  assign n69986 = \u0_L1_reg[28]/NET0131  & n69984 ;
  assign n69987 = ~n69985 & ~n69986 ;
  assign n69988 = ~n69388 & ~n69406 ;
  assign n69989 = n69375 & ~n69988 ;
  assign n69990 = ~n69395 & ~n69989 ;
  assign n69991 = n69402 & ~n69990 ;
  assign n69992 = ~n69375 & ~n69382 ;
  assign n69993 = n69404 & n69992 ;
  assign n69994 = ~n69991 & ~n69993 ;
  assign n69995 = ~n69363 & ~n69994 ;
  assign n69997 = n69376 & ~n69388 ;
  assign n69998 = ~n69382 & n69997 ;
  assign n70015 = n69425 & n69430 ;
  assign n70016 = ~n69392 & ~n70015 ;
  assign n70017 = ~n69433 & n70016 ;
  assign n70018 = ~n69998 & n70017 ;
  assign n70019 = ~n69402 & ~n70018 ;
  assign n69996 = n69375 & n69404 ;
  assign n70002 = n69369 & ~n69402 ;
  assign n70003 = n69394 & n70002 ;
  assign n70004 = ~n69996 & ~n70003 ;
  assign n70005 = ~n69998 & n70004 ;
  assign n69999 = ~n69388 & n69992 ;
  assign n70000 = n69402 & n69999 ;
  assign n70001 = n69382 & n69392 ;
  assign n70006 = ~n70000 & ~n70001 ;
  assign n70007 = n70005 & n70006 ;
  assign n70008 = n69363 & ~n70007 ;
  assign n70009 = n69382 & n69418 ;
  assign n70010 = ~n69388 & n70009 ;
  assign n70011 = ~n69427 & ~n70010 ;
  assign n70012 = n69402 & ~n70011 ;
  assign n70013 = ~n69363 & ~n69402 ;
  assign n70014 = n69391 & n70013 ;
  assign n70020 = ~n70012 & ~n70014 ;
  assign n70021 = ~n70008 & n70020 ;
  assign n70022 = ~n70019 & n70021 ;
  assign n70023 = ~n69995 & n70022 ;
  assign n70024 = \u0_L1_reg[15]/P0001  & n70023 ;
  assign n70025 = ~\u0_L1_reg[15]/P0001  & ~n70023 ;
  assign n70026 = ~n70024 & ~n70025 ;
  assign n70031 = ~n69465 & n69512 ;
  assign n70032 = ~n69493 & ~n69515 ;
  assign n70033 = ~n70031 & n70032 ;
  assign n70034 = n69475 & ~n70033 ;
  assign n70027 = n69492 & n69512 ;
  assign n70028 = n69452 & n69495 ;
  assign n70029 = ~n70027 & ~n70028 ;
  assign n70030 = ~n69475 & ~n70029 ;
  assign n70035 = ~n69523 & ~n69527 ;
  assign n70036 = ~n70030 & n70035 ;
  assign n70037 = ~n70034 & n70036 ;
  assign n70038 = ~n69507 & ~n70037 ;
  assign n70050 = ~n69484 & n69488 ;
  assign n70049 = ~n69465 & n70028 ;
  assign n70047 = ~n69465 & n69475 ;
  assign n70048 = n69491 & n70047 ;
  assign n70051 = n69465 & n69529 ;
  assign n70052 = ~n70048 & ~n70051 ;
  assign n70053 = ~n70049 & n70052 ;
  assign n70054 = ~n70050 & n70053 ;
  assign n70055 = n69507 & ~n70054 ;
  assign n70041 = ~n69509 & ~n69530 ;
  assign n70042 = n69475 & ~n69515 ;
  assign n70043 = n70041 & n70042 ;
  assign n70039 = ~n69521 & ~n69522 ;
  assign n70040 = ~n69475 & n70039 ;
  assign n70044 = n69465 & ~n70040 ;
  assign n70045 = ~n70043 & n70044 ;
  assign n70046 = n69488 & n69495 ;
  assign n70056 = ~n70045 & ~n70046 ;
  assign n70057 = ~n70055 & n70056 ;
  assign n70058 = ~n70038 & n70057 ;
  assign n70059 = ~\u0_L1_reg[4]/NET0131  & ~n70058 ;
  assign n70060 = \u0_L1_reg[4]/NET0131  & n70058 ;
  assign n70061 = ~n70059 & ~n70060 ;
  assign n70063 = ~n69375 & n69402 ;
  assign n70064 = n69382 & n69404 ;
  assign n70065 = ~n70063 & n70064 ;
  assign n70073 = ~n69393 & ~n69433 ;
  assign n70074 = ~n70065 & n70073 ;
  assign n70066 = ~n69392 & ~n69412 ;
  assign n70067 = n69402 & ~n70066 ;
  assign n70070 = ~n69363 & ~n69997 ;
  assign n70062 = n69425 & n70002 ;
  assign n70068 = ~n69388 & ~n69402 ;
  assign n70069 = n69411 & n70068 ;
  assign n70071 = ~n70062 & ~n70069 ;
  assign n70072 = n70070 & n70071 ;
  assign n70075 = ~n70067 & n70072 ;
  assign n70076 = n70074 & n70075 ;
  assign n70078 = n69402 & ~n69426 ;
  assign n70077 = n69376 & n69388 ;
  assign n70079 = ~n70009 & ~n70077 ;
  assign n70080 = n70078 & n70079 ;
  assign n70081 = n69388 & n69406 ;
  assign n70082 = ~n69402 & ~n70081 ;
  assign n70083 = ~n70001 & n70082 ;
  assign n70084 = ~n70080 & ~n70083 ;
  assign n70085 = ~n69412 & ~n69999 ;
  assign n70086 = n69369 & ~n70085 ;
  assign n70087 = n69363 & ~n70010 ;
  assign n70088 = ~n70086 & n70087 ;
  assign n70089 = ~n70084 & n70088 ;
  assign n70090 = ~n70076 & ~n70089 ;
  assign n70091 = n69402 & ~n69419 ;
  assign n70092 = n69389 & n69430 ;
  assign n70093 = ~n69402 & ~n70092 ;
  assign n70094 = ~n70091 & ~n70093 ;
  assign n70095 = ~n70090 & ~n70094 ;
  assign n70096 = ~\u0_L1_reg[21]/NET0131  & ~n70095 ;
  assign n70097 = \u0_L1_reg[21]/NET0131  & n70095 ;
  assign n70098 = ~n70096 & ~n70097 ;
  assign n70115 = ~n69466 & ~n69511 ;
  assign n70116 = ~n69482 & ~n70115 ;
  assign n70117 = n70039 & ~n70116 ;
  assign n70118 = n69475 & ~n70117 ;
  assign n70103 = n69465 & n69515 ;
  assign n70119 = ~n69465 & ~n69532 ;
  assign n70120 = ~n70103 & ~n70119 ;
  assign n70121 = ~n69475 & ~n70120 ;
  assign n70122 = ~n70027 & ~n70121 ;
  assign n70123 = ~n70118 & n70122 ;
  assign n70124 = ~n69507 & ~n70123 ;
  assign n70104 = n69465 & ~n69482 ;
  assign n70105 = n69459 & ~n70104 ;
  assign n70106 = ~n70103 & ~n70105 ;
  assign n70107 = n69475 & ~n70106 ;
  assign n70099 = n69465 & ~n69489 ;
  assign n70100 = ~n69512 & n70099 ;
  assign n70101 = ~n69509 & ~n70100 ;
  assign n70102 = ~n69475 & ~n70101 ;
  assign n70108 = n69465 & n69509 ;
  assign n70109 = n69494 & ~n69513 ;
  assign n70110 = ~n70108 & n70109 ;
  assign n70111 = ~n70102 & n70110 ;
  assign n70112 = ~n70107 & n70111 ;
  assign n70113 = n69507 & ~n70112 ;
  assign n70114 = n69529 & n70047 ;
  assign n70125 = ~n69523 & ~n70114 ;
  assign n70126 = ~n70113 & n70125 ;
  assign n70127 = ~n70124 & n70126 ;
  assign n70128 = \u0_L1_reg[29]/NET0131  & ~n70127 ;
  assign n70129 = ~\u0_L1_reg[29]/NET0131  & n70127 ;
  assign n70130 = ~n70128 & ~n70129 ;
  assign n70135 = ~n69931 & ~n69968 ;
  assign n70136 = ~n69915 & n69961 ;
  assign n70137 = ~n69939 & ~n70136 ;
  assign n70138 = ~n70135 & n70137 ;
  assign n70146 = n69909 & n69939 ;
  assign n70147 = n70136 & n70146 ;
  assign n70148 = ~n69946 & ~n70147 ;
  assign n70149 = ~n70138 & n70148 ;
  assign n70139 = ~n69915 & ~n69939 ;
  assign n70140 = ~n69909 & n69929 ;
  assign n70141 = n70139 & n70140 ;
  assign n70142 = n69909 & n69950 ;
  assign n70143 = ~n70141 & ~n70142 ;
  assign n70144 = ~n69961 & ~n69973 ;
  assign n70145 = ~n69909 & n70144 ;
  assign n70150 = n70143 & ~n70145 ;
  assign n70151 = n70149 & n70150 ;
  assign n70157 = n69909 & n69954 ;
  assign n70158 = ~n69962 & n70157 ;
  assign n70153 = ~n69909 & n69915 ;
  assign n70154 = ~n69953 & ~n70153 ;
  assign n70155 = n69939 & ~n70154 ;
  assign n70152 = n69955 & n69973 ;
  assign n70156 = n69947 & n70139 ;
  assign n70159 = n69946 & ~n70156 ;
  assign n70160 = ~n70152 & n70159 ;
  assign n70161 = ~n70155 & n70160 ;
  assign n70162 = ~n70158 & n70161 ;
  assign n70163 = ~n70151 & ~n70162 ;
  assign n70131 = n69923 & ~n69929 ;
  assign n70132 = n69915 & n69955 ;
  assign n70133 = ~n70131 & ~n70132 ;
  assign n70134 = n69939 & ~n70133 ;
  assign n70164 = ~n69916 & ~n70153 ;
  assign n70165 = ~n69939 & n69949 ;
  assign n70166 = n70164 & n70165 ;
  assign n70167 = ~n70134 & ~n70166 ;
  assign n70168 = ~n70163 & n70167 ;
  assign n70169 = \u0_L1_reg[2]/NET0131  & n70168 ;
  assign n70170 = ~\u0_L1_reg[2]/NET0131  & ~n70168 ;
  assign n70171 = ~n70169 & ~n70170 ;
  assign n70183 = ~n69590 & ~n69601 ;
  assign n70184 = n69551 & ~n70183 ;
  assign n70185 = ~n69596 & n69758 ;
  assign n70186 = ~n70184 & n70185 ;
  assign n70187 = n69579 & ~n70186 ;
  assign n70172 = ~n69563 & n69603 ;
  assign n70173 = ~n69614 & ~n70172 ;
  assign n70174 = n69579 & ~n70173 ;
  assign n70178 = ~n69588 & ~n69878 ;
  assign n70175 = ~n69590 & ~n69603 ;
  assign n70176 = n69563 & ~n69579 ;
  assign n70177 = ~n70175 & n70176 ;
  assign n70179 = ~n69624 & ~n70177 ;
  assign n70180 = ~n70178 & n70179 ;
  assign n70181 = ~n70174 & n70180 ;
  assign n70182 = ~n69551 & ~n70181 ;
  assign n70188 = ~n69551 & ~n69626 ;
  assign n70189 = ~n69564 & n69588 ;
  assign n70190 = n69622 & n70189 ;
  assign n70191 = ~n70188 & n70190 ;
  assign n70192 = ~n69612 & ~n69746 ;
  assign n70193 = n69551 & ~n69579 ;
  assign n70194 = ~n69582 & n70193 ;
  assign n70195 = ~n70192 & n70194 ;
  assign n70196 = ~n70191 & ~n70195 ;
  assign n70197 = ~n70182 & n70196 ;
  assign n70198 = ~n70187 & n70197 ;
  assign n70199 = ~\u0_L1_reg[1]/NET0131  & ~n70198 ;
  assign n70200 = \u0_L1_reg[1]/NET0131  & n70198 ;
  assign n70201 = ~n70199 & ~n70200 ;
  assign n70204 = ~n69475 & ~n69529 ;
  assign n70203 = ~n69458 & ~n69483 ;
  assign n70205 = ~n69468 & ~n70203 ;
  assign n70206 = ~n70204 & n70205 ;
  assign n70202 = ~n69475 & ~n70041 ;
  assign n70207 = ~n69507 & ~n70202 ;
  assign n70208 = ~n70206 & n70207 ;
  assign n70210 = n69465 & ~n70041 ;
  assign n70214 = n69507 & ~n69513 ;
  assign n70215 = ~n69518 & n70214 ;
  assign n70209 = n69468 & n69475 ;
  assign n70211 = n69475 & ~n69512 ;
  assign n70212 = ~n69452 & ~n69485 ;
  assign n70213 = ~n70211 & n70212 ;
  assign n70216 = ~n70209 & ~n70213 ;
  assign n70217 = n70215 & n70216 ;
  assign n70218 = ~n70210 & n70217 ;
  assign n70219 = ~n70208 & ~n70218 ;
  assign n70220 = n69517 & ~n69528 ;
  assign n70221 = ~n70219 & n70220 ;
  assign n70222 = ~\u0_L1_reg[19]/NET0131  & ~n70221 ;
  assign n70223 = \u0_L1_reg[19]/NET0131  & n70221 ;
  assign n70224 = ~n70222 & ~n70223 ;
  assign n70225 = n69200 & ~n69215 ;
  assign n70226 = ~n69180 & ~n69248 ;
  assign n70227 = ~n69820 & n70226 ;
  assign n70228 = ~n70225 & n70227 ;
  assign n70229 = n69193 & ~n69214 ;
  assign n70230 = ~n69237 & ~n70229 ;
  assign n70231 = n69180 & ~n69218 ;
  assign n70232 = ~n70230 & n70231 ;
  assign n70233 = ~n70228 & ~n70232 ;
  assign n70234 = n69193 & n69214 ;
  assign n70235 = n69199 & n70234 ;
  assign n70236 = ~n70233 & ~n70235 ;
  assign n70237 = n69174 & ~n70236 ;
  assign n70238 = n69215 & n69236 ;
  assign n70239 = ~n69193 & n69214 ;
  assign n70240 = n69819 & ~n70239 ;
  assign n70246 = ~n70238 & ~n70240 ;
  assign n70241 = ~n69229 & ~n70239 ;
  assign n70242 = n69180 & ~n70241 ;
  assign n70243 = ~n69200 & ~n69236 ;
  assign n70244 = ~n69215 & n69818 ;
  assign n70245 = n70243 & n70244 ;
  assign n70247 = ~n70242 & ~n70245 ;
  assign n70248 = n70246 & n70247 ;
  assign n70249 = ~n69174 & ~n70248 ;
  assign n70250 = n69180 & n69235 ;
  assign n70251 = ~n69214 & n69244 ;
  assign n70252 = n69211 & n70251 ;
  assign n70253 = ~n70250 & ~n70252 ;
  assign n70254 = ~n70249 & n70253 ;
  assign n70255 = ~n70237 & n70254 ;
  assign n70256 = \u0_L1_reg[32]/NET0131  & n70255 ;
  assign n70257 = ~\u0_L1_reg[32]/NET0131  & ~n70255 ;
  assign n70258 = ~n70256 & ~n70257 ;
  assign n70263 = ~n69186 & ~n70243 ;
  assign n70259 = n69199 & ~n69215 ;
  assign n70264 = ~n70234 & ~n70259 ;
  assign n70265 = ~n70263 & n70264 ;
  assign n70266 = ~n69180 & ~n70265 ;
  assign n70260 = ~n69229 & ~n70259 ;
  assign n70261 = n69193 & ~n70260 ;
  assign n70267 = ~n69193 & ~n69217 ;
  assign n70268 = n69215 & n70267 ;
  assign n70269 = n69180 & n70268 ;
  assign n70270 = ~n70261 & ~n70269 ;
  assign n70271 = ~n70266 & n70270 ;
  assign n70272 = n69174 & ~n70271 ;
  assign n70275 = ~n69215 & n69236 ;
  assign n70273 = n69193 & ~n69228 ;
  assign n70274 = n69215 & ~n70273 ;
  assign n70276 = ~n69174 & ~n70274 ;
  assign n70277 = ~n70275 & n70276 ;
  assign n70278 = ~n69219 & ~n70277 ;
  assign n70279 = n69180 & ~n70278 ;
  assign n70262 = ~n69180 & n70261 ;
  assign n70280 = ~n69180 & n70268 ;
  assign n70281 = ~n69219 & ~n70280 ;
  assign n70282 = ~n69174 & ~n70281 ;
  assign n70283 = ~n70262 & ~n70282 ;
  assign n70284 = ~n70279 & n70283 ;
  assign n70285 = ~n70272 & n70284 ;
  assign n70286 = ~\u0_L1_reg[7]/NET0131  & ~n70285 ;
  assign n70287 = \u0_L1_reg[7]/NET0131  & n70285 ;
  assign n70288 = ~n70286 & ~n70287 ;
  assign n70323 = decrypt_pad & ~\u0_uk_K_r1_reg[6]/NET0131  ;
  assign n70324 = ~decrypt_pad & ~\u0_uk_K_r1_reg[55]/NET0131  ;
  assign n70325 = ~n70323 & ~n70324 ;
  assign n70326 = \u0_R1_reg[11]/NET0131  & ~n70325 ;
  assign n70327 = ~\u0_R1_reg[11]/NET0131  & n70325 ;
  assign n70328 = ~n70326 & ~n70327 ;
  assign n70289 = decrypt_pad & ~\u0_uk_K_r1_reg[46]/NET0131  ;
  assign n70290 = ~decrypt_pad & ~\u0_uk_K_r1_reg[13]/NET0131  ;
  assign n70291 = ~n70289 & ~n70290 ;
  assign n70292 = \u0_R1_reg[12]/NET0131  & ~n70291 ;
  assign n70293 = ~\u0_R1_reg[12]/NET0131  & n70291 ;
  assign n70294 = ~n70292 & ~n70293 ;
  assign n70302 = decrypt_pad & ~\u0_uk_K_r1_reg[54]/NET0131  ;
  assign n70303 = ~decrypt_pad & ~\u0_uk_K_r1_reg[46]/NET0131  ;
  assign n70304 = ~n70302 & ~n70303 ;
  assign n70305 = \u0_R1_reg[9]/NET0131  & ~n70304 ;
  assign n70306 = ~\u0_R1_reg[9]/NET0131  & n70304 ;
  assign n70307 = ~n70305 & ~n70306 ;
  assign n70308 = decrypt_pad & ~\u0_uk_K_r1_reg[34]/NET0131  ;
  assign n70309 = ~decrypt_pad & ~\u0_uk_K_r1_reg[26]/NET0131  ;
  assign n70310 = ~n70308 & ~n70309 ;
  assign n70311 = \u0_R1_reg[13]/NET0131  & ~n70310 ;
  assign n70312 = ~\u0_R1_reg[13]/NET0131  & n70310 ;
  assign n70313 = ~n70311 & ~n70312 ;
  assign n70332 = ~n70307 & n70313 ;
  assign n70295 = decrypt_pad & ~\u0_uk_K_r1_reg[5]/NET0131  ;
  assign n70296 = ~decrypt_pad & ~\u0_uk_K_r1_reg[54]/NET0131  ;
  assign n70297 = ~n70295 & ~n70296 ;
  assign n70298 = \u0_R1_reg[10]/NET0131  & ~n70297 ;
  assign n70299 = ~\u0_R1_reg[10]/NET0131  & n70297 ;
  assign n70300 = ~n70298 & ~n70299 ;
  assign n70315 = decrypt_pad & ~\u0_uk_K_r1_reg[25]/NET0131  ;
  assign n70316 = ~decrypt_pad & ~\u0_uk_K_r1_reg[17]/NET0131  ;
  assign n70317 = ~n70315 & ~n70316 ;
  assign n70318 = \u0_R1_reg[8]/NET0131  & ~n70317 ;
  assign n70319 = ~\u0_R1_reg[8]/NET0131  & n70317 ;
  assign n70320 = ~n70318 & ~n70319 ;
  assign n70333 = n70313 & ~n70320 ;
  assign n70334 = n70300 & n70333 ;
  assign n70314 = n70307 & ~n70313 ;
  assign n70335 = n70314 & n70320 ;
  assign n70336 = ~n70334 & ~n70335 ;
  assign n70337 = ~n70332 & n70336 ;
  assign n70338 = n70294 & ~n70337 ;
  assign n70329 = ~n70313 & ~n70320 ;
  assign n70330 = ~n70300 & ~n70307 ;
  assign n70331 = n70329 & n70330 ;
  assign n70339 = n70300 & ~n70307 ;
  assign n70340 = n70313 & n70339 ;
  assign n70341 = ~n70331 & ~n70340 ;
  assign n70342 = ~n70338 & n70341 ;
  assign n70343 = n70328 & ~n70342 ;
  assign n70344 = ~n70300 & n70307 ;
  assign n70347 = ~n70339 & ~n70344 ;
  assign n70345 = ~n70320 & n70328 ;
  assign n70348 = n70313 & n70320 ;
  assign n70349 = ~n70329 & ~n70348 ;
  assign n70350 = ~n70345 & n70349 ;
  assign n70351 = n70347 & n70350 ;
  assign n70346 = n70344 & n70345 ;
  assign n70352 = ~n70347 & ~n70349 ;
  assign n70353 = ~n70346 & ~n70352 ;
  assign n70354 = ~n70351 & n70353 ;
  assign n70355 = ~n70294 & ~n70354 ;
  assign n70301 = n70294 & n70300 ;
  assign n70321 = n70314 & ~n70320 ;
  assign n70322 = n70301 & n70321 ;
  assign n70356 = n70320 & ~n70332 ;
  assign n70357 = ~n70344 & ~n70356 ;
  assign n70358 = ~n70314 & ~n70328 ;
  assign n70359 = n70294 & n70358 ;
  assign n70360 = ~n70357 & n70359 ;
  assign n70361 = ~n70322 & ~n70360 ;
  assign n70362 = ~n70355 & n70361 ;
  assign n70363 = ~n70343 & n70362 ;
  assign n70364 = ~\u0_L1_reg[6]/NET0131  & ~n70363 ;
  assign n70365 = \u0_L1_reg[6]/NET0131  & n70363 ;
  assign n70366 = ~n70364 & ~n70365 ;
  assign n70381 = ~n69405 & n69989 ;
  assign n70382 = n69402 & ~n70381 ;
  assign n70383 = ~n69412 & ~n69426 ;
  assign n70384 = n69420 & n70383 ;
  assign n70385 = ~n70382 & ~n70384 ;
  assign n70386 = ~n69393 & ~n70009 ;
  assign n70387 = ~n69427 & n70386 ;
  assign n70388 = ~n70385 & n70387 ;
  assign n70389 = n69363 & ~n70388 ;
  assign n70370 = n69402 & ~n69997 ;
  assign n70368 = n69382 & ~n69430 ;
  assign n70369 = ~n69382 & n69430 ;
  assign n70371 = ~n70368 & ~n70369 ;
  assign n70372 = n70370 & n70371 ;
  assign n70367 = n69389 & n70002 ;
  assign n70373 = ~n70069 & ~n70367 ;
  assign n70374 = ~n69434 & n70373 ;
  assign n70375 = ~n70372 & n70374 ;
  assign n70376 = ~n69363 & ~n70375 ;
  assign n70377 = ~n69413 & ~n69432 ;
  assign n70378 = ~n69402 & ~n70377 ;
  assign n70379 = n69369 & n69402 ;
  assign n70380 = n69992 & n70379 ;
  assign n70390 = ~n70378 & ~n70380 ;
  assign n70391 = ~n70376 & n70390 ;
  assign n70392 = ~n70389 & n70391 ;
  assign n70393 = ~\u0_L1_reg[27]/NET0131  & ~n70392 ;
  assign n70394 = \u0_L1_reg[27]/NET0131  & n70392 ;
  assign n70395 = ~n70393 & ~n70394 ;
  assign n70400 = ~n69326 & n69346 ;
  assign n70401 = n69345 & ~n70400 ;
  assign n70403 = ~n69266 & n69272 ;
  assign n70404 = ~n69286 & n70403 ;
  assign n70405 = ~n69294 & n70404 ;
  assign n70402 = ~n69293 & n69846 ;
  assign n70406 = ~n69307 & ~n70402 ;
  assign n70407 = ~n70405 & n70406 ;
  assign n70408 = ~n70401 & n70407 ;
  assign n70410 = n69307 & ~n69858 ;
  assign n70411 = ~n69330 & n70410 ;
  assign n70409 = n69293 & n69846 ;
  assign n70412 = ~n69336 & ~n70409 ;
  assign n70413 = n70411 & n70412 ;
  assign n70414 = ~n70408 & ~n70413 ;
  assign n70397 = ~n69285 & n69853 ;
  assign n70398 = ~n69342 & ~n70397 ;
  assign n70399 = ~n69266 & ~n70398 ;
  assign n70415 = n69279 & n69848 ;
  assign n70416 = ~n69849 & ~n70415 ;
  assign n70417 = n69272 & ~n69344 ;
  assign n70418 = ~n69266 & n69307 ;
  assign n70419 = ~n70417 & n70418 ;
  assign n70420 = n70416 & n70419 ;
  assign n70396 = n69266 & n69325 ;
  assign n70421 = ~n69287 & ~n70396 ;
  assign n70422 = ~n70420 & n70421 ;
  assign n70423 = ~n70399 & n70422 ;
  assign n70424 = ~n70414 & n70423 ;
  assign n70425 = \u0_L1_reg[23]/NET0131  & ~n70424 ;
  assign n70426 = ~\u0_L1_reg[23]/NET0131  & n70424 ;
  assign n70427 = ~n70425 & ~n70426 ;
  assign n70435 = ~n69915 & n69956 ;
  assign n70436 = ~n69971 & ~n69978 ;
  assign n70437 = ~n70435 & n70436 ;
  assign n70438 = ~n69939 & ~n70437 ;
  assign n70428 = n69939 & ~n69949 ;
  assign n70429 = ~n69955 & n70428 ;
  assign n70430 = ~n69930 & n70429 ;
  assign n70431 = n69939 & ~n69947 ;
  assign n70432 = ~n69973 & n70431 ;
  assign n70433 = ~n69950 & ~n70432 ;
  assign n70434 = ~n69909 & ~n70433 ;
  assign n70439 = ~n70430 & ~n70434 ;
  assign n70440 = ~n70438 & n70439 ;
  assign n70441 = ~n69946 & ~n70440 ;
  assign n70442 = n69961 & n70153 ;
  assign n70443 = ~n69932 & ~n70442 ;
  assign n70444 = ~n69939 & ~n70443 ;
  assign n70445 = ~n69915 & ~n69929 ;
  assign n70446 = n69909 & n70445 ;
  assign n70447 = n70137 & ~n70446 ;
  assign n70448 = ~n69909 & n70445 ;
  assign n70449 = n69939 & ~n69977 ;
  assign n70450 = ~n70448 & n70449 ;
  assign n70451 = ~n70447 & ~n70450 ;
  assign n70452 = n69915 & n69948 ;
  assign n70453 = n70443 & ~n70452 ;
  assign n70454 = n70143 & n70453 ;
  assign n70455 = ~n70451 & n70454 ;
  assign n70456 = n69946 & ~n70455 ;
  assign n70457 = ~n70444 & ~n70456 ;
  assign n70458 = ~n70441 & n70457 ;
  assign n70459 = ~\u0_L1_reg[13]/NET0131  & n70458 ;
  assign n70460 = \u0_L1_reg[13]/NET0131  & ~n70458 ;
  assign n70461 = ~n70459 & ~n70460 ;
  assign n70474 = ~n69665 & n69688 ;
  assign n70475 = ~n69796 & ~n70474 ;
  assign n70476 = n69646 & ~n70475 ;
  assign n70477 = ~n69665 & n69716 ;
  assign n70478 = ~n69728 & ~n70477 ;
  assign n70479 = ~n70476 & n70478 ;
  assign n70480 = n69705 & ~n70479 ;
  assign n70463 = n69646 & ~n69673 ;
  assign n70464 = ~n69800 & n70463 ;
  assign n70465 = n69676 & ~n69695 ;
  assign n70466 = n69797 & ~n70465 ;
  assign n70467 = ~n70464 & ~n70466 ;
  assign n70468 = ~n69685 & n69778 ;
  assign n70469 = ~n70467 & n70468 ;
  assign n70470 = ~n69705 & ~n70469 ;
  assign n70462 = ~n69658 & n69782 ;
  assign n70471 = n69676 & n69707 ;
  assign n70472 = ~n69675 & ~n70471 ;
  assign n70473 = n69646 & ~n70472 ;
  assign n70481 = ~n70462 & ~n70473 ;
  assign n70482 = ~n70470 & n70481 ;
  assign n70483 = ~n70480 & n70482 ;
  assign n70484 = ~\u0_L1_reg[8]/NET0131  & ~n70483 ;
  assign n70485 = \u0_L1_reg[8]/NET0131  & n70483 ;
  assign n70486 = ~n70484 & ~n70485 ;
  assign n70489 = n70300 & n70320 ;
  assign n70499 = ~n70307 & n70489 ;
  assign n70500 = ~n70313 & n70499 ;
  assign n70501 = n70300 & n70329 ;
  assign n70502 = ~n70300 & n70333 ;
  assign n70503 = ~n70501 & ~n70502 ;
  assign n70504 = ~n70321 & ~n70499 ;
  assign n70505 = n70503 & n70504 ;
  assign n70506 = n70328 & ~n70505 ;
  assign n70507 = ~n70500 & ~n70506 ;
  assign n70508 = ~n70294 & ~n70507 ;
  assign n70490 = n70307 & n70489 ;
  assign n70488 = n70330 & ~n70333 ;
  assign n70491 = ~n70334 & ~n70488 ;
  assign n70492 = ~n70490 & n70491 ;
  assign n70493 = n70328 & ~n70492 ;
  assign n70487 = n70330 & n70350 ;
  assign n70494 = ~n70328 & ~n70330 ;
  assign n70495 = ~n70349 & n70494 ;
  assign n70496 = ~n70487 & ~n70495 ;
  assign n70497 = ~n70493 & n70496 ;
  assign n70498 = n70294 & ~n70497 ;
  assign n70517 = n70330 & ~n70349 ;
  assign n70518 = n70336 & ~n70517 ;
  assign n70519 = ~n70294 & ~n70328 ;
  assign n70520 = ~n70518 & n70519 ;
  assign n70513 = ~n70300 & ~n70313 ;
  assign n70514 = n70320 & n70513 ;
  assign n70515 = ~n70307 & n70328 ;
  assign n70516 = n70514 & n70515 ;
  assign n70509 = n70307 & n70348 ;
  assign n70510 = n70300 & ~n70328 ;
  assign n70511 = n70509 & n70510 ;
  assign n70512 = n70313 & n70346 ;
  assign n70521 = ~n70511 & ~n70512 ;
  assign n70522 = ~n70516 & n70521 ;
  assign n70523 = ~n70520 & n70522 ;
  assign n70524 = ~n70498 & n70523 ;
  assign n70525 = ~n70508 & n70524 ;
  assign n70526 = ~\u0_L1_reg[24]/NET0131  & ~n70525 ;
  assign n70527 = \u0_L1_reg[24]/NET0131  & n70525 ;
  assign n70528 = ~n70526 & ~n70527 ;
  assign n70531 = ~n70314 & n70489 ;
  assign n70532 = n70307 & n70513 ;
  assign n70533 = ~n70531 & ~n70532 ;
  assign n70534 = n70328 & ~n70533 ;
  assign n70535 = ~n70307 & ~n70320 ;
  assign n70536 = ~n70489 & ~n70535 ;
  assign n70537 = n70358 & n70536 ;
  assign n70538 = n70333 & n70339 ;
  assign n70539 = ~n70294 & ~n70538 ;
  assign n70540 = ~n70517 & n70539 ;
  assign n70541 = ~n70537 & n70540 ;
  assign n70542 = ~n70534 & n70541 ;
  assign n70544 = ~n70321 & ~n70489 ;
  assign n70545 = ~n70328 & ~n70544 ;
  assign n70543 = n70328 & ~n70503 ;
  assign n70546 = n70294 & ~n70516 ;
  assign n70547 = ~n70543 & n70546 ;
  assign n70548 = ~n70545 & n70547 ;
  assign n70549 = ~n70542 & ~n70548 ;
  assign n70529 = n70307 & ~n70348 ;
  assign n70530 = n70301 & n70529 ;
  assign n70550 = ~n70307 & n70348 ;
  assign n70551 = n70328 & ~n70550 ;
  assign n70552 = n70300 & ~n70358 ;
  assign n70553 = ~n70551 & n70552 ;
  assign n70554 = ~n70530 & ~n70553 ;
  assign n70555 = ~n70549 & n70554 ;
  assign n70556 = \u0_L1_reg[30]/NET0131  & ~n70555 ;
  assign n70557 = ~\u0_L1_reg[30]/NET0131  & n70555 ;
  assign n70558 = ~n70556 & ~n70557 ;
  assign n70562 = ~n69665 & n69676 ;
  assign n70563 = ~n69712 & ~n70562 ;
  assign n70564 = n69646 & ~n70563 ;
  assign n70559 = ~n69687 & ~n69689 ;
  assign n70560 = ~n69796 & n70559 ;
  assign n70561 = ~n69646 & ~n70560 ;
  assign n70565 = ~n69659 & n69695 ;
  assign n70566 = ~n69705 & ~n70565 ;
  assign n70567 = ~n70561 & n70566 ;
  assign n70568 = ~n70564 & n70567 ;
  assign n70570 = ~n69709 & ~n69726 ;
  assign n70571 = n69646 & ~n70570 ;
  assign n70573 = ~n69680 & n69705 ;
  assign n70569 = n69665 & n69784 ;
  assign n70572 = ~n69646 & n69722 ;
  assign n70574 = ~n70569 & ~n70572 ;
  assign n70575 = n70573 & n70574 ;
  assign n70576 = ~n70571 & n70575 ;
  assign n70577 = ~n70568 & ~n70576 ;
  assign n70578 = n69676 & n69695 ;
  assign n70579 = n70463 & ~n70578 ;
  assign n70580 = ~n69646 & ~n69696 ;
  assign n70581 = ~n69733 & n70580 ;
  assign n70582 = ~n70474 & n70581 ;
  assign n70583 = ~n70579 & ~n70582 ;
  assign n70584 = ~n70577 & ~n70583 ;
  assign n70585 = ~\u0_L1_reg[3]/NET0131  & ~n70584 ;
  assign n70586 = \u0_L1_reg[3]/NET0131  & n70584 ;
  assign n70587 = ~n70585 & ~n70586 ;
  assign n70589 = ~n70529 & ~n70550 ;
  assign n70590 = ~n70329 & n70589 ;
  assign n70591 = n70314 & n70345 ;
  assign n70592 = ~n70590 & ~n70591 ;
  assign n70593 = ~n70300 & ~n70592 ;
  assign n70588 = n70307 & n70334 ;
  assign n70594 = ~n70501 & ~n70514 ;
  assign n70595 = ~n70328 & ~n70594 ;
  assign n70596 = ~n70588 & ~n70595 ;
  assign n70597 = ~n70593 & n70596 ;
  assign n70598 = n70294 & ~n70597 ;
  assign n70599 = ~n70332 & ~n70513 ;
  assign n70600 = ~n70320 & ~n70599 ;
  assign n70601 = ~n70509 & ~n70600 ;
  assign n70602 = ~n70294 & ~n70601 ;
  assign n70611 = ~n70499 & ~n70602 ;
  assign n70612 = ~n70328 & ~n70611 ;
  assign n70603 = n70331 & n70602 ;
  assign n70604 = ~n70313 & n70535 ;
  assign n70605 = ~n70335 & ~n70604 ;
  assign n70606 = n70300 & ~n70605 ;
  assign n70607 = ~n70294 & ~n70329 ;
  assign n70608 = ~n70589 & n70607 ;
  assign n70609 = ~n70606 & ~n70608 ;
  assign n70610 = n70328 & ~n70609 ;
  assign n70613 = ~n70603 & ~n70610 ;
  assign n70614 = ~n70612 & n70613 ;
  assign n70615 = ~n70598 & n70614 ;
  assign n70616 = ~\u0_L1_reg[16]/NET0131  & ~n70615 ;
  assign n70617 = \u0_L1_reg[16]/NET0131  & n70615 ;
  assign n70618 = ~n70616 & ~n70617 ;
  assign n70621 = ~n69321 & ~n69849 ;
  assign n70622 = ~n69286 & ~n70621 ;
  assign n70623 = ~n69293 & n69295 ;
  assign n70624 = n69266 & n69346 ;
  assign n70625 = ~n70623 & n70624 ;
  assign n70619 = ~n69320 & ~n69346 ;
  assign n70620 = ~n69266 & n70619 ;
  assign n70626 = ~n69307 & ~n70620 ;
  assign n70627 = ~n70625 & n70626 ;
  assign n70628 = ~n70622 & n70627 ;
  assign n70630 = n69285 & n70416 ;
  assign n70629 = n69312 & n70619 ;
  assign n70631 = n69863 & ~n70629 ;
  assign n70632 = ~n70630 & n70631 ;
  assign n70633 = ~n70628 & ~n70632 ;
  assign n70634 = ~n69266 & n69308 ;
  assign n70635 = ~n69337 & n70634 ;
  assign n70636 = ~n70633 & ~n70635 ;
  assign n70637 = ~\u0_L1_reg[9]/NET0131  & ~n70636 ;
  assign n70638 = \u0_L1_reg[9]/NET0131  & n70636 ;
  assign n70639 = ~n70637 & ~n70638 ;
  assign n70642 = n69939 & n70144 ;
  assign n70643 = ~n70140 & ~n70445 ;
  assign n70644 = n69922 & ~n69939 ;
  assign n70645 = ~n70643 & n70644 ;
  assign n70646 = n69946 & ~n70131 ;
  assign n70647 = ~n70645 & n70646 ;
  assign n70648 = ~n70642 & n70647 ;
  assign n70649 = n69929 & n69939 ;
  assign n70650 = n69953 & n70649 ;
  assign n70654 = ~n69946 & ~n70448 ;
  assign n70655 = ~n70650 & n70654 ;
  assign n70651 = n69931 & ~n69973 ;
  assign n70652 = ~n69922 & ~n70146 ;
  assign n70653 = n70164 & n70652 ;
  assign n70656 = ~n70651 & ~n70653 ;
  assign n70657 = n70655 & n70656 ;
  assign n70658 = ~n70648 & ~n70657 ;
  assign n70640 = ~n69929 & ~n70153 ;
  assign n70641 = n70429 & ~n70640 ;
  assign n70659 = ~n69939 & n69950 ;
  assign n70660 = ~n70641 & ~n70659 ;
  assign n70661 = ~n70658 & n70660 ;
  assign n70662 = \u0_L1_reg[18]/NET0131  & n70661 ;
  assign n70663 = ~\u0_L1_reg[18]/NET0131  & ~n70661 ;
  assign n70664 = ~n70662 & ~n70663 ;
  assign n70702 = decrypt_pad & ~\u0_uk_K_r0_reg[24]/P0001  ;
  assign n70703 = ~decrypt_pad & ~\u0_uk_K_r0_reg[20]/NET0131  ;
  assign n70704 = ~n70702 & ~n70703 ;
  assign n70705 = \u0_R0_reg[4]/NET0131  & ~n70704 ;
  assign n70706 = ~\u0_R0_reg[4]/NET0131  & n70704 ;
  assign n70707 = ~n70705 & ~n70706 ;
  assign n70685 = decrypt_pad & ~\u0_uk_K_r0_reg[54]/NET0131  ;
  assign n70686 = ~decrypt_pad & ~\u0_uk_K_r0_reg[18]/NET0131  ;
  assign n70687 = ~n70685 & ~n70686 ;
  assign n70688 = \u0_R0_reg[1]/NET0131  & ~n70687 ;
  assign n70689 = ~\u0_R0_reg[1]/NET0131  & n70687 ;
  assign n70690 = ~n70688 & ~n70689 ;
  assign n70665 = decrypt_pad & ~\u0_uk_K_r0_reg[33]/NET0131  ;
  assign n70666 = ~decrypt_pad & ~\u0_uk_K_r0_reg[54]/NET0131  ;
  assign n70667 = ~n70665 & ~n70666 ;
  assign n70668 = \u0_R0_reg[32]/NET0131  & ~n70667 ;
  assign n70669 = ~\u0_R0_reg[32]/NET0131  & n70667 ;
  assign n70670 = ~n70668 & ~n70669 ;
  assign n70671 = decrypt_pad & ~\u0_uk_K_r0_reg[12]/NET0131  ;
  assign n70672 = ~decrypt_pad & ~\u0_uk_K_r0_reg[33]/NET0131  ;
  assign n70673 = ~n70671 & ~n70672 ;
  assign n70674 = \u0_R0_reg[2]/NET0131  & ~n70673 ;
  assign n70675 = ~\u0_R0_reg[2]/NET0131  & n70673 ;
  assign n70676 = ~n70674 & ~n70675 ;
  assign n70677 = ~n70670 & n70676 ;
  assign n70678 = decrypt_pad & ~\u0_uk_K_r0_reg[46]/NET0131  ;
  assign n70679 = ~decrypt_pad & ~\u0_uk_K_r0_reg[10]/NET0131  ;
  assign n70680 = ~n70678 & ~n70679 ;
  assign n70681 = \u0_R0_reg[3]/NET0131  & ~n70680 ;
  assign n70682 = ~\u0_R0_reg[3]/NET0131  & n70680 ;
  assign n70683 = ~n70681 & ~n70682 ;
  assign n70684 = n70677 & n70683 ;
  assign n70691 = decrypt_pad & ~\u0_uk_K_r0_reg[27]/NET0131  ;
  assign n70692 = ~decrypt_pad & ~\u0_uk_K_r0_reg[48]/NET0131  ;
  assign n70693 = ~n70691 & ~n70692 ;
  assign n70694 = \u0_R0_reg[5]/NET0131  & ~n70693 ;
  assign n70695 = ~\u0_R0_reg[5]/NET0131  & n70693 ;
  assign n70696 = ~n70694 & ~n70695 ;
  assign n70721 = n70684 & n70696 ;
  assign n70722 = ~n70670 & ~n70696 ;
  assign n70723 = ~n70676 & n70722 ;
  assign n70724 = ~n70721 & ~n70723 ;
  assign n70725 = n70690 & ~n70724 ;
  assign n70715 = n70670 & ~n70676 ;
  assign n70716 = ~n70677 & ~n70715 ;
  assign n70717 = ~n70683 & n70716 ;
  assign n70708 = n70670 & n70690 ;
  assign n70718 = ~n70690 & n70696 ;
  assign n70719 = ~n70708 & ~n70718 ;
  assign n70720 = n70717 & n70719 ;
  assign n70709 = n70676 & ~n70696 ;
  assign n70710 = n70708 & n70709 ;
  assign n70711 = n70670 & n70696 ;
  assign n70712 = ~n70676 & n70711 ;
  assign n70713 = ~n70710 & ~n70712 ;
  assign n70714 = n70683 & ~n70713 ;
  assign n70726 = n70715 & n70718 ;
  assign n70727 = ~n70714 & ~n70726 ;
  assign n70728 = ~n70720 & n70727 ;
  assign n70729 = ~n70725 & n70728 ;
  assign n70730 = ~n70707 & ~n70729 ;
  assign n70731 = n70676 & n70722 ;
  assign n70732 = ~n70718 & ~n70731 ;
  assign n70733 = n70683 & ~n70732 ;
  assign n70739 = ~n70676 & n70683 ;
  assign n70740 = n70690 & ~n70739 ;
  assign n70741 = ~n70670 & n70696 ;
  assign n70742 = ~n70740 & n70741 ;
  assign n70734 = ~n70670 & n70690 ;
  assign n70735 = ~n70683 & n70690 ;
  assign n70736 = ~n70677 & ~n70735 ;
  assign n70737 = ~n70734 & ~n70736 ;
  assign n70697 = ~n70690 & ~n70696 ;
  assign n70738 = n70697 & n70715 ;
  assign n70743 = ~n70737 & ~n70738 ;
  assign n70744 = ~n70742 & n70743 ;
  assign n70745 = ~n70733 & n70744 ;
  assign n70746 = n70707 & ~n70745 ;
  assign n70749 = n70676 & n70711 ;
  assign n70750 = n70690 & n70749 ;
  assign n70747 = n70690 & ~n70696 ;
  assign n70748 = ~n70676 & n70747 ;
  assign n70751 = n70677 & n70718 ;
  assign n70752 = ~n70748 & ~n70751 ;
  assign n70753 = ~n70750 & n70752 ;
  assign n70754 = ~n70683 & ~n70753 ;
  assign n70698 = n70684 & n70697 ;
  assign n70699 = ~n70676 & ~n70690 ;
  assign n70700 = n70670 & n70683 ;
  assign n70701 = n70699 & n70700 ;
  assign n70755 = ~n70698 & ~n70701 ;
  assign n70756 = ~n70754 & n70755 ;
  assign n70757 = ~n70746 & n70756 ;
  assign n70758 = ~n70730 & n70757 ;
  assign n70759 = ~\u0_L0_reg[31]/NET0131  & ~n70758 ;
  assign n70760 = \u0_L0_reg[31]/NET0131  & n70758 ;
  assign n70761 = ~n70759 & ~n70760 ;
  assign n70817 = decrypt_pad & ~\u0_uk_K_r0_reg[21]/NET0131  ;
  assign n70818 = ~decrypt_pad & ~\u0_uk_K_r0_reg[42]/NET0131  ;
  assign n70819 = ~n70817 & ~n70818 ;
  assign n70820 = \u0_R0_reg[24]/NET0131  & ~n70819 ;
  assign n70821 = ~\u0_R0_reg[24]/NET0131  & n70819 ;
  assign n70822 = ~n70820 & ~n70821 ;
  assign n70775 = decrypt_pad & ~\u0_uk_K_r0_reg[37]/NET0131  ;
  assign n70776 = ~decrypt_pad & ~\u0_uk_K_r0_reg[31]/NET0131  ;
  assign n70777 = ~n70775 & ~n70776 ;
  assign n70778 = \u0_R0_reg[22]/NET0131  & ~n70777 ;
  assign n70779 = ~\u0_R0_reg[22]/NET0131  & n70777 ;
  assign n70780 = ~n70778 & ~n70779 ;
  assign n70762 = decrypt_pad & ~\u0_uk_K_r0_reg[15]/NET0131  ;
  assign n70763 = ~decrypt_pad & ~\u0_uk_K_r0_reg[36]/NET0131  ;
  assign n70764 = ~n70762 & ~n70763 ;
  assign n70765 = \u0_R0_reg[21]/NET0131  & ~n70764 ;
  assign n70766 = ~\u0_R0_reg[21]/NET0131  & n70764 ;
  assign n70767 = ~n70765 & ~n70766 ;
  assign n70768 = decrypt_pad & ~\u0_uk_K_r0_reg[0]/NET0131  ;
  assign n70769 = ~decrypt_pad & ~\u0_uk_K_r0_reg[21]/NET0131  ;
  assign n70770 = ~n70768 & ~n70769 ;
  assign n70771 = \u0_R0_reg[20]/NET0131  & ~n70770 ;
  assign n70772 = ~\u0_R0_reg[20]/NET0131  & n70770 ;
  assign n70773 = ~n70771 & ~n70772 ;
  assign n70774 = n70767 & ~n70773 ;
  assign n70792 = decrypt_pad & ~\u0_uk_K_r0_reg[16]/NET0131  ;
  assign n70793 = ~decrypt_pad & ~\u0_uk_K_r0_reg[37]/NET0131  ;
  assign n70794 = ~n70792 & ~n70793 ;
  assign n70795 = \u0_R0_reg[25]/NET0131  & ~n70794 ;
  assign n70796 = ~\u0_R0_reg[25]/NET0131  & n70794 ;
  assign n70797 = ~n70795 & ~n70796 ;
  assign n70806 = n70773 & n70797 ;
  assign n70847 = ~n70774 & ~n70806 ;
  assign n70848 = n70780 & ~n70847 ;
  assign n70785 = decrypt_pad & ~\u0_uk_K_r0_reg[50]/NET0131  ;
  assign n70786 = ~decrypt_pad & ~\u0_uk_K_r0_reg[16]/NET0131  ;
  assign n70787 = ~n70785 & ~n70786 ;
  assign n70788 = \u0_R0_reg[23]/NET0131  & ~n70787 ;
  assign n70789 = ~\u0_R0_reg[23]/NET0131  & n70787 ;
  assign n70790 = ~n70788 & ~n70789 ;
  assign n70844 = n70767 & n70797 ;
  assign n70845 = ~n70773 & n70844 ;
  assign n70846 = ~n70780 & ~n70845 ;
  assign n70849 = ~n70790 & ~n70846 ;
  assign n70850 = ~n70848 & n70849 ;
  assign n70804 = n70773 & ~n70797 ;
  assign n70837 = ~n70767 & n70804 ;
  assign n70838 = ~n70780 & n70837 ;
  assign n70781 = n70774 & n70780 ;
  assign n70836 = n70767 & n70806 ;
  assign n70839 = ~n70781 & ~n70836 ;
  assign n70840 = ~n70838 & n70839 ;
  assign n70841 = n70790 & ~n70840 ;
  assign n70803 = ~n70780 & ~n70790 ;
  assign n70842 = n70803 & n70806 ;
  assign n70843 = ~n70767 & n70842 ;
  assign n70851 = ~n70841 & ~n70843 ;
  assign n70852 = ~n70850 & n70851 ;
  assign n70853 = n70822 & ~n70852 ;
  assign n70782 = n70773 & ~n70780 ;
  assign n70783 = n70767 & n70782 ;
  assign n70784 = ~n70781 & ~n70783 ;
  assign n70791 = ~n70784 & ~n70790 ;
  assign n70811 = ~n70782 & n70790 ;
  assign n70810 = ~n70773 & ~n70797 ;
  assign n70812 = ~n70767 & ~n70810 ;
  assign n70813 = n70811 & n70812 ;
  assign n70798 = n70767 & ~n70797 ;
  assign n70799 = n70773 & ~n70798 ;
  assign n70800 = ~n70773 & ~n70790 ;
  assign n70801 = ~n70780 & ~n70800 ;
  assign n70802 = ~n70799 & n70801 ;
  assign n70805 = n70803 & n70804 ;
  assign n70807 = ~n70767 & n70780 ;
  assign n70808 = n70806 & n70807 ;
  assign n70809 = ~n70805 & ~n70808 ;
  assign n70814 = ~n70802 & n70809 ;
  assign n70815 = ~n70813 & n70814 ;
  assign n70816 = ~n70791 & n70815 ;
  assign n70823 = ~n70816 & ~n70822 ;
  assign n70833 = ~n70780 & n70798 ;
  assign n70834 = ~n70806 & ~n70833 ;
  assign n70835 = n70811 & ~n70834 ;
  assign n70824 = ~n70767 & n70810 ;
  assign n70825 = n70803 & n70824 ;
  assign n70826 = ~n70767 & ~n70780 ;
  assign n70827 = ~n70773 & n70797 ;
  assign n70828 = n70826 & n70827 ;
  assign n70829 = n70790 & n70828 ;
  assign n70830 = n70767 & n70804 ;
  assign n70831 = n70803 & n70830 ;
  assign n70832 = ~n70829 & ~n70831 ;
  assign n70854 = ~n70825 & n70832 ;
  assign n70855 = ~n70835 & n70854 ;
  assign n70856 = ~n70823 & n70855 ;
  assign n70857 = ~n70853 & n70856 ;
  assign n70858 = \u0_L0_reg[11]/NET0131  & ~n70857 ;
  assign n70859 = ~\u0_L0_reg[11]/NET0131  & n70857 ;
  assign n70860 = ~n70858 & ~n70859 ;
  assign n70861 = decrypt_pad & ~\u0_uk_K_r0_reg[28]/NET0131  ;
  assign n70862 = ~decrypt_pad & ~\u0_uk_K_r0_reg[49]/NET0131  ;
  assign n70863 = ~n70861 & ~n70862 ;
  assign n70864 = \u0_R0_reg[28]/NET0131  & ~n70863 ;
  assign n70865 = ~\u0_R0_reg[28]/NET0131  & n70863 ;
  assign n70866 = ~n70864 & ~n70865 ;
  assign n70897 = decrypt_pad & ~\u0_uk_K_r0_reg[45]/NET0131  ;
  assign n70898 = ~decrypt_pad & ~\u0_uk_K_r0_reg[7]/NET0131  ;
  assign n70899 = ~n70897 & ~n70898 ;
  assign n70900 = \u0_R0_reg[27]/NET0131  & ~n70899 ;
  assign n70901 = ~\u0_R0_reg[27]/NET0131  & n70899 ;
  assign n70902 = ~n70900 & ~n70901 ;
  assign n70867 = decrypt_pad & ~\u0_uk_K_r0_reg[8]/NET0131  ;
  assign n70868 = ~decrypt_pad & ~\u0_uk_K_r0_reg[29]/NET0131  ;
  assign n70869 = ~n70867 & ~n70868 ;
  assign n70870 = \u0_R0_reg[26]/NET0131  & ~n70869 ;
  assign n70871 = ~\u0_R0_reg[26]/NET0131  & n70869 ;
  assign n70872 = ~n70870 & ~n70871 ;
  assign n70873 = decrypt_pad & ~\u0_uk_K_r0_reg[43]/NET0131  ;
  assign n70874 = ~decrypt_pad & ~\u0_uk_K_r0_reg[9]/NET0131  ;
  assign n70875 = ~n70873 & ~n70874 ;
  assign n70876 = \u0_R0_reg[24]/NET0131  & ~n70875 ;
  assign n70877 = ~\u0_R0_reg[24]/NET0131  & n70875 ;
  assign n70878 = ~n70876 & ~n70877 ;
  assign n70882 = decrypt_pad & ~\u0_uk_K_r0_reg[51]/NET0131  ;
  assign n70883 = ~decrypt_pad & ~\u0_uk_K_r0_reg[45]/NET0131  ;
  assign n70884 = ~n70882 & ~n70883 ;
  assign n70885 = \u0_R0_reg[29]/NET0131  & ~n70884 ;
  assign n70886 = ~\u0_R0_reg[29]/NET0131  & n70884 ;
  assign n70887 = ~n70885 & ~n70886 ;
  assign n70910 = n70878 & ~n70887 ;
  assign n70911 = n70872 & ~n70910 ;
  assign n70888 = decrypt_pad & ~\u0_uk_K_r0_reg[23]/NET0131  ;
  assign n70889 = ~decrypt_pad & ~\u0_uk_K_r0_reg[44]/NET0131  ;
  assign n70890 = ~n70888 & ~n70889 ;
  assign n70891 = \u0_R0_reg[25]/NET0131  & ~n70890 ;
  assign n70892 = ~\u0_R0_reg[25]/NET0131  & n70890 ;
  assign n70893 = ~n70891 & ~n70892 ;
  assign n70904 = ~n70887 & ~n70893 ;
  assign n70912 = ~n70878 & ~n70904 ;
  assign n70913 = n70911 & ~n70912 ;
  assign n70914 = n70878 & n70893 ;
  assign n70915 = ~n70887 & n70914 ;
  assign n70916 = ~n70913 & ~n70915 ;
  assign n70917 = ~n70902 & ~n70916 ;
  assign n70879 = n70872 & n70878 ;
  assign n70880 = ~n70872 & ~n70878 ;
  assign n70881 = ~n70879 & ~n70880 ;
  assign n70894 = n70887 & n70893 ;
  assign n70895 = ~n70881 & n70894 ;
  assign n70896 = ~n70878 & n70887 ;
  assign n70903 = n70896 & ~n70902 ;
  assign n70905 = ~n70893 & n70902 ;
  assign n70906 = ~n70904 & ~n70905 ;
  assign n70907 = n70878 & ~n70906 ;
  assign n70908 = ~n70903 & ~n70907 ;
  assign n70909 = ~n70872 & ~n70908 ;
  assign n70918 = ~n70895 & ~n70909 ;
  assign n70919 = ~n70917 & n70918 ;
  assign n70920 = ~n70866 & ~n70919 ;
  assign n70926 = n70887 & ~n70893 ;
  assign n70927 = n70878 & n70926 ;
  assign n70928 = ~n70872 & n70927 ;
  assign n70929 = ~n70878 & n70894 ;
  assign n70930 = ~n70928 & ~n70929 ;
  assign n70931 = ~n70902 & ~n70930 ;
  assign n70923 = ~n70872 & ~n70893 ;
  assign n70932 = n70872 & n70893 ;
  assign n70933 = ~n70923 & ~n70932 ;
  assign n70934 = ~n70872 & ~n70887 ;
  assign n70935 = n70878 & n70902 ;
  assign n70936 = ~n70934 & n70935 ;
  assign n70937 = n70933 & n70936 ;
  assign n70921 = n70872 & ~n70893 ;
  assign n70922 = n70896 & n70921 ;
  assign n70924 = ~n70878 & ~n70887 ;
  assign n70925 = n70923 & n70924 ;
  assign n70938 = ~n70922 & ~n70925 ;
  assign n70939 = ~n70937 & n70938 ;
  assign n70940 = ~n70931 & n70939 ;
  assign n70941 = n70866 & ~n70940 ;
  assign n70944 = n70924 & n70932 ;
  assign n70945 = ~n70922 & ~n70944 ;
  assign n70946 = ~n70893 & n70910 ;
  assign n70947 = n70945 & ~n70946 ;
  assign n70948 = n70902 & ~n70947 ;
  assign n70942 = n70893 & ~n70902 ;
  assign n70943 = ~n70881 & n70942 ;
  assign n70949 = n70905 & n70934 ;
  assign n70950 = ~n70943 & ~n70949 ;
  assign n70951 = ~n70948 & n70950 ;
  assign n70952 = ~n70941 & n70951 ;
  assign n70953 = ~n70920 & n70952 ;
  assign n70954 = ~\u0_L0_reg[22]/NET0131  & ~n70953 ;
  assign n70955 = \u0_L0_reg[22]/NET0131  & n70953 ;
  assign n70956 = ~n70954 & ~n70955 ;
  assign n70957 = ~n70676 & n70696 ;
  assign n70958 = ~n70709 & ~n70957 ;
  assign n70959 = n70683 & n70734 ;
  assign n70960 = ~n70958 & n70959 ;
  assign n70966 = n70717 & ~n70734 ;
  assign n70961 = ~n70670 & ~n70699 ;
  assign n70962 = ~n70726 & ~n70961 ;
  assign n70963 = n70683 & ~n70962 ;
  assign n70964 = n70690 & ~n70722 ;
  assign n70965 = n70958 & n70964 ;
  assign n70967 = n70707 & ~n70965 ;
  assign n70968 = ~n70963 & n70967 ;
  assign n70969 = ~n70966 & n70968 ;
  assign n70972 = ~n70711 & ~n70722 ;
  assign n70973 = ~n70690 & ~n70972 ;
  assign n70974 = ~n70723 & ~n70973 ;
  assign n70975 = ~n70683 & ~n70974 ;
  assign n70970 = ~n70718 & ~n70747 ;
  assign n70971 = n70700 & n70970 ;
  assign n70976 = ~n70707 & ~n70710 ;
  assign n70977 = ~n70751 & n70976 ;
  assign n70978 = ~n70971 & n70977 ;
  assign n70979 = ~n70975 & n70978 ;
  assign n70980 = ~n70969 & ~n70979 ;
  assign n70981 = ~n70960 & ~n70980 ;
  assign n70982 = ~\u0_L0_reg[17]/NET0131  & ~n70981 ;
  assign n70983 = \u0_L0_reg[17]/NET0131  & n70981 ;
  assign n70984 = ~n70982 & ~n70983 ;
  assign n70989 = ~n70780 & n70827 ;
  assign n70990 = ~n70808 & ~n70830 ;
  assign n70991 = ~n70989 & n70990 ;
  assign n70992 = n70790 & ~n70991 ;
  assign n70985 = n70807 & n70827 ;
  assign n70986 = n70767 & n70810 ;
  assign n70987 = ~n70985 & ~n70986 ;
  assign n70988 = ~n70790 & ~n70987 ;
  assign n70993 = ~n70838 & ~n70842 ;
  assign n70994 = ~n70988 & n70993 ;
  assign n70995 = ~n70992 & n70994 ;
  assign n70996 = ~n70822 & ~n70995 ;
  assign n71008 = ~n70799 & n70803 ;
  assign n71007 = ~n70780 & n70986 ;
  assign n71005 = ~n70780 & n70790 ;
  assign n71006 = n70806 & n71005 ;
  assign n71009 = n70780 & n70844 ;
  assign n71010 = ~n71006 & ~n71009 ;
  assign n71011 = ~n71007 & n71010 ;
  assign n71012 = ~n71008 & n71011 ;
  assign n71013 = n70822 & ~n71012 ;
  assign n70999 = ~n70824 & ~n70845 ;
  assign n71000 = n70790 & ~n70830 ;
  assign n71001 = n70999 & n71000 ;
  assign n70997 = ~n70836 & ~n70837 ;
  assign n70998 = ~n70790 & n70997 ;
  assign n71002 = n70780 & ~n70998 ;
  assign n71003 = ~n71001 & n71002 ;
  assign n71004 = n70803 & n70810 ;
  assign n71014 = ~n71003 & ~n71004 ;
  assign n71015 = ~n71013 & n71014 ;
  assign n71016 = ~n70996 & n71015 ;
  assign n71017 = ~\u0_L0_reg[4]/NET0131  & ~n71016 ;
  assign n71018 = \u0_L0_reg[4]/NET0131  & n71016 ;
  assign n71019 = ~n71017 & ~n71018 ;
  assign n71033 = decrypt_pad & ~\u0_uk_K_r0_reg[18]/NET0131  ;
  assign n71034 = ~decrypt_pad & ~\u0_uk_K_r0_reg[39]/NET0131  ;
  assign n71035 = ~n71033 & ~n71034 ;
  assign n71036 = \u0_R0_reg[15]/NET0131  & ~n71035 ;
  assign n71037 = ~\u0_R0_reg[15]/NET0131  & n71035 ;
  assign n71038 = ~n71036 & ~n71037 ;
  assign n71020 = decrypt_pad & ~\u0_uk_K_r0_reg[6]/NET0131  ;
  assign n71021 = ~decrypt_pad & ~\u0_uk_K_r0_reg[27]/NET0131  ;
  assign n71022 = ~n71020 & ~n71021 ;
  assign n71023 = \u0_R0_reg[17]/NET0131  & ~n71022 ;
  assign n71024 = ~\u0_R0_reg[17]/NET0131  & n71022 ;
  assign n71025 = ~n71023 & ~n71024 ;
  assign n71047 = decrypt_pad & ~\u0_uk_K_r0_reg[10]/NET0131  ;
  assign n71048 = ~decrypt_pad & ~\u0_uk_K_r0_reg[6]/NET0131  ;
  assign n71049 = ~n71047 & ~n71048 ;
  assign n71050 = \u0_R0_reg[14]/NET0131  & ~n71049 ;
  assign n71051 = ~\u0_R0_reg[14]/NET0131  & n71049 ;
  assign n71052 = ~n71050 & ~n71051 ;
  assign n71026 = decrypt_pad & ~\u0_uk_K_r0_reg[47]/NET0131  ;
  assign n71027 = ~decrypt_pad & ~\u0_uk_K_r0_reg[11]/NET0131  ;
  assign n71028 = ~n71026 & ~n71027 ;
  assign n71029 = \u0_R0_reg[12]/NET0131  & ~n71028 ;
  assign n71030 = ~\u0_R0_reg[12]/NET0131  & n71028 ;
  assign n71031 = ~n71029 & ~n71030 ;
  assign n71040 = decrypt_pad & ~\u0_uk_K_r0_reg[41]/NET0131  ;
  assign n71041 = ~decrypt_pad & ~\u0_uk_K_r0_reg[5]/NET0131  ;
  assign n71042 = ~n71040 & ~n71041 ;
  assign n71043 = \u0_R0_reg[13]/NET0131  & ~n71042 ;
  assign n71044 = ~\u0_R0_reg[13]/NET0131  & n71042 ;
  assign n71045 = ~n71043 & ~n71044 ;
  assign n71068 = ~n71031 & ~n71045 ;
  assign n71069 = n71052 & n71068 ;
  assign n71070 = ~n71025 & n71069 ;
  assign n71071 = ~n71031 & n71045 ;
  assign n71072 = n71031 & ~n71045 ;
  assign n71073 = ~n71071 & ~n71072 ;
  assign n71074 = ~n71052 & ~n71073 ;
  assign n71075 = ~n71070 & ~n71074 ;
  assign n71076 = ~n71038 & ~n71075 ;
  assign n71032 = n71025 & ~n71031 ;
  assign n71053 = n71032 & n71045 ;
  assign n71054 = ~n71052 & n71053 ;
  assign n71055 = ~n71025 & n71031 ;
  assign n71056 = n71038 & n71045 ;
  assign n71057 = n71055 & n71056 ;
  assign n71058 = ~n71054 & ~n71057 ;
  assign n71059 = n71025 & n71031 ;
  assign n71060 = n71052 & n71059 ;
  assign n71061 = n71045 & n71060 ;
  assign n71039 = n71032 & n71038 ;
  assign n71046 = n71039 & ~n71045 ;
  assign n71062 = decrypt_pad & ~\u0_uk_K_r0_reg[26]/NET0131  ;
  assign n71063 = ~decrypt_pad & ~\u0_uk_K_r0_reg[47]/NET0131  ;
  assign n71064 = ~n71062 & ~n71063 ;
  assign n71065 = \u0_R0_reg[16]/NET0131  & ~n71064 ;
  assign n71066 = ~\u0_R0_reg[16]/NET0131  & n71064 ;
  assign n71067 = ~n71065 & ~n71066 ;
  assign n71077 = ~n71046 & n71067 ;
  assign n71078 = ~n71061 & n71077 ;
  assign n71079 = n71058 & n71078 ;
  assign n71080 = ~n71076 & n71079 ;
  assign n71081 = ~n71025 & ~n71031 ;
  assign n71095 = ~n71052 & n71081 ;
  assign n71096 = ~n71045 & n71095 ;
  assign n71091 = ~n71052 & n71072 ;
  assign n71092 = n71025 & n71091 ;
  assign n71093 = n71045 & n71081 ;
  assign n71094 = n71052 & n71093 ;
  assign n71100 = ~n71092 & ~n71094 ;
  assign n71101 = ~n71096 & n71100 ;
  assign n71087 = n71052 & n71055 ;
  assign n71088 = n71025 & ~n71045 ;
  assign n71089 = ~n71087 & ~n71088 ;
  assign n71090 = ~n71038 & ~n71089 ;
  assign n71082 = n71038 & ~n71045 ;
  assign n71083 = n71081 & n71082 ;
  assign n71097 = ~n71067 & ~n71083 ;
  assign n71084 = n71056 & n71059 ;
  assign n71085 = n71038 & n71052 ;
  assign n71086 = n71071 & n71085 ;
  assign n71098 = ~n71084 & ~n71086 ;
  assign n71099 = n71097 & n71098 ;
  assign n71102 = ~n71090 & n71099 ;
  assign n71103 = n71101 & n71102 ;
  assign n71104 = ~n71080 & ~n71103 ;
  assign n71108 = ~n71087 & ~n71095 ;
  assign n71109 = n71082 & ~n71108 ;
  assign n71105 = n71025 & ~n71052 ;
  assign n71106 = ~n71038 & n71105 ;
  assign n71107 = n71071 & n71106 ;
  assign n71110 = ~n71052 & n71057 ;
  assign n71111 = ~n71107 & ~n71110 ;
  assign n71112 = ~n71109 & n71111 ;
  assign n71113 = ~n71104 & n71112 ;
  assign n71114 = ~\u0_L0_reg[20]/NET0131  & ~n71113 ;
  assign n71115 = \u0_L0_reg[20]/NET0131  & n71113 ;
  assign n71116 = ~n71114 & ~n71115 ;
  assign n71133 = ~n70781 & ~n70826 ;
  assign n71134 = ~n70797 & ~n71133 ;
  assign n71135 = n70997 & ~n71134 ;
  assign n71136 = n70790 & ~n71135 ;
  assign n71121 = n70780 & n70830 ;
  assign n71137 = ~n70780 & ~n70847 ;
  assign n71138 = ~n71121 & ~n71137 ;
  assign n71139 = ~n70790 & ~n71138 ;
  assign n71140 = ~n70985 & ~n71139 ;
  assign n71141 = ~n71136 & n71140 ;
  assign n71142 = ~n70822 & ~n71141 ;
  assign n71122 = n70780 & ~n70797 ;
  assign n71123 = n70774 & ~n71122 ;
  assign n71124 = ~n71121 & ~n71123 ;
  assign n71125 = n70790 & ~n71124 ;
  assign n71117 = n70780 & ~n70804 ;
  assign n71118 = ~n70827 & n71117 ;
  assign n71119 = ~n70824 & ~n71118 ;
  assign n71120 = ~n70790 & ~n71119 ;
  assign n71126 = n70780 & n70824 ;
  assign n71127 = n70809 & ~n70828 ;
  assign n71128 = ~n71126 & n71127 ;
  assign n71129 = ~n71120 & n71128 ;
  assign n71130 = ~n71125 & n71129 ;
  assign n71131 = n70822 & ~n71130 ;
  assign n71132 = n70844 & n71005 ;
  assign n71143 = ~n70838 & ~n71132 ;
  assign n71144 = ~n71131 & n71143 ;
  assign n71145 = ~n71142 & n71144 ;
  assign n71146 = \u0_L0_reg[29]/NET0131  & ~n71145 ;
  assign n71147 = ~\u0_L0_reg[29]/NET0131  & n71145 ;
  assign n71148 = ~n71146 & ~n71147 ;
  assign n71149 = decrypt_pad & ~\u0_uk_K_r0_reg[34]/NET0131  ;
  assign n71150 = ~decrypt_pad & ~\u0_uk_K_r0_reg[55]/NET0131  ;
  assign n71151 = ~n71149 & ~n71150 ;
  assign n71152 = \u0_R0_reg[7]/NET0131  & ~n71151 ;
  assign n71153 = ~\u0_R0_reg[7]/NET0131  & n71151 ;
  assign n71154 = ~n71152 & ~n71153 ;
  assign n71161 = decrypt_pad & ~\u0_uk_K_r0_reg[17]/NET0131  ;
  assign n71162 = ~decrypt_pad & ~\u0_uk_K_r0_reg[13]/NET0131  ;
  assign n71163 = ~n71161 & ~n71162 ;
  assign n71164 = \u0_R0_reg[5]/NET0131  & ~n71163 ;
  assign n71165 = ~\u0_R0_reg[5]/NET0131  & n71163 ;
  assign n71166 = ~n71164 & ~n71165 ;
  assign n71167 = decrypt_pad & ~\u0_uk_K_r0_reg[40]/NET0131  ;
  assign n71168 = ~decrypt_pad & ~\u0_uk_K_r0_reg[4]/NET0131  ;
  assign n71169 = ~n71167 & ~n71168 ;
  assign n71170 = \u0_R0_reg[6]/NET0131  & ~n71169 ;
  assign n71171 = ~\u0_R0_reg[6]/NET0131  & n71169 ;
  assign n71172 = ~n71170 & ~n71171 ;
  assign n71173 = ~n71166 & n71172 ;
  assign n71155 = decrypt_pad & ~\u0_uk_K_r0_reg[5]/NET0131  ;
  assign n71156 = ~decrypt_pad & ~\u0_uk_K_r0_reg[26]/NET0131  ;
  assign n71157 = ~n71155 & ~n71156 ;
  assign n71158 = \u0_R0_reg[9]/NET0131  & ~n71157 ;
  assign n71159 = ~\u0_R0_reg[9]/NET0131  & n71157 ;
  assign n71160 = ~n71158 & ~n71159 ;
  assign n71174 = decrypt_pad & ~\u0_uk_K_r0_reg[13]/NET0131  ;
  assign n71175 = ~decrypt_pad & ~\u0_uk_K_r0_reg[34]/NET0131  ;
  assign n71176 = ~n71174 & ~n71175 ;
  assign n71177 = \u0_R0_reg[4]/NET0131  & ~n71176 ;
  assign n71178 = ~\u0_R0_reg[4]/NET0131  & n71176 ;
  assign n71179 = ~n71177 & ~n71178 ;
  assign n71199 = n71160 & n71179 ;
  assign n71200 = n71173 & n71199 ;
  assign n71201 = n71154 & n71200 ;
  assign n71186 = n71172 & ~n71179 ;
  assign n71187 = n71160 & n71166 ;
  assign n71188 = n71186 & n71187 ;
  assign n71189 = n71160 & ~n71166 ;
  assign n71190 = ~n71154 & ~n71172 ;
  assign n71191 = n71189 & n71190 ;
  assign n71192 = ~n71188 & ~n71191 ;
  assign n71193 = decrypt_pad & ~\u0_uk_K_r0_reg[25]/P0001  ;
  assign n71194 = ~decrypt_pad & ~\u0_uk_K_r0_reg[46]/NET0131  ;
  assign n71195 = ~n71193 & ~n71194 ;
  assign n71196 = \u0_R0_reg[8]/NET0131  & ~n71195 ;
  assign n71197 = ~\u0_R0_reg[8]/NET0131  & n71195 ;
  assign n71198 = ~n71196 & ~n71197 ;
  assign n71211 = n71192 & ~n71198 ;
  assign n71212 = ~n71201 & n71211 ;
  assign n71202 = n71172 & n71179 ;
  assign n71203 = ~n71189 & n71202 ;
  assign n71204 = n71160 & ~n71179 ;
  assign n71205 = ~n71166 & n71204 ;
  assign n71206 = ~n71203 & ~n71205 ;
  assign n71207 = ~n71154 & ~n71206 ;
  assign n71208 = ~n71160 & n71166 ;
  assign n71209 = ~n71205 & ~n71208 ;
  assign n71210 = ~n71172 & ~n71209 ;
  assign n71213 = ~n71207 & ~n71210 ;
  assign n71214 = n71212 & n71213 ;
  assign n71216 = ~n71160 & ~n71172 ;
  assign n71217 = ~n71166 & n71216 ;
  assign n71218 = n71179 & n71217 ;
  assign n71182 = ~n71172 & n71179 ;
  assign n71183 = n71166 & n71182 ;
  assign n71215 = n71160 & n71183 ;
  assign n71219 = n71154 & n71166 ;
  assign n71220 = ~n71186 & n71219 ;
  assign n71221 = n71198 & ~n71220 ;
  assign n71222 = ~n71215 & n71221 ;
  assign n71223 = ~n71218 & n71222 ;
  assign n71224 = ~n71214 & ~n71223 ;
  assign n71180 = n71173 & ~n71179 ;
  assign n71181 = ~n71160 & n71180 ;
  assign n71184 = ~n71181 & ~n71183 ;
  assign n71185 = n71154 & ~n71184 ;
  assign n71225 = ~n71173 & n71204 ;
  assign n71228 = ~n71173 & n71179 ;
  assign n71226 = ~n71160 & ~n71179 ;
  assign n71227 = ~n71199 & ~n71226 ;
  assign n71229 = n71198 & ~n71227 ;
  assign n71230 = ~n71228 & n71229 ;
  assign n71231 = ~n71225 & ~n71230 ;
  assign n71232 = n71166 & ~n71172 ;
  assign n71233 = ~n71154 & ~n71232 ;
  assign n71234 = ~n71231 & n71233 ;
  assign n71235 = ~n71185 & ~n71234 ;
  assign n71236 = ~n71224 & n71235 ;
  assign n71237 = \u0_L0_reg[2]/NET0131  & n71236 ;
  assign n71238 = ~\u0_L0_reg[2]/NET0131  & ~n71236 ;
  assign n71239 = ~n71237 & ~n71238 ;
  assign n71286 = decrypt_pad & ~\u0_uk_K_r0_reg[52]/NET0131  ;
  assign n71287 = ~decrypt_pad & ~\u0_uk_K_r0_reg[14]/NET0131  ;
  assign n71288 = ~n71286 & ~n71287 ;
  assign n71289 = \u0_R0_reg[32]/NET0131  & ~n71288 ;
  assign n71290 = ~\u0_R0_reg[32]/NET0131  & n71288 ;
  assign n71291 = ~n71289 & ~n71290 ;
  assign n71260 = decrypt_pad & ~\u0_uk_K_r0_reg[42]/NET0131  ;
  assign n71261 = ~decrypt_pad & ~\u0_uk_K_r0_reg[8]/NET0131  ;
  assign n71262 = ~n71260 & ~n71261 ;
  assign n71263 = \u0_R0_reg[31]/NET0131  & ~n71262 ;
  assign n71264 = ~\u0_R0_reg[31]/NET0131  & n71262 ;
  assign n71265 = ~n71263 & ~n71264 ;
  assign n71240 = decrypt_pad & ~\u0_uk_K_r0_reg[30]/NET0131  ;
  assign n71241 = ~decrypt_pad & ~\u0_uk_K_r0_reg[51]/NET0131  ;
  assign n71242 = ~n71240 & ~n71241 ;
  assign n71243 = \u0_R0_reg[30]/NET0131  & ~n71242 ;
  assign n71244 = ~\u0_R0_reg[30]/NET0131  & n71242 ;
  assign n71245 = ~n71243 & ~n71244 ;
  assign n71253 = decrypt_pad & ~\u0_uk_K_r0_reg[2]/NET0131  ;
  assign n71254 = ~decrypt_pad & ~\u0_uk_K_r0_reg[23]/NET0131  ;
  assign n71255 = ~n71253 & ~n71254 ;
  assign n71256 = \u0_R0_reg[28]/NET0131  & ~n71255 ;
  assign n71257 = ~\u0_R0_reg[28]/NET0131  & n71255 ;
  assign n71258 = ~n71256 & ~n71257 ;
  assign n71267 = ~n71245 & n71258 ;
  assign n71268 = decrypt_pad & ~\u0_uk_K_r0_reg[14]/NET0131  ;
  assign n71269 = ~decrypt_pad & ~\u0_uk_K_r0_reg[35]/NET0131  ;
  assign n71270 = ~n71268 & ~n71269 ;
  assign n71271 = \u0_R0_reg[1]/NET0131  & ~n71270 ;
  assign n71272 = ~\u0_R0_reg[1]/NET0131  & n71270 ;
  assign n71273 = ~n71271 & ~n71272 ;
  assign n71310 = ~n71245 & ~n71273 ;
  assign n71277 = n71258 & ~n71273 ;
  assign n71246 = decrypt_pad & ~\u0_uk_K_r0_reg[29]/NET0131  ;
  assign n71247 = ~decrypt_pad & ~\u0_uk_K_r0_reg[50]/NET0131  ;
  assign n71248 = ~n71246 & ~n71247 ;
  assign n71249 = \u0_R0_reg[29]/NET0131  & ~n71248 ;
  assign n71250 = ~\u0_R0_reg[29]/NET0131  & n71248 ;
  assign n71251 = ~n71249 & ~n71250 ;
  assign n71293 = ~n71251 & n71273 ;
  assign n71311 = ~n71277 & ~n71293 ;
  assign n71312 = ~n71310 & n71311 ;
  assign n71313 = ~n71267 & ~n71312 ;
  assign n71314 = ~n71265 & ~n71313 ;
  assign n71298 = ~n71258 & n71273 ;
  assign n71299 = ~n71251 & n71298 ;
  assign n71304 = n71245 & ~n71251 ;
  assign n71317 = n71277 & n71304 ;
  assign n71318 = ~n71299 & ~n71317 ;
  assign n71319 = n71265 & ~n71318 ;
  assign n71276 = ~n71245 & n71251 ;
  assign n71278 = n71276 & n71277 ;
  assign n71282 = n71245 & n71251 ;
  assign n71315 = n71258 & n71273 ;
  assign n71316 = n71282 & n71315 ;
  assign n71320 = ~n71278 & ~n71316 ;
  assign n71321 = ~n71319 & n71320 ;
  assign n71322 = ~n71314 & n71321 ;
  assign n71323 = ~n71291 & ~n71322 ;
  assign n71252 = ~n71245 & ~n71251 ;
  assign n71259 = n71252 & ~n71258 ;
  assign n71266 = ~n71259 & ~n71265 ;
  assign n71274 = n71251 & ~n71273 ;
  assign n71275 = ~n71267 & ~n71274 ;
  assign n71279 = ~n71275 & ~n71278 ;
  assign n71280 = n71265 & ~n71279 ;
  assign n71281 = ~n71266 & ~n71280 ;
  assign n71283 = ~n71258 & n71282 ;
  assign n71284 = n71273 & n71283 ;
  assign n71285 = ~n71281 & ~n71284 ;
  assign n71292 = ~n71285 & n71291 ;
  assign n71300 = n71245 & n71299 ;
  assign n71294 = n71267 & n71293 ;
  assign n71295 = ~n71258 & ~n71273 ;
  assign n71296 = ~n71252 & ~n71282 ;
  assign n71297 = n71295 & ~n71296 ;
  assign n71301 = ~n71294 & ~n71297 ;
  assign n71302 = ~n71300 & n71301 ;
  assign n71303 = n71265 & ~n71302 ;
  assign n71305 = n71291 & n71304 ;
  assign n71306 = ~n71245 & n71274 ;
  assign n71307 = ~n71305 & ~n71306 ;
  assign n71308 = n71258 & ~n71265 ;
  assign n71309 = ~n71307 & n71308 ;
  assign n71324 = ~n71303 & ~n71309 ;
  assign n71325 = ~n71292 & n71324 ;
  assign n71326 = ~n71323 & n71325 ;
  assign n71327 = \u0_L0_reg[5]/NET0131  & ~n71326 ;
  assign n71328 = ~\u0_L0_reg[5]/NET0131  & n71326 ;
  assign n71329 = ~n71327 & ~n71328 ;
  assign n71330 = n71251 & ~n71295 ;
  assign n71331 = ~n71252 & ~n71330 ;
  assign n71332 = n71267 & ~n71293 ;
  assign n71333 = ~n71331 & ~n71332 ;
  assign n71334 = n71265 & ~n71333 ;
  assign n71335 = n71296 & n71315 ;
  assign n71336 = n71267 & ~n71273 ;
  assign n71337 = ~n71265 & ~n71336 ;
  assign n71338 = ~n71335 & n71337 ;
  assign n71339 = ~n71334 & ~n71338 ;
  assign n71340 = ~n71251 & n71295 ;
  assign n71341 = n71258 & n71274 ;
  assign n71342 = ~n71340 & ~n71341 ;
  assign n71343 = n71245 & ~n71342 ;
  assign n71344 = n71259 & n71273 ;
  assign n71345 = n71291 & ~n71344 ;
  assign n71346 = ~n71343 & n71345 ;
  assign n71347 = ~n71339 & n71346 ;
  assign n71355 = n71258 & n71304 ;
  assign n71356 = ~n71259 & ~n71341 ;
  assign n71357 = ~n71355 & n71356 ;
  assign n71358 = n71265 & ~n71357 ;
  assign n71352 = ~n71265 & n71315 ;
  assign n71353 = ~n71340 & ~n71352 ;
  assign n71354 = ~n71245 & ~n71353 ;
  assign n71360 = ~n71283 & ~n71291 ;
  assign n71348 = n71245 & ~n71265 ;
  assign n71349 = n71298 & n71348 ;
  assign n71361 = ~n71317 & ~n71349 ;
  assign n71350 = ~n71258 & ~n71265 ;
  assign n71351 = n71274 & n71350 ;
  assign n71359 = n71276 & n71315 ;
  assign n71362 = ~n71351 & ~n71359 ;
  assign n71363 = n71361 & n71362 ;
  assign n71364 = n71360 & n71363 ;
  assign n71365 = ~n71354 & n71364 ;
  assign n71366 = ~n71358 & n71365 ;
  assign n71367 = ~n71347 & ~n71366 ;
  assign n71368 = ~\u0_L0_reg[21]/NET0131  & n71367 ;
  assign n71369 = \u0_L0_reg[21]/NET0131  & ~n71367 ;
  assign n71370 = ~n71368 & ~n71369 ;
  assign n71375 = n70880 & n70894 ;
  assign n71376 = n70866 & ~n70944 ;
  assign n71377 = ~n71375 & n71376 ;
  assign n71378 = ~n70928 & n71377 ;
  assign n71371 = ~n70903 & ~n70910 ;
  assign n71372 = n70921 & ~n71371 ;
  assign n71373 = ~n70914 & ~n70925 ;
  assign n71374 = n70902 & ~n71373 ;
  assign n71379 = ~n71372 & ~n71374 ;
  assign n71380 = n71378 & n71379 ;
  assign n71387 = ~n70878 & ~n70894 ;
  assign n71386 = ~n70926 & n70935 ;
  assign n71388 = n70872 & ~n71386 ;
  assign n71389 = ~n71387 & n71388 ;
  assign n71384 = n70896 & n70905 ;
  assign n71381 = n70910 & n70923 ;
  assign n71390 = ~n70866 & ~n71381 ;
  assign n71391 = ~n71384 & n71390 ;
  assign n71382 = ~n70894 & ~n70904 ;
  assign n71383 = ~n70902 & ~n71382 ;
  assign n71385 = n70924 & n70933 ;
  assign n71392 = ~n71383 & ~n71385 ;
  assign n71393 = n71391 & n71392 ;
  assign n71394 = ~n71389 & n71393 ;
  assign n71395 = ~n71380 & ~n71394 ;
  assign n71396 = \u0_L0_reg[12]/NET0131  & n71395 ;
  assign n71397 = ~\u0_L0_reg[12]/NET0131  & ~n71395 ;
  assign n71398 = ~n71396 & ~n71397 ;
  assign n71405 = ~n70708 & ~n70749 ;
  assign n71406 = ~n70683 & ~n71405 ;
  assign n71407 = ~n70707 & ~n70721 ;
  assign n71399 = ~n70696 & n70959 ;
  assign n71404 = n70958 & n70970 ;
  assign n71408 = ~n71399 & ~n71404 ;
  assign n71409 = n71407 & n71408 ;
  assign n71410 = ~n71406 & n71409 ;
  assign n71411 = ~n70711 & n70964 ;
  assign n71412 = ~n70973 & ~n71411 ;
  assign n71413 = n70670 & ~n70709 ;
  assign n71414 = ~n70683 & ~n71413 ;
  assign n71415 = n71412 & n71414 ;
  assign n71416 = n70683 & ~n70715 ;
  assign n71417 = n71411 & n71416 ;
  assign n71418 = n70707 & ~n70726 ;
  assign n71419 = ~n70698 & n71418 ;
  assign n71420 = ~n71417 & n71419 ;
  assign n71421 = ~n71415 & n71420 ;
  assign n71422 = ~n71410 & ~n71421 ;
  assign n71400 = ~n70683 & ~n70711 ;
  assign n71401 = ~n70719 & n71400 ;
  assign n71402 = ~n71399 & ~n71401 ;
  assign n71403 = ~n70676 & ~n71402 ;
  assign n71423 = n70735 & n70749 ;
  assign n71424 = ~n70701 & ~n71423 ;
  assign n71425 = ~n71403 & n71424 ;
  assign n71426 = ~n71422 & n71425 ;
  assign n71427 = \u0_L0_reg[23]/NET0131  & ~n71426 ;
  assign n71428 = ~\u0_L0_reg[23]/NET0131  & n71426 ;
  assign n71429 = ~n71427 & ~n71428 ;
  assign n71436 = n71045 & ~n71095 ;
  assign n71437 = n71038 & ~n71108 ;
  assign n71438 = ~n71436 & n71437 ;
  assign n71430 = ~n71052 & n71055 ;
  assign n71433 = ~n71059 & ~n71430 ;
  assign n71434 = ~n71038 & ~n71045 ;
  assign n71435 = ~n71433 & n71434 ;
  assign n71431 = ~n71060 & ~n71430 ;
  assign n71432 = n71045 & ~n71431 ;
  assign n71439 = ~n71054 & ~n71432 ;
  assign n71440 = ~n71435 & n71439 ;
  assign n71441 = ~n71438 & n71440 ;
  assign n71442 = ~n71067 & ~n71441 ;
  assign n71453 = n71045 & ~n71052 ;
  assign n71454 = ~n71055 & n71453 ;
  assign n71455 = ~n71053 & ~n71454 ;
  assign n71456 = ~n71038 & ~n71455 ;
  assign n71447 = n71045 & n71087 ;
  assign n71457 = ~n71069 & ~n71447 ;
  assign n71458 = ~n71456 & n71457 ;
  assign n71459 = n71067 & ~n71458 ;
  assign n71443 = n71025 & n71069 ;
  assign n71444 = ~n71061 & ~n71443 ;
  assign n71445 = ~n71094 & n71444 ;
  assign n71446 = n71038 & ~n71445 ;
  assign n71448 = ~n71070 & ~n71447 ;
  assign n71449 = ~n71038 & ~n71448 ;
  assign n71450 = ~n71088 & ~n71091 ;
  assign n71451 = n71038 & n71067 ;
  assign n71452 = ~n71450 & n71451 ;
  assign n71460 = ~n71449 & ~n71452 ;
  assign n71461 = ~n71446 & n71460 ;
  assign n71462 = ~n71459 & n71461 ;
  assign n71463 = ~n71442 & n71462 ;
  assign n71464 = ~\u0_L0_reg[1]/NET0131  & ~n71463 ;
  assign n71465 = \u0_L0_reg[1]/NET0131  & n71463 ;
  assign n71466 = ~n71464 & ~n71465 ;
  assign n71467 = ~n71187 & ~n71216 ;
  assign n71468 = ~n71179 & ~n71467 ;
  assign n71469 = n71154 & ~n71468 ;
  assign n71471 = ~n71189 & n71228 ;
  assign n71470 = ~n71154 & ~n71180 ;
  assign n71472 = ~n71205 & n71470 ;
  assign n71473 = ~n71471 & n71472 ;
  assign n71474 = ~n71469 & ~n71473 ;
  assign n71475 = n71179 & n71208 ;
  assign n71476 = ~n71166 & ~n71227 ;
  assign n71477 = ~n71475 & ~n71476 ;
  assign n71478 = n71172 & ~n71477 ;
  assign n71479 = ~n71198 & ~n71478 ;
  assign n71480 = ~n71474 & n71479 ;
  assign n71483 = n71179 & ~n71208 ;
  assign n71484 = ~n71189 & n71483 ;
  assign n71481 = ~n71179 & n71208 ;
  assign n71482 = n71172 & n71481 ;
  assign n71485 = n71154 & ~n71482 ;
  assign n71486 = ~n71484 & n71485 ;
  assign n71487 = n71172 & n71475 ;
  assign n71488 = ~n71468 & n71470 ;
  assign n71489 = ~n71487 & n71488 ;
  assign n71490 = ~n71486 & ~n71489 ;
  assign n71491 = ~n71154 & ~n71189 ;
  assign n71492 = n71182 & ~n71491 ;
  assign n71493 = n71173 & n71204 ;
  assign n71494 = n71198 & ~n71493 ;
  assign n71495 = ~n71492 & n71494 ;
  assign n71496 = ~n71490 & n71495 ;
  assign n71497 = ~n71480 & ~n71496 ;
  assign n71498 = \u0_L0_reg[28]/NET0131  & n71497 ;
  assign n71499 = ~\u0_L0_reg[28]/NET0131  & ~n71497 ;
  assign n71500 = ~n71498 & ~n71499 ;
  assign n71502 = ~n71258 & ~n71310 ;
  assign n71503 = n71251 & ~n71502 ;
  assign n71504 = ~n71299 & ~n71503 ;
  assign n71505 = n71265 & ~n71504 ;
  assign n71501 = n71252 & n71277 ;
  assign n71506 = ~n71291 & ~n71501 ;
  assign n71507 = ~n71505 & n71506 ;
  assign n71509 = ~n71251 & n71348 ;
  assign n71510 = ~n71355 & ~n71509 ;
  assign n71511 = n71273 & ~n71510 ;
  assign n71513 = ~n71273 & n71283 ;
  assign n71512 = n71265 & n71340 ;
  assign n71508 = n71258 & n71276 ;
  assign n71514 = n71291 & ~n71508 ;
  assign n71515 = ~n71512 & n71514 ;
  assign n71516 = ~n71513 & n71515 ;
  assign n71517 = ~n71511 & n71516 ;
  assign n71518 = ~n71507 & ~n71517 ;
  assign n71520 = ~n71245 & n71291 ;
  assign n71521 = ~n71251 & n71258 ;
  assign n71522 = ~n71520 & n71521 ;
  assign n71519 = n71276 & n71298 ;
  assign n71523 = ~n71265 & ~n71519 ;
  assign n71524 = ~n71522 & n71523 ;
  assign n71525 = ~n71297 & n71524 ;
  assign n71526 = n71265 & ~n71284 ;
  assign n71527 = ~n71344 & n71526 ;
  assign n71528 = ~n71525 & ~n71527 ;
  assign n71529 = ~n71518 & ~n71528 ;
  assign n71530 = \u0_L0_reg[15]/P0001  & n71529 ;
  assign n71531 = ~\u0_L0_reg[15]/P0001  & ~n71529 ;
  assign n71532 = ~n71530 & ~n71531 ;
  assign n71533 = decrypt_pad & ~\u0_uk_K_r0_reg[3]/NET0131  ;
  assign n71534 = ~decrypt_pad & ~\u0_uk_K_r0_reg[24]/P0001  ;
  assign n71535 = ~n71533 & ~n71534 ;
  assign n71536 = \u0_R0_reg[12]/NET0131  & ~n71535 ;
  assign n71537 = ~\u0_R0_reg[12]/NET0131  & n71535 ;
  assign n71538 = ~n71536 & ~n71537 ;
  assign n71539 = decrypt_pad & ~\u0_uk_K_r0_reg[11]/NET0131  ;
  assign n71540 = ~decrypt_pad & ~\u0_uk_K_r0_reg[32]/NET0131  ;
  assign n71541 = ~n71539 & ~n71540 ;
  assign n71542 = \u0_R0_reg[9]/NET0131  & ~n71541 ;
  assign n71543 = ~\u0_R0_reg[9]/NET0131  & n71541 ;
  assign n71544 = ~n71542 & ~n71543 ;
  assign n71553 = decrypt_pad & ~\u0_uk_K_r0_reg[39]/NET0131  ;
  assign n71554 = ~decrypt_pad & ~\u0_uk_K_r0_reg[3]/NET0131  ;
  assign n71555 = ~n71553 & ~n71554 ;
  assign n71556 = \u0_R0_reg[8]/NET0131  & ~n71555 ;
  assign n71557 = ~\u0_R0_reg[8]/NET0131  & n71555 ;
  assign n71558 = ~n71556 & ~n71557 ;
  assign n71545 = decrypt_pad & ~\u0_uk_K_r0_reg[19]/NET0131  ;
  assign n71546 = ~decrypt_pad & ~\u0_uk_K_r0_reg[40]/NET0131  ;
  assign n71547 = ~n71545 & ~n71546 ;
  assign n71548 = \u0_R0_reg[10]/NET0131  & ~n71547 ;
  assign n71549 = ~\u0_R0_reg[10]/NET0131  & n71547 ;
  assign n71550 = ~n71548 & ~n71549 ;
  assign n71559 = decrypt_pad & ~\u0_uk_K_r0_reg[48]/NET0131  ;
  assign n71560 = ~decrypt_pad & ~\u0_uk_K_r0_reg[12]/NET0131  ;
  assign n71561 = ~n71559 & ~n71560 ;
  assign n71562 = \u0_R0_reg[13]/NET0131  & ~n71561 ;
  assign n71563 = ~\u0_R0_reg[13]/NET0131  & n71561 ;
  assign n71564 = ~n71562 & ~n71563 ;
  assign n71582 = ~n71550 & ~n71564 ;
  assign n71583 = n71558 & n71582 ;
  assign n71584 = ~n71544 & n71583 ;
  assign n71576 = ~n71558 & n71564 ;
  assign n71585 = ~n71550 & n71576 ;
  assign n71570 = decrypt_pad & ~\u0_uk_K_r0_reg[20]/NET0131  ;
  assign n71571 = ~decrypt_pad & ~\u0_uk_K_r0_reg[41]/NET0131  ;
  assign n71572 = ~n71570 & ~n71571 ;
  assign n71573 = \u0_R0_reg[11]/NET0131  & ~n71572 ;
  assign n71574 = ~\u0_R0_reg[11]/NET0131  & n71572 ;
  assign n71575 = ~n71573 & ~n71574 ;
  assign n71586 = ~n71544 & ~n71575 ;
  assign n71587 = n71585 & n71586 ;
  assign n71588 = ~n71584 & ~n71587 ;
  assign n71551 = n71544 & n71550 ;
  assign n71552 = ~n71544 & ~n71550 ;
  assign n71565 = ~n71558 & ~n71564 ;
  assign n71566 = n71558 & n71564 ;
  assign n71567 = ~n71565 & ~n71566 ;
  assign n71568 = ~n71552 & ~n71567 ;
  assign n71569 = ~n71551 & n71568 ;
  assign n71577 = n71551 & n71576 ;
  assign n71578 = ~n71575 & n71577 ;
  assign n71579 = n71544 & ~n71564 ;
  assign n71580 = n71550 & n71558 ;
  assign n71581 = n71579 & n71580 ;
  assign n71589 = n71544 & ~n71550 ;
  assign n71590 = ~n71558 & n71575 ;
  assign n71591 = n71589 & n71590 ;
  assign n71592 = ~n71581 & ~n71591 ;
  assign n71593 = ~n71578 & n71592 ;
  assign n71594 = ~n71569 & n71593 ;
  assign n71595 = n71588 & n71594 ;
  assign n71596 = ~n71538 & ~n71595 ;
  assign n71597 = ~n71544 & n71564 ;
  assign n71609 = n71558 & n71579 ;
  assign n71610 = n71550 & n71576 ;
  assign n71611 = ~n71609 & ~n71610 ;
  assign n71612 = ~n71597 & n71611 ;
  assign n71613 = n71538 & n71575 ;
  assign n71614 = ~n71612 & n71613 ;
  assign n71605 = ~n71575 & ~n71579 ;
  assign n71604 = ~n71558 & ~n71589 ;
  assign n71606 = n71538 & ~n71597 ;
  assign n71607 = ~n71604 & n71606 ;
  assign n71608 = n71605 & n71607 ;
  assign n71598 = n71550 & n71597 ;
  assign n71599 = n71552 & n71565 ;
  assign n71600 = ~n71598 & ~n71599 ;
  assign n71601 = n71575 & ~n71600 ;
  assign n71602 = n71538 & n71551 ;
  assign n71603 = n71565 & n71602 ;
  assign n71615 = ~n71601 & ~n71603 ;
  assign n71616 = ~n71608 & n71615 ;
  assign n71617 = ~n71614 & n71616 ;
  assign n71618 = ~n71596 & n71617 ;
  assign n71619 = ~\u0_L0_reg[6]/NET0131  & ~n71618 ;
  assign n71620 = \u0_L0_reg[6]/NET0131  & n71618 ;
  assign n71621 = ~n71619 & ~n71620 ;
  assign n71622 = decrypt_pad & ~\u0_uk_K_r0_reg[9]/NET0131  ;
  assign n71623 = ~decrypt_pad & ~\u0_uk_K_r0_reg[30]/NET0131  ;
  assign n71624 = ~n71622 & ~n71623 ;
  assign n71625 = \u0_R0_reg[20]/NET0131  & ~n71624 ;
  assign n71626 = ~\u0_R0_reg[20]/NET0131  & n71624 ;
  assign n71627 = ~n71625 & ~n71626 ;
  assign n71628 = decrypt_pad & ~\u0_uk_K_r0_reg[7]/NET0131  ;
  assign n71629 = ~decrypt_pad & ~\u0_uk_K_r0_reg[28]/NET0131  ;
  assign n71630 = ~n71628 & ~n71629 ;
  assign n71631 = \u0_R0_reg[18]/NET0131  & ~n71630 ;
  assign n71632 = ~\u0_R0_reg[18]/NET0131  & n71630 ;
  assign n71633 = ~n71631 & ~n71632 ;
  assign n71648 = decrypt_pad & ~\u0_uk_K_r0_reg[38]/NET0131  ;
  assign n71649 = ~decrypt_pad & ~\u0_uk_K_r0_reg[0]/NET0131  ;
  assign n71650 = ~n71648 & ~n71649 ;
  assign n71651 = \u0_R0_reg[21]/NET0131  & ~n71650 ;
  assign n71652 = ~\u0_R0_reg[21]/NET0131  & n71650 ;
  assign n71653 = ~n71651 & ~n71652 ;
  assign n71655 = decrypt_pad & ~\u0_uk_K_r0_reg[49]/NET0131  ;
  assign n71656 = ~decrypt_pad & ~\u0_uk_K_r0_reg[15]/NET0131  ;
  assign n71657 = ~n71655 & ~n71656 ;
  assign n71658 = \u0_R0_reg[19]/NET0131  & ~n71657 ;
  assign n71659 = ~\u0_R0_reg[19]/NET0131  & n71657 ;
  assign n71660 = ~n71658 & ~n71659 ;
  assign n71634 = decrypt_pad & ~\u0_uk_K_r0_reg[44]/NET0131  ;
  assign n71635 = ~decrypt_pad & ~\u0_uk_K_r0_reg[38]/NET0131  ;
  assign n71636 = ~n71634 & ~n71635 ;
  assign n71637 = \u0_R0_reg[17]/NET0131  & ~n71636 ;
  assign n71638 = ~\u0_R0_reg[17]/NET0131  & n71636 ;
  assign n71639 = ~n71637 & ~n71638 ;
  assign n71641 = decrypt_pad & ~\u0_uk_K_r0_reg[22]/NET0131  ;
  assign n71642 = ~decrypt_pad & ~\u0_uk_K_r0_reg[43]/NET0131  ;
  assign n71643 = ~n71641 & ~n71642 ;
  assign n71644 = \u0_R0_reg[16]/NET0131  & ~n71643 ;
  assign n71645 = ~\u0_R0_reg[16]/NET0131  & n71643 ;
  assign n71646 = ~n71644 & ~n71645 ;
  assign n71669 = ~n71639 & ~n71646 ;
  assign n71698 = ~n71660 & n71669 ;
  assign n71699 = ~n71653 & n71698 ;
  assign n71661 = n71646 & n71653 ;
  assign n71702 = ~n71639 & n71661 ;
  assign n71667 = n71639 & ~n71653 ;
  assign n71694 = n71646 & n71667 ;
  assign n71692 = ~n71646 & n71653 ;
  assign n71700 = n71639 & ~n71660 ;
  assign n71701 = n71692 & n71700 ;
  assign n71703 = ~n71694 & ~n71701 ;
  assign n71704 = ~n71702 & n71703 ;
  assign n71705 = ~n71699 & n71704 ;
  assign n71706 = ~n71633 & ~n71705 ;
  assign n71664 = n71646 & ~n71653 ;
  assign n71665 = ~n71639 & n71664 ;
  assign n71688 = n71639 & n71661 ;
  assign n71689 = ~n71660 & n71688 ;
  assign n71690 = ~n71665 & ~n71689 ;
  assign n71691 = n71633 & ~n71690 ;
  assign n71662 = ~n71633 & n71661 ;
  assign n71640 = ~n71633 & n71639 ;
  assign n71693 = ~n71640 & n71692 ;
  assign n71695 = ~n71662 & ~n71693 ;
  assign n71696 = ~n71694 & n71695 ;
  assign n71697 = n71660 & ~n71696 ;
  assign n71707 = ~n71691 & ~n71697 ;
  assign n71708 = ~n71706 & n71707 ;
  assign n71709 = n71627 & ~n71708 ;
  assign n71666 = ~n71633 & n71665 ;
  assign n71663 = n71639 & n71662 ;
  assign n71668 = n71633 & n71667 ;
  assign n71670 = n71653 & n71669 ;
  assign n71671 = ~n71668 & ~n71670 ;
  assign n71672 = ~n71663 & n71671 ;
  assign n71673 = ~n71666 & n71672 ;
  assign n71674 = ~n71660 & ~n71673 ;
  assign n71677 = n71633 & n71653 ;
  assign n71678 = n71646 & n71677 ;
  assign n71647 = n71640 & ~n71646 ;
  assign n71675 = ~n71646 & ~n71653 ;
  assign n71676 = ~n71639 & n71675 ;
  assign n71679 = ~n71647 & ~n71676 ;
  assign n71680 = ~n71678 & n71679 ;
  assign n71681 = n71660 & ~n71680 ;
  assign n71654 = n71647 & ~n71653 ;
  assign n71682 = n71633 & ~n71639 ;
  assign n71683 = n71661 & n71682 ;
  assign n71684 = ~n71654 & ~n71683 ;
  assign n71685 = ~n71681 & n71684 ;
  assign n71686 = ~n71674 & n71685 ;
  assign n71687 = ~n71627 & ~n71686 ;
  assign n71710 = ~n71646 & n71667 ;
  assign n71711 = ~n71670 & ~n71710 ;
  assign n71712 = n71633 & ~n71711 ;
  assign n71713 = ~n71660 & n71712 ;
  assign n71714 = ~n71633 & n71694 ;
  assign n71715 = n71675 & n71682 ;
  assign n71716 = ~n71714 & ~n71715 ;
  assign n71717 = n71660 & ~n71716 ;
  assign n71718 = ~n71713 & ~n71717 ;
  assign n71719 = ~n71687 & n71718 ;
  assign n71720 = ~n71709 & n71719 ;
  assign n71721 = ~\u0_L0_reg[14]/NET0131  & ~n71720 ;
  assign n71722 = \u0_L0_reg[14]/NET0131  & n71720 ;
  assign n71723 = ~n71721 & ~n71722 ;
  assign n71726 = ~n70790 & ~n70844 ;
  assign n71725 = ~n70773 & ~n70798 ;
  assign n71727 = ~n70783 & ~n71725 ;
  assign n71728 = ~n71726 & n71727 ;
  assign n71724 = ~n70790 & ~n70999 ;
  assign n71729 = ~n70822 & ~n71724 ;
  assign n71730 = ~n71728 & n71729 ;
  assign n71732 = n70780 & ~n70999 ;
  assign n71736 = n70822 & ~n70828 ;
  assign n71737 = ~n70833 & n71736 ;
  assign n71731 = n70783 & n70790 ;
  assign n71733 = n70790 & ~n70827 ;
  assign n71734 = ~n70767 & ~n70800 ;
  assign n71735 = ~n71733 & n71734 ;
  assign n71738 = ~n71731 & ~n71735 ;
  assign n71739 = n71737 & n71738 ;
  assign n71740 = ~n71732 & n71739 ;
  assign n71741 = ~n71730 & ~n71740 ;
  assign n71742 = n70832 & ~n70843 ;
  assign n71743 = ~n71741 & n71742 ;
  assign n71744 = ~\u0_L0_reg[19]/P0001  & ~n71743 ;
  assign n71745 = \u0_L0_reg[19]/P0001  & n71743 ;
  assign n71746 = ~n71744 & ~n71745 ;
  assign n71750 = ~n71633 & ~n71639 ;
  assign n71751 = n71633 & ~n71646 ;
  assign n71752 = ~n71750 & ~n71751 ;
  assign n71753 = ~n71653 & ~n71752 ;
  assign n71754 = ~n71669 & ~n71688 ;
  assign n71755 = ~n71753 & n71754 ;
  assign n71756 = n71660 & ~n71755 ;
  assign n71747 = ~n71647 & ~n71702 ;
  assign n71748 = ~n71660 & ~n71747 ;
  assign n71749 = n71640 & n71653 ;
  assign n71757 = n71633 & n71694 ;
  assign n71758 = ~n71749 & ~n71757 ;
  assign n71759 = ~n71748 & n71758 ;
  assign n71760 = ~n71756 & n71759 ;
  assign n71761 = n71627 & ~n71760 ;
  assign n71769 = n71660 & n71667 ;
  assign n71770 = ~n71698 & ~n71769 ;
  assign n71771 = ~n71633 & ~n71770 ;
  assign n71768 = ~n71660 & n71665 ;
  assign n71772 = ~n71653 & n71660 ;
  assign n71773 = n71639 & n71751 ;
  assign n71774 = ~n71772 & n71773 ;
  assign n71775 = ~n71768 & ~n71774 ;
  assign n71776 = ~n71771 & n71775 ;
  assign n71777 = ~n71627 & ~n71776 ;
  assign n71762 = ~n71715 & ~n71757 ;
  assign n71763 = n71692 & n71750 ;
  assign n71764 = n71762 & ~n71763 ;
  assign n71765 = n71660 & ~n71764 ;
  assign n71766 = n71646 & ~n71660 ;
  assign n71767 = n71682 & n71766 ;
  assign n71778 = ~n71663 & ~n71767 ;
  assign n71779 = ~n71765 & n71778 ;
  assign n71780 = ~n71777 & n71779 ;
  assign n71781 = ~n71761 & n71780 ;
  assign n71782 = ~\u0_L0_reg[25]/NET0131  & ~n71781 ;
  assign n71783 = \u0_L0_reg[25]/NET0131  & n71781 ;
  assign n71784 = ~n71782 & ~n71783 ;
  assign n71789 = ~n71032 & n71045 ;
  assign n71790 = ~n71055 & ~n71789 ;
  assign n71788 = n71045 & n71055 ;
  assign n71791 = ~n71052 & ~n71788 ;
  assign n71792 = ~n71790 & n71791 ;
  assign n71785 = ~n71025 & ~n71045 ;
  assign n71786 = ~n71069 & ~n71785 ;
  assign n71787 = ~n71067 & ~n71786 ;
  assign n71793 = ~n71038 & ~n71787 ;
  assign n71794 = ~n71792 & n71793 ;
  assign n71795 = n71038 & ~n71054 ;
  assign n71796 = ~n71092 & n71795 ;
  assign n71797 = ~n71794 & ~n71796 ;
  assign n71798 = n71045 & ~n71108 ;
  assign n71804 = n71067 & ~n71083 ;
  assign n71805 = ~n71798 & n71804 ;
  assign n71799 = n71068 & n71105 ;
  assign n71800 = ~n71060 & ~n71799 ;
  assign n71801 = ~n71038 & ~n71800 ;
  assign n71802 = ~n71039 & ~n71053 ;
  assign n71803 = n71052 & ~n71802 ;
  assign n71806 = ~n71801 & ~n71803 ;
  assign n71807 = n71805 & n71806 ;
  assign n71808 = n71085 & n71789 ;
  assign n71809 = ~n71067 & ~n71091 ;
  assign n71810 = ~n71808 & n71809 ;
  assign n71811 = n71058 & n71810 ;
  assign n71812 = ~n71807 & ~n71811 ;
  assign n71813 = ~n71797 & ~n71812 ;
  assign n71814 = ~\u0_L0_reg[26]/NET0131  & ~n71813 ;
  assign n71815 = \u0_L0_reg[26]/NET0131  & n71813 ;
  assign n71816 = ~n71814 & ~n71815 ;
  assign n71821 = n71202 & ~n71208 ;
  assign n71820 = n71182 & n71208 ;
  assign n71822 = n71154 & ~n71820 ;
  assign n71823 = ~n71821 & n71822 ;
  assign n71824 = ~n71476 & n71823 ;
  assign n71825 = ~n71215 & ~n71487 ;
  assign n71826 = ~n71154 & ~n71481 ;
  assign n71827 = ~n71493 & n71826 ;
  assign n71828 = ~n71218 & n71827 ;
  assign n71829 = n71825 & n71828 ;
  assign n71830 = ~n71824 & ~n71829 ;
  assign n71817 = ~n71154 & ~n71166 ;
  assign n71818 = ~n71172 & n71204 ;
  assign n71819 = ~n71817 & n71818 ;
  assign n71831 = ~n71198 & ~n71819 ;
  assign n71832 = ~n71830 & n71831 ;
  assign n71839 = n71192 & n71198 ;
  assign n71833 = ~n71172 & n71481 ;
  assign n71837 = ~n71204 & ~n71216 ;
  assign n71838 = n71817 & n71837 ;
  assign n71840 = ~n71833 & ~n71838 ;
  assign n71841 = n71839 & n71840 ;
  assign n71834 = n71172 & n71204 ;
  assign n71835 = ~n71217 & ~n71834 ;
  assign n71836 = n71154 & ~n71835 ;
  assign n71842 = n71825 & ~n71836 ;
  assign n71843 = n71841 & n71842 ;
  assign n71844 = ~n71832 & ~n71843 ;
  assign n71845 = ~\u0_L0_reg[13]/NET0131  & ~n71844 ;
  assign n71846 = \u0_L0_reg[13]/NET0131  & n71844 ;
  assign n71847 = ~n71845 & ~n71846 ;
  assign n71849 = ~n71633 & n71676 ;
  assign n71850 = ~n71702 & ~n71849 ;
  assign n71851 = n71660 & ~n71850 ;
  assign n71848 = ~n71633 & n71766 ;
  assign n71852 = n71627 & ~n71848 ;
  assign n71853 = ~n71712 & n71852 ;
  assign n71854 = ~n71851 & n71853 ;
  assign n71855 = n71660 & ~n71666 ;
  assign n71856 = ~n71688 & n71855 ;
  assign n71857 = ~n71682 & n71692 ;
  assign n71858 = ~n71660 & ~n71702 ;
  assign n71859 = ~n71857 & n71858 ;
  assign n71860 = ~n71856 & ~n71859 ;
  assign n71861 = ~n71627 & ~n71647 ;
  assign n71862 = n71762 & n71861 ;
  assign n71863 = ~n71860 & n71862 ;
  assign n71864 = ~n71854 & ~n71863 ;
  assign n71865 = ~n71653 & n71767 ;
  assign n71866 = ~n71640 & ~n71682 ;
  assign n71867 = n71692 & ~n71866 ;
  assign n71868 = ~n71668 & ~n71867 ;
  assign n71869 = n71660 & ~n71868 ;
  assign n71870 = ~n71865 & ~n71869 ;
  assign n71871 = ~n71864 & n71870 ;
  assign n71872 = ~\u0_L0_reg[8]/NET0131  & ~n71871 ;
  assign n71873 = \u0_L0_reg[8]/NET0131  & n71871 ;
  assign n71874 = ~n71872 & ~n71873 ;
  assign n71875 = n71544 & n71565 ;
  assign n71876 = n71575 & n71875 ;
  assign n71877 = n71544 & n71566 ;
  assign n71878 = ~n71544 & ~n71566 ;
  assign n71879 = ~n71877 & ~n71878 ;
  assign n71880 = ~n71565 & ~n71879 ;
  assign n71881 = ~n71876 & ~n71880 ;
  assign n71882 = ~n71550 & ~n71881 ;
  assign n71883 = n71550 & n71565 ;
  assign n71884 = ~n71583 & ~n71883 ;
  assign n71885 = ~n71575 & ~n71884 ;
  assign n71886 = n71538 & ~n71577 ;
  assign n71887 = ~n71885 & n71886 ;
  assign n71888 = ~n71882 & n71887 ;
  assign n71889 = ~n71582 & ~n71597 ;
  assign n71890 = ~n71558 & ~n71889 ;
  assign n71891 = ~n71877 & ~n71890 ;
  assign n71892 = ~n71575 & ~n71891 ;
  assign n71893 = ~n71565 & n71575 ;
  assign n71894 = n71879 & n71893 ;
  assign n71895 = ~n71538 & ~n71599 ;
  assign n71896 = ~n71894 & n71895 ;
  assign n71897 = ~n71892 & n71896 ;
  assign n71898 = ~n71888 & ~n71897 ;
  assign n71899 = ~n71544 & n71580 ;
  assign n71900 = ~n71575 & ~n71899 ;
  assign n71901 = ~n71544 & n71883 ;
  assign n71902 = n71575 & ~n71581 ;
  assign n71903 = ~n71901 & n71902 ;
  assign n71904 = ~n71900 & ~n71903 ;
  assign n71905 = ~n71898 & ~n71904 ;
  assign n71906 = ~\u0_L0_reg[16]/NET0131  & ~n71905 ;
  assign n71907 = \u0_L0_reg[16]/NET0131  & n71905 ;
  assign n71908 = ~n71906 & ~n71907 ;
  assign n71914 = ~n70878 & ~n70933 ;
  assign n71909 = ~n70896 & ~n70910 ;
  assign n71910 = n70893 & ~n71909 ;
  assign n71915 = n70879 & ~n70887 ;
  assign n71916 = ~n71910 & ~n71915 ;
  assign n71917 = ~n71914 & n71916 ;
  assign n71918 = ~n70902 & ~n71917 ;
  assign n71911 = ~n70927 & ~n71910 ;
  assign n71912 = n70872 & ~n71911 ;
  assign n71919 = ~n70872 & ~n70904 ;
  assign n71920 = n71909 & n71919 ;
  assign n71921 = n70902 & n71920 ;
  assign n71922 = ~n71912 & ~n71921 ;
  assign n71923 = ~n71918 & n71922 ;
  assign n71924 = n70866 & ~n71923 ;
  assign n71925 = n70866 & ~n70902 ;
  assign n71926 = ~n70902 & n71920 ;
  assign n71927 = n70921 & n70924 ;
  assign n71928 = ~n71926 & ~n71927 ;
  assign n71929 = ~n71925 & ~n71928 ;
  assign n71913 = ~n70902 & n71912 ;
  assign n71931 = n70872 & ~n70926 ;
  assign n71932 = n71909 & ~n71931 ;
  assign n71930 = n70932 & ~n71909 ;
  assign n71933 = ~n70866 & n70902 ;
  assign n71934 = ~n71930 & n71933 ;
  assign n71935 = ~n71932 & n71934 ;
  assign n71936 = ~n71913 & ~n71935 ;
  assign n71937 = ~n71929 & n71936 ;
  assign n71938 = ~n71924 & n71937 ;
  assign n71939 = ~\u0_L0_reg[7]/NET0131  & ~n71938 ;
  assign n71940 = \u0_L0_reg[7]/NET0131  & n71938 ;
  assign n71941 = ~n71939 & ~n71940 ;
  assign n71944 = ~n70712 & ~n70973 ;
  assign n71945 = ~n70699 & ~n71944 ;
  assign n71946 = n70690 & n70715 ;
  assign n71947 = n70683 & ~n70970 ;
  assign n71948 = ~n71946 & n71947 ;
  assign n71942 = n70719 & ~n70747 ;
  assign n71943 = ~n70683 & n71942 ;
  assign n71949 = ~n70707 & ~n71943 ;
  assign n71950 = ~n71948 & n71949 ;
  assign n71951 = ~n71945 & n71950 ;
  assign n71953 = n70676 & n71412 ;
  assign n71954 = n70739 & n71942 ;
  assign n71952 = n70715 & n70747 ;
  assign n71955 = n70707 & ~n71952 ;
  assign n71956 = ~n71954 & n71955 ;
  assign n71957 = ~n71953 & n71956 ;
  assign n71958 = ~n71951 & ~n71957 ;
  assign n71959 = n70696 & n70735 ;
  assign n71960 = ~n70716 & n71959 ;
  assign n71961 = ~n71958 & ~n71960 ;
  assign n71962 = ~\u0_L0_reg[9]/NET0131  & ~n71961 ;
  assign n71963 = \u0_L0_reg[9]/NET0131  & n71961 ;
  assign n71964 = ~n71962 & ~n71963 ;
  assign n71971 = ~n70923 & n71382 ;
  assign n71972 = n71909 & ~n71971 ;
  assign n71973 = ~n70923 & ~n71909 ;
  assign n71974 = ~n70902 & ~n71973 ;
  assign n71975 = ~n71972 & n71974 ;
  assign n71965 = n70910 & n70932 ;
  assign n71966 = ~n70926 & ~n70934 ;
  assign n71967 = ~n70911 & n71966 ;
  assign n71968 = ~n70893 & n70924 ;
  assign n71969 = ~n71967 & ~n71968 ;
  assign n71970 = n70902 & ~n71969 ;
  assign n71976 = ~n71965 & ~n71970 ;
  assign n71977 = ~n71975 & n71976 ;
  assign n71978 = n70866 & ~n71977 ;
  assign n71980 = ~n70872 & n70910 ;
  assign n71981 = n71383 & ~n71980 ;
  assign n71982 = n70935 & ~n71966 ;
  assign n71979 = n70914 & n70934 ;
  assign n71983 = n70879 & n70894 ;
  assign n71984 = ~n71979 & ~n71983 ;
  assign n71985 = n70945 & n71984 ;
  assign n71986 = ~n71982 & n71985 ;
  assign n71987 = ~n71981 & n71986 ;
  assign n71988 = ~n70866 & ~n71987 ;
  assign n71989 = n70872 & n71384 ;
  assign n71990 = ~n70934 & n70942 ;
  assign n71991 = n70881 & n71990 ;
  assign n71992 = ~n71989 & ~n71991 ;
  assign n71993 = ~n71988 & n71992 ;
  assign n71994 = ~n71978 & n71993 ;
  assign n71995 = \u0_L0_reg[32]/NET0131  & n71994 ;
  assign n71996 = ~\u0_L0_reg[32]/NET0131  & ~n71994 ;
  assign n71997 = ~n71995 & ~n71996 ;
  assign n71999 = ~n71277 & n71503 ;
  assign n72000 = n71265 & ~n71999 ;
  assign n72001 = ~n71315 & n71330 ;
  assign n72002 = n71266 & ~n72001 ;
  assign n72003 = ~n72000 & ~n72002 ;
  assign n71998 = ~n71245 & n71293 ;
  assign n72004 = n71291 & ~n71317 ;
  assign n72005 = ~n71998 & n72004 ;
  assign n72006 = ~n71284 & n72005 ;
  assign n72007 = ~n72003 & n72006 ;
  assign n72011 = n71265 & ~n71283 ;
  assign n72010 = n71273 & ~n71276 ;
  assign n72012 = ~n71306 & ~n72010 ;
  assign n72013 = n72011 & n72012 ;
  assign n72008 = ~n71299 & ~n71352 ;
  assign n72009 = n71245 & ~n72008 ;
  assign n72014 = ~n71291 & ~n71351 ;
  assign n72015 = ~n72009 & n72014 ;
  assign n72016 = ~n72013 & n72015 ;
  assign n72017 = ~n72007 & ~n72016 ;
  assign n72018 = ~n71278 & ~n71294 ;
  assign n72019 = ~n71513 & n72018 ;
  assign n72020 = ~n71265 & ~n72019 ;
  assign n72021 = n71265 & ~n71273 ;
  assign n72022 = n71304 & n72021 ;
  assign n72023 = ~n72020 & ~n72022 ;
  assign n72024 = ~n72017 & n72023 ;
  assign n72025 = ~\u0_L0_reg[27]/NET0131  & ~n72024 ;
  assign n72026 = \u0_L0_reg[27]/NET0131  & n72024 ;
  assign n72027 = ~n72025 & ~n72026 ;
  assign n72028 = ~n71579 & n71580 ;
  assign n72029 = n71544 & n71582 ;
  assign n72030 = ~n72028 & ~n72029 ;
  assign n72031 = n71575 & ~n72030 ;
  assign n72032 = ~n71544 & ~n71558 ;
  assign n72033 = ~n71580 & ~n72032 ;
  assign n72034 = n71605 & n72033 ;
  assign n72037 = ~n71538 & ~n72034 ;
  assign n72035 = n71552 & ~n71567 ;
  assign n72036 = ~n71544 & n71610 ;
  assign n72038 = ~n72035 & ~n72036 ;
  assign n72039 = n72037 & n72038 ;
  assign n72040 = ~n72031 & n72039 ;
  assign n72043 = ~n71585 & ~n71883 ;
  assign n72044 = ~n71584 & n72043 ;
  assign n72045 = n71575 & ~n72044 ;
  assign n72041 = ~n71580 & ~n71875 ;
  assign n72042 = ~n71575 & ~n72041 ;
  assign n72046 = n71538 & ~n72042 ;
  assign n72047 = ~n72045 & n72046 ;
  assign n72048 = ~n72040 & ~n72047 ;
  assign n72052 = n71564 & n71575 ;
  assign n72053 = n71899 & n72052 ;
  assign n72049 = ~n71566 & n71602 ;
  assign n72050 = n71550 & ~n71575 ;
  assign n72051 = n71579 & n72050 ;
  assign n72054 = ~n72049 & ~n72051 ;
  assign n72055 = ~n72053 & n72054 ;
  assign n72056 = ~n72048 & n72055 ;
  assign n72057 = \u0_L0_reg[30]/P0001  & ~n72056 ;
  assign n72058 = ~\u0_L0_reg[30]/P0001  & n72056 ;
  assign n72059 = ~n72057 & ~n72058 ;
  assign n72074 = n71154 & ~n71209 ;
  assign n72075 = n71160 & n71172 ;
  assign n72076 = ~n71154 & ~n72075 ;
  assign n72077 = n71483 & n72076 ;
  assign n72078 = ~n71181 & ~n72077 ;
  assign n72079 = ~n72074 & n72078 ;
  assign n72080 = n71198 & ~n72079 ;
  assign n72061 = ~n71179 & ~n71219 ;
  assign n72062 = ~n71216 & ~n72061 ;
  assign n72063 = ~n71173 & ~n71232 ;
  assign n72064 = ~n72062 & n72063 ;
  assign n72060 = n71199 & n71219 ;
  assign n72065 = ~n71200 & ~n72060 ;
  assign n72066 = ~n71487 & n72065 ;
  assign n72067 = ~n72064 & n72066 ;
  assign n72068 = ~n71198 & ~n72067 ;
  assign n72069 = n71160 & n71202 ;
  assign n72070 = ~n71833 & ~n72069 ;
  assign n72071 = n71154 & ~n72070 ;
  assign n72072 = ~n71154 & n71166 ;
  assign n72073 = n71204 & n72072 ;
  assign n72081 = ~n72071 & ~n72073 ;
  assign n72082 = ~n72068 & n72081 ;
  assign n72083 = ~n72080 & n72082 ;
  assign n72084 = ~\u0_L0_reg[18]/NET0131  & ~n72083 ;
  assign n72085 = \u0_L0_reg[18]/NET0131  & n72083 ;
  assign n72086 = ~n72084 & ~n72085 ;
  assign n72098 = ~n71564 & n71899 ;
  assign n72099 = ~n71875 & ~n71899 ;
  assign n72100 = n72043 & n72099 ;
  assign n72101 = n71575 & ~n72100 ;
  assign n72102 = ~n72098 & ~n72101 ;
  assign n72103 = ~n71538 & ~n72102 ;
  assign n72088 = n71552 & n71575 ;
  assign n72089 = ~n71576 & n72088 ;
  assign n72094 = n71588 & ~n72089 ;
  assign n72090 = n71544 & n71580 ;
  assign n72091 = ~n71610 & ~n72090 ;
  assign n72092 = n71575 & ~n72091 ;
  assign n72093 = n71568 & ~n71575 ;
  assign n72095 = ~n72092 & ~n72093 ;
  assign n72096 = n72094 & n72095 ;
  assign n72097 = n71538 & ~n72096 ;
  assign n72104 = n71611 & ~n72035 ;
  assign n72105 = ~n71538 & ~n71575 ;
  assign n72106 = ~n72104 & n72105 ;
  assign n72108 = n71575 & n71584 ;
  assign n72087 = n71877 & n72050 ;
  assign n72107 = n71564 & n71591 ;
  assign n72109 = ~n72087 & ~n72107 ;
  assign n72110 = ~n72108 & n72109 ;
  assign n72111 = ~n72106 & n72110 ;
  assign n72112 = ~n72097 & n72111 ;
  assign n72113 = ~n72103 & n72112 ;
  assign n72114 = ~\u0_L0_reg[24]/NET0131  & ~n72113 ;
  assign n72115 = \u0_L0_reg[24]/NET0131  & n72113 ;
  assign n72116 = ~n72114 & ~n72115 ;
  assign n72118 = ~n71662 & ~n71710 ;
  assign n72119 = n71660 & ~n72118 ;
  assign n72117 = n71633 & n71665 ;
  assign n72120 = ~n71663 & ~n71701 ;
  assign n72121 = ~n72117 & n72120 ;
  assign n72122 = ~n72119 & n72121 ;
  assign n72123 = n71627 & ~n72122 ;
  assign n72125 = ~n71633 & n71692 ;
  assign n72126 = ~n71664 & ~n71682 ;
  assign n72127 = ~n71665 & ~n72126 ;
  assign n72128 = ~n72125 & ~n72127 ;
  assign n72129 = ~n71627 & ~n72128 ;
  assign n72124 = n71633 & n71670 ;
  assign n72130 = n71855 & ~n72124 ;
  assign n72131 = ~n72129 & n72130 ;
  assign n72132 = n71627 & ~n71683 ;
  assign n72133 = ~n71675 & ~n71677 ;
  assign n72134 = ~n71702 & n72133 ;
  assign n72135 = ~n72132 & ~n72134 ;
  assign n72136 = ~n71660 & ~n71714 ;
  assign n72137 = ~n71849 & n72136 ;
  assign n72138 = ~n72135 & n72137 ;
  assign n72139 = ~n72131 & ~n72138 ;
  assign n72140 = ~n72123 & ~n72139 ;
  assign n72141 = ~\u0_L0_reg[3]/NET0131  & ~n72140 ;
  assign n72142 = \u0_L0_reg[3]/NET0131  & n72140 ;
  assign n72143 = ~n72141 & ~n72142 ;
  assign n72144 = decrypt_pad & ~\u0_key_r_reg[35]/P0001  ;
  assign n72145 = ~decrypt_pad & ~\u0_key_r_reg[42]/P0001  ;
  assign n72146 = ~n72144 & ~n72145 ;
  assign n72147 = \u0_desIn_r_reg[25]/NET0131  & ~n72146 ;
  assign n72148 = ~\u0_desIn_r_reg[25]/NET0131  & n72146 ;
  assign n72149 = ~n72147 & ~n72148 ;
  assign n72169 = decrypt_pad & ~\u0_key_r_reg[15]/NET0131  ;
  assign n72170 = ~decrypt_pad & ~\u0_key_r_reg[22]/NET0131  ;
  assign n72171 = ~n72169 & ~n72170 ;
  assign n72172 = \u0_desIn_r_reg[9]/NET0131  & ~n72171 ;
  assign n72173 = ~\u0_desIn_r_reg[9]/NET0131  & n72171 ;
  assign n72174 = ~n72172 & ~n72173 ;
  assign n72150 = decrypt_pad & ~\u0_key_r_reg[50]/NET0131  ;
  assign n72151 = ~decrypt_pad & ~\u0_key_r_reg[2]/NET0131  ;
  assign n72152 = ~n72150 & ~n72151 ;
  assign n72153 = \u0_desIn_r_reg[59]/NET0131  & ~n72152 ;
  assign n72154 = ~\u0_desIn_r_reg[59]/NET0131  & n72152 ;
  assign n72155 = ~n72153 & ~n72154 ;
  assign n72156 = decrypt_pad & ~\u0_key_r_reg[31]/NET0131  ;
  assign n72157 = ~decrypt_pad & ~\u0_key_r_reg[38]/NET0131  ;
  assign n72158 = ~n72156 & ~n72157 ;
  assign n72159 = \u0_desIn_r_reg[33]/NET0131  & ~n72158 ;
  assign n72160 = ~\u0_desIn_r_reg[33]/NET0131  & n72158 ;
  assign n72161 = ~n72159 & ~n72160 ;
  assign n72177 = decrypt_pad & ~\u0_key_r_reg[30]/NET0131  ;
  assign n72178 = ~decrypt_pad & ~\u0_key_r_reg[37]/NET0131  ;
  assign n72179 = ~n72177 & ~n72178 ;
  assign n72180 = \u0_desIn_r_reg[1]/NET0131  & ~n72179 ;
  assign n72181 = ~\u0_desIn_r_reg[1]/NET0131  & n72179 ;
  assign n72182 = ~n72180 & ~n72181 ;
  assign n72193 = n72161 & n72182 ;
  assign n72225 = ~n72155 & n72193 ;
  assign n72227 = n72174 & ~n72225 ;
  assign n72163 = decrypt_pad & ~\u0_key_r_reg[52]/NET0131  ;
  assign n72164 = ~decrypt_pad & ~\u0_key_r_reg[0]/NET0131  ;
  assign n72165 = ~n72163 & ~n72164 ;
  assign n72166 = \u0_desIn_r_reg[17]/NET0131  & ~n72165 ;
  assign n72167 = ~\u0_desIn_r_reg[17]/NET0131  & n72165 ;
  assign n72168 = ~n72166 & ~n72167 ;
  assign n72188 = n72155 & n72161 ;
  assign n72224 = ~n72182 & n72188 ;
  assign n72226 = ~n72224 & ~n72225 ;
  assign n72228 = ~n72168 & ~n72226 ;
  assign n72229 = ~n72227 & n72228 ;
  assign n72219 = n72155 & n72174 ;
  assign n72220 = ~n72182 & n72219 ;
  assign n72195 = n72155 & ~n72174 ;
  assign n72221 = n72193 & n72195 ;
  assign n72222 = ~n72220 & ~n72221 ;
  assign n72223 = n72168 & ~n72222 ;
  assign n72162 = ~n72155 & n72161 ;
  assign n72207 = n72162 & ~n72182 ;
  assign n72208 = n72174 & n72207 ;
  assign n72198 = ~n72174 & ~n72182 ;
  assign n72217 = ~n72155 & n72198 ;
  assign n72218 = ~n72161 & n72217 ;
  assign n72230 = ~n72208 & ~n72218 ;
  assign n72231 = ~n72223 & n72230 ;
  assign n72232 = ~n72229 & n72231 ;
  assign n72233 = n72149 & ~n72232 ;
  assign n72183 = ~n72161 & ~n72182 ;
  assign n72184 = ~n72155 & n72183 ;
  assign n72185 = n72174 & n72184 ;
  assign n72186 = n72155 & n72182 ;
  assign n72187 = ~n72161 & n72186 ;
  assign n72189 = n72174 & n72188 ;
  assign n72190 = ~n72187 & ~n72189 ;
  assign n72191 = ~n72185 & n72190 ;
  assign n72192 = ~n72168 & ~n72191 ;
  assign n72199 = n72161 & ~n72168 ;
  assign n72200 = n72155 & n72198 ;
  assign n72201 = ~n72199 & n72200 ;
  assign n72175 = ~n72168 & ~n72174 ;
  assign n72176 = n72162 & n72175 ;
  assign n72194 = ~n72155 & n72174 ;
  assign n72196 = ~n72194 & ~n72195 ;
  assign n72197 = n72193 & n72196 ;
  assign n72202 = ~n72176 & ~n72197 ;
  assign n72203 = ~n72201 & n72202 ;
  assign n72204 = ~n72192 & n72203 ;
  assign n72205 = ~n72149 & ~n72204 ;
  assign n72209 = ~n72155 & ~n72161 ;
  assign n72210 = n72182 & n72209 ;
  assign n72211 = n72174 & n72210 ;
  assign n72206 = n72183 & ~n72194 ;
  assign n72212 = ~n72206 & ~n72208 ;
  assign n72213 = ~n72211 & n72212 ;
  assign n72214 = n72168 & ~n72213 ;
  assign n72215 = ~n72168 & n72182 ;
  assign n72216 = n72196 & n72215 ;
  assign n72234 = ~n72214 & ~n72216 ;
  assign n72235 = ~n72205 & n72234 ;
  assign n72236 = ~n72233 & n72235 ;
  assign n72237 = ~\u0_desIn_r_reg[42]/NET0131  & ~n72236 ;
  assign n72238 = \u0_desIn_r_reg[42]/NET0131  & n72236 ;
  assign n72239 = ~n72237 & ~n72238 ;
  assign n72259 = decrypt_pad & ~\u0_key_r_reg[40]/NET0131  ;
  assign n72260 = ~decrypt_pad & ~\u0_key_r_reg[47]/NET0131  ;
  assign n72261 = ~n72259 & ~n72260 ;
  assign n72262 = \u0_desIn_r_reg[57]/NET0131  & ~n72261 ;
  assign n72263 = ~\u0_desIn_r_reg[57]/NET0131  & n72261 ;
  assign n72264 = ~n72262 & ~n72263 ;
  assign n72240 = decrypt_pad & ~\u0_key_r_reg[53]/NET0131  ;
  assign n72241 = ~decrypt_pad & ~\u0_key_r_reg[3]/NET0131  ;
  assign n72242 = ~n72240 & ~n72241 ;
  assign n72243 = \u0_desIn_r_reg[23]/NET0131  & ~n72242 ;
  assign n72244 = ~\u0_desIn_r_reg[23]/NET0131  & n72242 ;
  assign n72245 = ~n72243 & ~n72244 ;
  assign n72253 = decrypt_pad & ~\u0_key_r_reg[4]/NET0131  ;
  assign n72254 = ~decrypt_pad & ~\u0_key_r_reg[11]/NET0131  ;
  assign n72255 = ~n72253 & ~n72254 ;
  assign n72256 = \u0_desIn_r_reg[7]/NET0131  & ~n72255 ;
  assign n72257 = ~\u0_desIn_r_reg[7]/NET0131  & n72255 ;
  assign n72258 = ~n72256 & ~n72257 ;
  assign n72308 = ~n72245 & n72258 ;
  assign n72267 = decrypt_pad & ~\u0_key_r_reg[34]/NET0131  ;
  assign n72268 = ~decrypt_pad & ~\u0_key_r_reg[41]/NET0131  ;
  assign n72269 = ~n72267 & ~n72268 ;
  assign n72270 = \u0_desIn_r_reg[39]/NET0131  & ~n72269 ;
  assign n72271 = ~\u0_desIn_r_reg[39]/NET0131  & n72269 ;
  assign n72272 = ~n72270 & ~n72271 ;
  assign n72246 = decrypt_pad & ~\u0_key_r_reg[19]/NET0131  ;
  assign n72247 = ~decrypt_pad & ~\u0_key_r_reg[26]/NET0131  ;
  assign n72248 = ~n72246 & ~n72247 ;
  assign n72249 = \u0_desIn_r_reg[15]/NET0131  & ~n72248 ;
  assign n72250 = ~\u0_desIn_r_reg[15]/NET0131  & n72248 ;
  assign n72251 = ~n72249 & ~n72250 ;
  assign n72309 = ~n72251 & ~n72258 ;
  assign n72310 = ~n72272 & n72309 ;
  assign n72311 = ~n72308 & ~n72310 ;
  assign n72312 = n72264 & ~n72311 ;
  assign n72280 = ~n72258 & n72272 ;
  assign n72300 = ~n72264 & ~n72272 ;
  assign n72301 = n72251 & n72300 ;
  assign n72302 = ~n72280 & ~n72301 ;
  assign n72303 = n72245 & ~n72302 ;
  assign n72287 = decrypt_pad & ~\u0_key_r_reg[6]/NET0131  ;
  assign n72288 = ~decrypt_pad & ~\u0_key_r_reg[13]/NET0131  ;
  assign n72289 = ~n72287 & ~n72288 ;
  assign n72290 = \u0_desIn_r_reg[31]/NET0131  & ~n72289 ;
  assign n72291 = ~\u0_desIn_r_reg[31]/NET0131  & n72289 ;
  assign n72292 = ~n72290 & ~n72291 ;
  assign n72252 = n72245 & ~n72251 ;
  assign n72304 = ~n72252 & n72258 ;
  assign n72274 = n72251 & ~n72264 ;
  assign n72305 = ~n72264 & n72272 ;
  assign n72306 = ~n72274 & ~n72305 ;
  assign n72307 = ~n72304 & ~n72306 ;
  assign n72313 = n72292 & ~n72307 ;
  assign n72314 = ~n72303 & n72313 ;
  assign n72315 = ~n72312 & n72314 ;
  assign n72277 = n72264 & n72272 ;
  assign n72319 = n72277 & ~n72308 ;
  assign n72316 = n72258 & ~n72272 ;
  assign n72320 = ~n72264 & n72316 ;
  assign n72321 = ~n72319 & ~n72320 ;
  assign n72322 = ~n72251 & ~n72321 ;
  assign n72275 = n72245 & n72274 ;
  assign n72323 = n72258 & n72272 ;
  assign n72324 = n72275 & n72323 ;
  assign n72284 = n72251 & n72264 ;
  assign n72317 = n72284 & n72316 ;
  assign n72318 = n72245 & n72317 ;
  assign n72325 = ~n72292 & ~n72318 ;
  assign n72326 = ~n72324 & n72325 ;
  assign n72327 = ~n72322 & n72326 ;
  assign n72328 = ~n72315 & ~n72327 ;
  assign n72282 = ~n72251 & ~n72264 ;
  assign n72283 = ~n72280 & n72282 ;
  assign n72273 = ~n72258 & ~n72272 ;
  assign n72285 = n72273 & n72284 ;
  assign n72286 = ~n72283 & ~n72285 ;
  assign n72293 = ~n72286 & ~n72292 ;
  assign n72278 = n72251 & n72277 ;
  assign n72279 = n72258 & n72278 ;
  assign n72281 = n72274 & n72280 ;
  assign n72294 = ~n72251 & n72258 ;
  assign n72295 = ~n72272 & n72294 ;
  assign n72296 = ~n72281 & ~n72295 ;
  assign n72297 = ~n72279 & n72296 ;
  assign n72298 = ~n72293 & n72297 ;
  assign n72299 = ~n72245 & ~n72298 ;
  assign n72265 = ~n72258 & n72264 ;
  assign n72266 = n72252 & n72265 ;
  assign n72276 = n72273 & n72275 ;
  assign n72329 = ~n72266 & ~n72276 ;
  assign n72330 = ~n72299 & n72329 ;
  assign n72331 = ~n72328 & n72330 ;
  assign n72332 = ~\u0_desIn_r_reg[48]/NET0131  & ~n72331 ;
  assign n72333 = \u0_desIn_r_reg[48]/NET0131  & n72331 ;
  assign n72334 = ~n72332 & ~n72333 ;
  assign n72335 = decrypt_pad & ~\u0_key_r_reg[54]/NET0131  ;
  assign n72336 = ~decrypt_pad & ~\u0_key_r_reg[4]/NET0131  ;
  assign n72337 = ~n72335 & ~n72336 ;
  assign n72338 = \u0_desIn_r_reg[29]/NET0131  & ~n72337 ;
  assign n72339 = ~\u0_desIn_r_reg[29]/NET0131  & n72337 ;
  assign n72340 = ~n72338 & ~n72339 ;
  assign n72341 = decrypt_pad & ~\u0_key_r_reg[13]/NET0131  ;
  assign n72342 = ~decrypt_pad & ~\u0_key_r_reg[20]/NET0131  ;
  assign n72343 = ~n72341 & ~n72342 ;
  assign n72344 = \u0_desIn_r_reg[3]/NET0131  & ~n72343 ;
  assign n72345 = ~\u0_desIn_r_reg[3]/NET0131  & n72343 ;
  assign n72346 = ~n72344 & ~n72345 ;
  assign n72347 = ~n72340 & n72346 ;
  assign n72354 = decrypt_pad & ~\u0_key_r_reg[48]/NET0131  ;
  assign n72355 = ~decrypt_pad & ~\u0_key_r_reg[55]/NET0131  ;
  assign n72356 = ~n72354 & ~n72355 ;
  assign n72357 = \u0_desIn_r_reg[37]/NET0131  & ~n72356 ;
  assign n72358 = ~\u0_desIn_r_reg[37]/NET0131  & n72356 ;
  assign n72359 = ~n72357 & ~n72358 ;
  assign n72362 = decrypt_pad & ~\u0_key_r_reg[17]/NET0131  ;
  assign n72363 = ~decrypt_pad & ~\u0_key_r_reg[24]/NET0131  ;
  assign n72364 = ~n72362 & ~n72363 ;
  assign n72365 = \u0_desIn_r_reg[45]/NET0131  & ~n72364 ;
  assign n72366 = ~\u0_desIn_r_reg[45]/NET0131  & n72364 ;
  assign n72367 = ~n72365 & ~n72366 ;
  assign n72368 = n72359 & ~n72367 ;
  assign n72369 = n72347 & n72368 ;
  assign n72370 = n72340 & n72346 ;
  assign n72371 = n72359 & n72370 ;
  assign n72372 = n72367 & n72371 ;
  assign n72373 = ~n72369 & ~n72372 ;
  assign n72382 = n72340 & ~n72346 ;
  assign n72348 = decrypt_pad & ~\u0_key_r_reg[25]/NET0131  ;
  assign n72349 = ~decrypt_pad & ~\u0_key_r_reg[32]/NET0131  ;
  assign n72350 = ~n72348 & ~n72349 ;
  assign n72351 = \u0_desIn_r_reg[53]/NET0131  & ~n72350 ;
  assign n72352 = ~\u0_desIn_r_reg[53]/NET0131  & n72350 ;
  assign n72353 = ~n72351 & ~n72352 ;
  assign n72383 = n72353 & n72359 ;
  assign n72384 = n72382 & n72383 ;
  assign n72360 = n72353 & ~n72359 ;
  assign n72361 = n72347 & n72360 ;
  assign n72385 = decrypt_pad & ~\u0_key_r_reg[33]/NET0131  ;
  assign n72386 = ~decrypt_pad & ~\u0_key_r_reg[40]/NET0131  ;
  assign n72387 = ~n72385 & ~n72386 ;
  assign n72388 = \u0_desIn_r_reg[61]/NET0131  & ~n72387 ;
  assign n72389 = ~\u0_desIn_r_reg[61]/NET0131  & n72387 ;
  assign n72390 = ~n72388 & ~n72389 ;
  assign n72391 = ~n72361 & n72390 ;
  assign n72392 = ~n72384 & n72391 ;
  assign n72374 = ~n72353 & ~n72367 ;
  assign n72375 = n72340 & n72359 ;
  assign n72376 = ~n72340 & ~n72359 ;
  assign n72377 = ~n72375 & ~n72376 ;
  assign n72378 = n72374 & n72377 ;
  assign n72379 = ~n72353 & n72367 ;
  assign n72380 = ~n72346 & n72376 ;
  assign n72381 = n72379 & n72380 ;
  assign n72393 = ~n72378 & ~n72381 ;
  assign n72394 = n72392 & n72393 ;
  assign n72395 = n72373 & n72394 ;
  assign n72401 = n72346 & ~n72359 ;
  assign n72407 = ~n72367 & n72401 ;
  assign n72408 = n72340 & n72407 ;
  assign n72397 = ~n72340 & n72367 ;
  assign n72398 = ~n72370 & ~n72397 ;
  assign n72399 = n72383 & ~n72398 ;
  assign n72404 = ~n72346 & n72359 ;
  assign n72405 = ~n72340 & n72404 ;
  assign n72406 = n72367 & n72405 ;
  assign n72410 = ~n72399 & ~n72406 ;
  assign n72411 = ~n72408 & n72410 ;
  assign n72400 = n72367 & n72382 ;
  assign n72402 = ~n72400 & ~n72401 ;
  assign n72403 = ~n72353 & ~n72402 ;
  assign n72396 = ~n72379 & n72380 ;
  assign n72409 = ~n72390 & ~n72396 ;
  assign n72412 = ~n72403 & n72409 ;
  assign n72413 = n72411 & n72412 ;
  assign n72414 = ~n72395 & ~n72413 ;
  assign n72415 = ~n72353 & ~n72369 ;
  assign n72416 = n72340 & ~n72367 ;
  assign n72417 = n72404 & n72416 ;
  assign n72418 = n72353 & ~n72417 ;
  assign n72419 = ~n72415 & ~n72418 ;
  assign n72420 = ~n72346 & ~n72367 ;
  assign n72421 = ~n72340 & n72420 ;
  assign n72422 = ~n72400 & ~n72421 ;
  assign n72423 = n72360 & ~n72422 ;
  assign n72424 = ~n72419 & ~n72423 ;
  assign n72425 = ~n72414 & n72424 ;
  assign n72426 = ~\u0_desIn_r_reg[26]/NET0131  & ~n72425 ;
  assign n72427 = \u0_desIn_r_reg[26]/NET0131  & n72425 ;
  assign n72428 = ~n72426 & ~n72427 ;
  assign n72435 = decrypt_pad & ~\u0_key_r_reg[9]/NET0131  ;
  assign n72436 = ~decrypt_pad & ~\u0_key_r_reg[16]/NET0131  ;
  assign n72437 = ~n72435 & ~n72436 ;
  assign n72438 = \u0_desIn_r_reg[25]/NET0131  & ~n72437 ;
  assign n72439 = ~\u0_desIn_r_reg[25]/NET0131  & n72437 ;
  assign n72440 = ~n72438 & ~n72439 ;
  assign n72441 = decrypt_pad & ~\u0_key_r_reg[21]/NET0131  ;
  assign n72442 = ~decrypt_pad & ~\u0_key_r_reg[28]/NET0131  ;
  assign n72443 = ~n72441 & ~n72442 ;
  assign n72444 = \u0_desIn_r_reg[7]/NET0131  & ~n72443 ;
  assign n72445 = ~\u0_desIn_r_reg[7]/NET0131  & n72443 ;
  assign n72446 = ~n72444 & ~n72445 ;
  assign n72448 = decrypt_pad & ~\u0_key_r_reg[36]/NET0131  ;
  assign n72449 = ~decrypt_pad & ~\u0_key_r_reg[43]/NET0131  ;
  assign n72450 = ~n72448 & ~n72449 ;
  assign n72451 = \u0_desIn_r_reg[33]/NET0131  & ~n72450 ;
  assign n72452 = ~\u0_desIn_r_reg[33]/NET0131  & n72450 ;
  assign n72453 = ~n72451 & ~n72452 ;
  assign n72456 = decrypt_pad & ~\u0_key_r_reg[37]/NET0131  ;
  assign n72457 = ~decrypt_pad & ~\u0_key_r_reg[44]/NET0131  ;
  assign n72458 = ~n72456 & ~n72457 ;
  assign n72459 = \u0_desIn_r_reg[41]/NET0131  & ~n72458 ;
  assign n72460 = ~\u0_desIn_r_reg[41]/NET0131  & n72458 ;
  assign n72461 = ~n72459 & ~n72460 ;
  assign n72472 = n72453 & n72461 ;
  assign n72473 = n72446 & n72472 ;
  assign n72465 = decrypt_pad & ~\u0_key_r_reg[49]/NET0131  ;
  assign n72466 = ~decrypt_pad & ~\u0_key_r_reg[1]/NET0131  ;
  assign n72467 = ~n72465 & ~n72466 ;
  assign n72468 = \u0_desIn_r_reg[49]/NET0131  & ~n72467 ;
  assign n72469 = ~\u0_desIn_r_reg[49]/NET0131  & n72467 ;
  assign n72470 = ~n72468 & ~n72469 ;
  assign n72474 = ~n72446 & n72453 ;
  assign n72475 = n72470 & ~n72474 ;
  assign n72476 = ~n72461 & ~n72475 ;
  assign n72477 = ~n72473 & ~n72476 ;
  assign n72478 = n72440 & ~n72477 ;
  assign n72447 = ~n72440 & n72446 ;
  assign n72454 = n72447 & ~n72453 ;
  assign n72455 = n72440 & ~n72453 ;
  assign n72462 = ~n72446 & n72461 ;
  assign n72463 = n72455 & n72462 ;
  assign n72464 = ~n72454 & ~n72463 ;
  assign n72471 = ~n72464 & n72470 ;
  assign n72429 = decrypt_pad & ~\u0_key_r_reg[0]/NET0131  ;
  assign n72430 = ~decrypt_pad & ~\u0_key_r_reg[7]/NET0131  ;
  assign n72431 = ~n72429 & ~n72430 ;
  assign n72432 = \u0_desIn_r_reg[57]/NET0131  & ~n72431 ;
  assign n72433 = ~\u0_desIn_r_reg[57]/NET0131  & n72431 ;
  assign n72434 = ~n72432 & ~n72433 ;
  assign n72479 = n72446 & ~n72453 ;
  assign n72482 = ~n72470 & ~n72479 ;
  assign n72480 = n72440 & ~n72446 ;
  assign n72481 = ~n72446 & ~n72461 ;
  assign n72483 = ~n72480 & ~n72481 ;
  assign n72484 = n72482 & n72483 ;
  assign n72485 = ~n72434 & ~n72484 ;
  assign n72486 = ~n72471 & n72485 ;
  assign n72487 = ~n72478 & n72486 ;
  assign n72490 = n72440 & ~n72461 ;
  assign n72492 = n72474 & n72490 ;
  assign n72491 = ~n72474 & ~n72490 ;
  assign n72493 = n72470 & ~n72491 ;
  assign n72494 = ~n72492 & n72493 ;
  assign n72495 = ~n72453 & ~n72461 ;
  assign n72496 = ~n72440 & n72495 ;
  assign n72497 = ~n72470 & n72496 ;
  assign n72488 = ~n72440 & n72472 ;
  assign n72489 = n72446 & n72488 ;
  assign n72498 = n72434 & ~n72489 ;
  assign n72499 = ~n72497 & n72498 ;
  assign n72500 = ~n72494 & n72499 ;
  assign n72501 = ~n72487 & ~n72500 ;
  assign n72502 = ~n72446 & n72496 ;
  assign n72507 = n72470 & ~n72502 ;
  assign n72503 = n72454 & n72461 ;
  assign n72504 = n72453 & ~n72461 ;
  assign n72505 = ~n72480 & ~n72504 ;
  assign n72506 = ~n72491 & n72505 ;
  assign n72508 = ~n72503 & ~n72506 ;
  assign n72509 = n72507 & n72508 ;
  assign n72510 = n72455 & n72461 ;
  assign n72511 = n72434 & n72510 ;
  assign n72512 = ~n72470 & ~n72492 ;
  assign n72513 = ~n72511 & n72512 ;
  assign n72514 = ~n72509 & ~n72513 ;
  assign n72515 = ~n72501 & ~n72514 ;
  assign n72516 = \u0_desIn_r_reg[38]/NET0131  & ~n72515 ;
  assign n72517 = ~\u0_desIn_r_reg[38]/NET0131  & n72515 ;
  assign n72518 = ~n72516 & ~n72517 ;
  assign n72519 = decrypt_pad & ~\u0_key_r_reg[10]/P0001  ;
  assign n72520 = ~decrypt_pad & ~\u0_key_r_reg[17]/NET0131  ;
  assign n72521 = ~n72519 & ~n72520 ;
  assign n72522 = \u0_desIn_r_reg[29]/NET0131  & ~n72521 ;
  assign n72523 = ~\u0_desIn_r_reg[29]/NET0131  & n72521 ;
  assign n72524 = ~n72522 & ~n72523 ;
  assign n72525 = decrypt_pad & ~\u0_key_r_reg[55]/NET0131  ;
  assign n72526 = ~decrypt_pad & ~\u0_key_r_reg[5]/NET0131  ;
  assign n72527 = ~n72525 & ~n72526 ;
  assign n72528 = \u0_desIn_r_reg[37]/NET0131  & ~n72527 ;
  assign n72529 = ~\u0_desIn_r_reg[37]/NET0131  & n72527 ;
  assign n72530 = ~n72528 & ~n72529 ;
  assign n72531 = decrypt_pad & ~\u0_key_r_reg[46]/NET0131  ;
  assign n72532 = ~decrypt_pad & ~\u0_key_r_reg[53]/NET0131  ;
  assign n72533 = ~n72531 & ~n72532 ;
  assign n72534 = \u0_desIn_r_reg[63]/NET0131  & ~n72533 ;
  assign n72535 = ~\u0_desIn_r_reg[63]/NET0131  & n72533 ;
  assign n72536 = ~n72534 & ~n72535 ;
  assign n72537 = n72530 & ~n72536 ;
  assign n72538 = decrypt_pad & ~\u0_key_r_reg[26]/NET0131  ;
  assign n72539 = ~decrypt_pad & ~\u0_key_r_reg[33]/NET0131  ;
  assign n72540 = ~n72538 & ~n72539 ;
  assign n72541 = \u0_desIn_r_reg[13]/NET0131  & ~n72540 ;
  assign n72542 = ~\u0_desIn_r_reg[13]/NET0131  & n72540 ;
  assign n72543 = ~n72541 & ~n72542 ;
  assign n72544 = n72537 & n72543 ;
  assign n72545 = decrypt_pad & ~\u0_key_r_reg[18]/NET0131  ;
  assign n72546 = ~decrypt_pad & ~\u0_key_r_reg[25]/NET0131  ;
  assign n72547 = ~n72545 & ~n72546 ;
  assign n72548 = \u0_desIn_r_reg[5]/NET0131  & ~n72547 ;
  assign n72549 = ~\u0_desIn_r_reg[5]/NET0131  & n72547 ;
  assign n72550 = ~n72548 & ~n72549 ;
  assign n72551 = n72544 & n72550 ;
  assign n72552 = decrypt_pad & ~\u0_key_r_reg[27]/NET0131  ;
  assign n72553 = ~decrypt_pad & ~\u0_key_r_reg[34]/NET0131  ;
  assign n72554 = ~n72552 & ~n72553 ;
  assign n72555 = \u0_desIn_r_reg[21]/NET0131  & ~n72554 ;
  assign n72556 = ~\u0_desIn_r_reg[21]/NET0131  & n72554 ;
  assign n72557 = ~n72555 & ~n72556 ;
  assign n72558 = n72551 & ~n72557 ;
  assign n72559 = n72543 & ~n72550 ;
  assign n72560 = ~n72530 & ~n72536 ;
  assign n72561 = n72530 & n72536 ;
  assign n72562 = ~n72560 & ~n72561 ;
  assign n72563 = n72559 & ~n72562 ;
  assign n72570 = ~n72530 & n72550 ;
  assign n72571 = n72543 & n72570 ;
  assign n72572 = n72536 & n72571 ;
  assign n72573 = ~n72563 & ~n72572 ;
  assign n72574 = ~n72558 & n72573 ;
  assign n72564 = n72530 & n72557 ;
  assign n72565 = n72562 & ~n72564 ;
  assign n72566 = ~n72543 & n72550 ;
  assign n72567 = ~n72565 & n72566 ;
  assign n72568 = ~n72543 & ~n72550 ;
  assign n72569 = n72565 & n72568 ;
  assign n72575 = ~n72567 & ~n72569 ;
  assign n72576 = n72574 & n72575 ;
  assign n72577 = ~n72524 & ~n72576 ;
  assign n72586 = n72530 & ~n72550 ;
  assign n72592 = ~n72530 & n72536 ;
  assign n72593 = n72550 & n72592 ;
  assign n72594 = ~n72544 & ~n72593 ;
  assign n72595 = ~n72586 & n72594 ;
  assign n72596 = n72524 & n72557 ;
  assign n72597 = ~n72595 & n72596 ;
  assign n72581 = ~n72543 & n72560 ;
  assign n72582 = ~n72550 & n72581 ;
  assign n72583 = n72530 & n72559 ;
  assign n72584 = ~n72582 & ~n72583 ;
  assign n72585 = n72557 & ~n72584 ;
  assign n72578 = n72543 & n72560 ;
  assign n72579 = n72524 & n72550 ;
  assign n72580 = n72578 & n72579 ;
  assign n72587 = ~n72536 & ~n72566 ;
  assign n72588 = n72524 & ~n72557 ;
  assign n72589 = ~n72570 & ~n72586 ;
  assign n72590 = n72588 & n72589 ;
  assign n72591 = ~n72587 & n72590 ;
  assign n72598 = ~n72580 & ~n72591 ;
  assign n72599 = ~n72585 & n72598 ;
  assign n72600 = ~n72597 & n72599 ;
  assign n72601 = ~n72577 & n72600 ;
  assign n72602 = ~\u0_desIn_r_reg[46]/NET0131  & ~n72601 ;
  assign n72603 = \u0_desIn_r_reg[46]/NET0131  & n72601 ;
  assign n72604 = ~n72602 & ~n72603 ;
  assign n72650 = decrypt_pad & ~\u0_key_r_reg[28]/NET0131  ;
  assign n72651 = ~decrypt_pad & ~\u0_key_r_reg[35]/P0001  ;
  assign n72652 = ~n72650 & ~n72651 ;
  assign n72653 = \u0_desIn_r_reg[59]/NET0131  & ~n72652 ;
  assign n72654 = ~\u0_desIn_r_reg[59]/NET0131  & n72652 ;
  assign n72655 = ~n72653 & ~n72654 ;
  assign n72633 = decrypt_pad & ~\u0_key_r_reg[2]/NET0131  ;
  assign n72634 = ~decrypt_pad & ~\u0_key_r_reg[9]/NET0131  ;
  assign n72635 = ~n72633 & ~n72634 ;
  assign n72636 = \u0_desIn_r_reg[51]/NET0131  & ~n72635 ;
  assign n72637 = ~\u0_desIn_r_reg[51]/NET0131  & n72635 ;
  assign n72638 = ~n72636 & ~n72637 ;
  assign n72618 = decrypt_pad & ~\u0_key_r_reg[22]/NET0131  ;
  assign n72619 = ~decrypt_pad & ~\u0_key_r_reg[29]/NET0131  ;
  assign n72620 = ~n72618 & ~n72619 ;
  assign n72621 = \u0_desIn_r_reg[35]/NET0131  & ~n72620 ;
  assign n72622 = ~\u0_desIn_r_reg[35]/NET0131  & n72620 ;
  assign n72623 = ~n72621 & ~n72622 ;
  assign n72605 = decrypt_pad & ~\u0_key_r_reg[7]/NET0131  ;
  assign n72606 = ~decrypt_pad & ~\u0_key_r_reg[14]/NET0131  ;
  assign n72607 = ~n72605 & ~n72606 ;
  assign n72608 = \u0_desIn_r_reg[27]/NET0131  & ~n72607 ;
  assign n72609 = ~\u0_desIn_r_reg[27]/NET0131  & n72607 ;
  assign n72610 = ~n72608 & ~n72609 ;
  assign n72625 = decrypt_pad & ~\u0_key_r_reg[23]/NET0131  ;
  assign n72626 = ~decrypt_pad & ~\u0_key_r_reg[30]/NET0131  ;
  assign n72627 = ~n72625 & ~n72626 ;
  assign n72628 = \u0_desIn_r_reg[1]/NET0131  & ~n72627 ;
  assign n72629 = ~\u0_desIn_r_reg[1]/NET0131  & n72627 ;
  assign n72630 = ~n72628 & ~n72629 ;
  assign n72657 = n72610 & ~n72630 ;
  assign n72658 = n72623 & n72657 ;
  assign n72611 = decrypt_pad & ~\u0_key_r_reg[44]/NET0131  ;
  assign n72612 = ~decrypt_pad & ~\u0_key_r_reg[51]/NET0131  ;
  assign n72613 = ~n72611 & ~n72612 ;
  assign n72614 = \u0_desIn_r_reg[43]/NET0131  & ~n72613 ;
  assign n72615 = ~\u0_desIn_r_reg[43]/NET0131  & n72613 ;
  assign n72616 = ~n72614 & ~n72615 ;
  assign n72617 = ~n72610 & ~n72616 ;
  assign n72674 = n72610 & ~n72623 ;
  assign n72675 = n72616 & n72674 ;
  assign n72676 = ~n72617 & ~n72675 ;
  assign n72677 = n72630 & ~n72676 ;
  assign n72678 = ~n72658 & ~n72677 ;
  assign n72679 = n72638 & ~n72678 ;
  assign n72680 = ~n72610 & ~n72623 ;
  assign n72681 = n72616 & n72630 ;
  assign n72682 = n72680 & n72681 ;
  assign n72644 = ~n72610 & ~n72630 ;
  assign n72683 = n72623 & n72644 ;
  assign n72684 = ~n72682 & ~n72683 ;
  assign n72685 = ~n72638 & ~n72684 ;
  assign n72640 = n72610 & n72630 ;
  assign n72672 = ~n72616 & ~n72638 ;
  assign n72673 = n72640 & n72672 ;
  assign n72667 = ~n72623 & n72657 ;
  assign n72686 = ~n72616 & n72667 ;
  assign n72687 = ~n72673 & ~n72686 ;
  assign n72688 = ~n72685 & n72687 ;
  assign n72689 = ~n72679 & n72688 ;
  assign n72690 = ~n72655 & ~n72689 ;
  assign n72624 = ~n72616 & n72623 ;
  assign n72631 = n72624 & ~n72630 ;
  assign n72632 = ~n72617 & ~n72631 ;
  assign n72639 = ~n72632 & ~n72638 ;
  assign n72641 = ~n72616 & n72638 ;
  assign n72642 = n72640 & n72641 ;
  assign n72645 = ~n72616 & ~n72644 ;
  assign n72643 = n72616 & ~n72630 ;
  assign n72646 = n72623 & ~n72643 ;
  assign n72647 = ~n72645 & n72646 ;
  assign n72648 = ~n72642 & ~n72647 ;
  assign n72649 = ~n72639 & n72648 ;
  assign n72656 = ~n72649 & n72655 ;
  assign n72659 = ~n72610 & n72623 ;
  assign n72660 = n72630 & n72659 ;
  assign n72661 = ~n72623 & n72644 ;
  assign n72662 = ~n72660 & ~n72661 ;
  assign n72663 = ~n72658 & n72662 ;
  assign n72664 = n72616 & n72638 ;
  assign n72665 = ~n72663 & n72664 ;
  assign n72666 = n72623 & n72640 ;
  assign n72668 = ~n72666 & ~n72667 ;
  assign n72669 = n72616 & n72668 ;
  assign n72670 = ~n72638 & ~n72645 ;
  assign n72671 = ~n72669 & n72670 ;
  assign n72691 = ~n72665 & ~n72671 ;
  assign n72692 = ~n72656 & n72691 ;
  assign n72693 = ~n72690 & n72692 ;
  assign n72694 = ~\u0_desIn_r_reg[30]/NET0131  & ~n72693 ;
  assign n72695 = \u0_desIn_r_reg[30]/NET0131  & n72693 ;
  assign n72696 = ~n72694 & ~n72695 ;
  assign n72697 = decrypt_pad & ~\u0_key_r_reg[1]/NET0131  ;
  assign n72698 = ~decrypt_pad & ~\u0_key_r_reg[8]/NET0131  ;
  assign n72699 = ~n72697 & ~n72698 ;
  assign n72700 = \u0_desIn_r_reg[19]/NET0131  & ~n72699 ;
  assign n72701 = ~\u0_desIn_r_reg[19]/NET0131  & n72699 ;
  assign n72702 = ~n72700 & ~n72701 ;
  assign n72723 = decrypt_pad & ~\u0_key_r_reg[29]/NET0131  ;
  assign n72724 = ~decrypt_pad & ~\u0_key_r_reg[36]/NET0131  ;
  assign n72725 = ~n72723 & ~n72724 ;
  assign n72726 = \u0_desIn_r_reg[61]/NET0131  & ~n72725 ;
  assign n72727 = ~\u0_desIn_r_reg[61]/NET0131  & n72725 ;
  assign n72728 = ~n72726 & ~n72727 ;
  assign n72703 = decrypt_pad & ~\u0_key_r_reg[45]/NET0131  ;
  assign n72704 = ~decrypt_pad & ~\u0_key_r_reg[52]/NET0131  ;
  assign n72705 = ~n72703 & ~n72704 ;
  assign n72706 = \u0_desIn_r_reg[35]/NET0131  & ~n72705 ;
  assign n72707 = ~\u0_desIn_r_reg[35]/NET0131  & n72705 ;
  assign n72708 = ~n72706 & ~n72707 ;
  assign n72709 = decrypt_pad & ~\u0_key_r_reg[51]/NET0131  ;
  assign n72710 = ~decrypt_pad & ~\u0_key_r_reg[31]/NET0131  ;
  assign n72711 = ~n72709 & ~n72710 ;
  assign n72712 = \u0_desIn_r_reg[3]/NET0131  & ~n72711 ;
  assign n72713 = ~\u0_desIn_r_reg[3]/NET0131  & n72711 ;
  assign n72714 = ~n72712 & ~n72713 ;
  assign n72716 = decrypt_pad & ~\u0_key_r_reg[14]/NET0131  ;
  assign n72717 = ~decrypt_pad & ~\u0_key_r_reg[21]/NET0131  ;
  assign n72718 = ~n72716 & ~n72717 ;
  assign n72719 = \u0_desIn_r_reg[11]/NET0131  & ~n72718 ;
  assign n72720 = ~\u0_desIn_r_reg[11]/NET0131  & n72718 ;
  assign n72721 = ~n72719 & ~n72720 ;
  assign n72734 = n72714 & ~n72721 ;
  assign n72735 = n72708 & n72734 ;
  assign n72736 = n72728 & n72735 ;
  assign n72731 = ~n72708 & n72728 ;
  assign n72732 = ~n72714 & ~n72721 ;
  assign n72733 = n72731 & n72732 ;
  assign n72715 = ~n72708 & n72714 ;
  assign n72722 = n72715 & n72721 ;
  assign n72729 = ~n72714 & ~n72728 ;
  assign n72730 = n72708 & n72729 ;
  assign n72737 = ~n72722 & ~n72730 ;
  assign n72738 = ~n72733 & n72737 ;
  assign n72739 = ~n72736 & n72738 ;
  assign n72740 = ~n72702 & ~n72739 ;
  assign n72748 = n72708 & n72721 ;
  assign n72749 = n72728 & n72748 ;
  assign n72744 = ~n72728 & n72734 ;
  assign n72746 = ~n72708 & ~n72728 ;
  assign n72747 = ~n72714 & n72746 ;
  assign n72750 = ~n72744 & ~n72747 ;
  assign n72751 = ~n72749 & n72750 ;
  assign n72752 = n72702 & ~n72751 ;
  assign n72741 = n72708 & n72728 ;
  assign n72742 = ~n72714 & n72741 ;
  assign n72743 = n72721 & n72742 ;
  assign n72745 = ~n72708 & n72744 ;
  assign n72753 = ~n72743 & ~n72745 ;
  assign n72754 = ~n72752 & n72753 ;
  assign n72755 = ~n72740 & n72754 ;
  assign n72756 = decrypt_pad & ~\u0_key_r_reg[16]/NET0131  ;
  assign n72757 = ~decrypt_pad & ~\u0_key_r_reg[23]/NET0131  ;
  assign n72758 = ~n72756 & ~n72757 ;
  assign n72759 = \u0_desIn_r_reg[27]/NET0131  & ~n72758 ;
  assign n72760 = ~\u0_desIn_r_reg[27]/NET0131  & n72758 ;
  assign n72761 = ~n72759 & ~n72760 ;
  assign n72762 = ~n72755 & ~n72761 ;
  assign n72769 = n72715 & n72728 ;
  assign n72766 = ~n72721 & n72741 ;
  assign n72767 = n72708 & ~n72728 ;
  assign n72768 = ~n72734 & n72767 ;
  assign n72770 = ~n72766 & ~n72768 ;
  assign n72771 = ~n72769 & n72770 ;
  assign n72772 = n72702 & ~n72771 ;
  assign n72773 = ~n72702 & ~n72721 ;
  assign n72774 = n72714 & n72767 ;
  assign n72775 = ~n72747 & ~n72774 ;
  assign n72776 = n72773 & ~n72775 ;
  assign n72763 = ~n72714 & n72721 ;
  assign n72764 = ~n72734 & ~n72763 ;
  assign n72765 = n72731 & ~n72764 ;
  assign n72777 = n72702 & n72714 ;
  assign n72778 = n72741 & ~n72777 ;
  assign n72779 = n72764 & n72778 ;
  assign n72780 = ~n72765 & ~n72779 ;
  assign n72781 = ~n72776 & n72780 ;
  assign n72782 = ~n72772 & n72781 ;
  assign n72783 = n72761 & ~n72782 ;
  assign n72784 = ~n72721 & n72769 ;
  assign n72785 = n72746 & n72763 ;
  assign n72786 = ~n72784 & ~n72785 ;
  assign n72787 = n72702 & ~n72786 ;
  assign n72788 = n72729 & n72748 ;
  assign n72789 = n72721 & ~n72728 ;
  assign n72790 = n72715 & n72789 ;
  assign n72791 = ~n72788 & ~n72790 ;
  assign n72792 = ~n72702 & ~n72791 ;
  assign n72793 = ~n72787 & ~n72792 ;
  assign n72794 = ~n72783 & n72793 ;
  assign n72795 = ~n72762 & n72794 ;
  assign n72796 = ~\u0_desIn_r_reg[44]/NET0131  & ~n72795 ;
  assign n72797 = \u0_desIn_r_reg[44]/NET0131  & n72795 ;
  assign n72798 = ~n72796 & ~n72797 ;
  assign n72825 = n72616 & ~n72659 ;
  assign n72826 = ~n72640 & n72825 ;
  assign n72827 = ~n72616 & n72630 ;
  assign n72828 = n72659 & n72827 ;
  assign n72829 = ~n72826 & ~n72828 ;
  assign n72830 = ~n72638 & ~n72829 ;
  assign n72801 = n72616 & n72659 ;
  assign n72822 = ~n72666 & ~n72801 ;
  assign n72823 = ~n72686 & n72822 ;
  assign n72824 = n72638 & ~n72823 ;
  assign n72831 = ~n72623 & n72673 ;
  assign n72832 = ~n72824 & ~n72831 ;
  assign n72833 = ~n72830 & n72832 ;
  assign n72834 = n72655 & ~n72833 ;
  assign n72799 = n72638 & n72676 ;
  assign n72800 = n72610 & n72624 ;
  assign n72802 = ~n72638 & ~n72800 ;
  assign n72803 = ~n72801 & n72802 ;
  assign n72804 = ~n72799 & ~n72803 ;
  assign n72807 = n72657 & n72672 ;
  assign n72808 = n72630 & n72675 ;
  assign n72809 = ~n72807 & ~n72808 ;
  assign n72805 = n72630 & n72638 ;
  assign n72806 = n72680 & n72805 ;
  assign n72810 = n72624 & n72657 ;
  assign n72811 = ~n72806 & ~n72810 ;
  assign n72812 = n72809 & n72811 ;
  assign n72813 = ~n72804 & n72812 ;
  assign n72814 = ~n72655 & ~n72813 ;
  assign n72819 = ~n72616 & n72806 ;
  assign n72820 = n72623 & n72807 ;
  assign n72821 = ~n72819 & ~n72820 ;
  assign n72815 = ~n72624 & ~n72640 ;
  assign n72816 = n72638 & ~n72645 ;
  assign n72817 = ~n72815 & n72816 ;
  assign n72818 = n72661 & n72672 ;
  assign n72835 = ~n72817 & ~n72818 ;
  assign n72836 = n72821 & n72835 ;
  assign n72837 = ~n72814 & n72836 ;
  assign n72838 = ~n72834 & n72837 ;
  assign n72839 = \u0_desIn_r_reg[20]/NET0131  & ~n72838 ;
  assign n72840 = ~\u0_desIn_r_reg[20]/NET0131  & n72838 ;
  assign n72841 = ~n72839 & ~n72840 ;
  assign n72842 = n72353 & ~n72408 ;
  assign n72843 = ~n72405 & n72842 ;
  assign n72844 = ~n72368 & n72382 ;
  assign n72845 = n72415 & ~n72844 ;
  assign n72846 = ~n72843 & ~n72845 ;
  assign n72847 = n72367 & ~n72377 ;
  assign n72848 = n72346 & n72847 ;
  assign n72849 = ~n72846 & ~n72848 ;
  assign n72850 = n72390 & ~n72849 ;
  assign n72861 = ~n72360 & ~n72368 ;
  assign n72862 = n72340 & ~n72407 ;
  assign n72863 = ~n72861 & n72862 ;
  assign n72856 = n72353 & n72367 ;
  assign n72857 = n72347 & n72353 ;
  assign n72858 = ~n72380 & ~n72857 ;
  assign n72859 = ~n72856 & ~n72858 ;
  assign n72860 = n72370 & n72374 ;
  assign n72864 = ~n72406 & ~n72860 ;
  assign n72865 = ~n72859 & n72864 ;
  assign n72866 = ~n72863 & n72865 ;
  assign n72867 = ~n72390 & ~n72866 ;
  assign n72851 = n72383 & n72397 ;
  assign n72852 = n72376 & n72420 ;
  assign n72853 = ~n72353 & ~n72852 ;
  assign n72854 = ~n72848 & n72853 ;
  assign n72855 = ~n72418 & ~n72854 ;
  assign n72868 = ~n72851 & ~n72855 ;
  assign n72869 = ~n72867 & n72868 ;
  assign n72870 = ~n72850 & n72869 ;
  assign n72871 = ~\u0_desIn_r_reg[12]/NET0131  & ~n72870 ;
  assign n72872 = \u0_desIn_r_reg[12]/NET0131  & n72870 ;
  assign n72873 = ~n72871 & ~n72872 ;
  assign n72887 = ~n72763 & n72767 ;
  assign n72888 = ~n72742 & ~n72887 ;
  assign n72889 = ~n72702 & ~n72888 ;
  assign n72895 = ~n72744 & ~n72889 ;
  assign n72890 = n72714 & n72741 ;
  assign n72891 = ~n72733 & ~n72890 ;
  assign n72892 = n72702 & ~n72891 ;
  assign n72893 = n72721 & n72769 ;
  assign n72894 = ~n72785 & ~n72893 ;
  assign n72896 = ~n72892 & n72894 ;
  assign n72897 = n72895 & n72896 ;
  assign n72898 = ~n72761 & ~n72897 ;
  assign n72877 = ~n72721 & n72747 ;
  assign n72878 = ~n72742 & ~n72877 ;
  assign n72879 = n72702 & ~n72878 ;
  assign n72880 = n72728 & n72773 ;
  assign n72881 = n72791 & ~n72880 ;
  assign n72882 = ~n72879 & n72881 ;
  assign n72883 = n72761 & ~n72882 ;
  assign n72874 = n72728 & n72763 ;
  assign n72875 = ~n72702 & n72874 ;
  assign n72876 = ~n72708 & n72875 ;
  assign n72884 = ~n72764 & n72767 ;
  assign n72885 = ~n72722 & ~n72884 ;
  assign n72886 = n72702 & ~n72885 ;
  assign n72899 = ~n72876 & ~n72886 ;
  assign n72900 = ~n72883 & n72899 ;
  assign n72901 = ~n72898 & n72900 ;
  assign n72902 = ~\u0_desIn_r_reg[62]/NET0131  & ~n72901 ;
  assign n72903 = \u0_desIn_r_reg[62]/NET0131  & n72901 ;
  assign n72904 = ~n72902 & ~n72903 ;
  assign n72905 = ~n72369 & n72842 ;
  assign n72909 = ~n72346 & n72377 ;
  assign n72910 = ~n72371 & ~n72909 ;
  assign n72911 = ~n72367 & ~n72910 ;
  assign n72906 = n72346 & ~n72397 ;
  assign n72907 = ~n72359 & ~n72390 ;
  assign n72908 = ~n72906 & n72907 ;
  assign n72912 = ~n72353 & ~n72908 ;
  assign n72913 = ~n72911 & n72912 ;
  assign n72914 = ~n72905 & ~n72913 ;
  assign n72915 = ~n72347 & n72367 ;
  assign n72916 = n72383 & n72915 ;
  assign n72917 = ~n72359 & n72416 ;
  assign n72918 = ~n72369 & ~n72384 ;
  assign n72919 = ~n72917 & n72918 ;
  assign n72920 = ~n72916 & n72919 ;
  assign n72921 = ~n72390 & ~n72920 ;
  assign n72922 = ~n72370 & ~n72407 ;
  assign n72923 = ~n72353 & ~n72922 ;
  assign n72924 = ~n72340 & n72353 ;
  assign n72925 = ~n72359 & ~n72924 ;
  assign n72926 = ~n72906 & ~n72925 ;
  assign n72927 = ~n72406 & n72926 ;
  assign n72928 = ~n72923 & ~n72927 ;
  assign n72929 = n72390 & ~n72416 ;
  assign n72930 = ~n72928 & n72929 ;
  assign n72931 = ~n72921 & ~n72930 ;
  assign n72932 = ~n72914 & n72931 ;
  assign n72933 = ~\u0_desIn_r_reg[8]/NET0131  & ~n72932 ;
  assign n72934 = \u0_desIn_r_reg[8]/NET0131  & n72932 ;
  assign n72935 = ~n72933 & ~n72934 ;
  assign n72936 = decrypt_pad & ~\u0_key_r_reg[41]/NET0131  ;
  assign n72937 = ~decrypt_pad & ~\u0_key_r_reg[48]/NET0131  ;
  assign n72938 = ~n72936 & ~n72937 ;
  assign n72939 = \u0_desIn_r_reg[55]/NET0131  & ~n72938 ;
  assign n72940 = ~\u0_desIn_r_reg[55]/NET0131  & n72938 ;
  assign n72941 = ~n72939 & ~n72940 ;
  assign n72948 = decrypt_pad & ~\u0_key_r_reg[24]/NET0131  ;
  assign n72949 = ~decrypt_pad & ~\u0_key_r_reg[6]/NET0131  ;
  assign n72950 = ~n72948 & ~n72949 ;
  assign n72951 = \u0_desIn_r_reg[39]/NET0131  & ~n72950 ;
  assign n72952 = ~\u0_desIn_r_reg[39]/NET0131  & n72950 ;
  assign n72953 = ~n72951 & ~n72952 ;
  assign n72973 = ~n72941 & ~n72953 ;
  assign n72942 = decrypt_pad & ~\u0_key_r_reg[12]/NET0131  ;
  assign n72943 = ~decrypt_pad & ~\u0_key_r_reg[19]/NET0131  ;
  assign n72944 = ~n72942 & ~n72943 ;
  assign n72945 = \u0_desIn_r_reg[5]/NET0131  & ~n72944 ;
  assign n72946 = ~\u0_desIn_r_reg[5]/NET0131  & n72944 ;
  assign n72947 = ~n72945 & ~n72946 ;
  assign n72961 = decrypt_pad & ~\u0_key_r_reg[47]/NET0131  ;
  assign n72962 = ~decrypt_pad & ~\u0_key_r_reg[54]/NET0131  ;
  assign n72963 = ~n72961 & ~n72962 ;
  assign n72964 = \u0_desIn_r_reg[47]/NET0131  & ~n72963 ;
  assign n72965 = ~\u0_desIn_r_reg[47]/NET0131  & n72963 ;
  assign n72966 = ~n72964 & ~n72965 ;
  assign n72974 = n72947 & ~n72966 ;
  assign n72975 = n72973 & n72974 ;
  assign n72955 = decrypt_pad & ~\u0_key_r_reg[20]/NET0131  ;
  assign n72956 = ~decrypt_pad & ~\u0_key_r_reg[27]/NET0131  ;
  assign n72957 = ~n72955 & ~n72956 ;
  assign n72958 = \u0_desIn_r_reg[31]/NET0131  & ~n72957 ;
  assign n72959 = ~\u0_desIn_r_reg[31]/NET0131  & n72957 ;
  assign n72960 = ~n72958 & ~n72959 ;
  assign n72976 = n72947 & ~n72960 ;
  assign n72977 = n72953 & n72976 ;
  assign n72978 = n72966 & n72977 ;
  assign n72979 = ~n72975 & ~n72978 ;
  assign n72980 = decrypt_pad & ~\u0_key_r_reg[32]/NET0131  ;
  assign n72981 = ~decrypt_pad & ~\u0_key_r_reg[39]/P0001  ;
  assign n72982 = ~n72980 & ~n72981 ;
  assign n72983 = \u0_desIn_r_reg[63]/NET0131  & ~n72982 ;
  assign n72984 = ~\u0_desIn_r_reg[63]/NET0131  & n72982 ;
  assign n72985 = ~n72983 & ~n72984 ;
  assign n72986 = n72947 & ~n72953 ;
  assign n72987 = n72960 & n72966 ;
  assign n72988 = n72941 & n72987 ;
  assign n72989 = n72986 & n72988 ;
  assign n72998 = ~n72985 & ~n72989 ;
  assign n72999 = n72979 & n72998 ;
  assign n72990 = ~n72947 & n72953 ;
  assign n72991 = ~n72960 & n72986 ;
  assign n72992 = ~n72990 & ~n72991 ;
  assign n72993 = ~n72966 & ~n72992 ;
  assign n72994 = n72960 & n72986 ;
  assign n72995 = ~n72941 & ~n72994 ;
  assign n72996 = ~n72986 & ~n72987 ;
  assign n72997 = n72995 & ~n72996 ;
  assign n73000 = ~n72993 & ~n72997 ;
  assign n73001 = n72999 & n73000 ;
  assign n73008 = ~n72941 & n72966 ;
  assign n73002 = ~n72947 & ~n72960 ;
  assign n73009 = ~n72994 & ~n73002 ;
  assign n73010 = n73008 & ~n73009 ;
  assign n72967 = ~n72960 & n72966 ;
  assign n73011 = n72941 & n72953 ;
  assign n73012 = ~n72967 & n73011 ;
  assign n73003 = n72973 & n73002 ;
  assign n73013 = n72985 & ~n73003 ;
  assign n73014 = ~n73012 & n73013 ;
  assign n73004 = n72960 & ~n72966 ;
  assign n73005 = ~n72947 & n73004 ;
  assign n73006 = ~n72953 & n73005 ;
  assign n72969 = n72953 & n72960 ;
  assign n72970 = ~n72966 & n72969 ;
  assign n73007 = n72947 & n72970 ;
  assign n73015 = ~n73006 & ~n73007 ;
  assign n73016 = n73014 & n73015 ;
  assign n73017 = ~n73010 & n73016 ;
  assign n73018 = ~n73001 & ~n73017 ;
  assign n72954 = ~n72947 & ~n72953 ;
  assign n72968 = n72954 & n72967 ;
  assign n72971 = ~n72968 & ~n72970 ;
  assign n72972 = n72941 & ~n72971 ;
  assign n73020 = ~n72973 & ~n73008 ;
  assign n73019 = ~n72953 & n72966 ;
  assign n73021 = n72976 & ~n73019 ;
  assign n73022 = ~n73020 & n73021 ;
  assign n73023 = ~n72972 & ~n73022 ;
  assign n73024 = ~n73018 & n73023 ;
  assign n73025 = \u0_desIn_r_reg[14]/NET0131  & n73024 ;
  assign n73026 = ~\u0_desIn_r_reg[14]/NET0131  & ~n73024 ;
  assign n73027 = ~n73025 & ~n73026 ;
  assign n73028 = ~n72966 & n73002 ;
  assign n73029 = ~n72977 & ~n73028 ;
  assign n73048 = n72941 & n73029 ;
  assign n73049 = ~n72941 & ~n72969 ;
  assign n73050 = ~n72991 & n73049 ;
  assign n73051 = ~n73005 & n73050 ;
  assign n73052 = ~n73048 & ~n73051 ;
  assign n73053 = n72987 & n72990 ;
  assign n73054 = ~n73009 & n73019 ;
  assign n73055 = ~n73053 & ~n73054 ;
  assign n73056 = ~n73052 & n73055 ;
  assign n73057 = ~n72985 & ~n73056 ;
  assign n73033 = n72960 & ~n72990 ;
  assign n73034 = ~n72986 & n73033 ;
  assign n73035 = ~n72960 & n72990 ;
  assign n73036 = n72966 & n73035 ;
  assign n73037 = ~n73034 & ~n73036 ;
  assign n73038 = n72941 & ~n73037 ;
  assign n73030 = ~n72941 & ~n73029 ;
  assign n73031 = ~n72941 & ~n72986 ;
  assign n73032 = n73004 & ~n73031 ;
  assign n73039 = n72967 & n72986 ;
  assign n73040 = ~n73032 & ~n73039 ;
  assign n73041 = ~n73030 & n73040 ;
  assign n73042 = ~n73038 & n73041 ;
  assign n73043 = n72985 & ~n73042 ;
  assign n73044 = ~n72960 & ~n73019 ;
  assign n73045 = ~n72941 & ~n73004 ;
  assign n73046 = ~n73033 & n73045 ;
  assign n73047 = ~n73044 & n73046 ;
  assign n73058 = ~n73043 & ~n73047 ;
  assign n73059 = ~n73057 & n73058 ;
  assign n73060 = ~\u0_desIn_r_reg[24]/NET0131  & ~n73059 ;
  assign n73061 = \u0_desIn_r_reg[24]/NET0131  & n73059 ;
  assign n73062 = ~n73060 & ~n73061 ;
  assign n73077 = ~n72732 & ~n72789 ;
  assign n73078 = ~n72708 & ~n73077 ;
  assign n73079 = ~n72729 & ~n72890 ;
  assign n73080 = ~n73078 & n73079 ;
  assign n73081 = n72702 & ~n73080 ;
  assign n73075 = ~n72742 & ~n72744 ;
  assign n73076 = ~n72702 & ~n73075 ;
  assign n73082 = ~n72735 & ~n72893 ;
  assign n73083 = ~n73076 & n73082 ;
  assign n73084 = ~n73081 & n73083 ;
  assign n73085 = n72761 & ~n73084 ;
  assign n73069 = n72702 & ~n72715 ;
  assign n73068 = ~n72702 & ~n72729 ;
  assign n73070 = ~n72721 & ~n73068 ;
  assign n73071 = ~n73069 & n73070 ;
  assign n73063 = n72721 & n72774 ;
  assign n73065 = ~n72714 & ~n72731 ;
  assign n73064 = n72714 & ~n72789 ;
  assign n73066 = ~n72702 & ~n73064 ;
  assign n73067 = ~n73065 & n73066 ;
  assign n73072 = ~n73063 & ~n73067 ;
  assign n73073 = ~n73071 & n73072 ;
  assign n73074 = ~n72761 & ~n73073 ;
  assign n73086 = n72732 & n72767 ;
  assign n73087 = n72894 & ~n73086 ;
  assign n73088 = n72702 & ~n73087 ;
  assign n73089 = ~n72736 & ~n72875 ;
  assign n73090 = ~n73088 & n73089 ;
  assign n73091 = ~n73074 & n73090 ;
  assign n73092 = ~n73085 & n73091 ;
  assign n73093 = ~\u0_desIn_r_reg[0]/NET0131  & ~n73092 ;
  assign n73094 = \u0_desIn_r_reg[0]/NET0131  & n73092 ;
  assign n73095 = ~n73093 & ~n73094 ;
  assign n73096 = ~n72186 & ~n72218 ;
  assign n73097 = n72168 & ~n73096 ;
  assign n73098 = n72174 & n72182 ;
  assign n73099 = ~n72155 & n73098 ;
  assign n73100 = ~n72220 & ~n73099 ;
  assign n73101 = ~n72161 & ~n73100 ;
  assign n73104 = n72149 & ~n73101 ;
  assign n73102 = ~n72168 & n72208 ;
  assign n73103 = ~n72174 & ~n72226 ;
  assign n73105 = ~n73102 & ~n73103 ;
  assign n73106 = n73104 & n73105 ;
  assign n73107 = ~n73097 & n73106 ;
  assign n73108 = n72161 & n73099 ;
  assign n73116 = ~n72149 & ~n73108 ;
  assign n73109 = n72168 & n72207 ;
  assign n73110 = n72183 & ~n72196 ;
  assign n73117 = ~n73109 & ~n73110 ;
  assign n73118 = n73116 & n73117 ;
  assign n73111 = ~n72189 & ~n72210 ;
  assign n73112 = ~n73098 & ~n73111 ;
  assign n73113 = ~n72183 & ~n72193 ;
  assign n73114 = ~n72219 & n73113 ;
  assign n73115 = ~n72168 & ~n73114 ;
  assign n73119 = ~n73112 & ~n73115 ;
  assign n73120 = n73118 & n73119 ;
  assign n73121 = ~n73107 & ~n73120 ;
  assign n73122 = \u0_desIn_r_reg[28]/NET0131  & n73121 ;
  assign n73123 = ~\u0_desIn_r_reg[28]/NET0131  & ~n73121 ;
  assign n73124 = ~n73122 & ~n73123 ;
  assign n73130 = n72616 & n72658 ;
  assign n73140 = ~n72643 & n72659 ;
  assign n73141 = ~n73130 & ~n73140 ;
  assign n73142 = n72638 & ~n73141 ;
  assign n73143 = n72616 & n72640 ;
  assign n73144 = ~n72624 & n72644 ;
  assign n73145 = ~n73143 & ~n73144 ;
  assign n73146 = ~n72638 & ~n73145 ;
  assign n73138 = ~n72643 & ~n72827 ;
  assign n73139 = n72680 & ~n73138 ;
  assign n73147 = n72809 & ~n73139 ;
  assign n73148 = ~n73146 & n73147 ;
  assign n73149 = ~n73142 & n73148 ;
  assign n73150 = n72655 & ~n73149 ;
  assign n73131 = ~n72616 & ~n72657 ;
  assign n73132 = ~n72680 & n73131 ;
  assign n73133 = ~n73130 & ~n73132 ;
  assign n73134 = ~n72638 & ~n73133 ;
  assign n73126 = ~n72624 & ~n72630 ;
  assign n73127 = ~n72825 & n73126 ;
  assign n73128 = n72668 & ~n73127 ;
  assign n73129 = n72638 & ~n73128 ;
  assign n73135 = ~n72682 & ~n73129 ;
  assign n73136 = ~n73134 & n73135 ;
  assign n73137 = ~n72655 & ~n73136 ;
  assign n73125 = n72624 & n72805 ;
  assign n73151 = ~n72686 & ~n73125 ;
  assign n73152 = ~n73137 & n73151 ;
  assign n73153 = ~n73150 & n73152 ;
  assign n73154 = \u0_desIn_r_reg[32]/NET0131  & ~n73153 ;
  assign n73155 = ~\u0_desIn_r_reg[32]/NET0131  & n73153 ;
  assign n73156 = ~n73154 & ~n73155 ;
  assign n73172 = ~n72401 & ~n72420 ;
  assign n73173 = n72340 & ~n73172 ;
  assign n73174 = ~n72353 & ~n73173 ;
  assign n73175 = ~n72359 & n72400 ;
  assign n73176 = n72353 & ~n72421 ;
  assign n73177 = ~n73175 & n73176 ;
  assign n73178 = ~n73174 & ~n73177 ;
  assign n73179 = n72373 & ~n72417 ;
  assign n73180 = ~n73178 & n73179 ;
  assign n73181 = ~n72390 & ~n73180 ;
  assign n73157 = n72346 & ~n72377 ;
  assign n73158 = ~n72405 & ~n73157 ;
  assign n73159 = n72367 & ~n73158 ;
  assign n73160 = ~n72401 & ~n72917 ;
  assign n73161 = n72390 & ~n73160 ;
  assign n73162 = ~n73159 & ~n73161 ;
  assign n73163 = n72353 & ~n73162 ;
  assign n73164 = ~n72370 & n72847 ;
  assign n73165 = ~n72353 & n72359 ;
  assign n73166 = ~n72382 & n73165 ;
  assign n73167 = ~n72915 & n73166 ;
  assign n73168 = ~n73164 & ~n73167 ;
  assign n73169 = n72390 & ~n73168 ;
  assign n73170 = ~n72346 & ~n72353 ;
  assign n73171 = n72847 & n73170 ;
  assign n73182 = ~n73169 & ~n73171 ;
  assign n73183 = ~n73163 & n73182 ;
  assign n73184 = ~n73181 & n73183 ;
  assign n73185 = ~\u0_desIn_r_reg[6]/NET0131  & ~n73184 ;
  assign n73186 = \u0_desIn_r_reg[6]/NET0131  & n73184 ;
  assign n73187 = ~n73185 & ~n73186 ;
  assign n73190 = ~n72264 & ~n72309 ;
  assign n73191 = ~n72251 & n72264 ;
  assign n73194 = n72280 & n73191 ;
  assign n73195 = ~n73190 & ~n73194 ;
  assign n73196 = n72245 & ~n73195 ;
  assign n73188 = n72264 & n72295 ;
  assign n73189 = n72292 & ~n73188 ;
  assign n73192 = ~n72245 & ~n73191 ;
  assign n73193 = ~n73190 & n73192 ;
  assign n73197 = n72251 & n72323 ;
  assign n73198 = ~n73193 & ~n73197 ;
  assign n73199 = n73189 & n73198 ;
  assign n73200 = ~n73196 & n73199 ;
  assign n73203 = ~n72251 & n72305 ;
  assign n73204 = ~n72301 & ~n73203 ;
  assign n73205 = n72258 & ~n73204 ;
  assign n73201 = ~n72280 & ~n72316 ;
  assign n73202 = n72264 & n73201 ;
  assign n73206 = n72245 & ~n73202 ;
  assign n73207 = ~n73205 & n73206 ;
  assign n73208 = ~n72277 & ~n72300 ;
  assign n73209 = ~n72258 & ~n73208 ;
  assign n73210 = ~n72272 & n72282 ;
  assign n73211 = ~n72245 & ~n73210 ;
  assign n73212 = ~n73209 & n73211 ;
  assign n73213 = ~n73207 & ~n73212 ;
  assign n73214 = ~n72281 & ~n72292 ;
  assign n73215 = ~n72317 & n73214 ;
  assign n73216 = ~n73213 & n73215 ;
  assign n73217 = ~n73200 & ~n73216 ;
  assign n73218 = \u0_desIn_r_reg[2]/NET0131  & ~n73217 ;
  assign n73219 = ~\u0_desIn_r_reg[2]/NET0131  & n73217 ;
  assign n73220 = ~n73218 & ~n73219 ;
  assign n73221 = n72988 & ~n72990 ;
  assign n73222 = ~n72966 & ~n72973 ;
  assign n73223 = n72976 & n73222 ;
  assign n73224 = ~n73221 & ~n73223 ;
  assign n73225 = ~n72941 & ~n72985 ;
  assign n73226 = ~n73035 & n73225 ;
  assign n73227 = ~n73039 & n73226 ;
  assign n73228 = ~n73006 & n73227 ;
  assign n73229 = n73224 & n73228 ;
  assign n73230 = n72954 & n72966 ;
  assign n73231 = n72995 & ~n73230 ;
  assign n73233 = n72966 & n72976 ;
  assign n73232 = n72954 & ~n72966 ;
  assign n73234 = n72941 & ~n73232 ;
  assign n73235 = ~n73233 & n73234 ;
  assign n73236 = ~n73231 & ~n73235 ;
  assign n73237 = n72953 & n73028 ;
  assign n73238 = n72985 & ~n73237 ;
  assign n73239 = n72979 & n73238 ;
  assign n73240 = ~n73236 & n73239 ;
  assign n73241 = ~n73229 & ~n73240 ;
  assign n73242 = ~n73007 & ~n73053 ;
  assign n73243 = ~n73241 & n73242 ;
  assign n73244 = ~n72953 & ~n73009 ;
  assign n73245 = n72953 & n73005 ;
  assign n73246 = n72941 & ~n72985 ;
  assign n73247 = ~n73245 & n73246 ;
  assign n73248 = n73224 & n73247 ;
  assign n73249 = ~n73244 & n73248 ;
  assign n73250 = ~n73243 & ~n73249 ;
  assign n73251 = ~\u0_desIn_r_reg[36]/NET0131  & ~n73250 ;
  assign n73252 = \u0_desIn_r_reg[36]/NET0131  & n73250 ;
  assign n73253 = ~n73251 & ~n73252 ;
  assign n73258 = ~n72638 & ~n72662 ;
  assign n73255 = n72610 & ~n72624 ;
  assign n73256 = ~n72683 & ~n73255 ;
  assign n73257 = n72638 & ~n73256 ;
  assign n73254 = n72623 & n73143 ;
  assign n73259 = ~n72655 & ~n73254 ;
  assign n73260 = ~n73257 & n73259 ;
  assign n73261 = ~n73258 & n73260 ;
  assign n73265 = ~n72631 & n72655 ;
  assign n73262 = ~n72638 & n72674 ;
  assign n73266 = ~n72806 & ~n73262 ;
  assign n73267 = n73265 & n73266 ;
  assign n73264 = n72638 & n72800 ;
  assign n73263 = n72630 & n72801 ;
  assign n73268 = ~n73139 & ~n73263 ;
  assign n73269 = ~n73264 & n73268 ;
  assign n73270 = n73267 & n73269 ;
  assign n73271 = ~n73261 & ~n73270 ;
  assign n73272 = n72821 & ~n72831 ;
  assign n73273 = ~n73271 & n73272 ;
  assign n73274 = \u0_desIn_r_reg[18]/NET0131  & n73273 ;
  assign n73275 = ~\u0_desIn_r_reg[18]/NET0131  & ~n73273 ;
  assign n73276 = ~n73274 & ~n73275 ;
  assign n73292 = n72258 & n72264 ;
  assign n73293 = ~n72278 & ~n73292 ;
  assign n73294 = ~n72245 & ~n73293 ;
  assign n73296 = n72272 & n72275 ;
  assign n73295 = n72245 & n72320 ;
  assign n73297 = ~n72310 & ~n73197 ;
  assign n73298 = ~n73295 & n73297 ;
  assign n73299 = ~n73296 & n73298 ;
  assign n73300 = ~n73294 & n73299 ;
  assign n73301 = ~n72292 & ~n73300 ;
  assign n73278 = ~n72264 & ~n73201 ;
  assign n73279 = ~n72285 & ~n73278 ;
  assign n73280 = n72292 & ~n73279 ;
  assign n73277 = ~n72258 & n73203 ;
  assign n73281 = ~n72279 & ~n73188 ;
  assign n73282 = ~n73277 & n73281 ;
  assign n73283 = ~n73280 & n73282 ;
  assign n73284 = ~n72245 & ~n73283 ;
  assign n73285 = ~n72265 & ~n72320 ;
  assign n73286 = n72252 & ~n73285 ;
  assign n73287 = n72245 & ~n72306 ;
  assign n73288 = n73201 & n73287 ;
  assign n73289 = ~n72318 & ~n73194 ;
  assign n73290 = ~n73288 & n73289 ;
  assign n73291 = n72292 & ~n73290 ;
  assign n73302 = ~n73286 & ~n73291 ;
  assign n73303 = ~n73284 & n73302 ;
  assign n73304 = ~n73301 & n73303 ;
  assign n73305 = \u0_desIn_r_reg[50]/NET0131  & ~n73304 ;
  assign n73306 = ~\u0_desIn_r_reg[50]/NET0131  & n73304 ;
  assign n73307 = ~n73305 & ~n73306 ;
  assign n73336 = n72446 & n72510 ;
  assign n73337 = ~n72461 & n72480 ;
  assign n73338 = ~n73336 & ~n73337 ;
  assign n73339 = ~n72470 & ~n73338 ;
  assign n73311 = ~n72440 & ~n72446 ;
  assign n73328 = n72453 & ~n73311 ;
  assign n73329 = ~n72490 & n73328 ;
  assign n73330 = n72446 & n72495 ;
  assign n73331 = ~n73329 & ~n73330 ;
  assign n73332 = n72470 & ~n73331 ;
  assign n73308 = n72440 & n72474 ;
  assign n73333 = ~n72453 & n73311 ;
  assign n73334 = ~n73308 & ~n73333 ;
  assign n73335 = n72461 & ~n73334 ;
  assign n73340 = n72454 & ~n72461 ;
  assign n73341 = ~n73335 & ~n73340 ;
  assign n73342 = ~n73332 & n73341 ;
  assign n73343 = ~n73339 & n73342 ;
  assign n73344 = n72434 & ~n73343 ;
  assign n73309 = ~n72510 & ~n73308 ;
  assign n73310 = n72470 & ~n73309 ;
  assign n73319 = ~n72463 & ~n72488 ;
  assign n73312 = n72453 & ~n72470 ;
  assign n73313 = n73311 & n73312 ;
  assign n73317 = n72461 & ~n72470 ;
  assign n73318 = n72447 & n73317 ;
  assign n73320 = ~n73313 & ~n73318 ;
  assign n73321 = n73319 & n73320 ;
  assign n73314 = ~n72453 & n72470 ;
  assign n73315 = n72446 & n72490 ;
  assign n73316 = ~n73314 & n73315 ;
  assign n73322 = ~n72502 & ~n73316 ;
  assign n73323 = n73321 & n73322 ;
  assign n73324 = ~n73310 & n73323 ;
  assign n73325 = ~n72434 & ~n73324 ;
  assign n73326 = n72470 & n72496 ;
  assign n73327 = n73312 & n73315 ;
  assign n73345 = ~n73326 & ~n73327 ;
  assign n73346 = ~n73325 & n73345 ;
  assign n73347 = ~n73344 & n73346 ;
  assign n73348 = ~\u0_desIn_r_reg[34]/NET0131  & ~n73347 ;
  assign n73349 = \u0_desIn_r_reg[34]/NET0131  & n73347 ;
  assign n73350 = ~n73348 & ~n73349 ;
  assign n73354 = n72550 & n72561 ;
  assign n73355 = ~n72550 & ~n72561 ;
  assign n73356 = ~n73354 & ~n73355 ;
  assign n73357 = ~n72560 & ~n73356 ;
  assign n73358 = n72550 & n72560 ;
  assign n73359 = n72557 & n73358 ;
  assign n73360 = ~n73357 & ~n73359 ;
  assign n73361 = ~n72543 & ~n73360 ;
  assign n73362 = ~n72543 & n72592 ;
  assign n73363 = ~n72578 & ~n73362 ;
  assign n73364 = ~n72557 & ~n73363 ;
  assign n73365 = ~n72551 & ~n73364 ;
  assign n73366 = ~n73361 & n73365 ;
  assign n73367 = n72524 & ~n73366 ;
  assign n73371 = ~n72536 & ~n72550 ;
  assign n73372 = n72530 & n73371 ;
  assign n73373 = ~n72581 & ~n73354 ;
  assign n73374 = ~n73372 & n73373 ;
  assign n73375 = ~n72557 & ~n73374 ;
  assign n73376 = n72557 & ~n72560 ;
  assign n73377 = n73356 & n73376 ;
  assign n73378 = ~n72582 & ~n73377 ;
  assign n73379 = ~n73375 & n73378 ;
  assign n73380 = ~n72524 & ~n73379 ;
  assign n73351 = n72536 & ~n72550 ;
  assign n73352 = n72543 & ~n72557 ;
  assign n73353 = n73351 & n73352 ;
  assign n73368 = ~n72550 & n72578 ;
  assign n73369 = ~n72572 & ~n73368 ;
  assign n73370 = n72557 & ~n73369 ;
  assign n73381 = ~n73353 & ~n73370 ;
  assign n73382 = ~n73380 & n73381 ;
  assign n73383 = ~n73367 & n73382 ;
  assign n73384 = ~\u0_desIn_r_reg[60]/NET0131  & ~n73383 ;
  assign n73385 = \u0_desIn_r_reg[60]/NET0131  & n73383 ;
  assign n73386 = ~n73384 & ~n73385 ;
  assign n73392 = ~n72496 & ~n73328 ;
  assign n73391 = n72440 & n72446 ;
  assign n73393 = ~n72470 & ~n73391 ;
  assign n73394 = ~n73392 & n73393 ;
  assign n73387 = ~n72440 & ~n72481 ;
  assign n73388 = n72453 & ~n73387 ;
  assign n73389 = n72470 & ~n72480 ;
  assign n73390 = n73388 & n73389 ;
  assign n73395 = ~n72463 & ~n73330 ;
  assign n73396 = ~n72489 & n73395 ;
  assign n73397 = ~n73390 & n73396 ;
  assign n73398 = ~n73394 & n73397 ;
  assign n73399 = n72434 & ~n73398 ;
  assign n73406 = n72470 & ~n72488 ;
  assign n73404 = ~n72446 & n72504 ;
  assign n73405 = n72446 & ~n72504 ;
  assign n73407 = ~n73404 & ~n73405 ;
  assign n73408 = n73406 & n73407 ;
  assign n73403 = n73317 & n73391 ;
  assign n73409 = ~n73313 & ~n73403 ;
  assign n73410 = ~n72503 & n73409 ;
  assign n73411 = ~n73408 & n73410 ;
  assign n73412 = ~n72434 & ~n73411 ;
  assign n73400 = ~n72492 & ~n72506 ;
  assign n73401 = ~n72470 & ~n73400 ;
  assign n73402 = n72462 & n73314 ;
  assign n73413 = ~n73401 & ~n73402 ;
  assign n73414 = ~n73412 & n73413 ;
  assign n73415 = ~n73399 & n73414 ;
  assign n73416 = ~\u0_desIn_r_reg[16]/NET0131  & ~n73415 ;
  assign n73417 = \u0_desIn_r_reg[16]/NET0131  & n73415 ;
  assign n73418 = ~n73416 & ~n73417 ;
  assign n73443 = n72174 & n72224 ;
  assign n73422 = ~n72188 & ~n72209 ;
  assign n73442 = n72198 & n73422 ;
  assign n73444 = ~n72210 & ~n73442 ;
  assign n73445 = ~n73443 & n73444 ;
  assign n73446 = ~n72168 & ~n73445 ;
  assign n73436 = ~n72161 & n72219 ;
  assign n73437 = n72182 & n73436 ;
  assign n73438 = ~n72174 & n72193 ;
  assign n73439 = ~n72184 & ~n73436 ;
  assign n73440 = ~n73438 & n73439 ;
  assign n73441 = n72168 & ~n73440 ;
  assign n73447 = ~n73437 & ~n73441 ;
  assign n73448 = ~n73446 & n73447 ;
  assign n73449 = n72149 & ~n73448 ;
  assign n73423 = ~n72196 & n73422 ;
  assign n73424 = n73113 & ~n73423 ;
  assign n73419 = ~n72161 & n72195 ;
  assign n73425 = ~n72168 & ~n73419 ;
  assign n73426 = ~n73113 & ~n73425 ;
  assign n73427 = ~n73424 & ~n73426 ;
  assign n73420 = ~n72224 & ~n73419 ;
  assign n73421 = n72168 & ~n73420 ;
  assign n73428 = n73098 & ~n73422 ;
  assign n73429 = ~n73421 & ~n73428 ;
  assign n73430 = ~n73427 & n73429 ;
  assign n73431 = ~n72149 & ~n73430 ;
  assign n73432 = n72168 & ~n72208 ;
  assign n73433 = ~n72168 & ~n72221 ;
  assign n73434 = ~n73099 & n73433 ;
  assign n73435 = ~n73432 & ~n73434 ;
  assign n73450 = ~n73431 & ~n73435 ;
  assign n73451 = ~n73449 & n73450 ;
  assign n73452 = \u0_desIn_r_reg[56]/NET0131  & n73451 ;
  assign n73453 = ~\u0_desIn_r_reg[56]/NET0131  & ~n73451 ;
  assign n73454 = ~n73452 & ~n73453 ;
  assign n73468 = ~n72746 & ~n72748 ;
  assign n73469 = ~n72742 & n73468 ;
  assign n73470 = ~n72702 & ~n73469 ;
  assign n73464 = n72721 & n73065 ;
  assign n73465 = ~n72721 & n72767 ;
  assign n73466 = ~n72769 & ~n73465 ;
  assign n73467 = n72702 & ~n73466 ;
  assign n73471 = ~n73464 & ~n73467 ;
  assign n73472 = ~n73470 & n73471 ;
  assign n73473 = ~n72761 & ~n73472 ;
  assign n73456 = n72715 & ~n72728 ;
  assign n73457 = ~n72766 & ~n73456 ;
  assign n73458 = n72702 & ~n73457 ;
  assign n73459 = ~n72702 & n72774 ;
  assign n73455 = ~n72708 & n72874 ;
  assign n73460 = ~n72736 & ~n73455 ;
  assign n73461 = ~n73459 & n73460 ;
  assign n73462 = ~n73458 & n73461 ;
  assign n73463 = n72761 & ~n73462 ;
  assign n73474 = ~n72702 & ~n72743 ;
  assign n73475 = ~n72784 & ~n72877 ;
  assign n73476 = n73474 & n73475 ;
  assign n73477 = n72702 & ~n72733 ;
  assign n73478 = ~n72788 & n73477 ;
  assign n73479 = ~n73476 & ~n73478 ;
  assign n73480 = ~n73463 & ~n73479 ;
  assign n73481 = ~n73473 & n73480 ;
  assign n73482 = ~\u0_desIn_r_reg[22]/NET0131  & ~n73481 ;
  assign n73483 = \u0_desIn_r_reg[22]/NET0131  & n73481 ;
  assign n73484 = ~n73482 & ~n73483 ;
  assign n73486 = n72536 & n72543 ;
  assign n73487 = ~n72570 & ~n73486 ;
  assign n73488 = n72557 & ~n72571 ;
  assign n73489 = ~n73487 & n73488 ;
  assign n73491 = ~n72557 & ~n73371 ;
  assign n73492 = n73487 & n73491 ;
  assign n73485 = n72537 & n72559 ;
  assign n73490 = ~n72562 & n72568 ;
  assign n73493 = ~n73485 & ~n73490 ;
  assign n73494 = ~n73492 & n73493 ;
  assign n73495 = ~n73489 & n73494 ;
  assign n73496 = ~n72524 & ~n73495 ;
  assign n73497 = n72537 & ~n72543 ;
  assign n73498 = ~n72578 & ~n73497 ;
  assign n73499 = n72557 & ~n73498 ;
  assign n73500 = n72557 & n72568 ;
  assign n73501 = n72592 & n73500 ;
  assign n73502 = ~n73499 & ~n73501 ;
  assign n73503 = n72524 & ~n73502 ;
  assign n73504 = ~n73358 & ~n73486 ;
  assign n73505 = n72588 & ~n73504 ;
  assign n73509 = n72543 & ~n72561 ;
  assign n73510 = n72579 & n73509 ;
  assign n73506 = ~n72550 & n73486 ;
  assign n73507 = n72564 & n73506 ;
  assign n73508 = n72570 & n73352 ;
  assign n73511 = ~n73507 & ~n73508 ;
  assign n73512 = ~n73510 & n73511 ;
  assign n73513 = ~n73505 & n73512 ;
  assign n73514 = ~n73503 & n73513 ;
  assign n73515 = ~n73496 & n73514 ;
  assign n73516 = \u0_desIn_r_reg[40]/NET0131  & ~n73515 ;
  assign n73517 = ~\u0_desIn_r_reg[40]/NET0131  & n73515 ;
  assign n73518 = ~n73516 & ~n73517 ;
  assign n73519 = n72182 & n73422 ;
  assign n73523 = ~n72217 & ~n73099 ;
  assign n73524 = ~n73436 & n73523 ;
  assign n73525 = ~n73519 & n73524 ;
  assign n73526 = ~n72168 & ~n73525 ;
  assign n73520 = ~n72224 & ~n73519 ;
  assign n73521 = n72174 & ~n73520 ;
  assign n73527 = ~n72183 & ~n73422 ;
  assign n73528 = n72168 & ~n72174 ;
  assign n73529 = n73527 & n73528 ;
  assign n73530 = ~n73521 & ~n73529 ;
  assign n73531 = ~n73526 & n73530 ;
  assign n73532 = n72149 & ~n73531 ;
  assign n73537 = ~n72194 & ~n73422 ;
  assign n73538 = ~n73098 & ~n73537 ;
  assign n73539 = ~n73428 & ~n73538 ;
  assign n73536 = n72149 & ~n72185 ;
  assign n73540 = n72168 & ~n73536 ;
  assign n73541 = ~n73539 & n73540 ;
  assign n73522 = ~n72168 & n73521 ;
  assign n73533 = n72175 & n73527 ;
  assign n73534 = ~n72185 & ~n73533 ;
  assign n73535 = ~n72149 & ~n73534 ;
  assign n73542 = ~n73522 & ~n73535 ;
  assign n73543 = ~n73541 & n73542 ;
  assign n73544 = ~n73532 & n73543 ;
  assign n73545 = ~\u0_desIn_r_reg[54]/NET0131  & ~n73544 ;
  assign n73546 = \u0_desIn_r_reg[54]/NET0131  & n73544 ;
  assign n73547 = ~n73545 & ~n73546 ;
  assign n73548 = n72272 & n73191 ;
  assign n73549 = ~n73209 & ~n73548 ;
  assign n73550 = ~n72309 & ~n73549 ;
  assign n73553 = n72294 & ~n72300 ;
  assign n73554 = n72245 & ~n73201 ;
  assign n73555 = ~n73553 & n73554 ;
  assign n73551 = ~n72277 & n73201 ;
  assign n73552 = ~n72245 & n73551 ;
  assign n73556 = ~n72292 & ~n73552 ;
  assign n73557 = ~n73555 & n73556 ;
  assign n73558 = ~n73550 & n73557 ;
  assign n73560 = ~n73202 & ~n73278 ;
  assign n73561 = n72251 & ~n73560 ;
  assign n73559 = n72252 & n73551 ;
  assign n73562 = n73189 & ~n73559 ;
  assign n73563 = ~n73561 & n73562 ;
  assign n73564 = ~n73558 & ~n73563 ;
  assign n73565 = n72272 & ~n72282 ;
  assign n73566 = ~n72284 & n72308 ;
  assign n73567 = n73565 & n73566 ;
  assign n73568 = ~n73564 & ~n73567 ;
  assign n73569 = ~\u0_desIn_r_reg[4]/NET0131  & ~n73568 ;
  assign n73570 = \u0_desIn_r_reg[4]/NET0131  & n73568 ;
  assign n73571 = ~n73569 & ~n73570 ;
  assign n73572 = ~n72454 & ~n73388 ;
  assign n73573 = n72470 & ~n73572 ;
  assign n73574 = ~n72453 & n73337 ;
  assign n73575 = ~n73573 & ~n73574 ;
  assign n73576 = ~n72434 & ~n73575 ;
  assign n73580 = ~n72470 & ~n72510 ;
  assign n73578 = ~n72434 & n72455 ;
  assign n73579 = n72447 & n72504 ;
  assign n73581 = ~n73578 & ~n73579 ;
  assign n73582 = n73580 & n73581 ;
  assign n73577 = ~n72446 & n72488 ;
  assign n73583 = ~n72502 & ~n73577 ;
  assign n73584 = n73582 & n73583 ;
  assign n73585 = n72470 & ~n72489 ;
  assign n73586 = ~n73340 & n73585 ;
  assign n73587 = ~n73584 & ~n73586 ;
  assign n73588 = n72453 & n72490 ;
  assign n73589 = n72479 & n73317 ;
  assign n73591 = ~n73588 & ~n73589 ;
  assign n73592 = ~n73336 & n73591 ;
  assign n73590 = n72470 & n73333 ;
  assign n73593 = ~n73577 & ~n73590 ;
  assign n73594 = n73592 & n73593 ;
  assign n73595 = n72434 & ~n73594 ;
  assign n73596 = ~n73587 & ~n73595 ;
  assign n73597 = ~n73576 & n73596 ;
  assign n73598 = ~\u0_desIn_r_reg[52]/NET0131  & ~n73597 ;
  assign n73599 = \u0_desIn_r_reg[52]/NET0131  & n73597 ;
  assign n73600 = ~n73598 & ~n73599 ;
  assign n73601 = decrypt_pad & \key3[51]_pad  ;
  assign n73602 = ~decrypt_pad & \key1[51]_pad  ;
  assign n73603 = ~n73601 & ~n73602 ;
  assign n73604 = decrypt_pad & \key1[33]_pad  ;
  assign n73605 = ~decrypt_pad & \key3[33]_pad  ;
  assign n73606 = ~n73604 & ~n73605 ;
  assign n73607 = decrypt_pad & \key1[35]_pad  ;
  assign n73608 = ~decrypt_pad & \key3[35]_pad  ;
  assign n73609 = ~n73607 & ~n73608 ;
  assign n73610 = decrypt_pad & \key1[45]_pad  ;
  assign n73611 = ~decrypt_pad & \key3[45]_pad  ;
  assign n73612 = ~n73610 & ~n73611 ;
  assign n73613 = decrypt_pad & \key1[7]_pad  ;
  assign n73614 = ~decrypt_pad & \key3[7]_pad  ;
  assign n73615 = ~n73613 & ~n73614 ;
  assign n73616 = decrypt_pad & \key1[38]_pad  ;
  assign n73617 = ~decrypt_pad & \key3[38]_pad  ;
  assign n73618 = ~n73616 & ~n73617 ;
  assign n73619 = decrypt_pad & \key3[23]_pad  ;
  assign n73620 = ~decrypt_pad & \key1[23]_pad  ;
  assign n73621 = ~n73619 & ~n73620 ;
  assign n73622 = decrypt_pad & \key1[11]_pad  ;
  assign n73623 = ~decrypt_pad & \key3[11]_pad  ;
  assign n73624 = ~n73622 & ~n73623 ;
  assign n73625 = decrypt_pad & \key1[27]_pad  ;
  assign n73626 = ~decrypt_pad & \key3[27]_pad  ;
  assign n73627 = ~n73625 & ~n73626 ;
  assign n73628 = decrypt_pad & \key1[32]_pad  ;
  assign n73629 = ~decrypt_pad & \key3[32]_pad  ;
  assign n73630 = ~n73628 & ~n73629 ;
  assign n73631 = decrypt_pad & \key3[10]_pad  ;
  assign n73632 = ~decrypt_pad & \key1[10]_pad  ;
  assign n73633 = ~n73631 & ~n73632 ;
  assign n73634 = decrypt_pad & \key3[19]_pad  ;
  assign n73635 = ~decrypt_pad & \key1[19]_pad  ;
  assign n73636 = ~n73634 & ~n73635 ;
  assign n73637 = decrypt_pad & \key3[14]_pad  ;
  assign n73638 = ~decrypt_pad & \key1[14]_pad  ;
  assign n73639 = ~n73637 & ~n73638 ;
  assign n73640 = decrypt_pad & \key3[12]_pad  ;
  assign n73641 = ~decrypt_pad & \key1[12]_pad  ;
  assign n73642 = ~n73640 & ~n73641 ;
  assign n73643 = decrypt_pad & \key3[30]_pad  ;
  assign n73644 = ~decrypt_pad & \key1[30]_pad  ;
  assign n73645 = ~n73643 & ~n73644 ;
  assign n73646 = decrypt_pad & \key3[17]_pad  ;
  assign n73647 = ~decrypt_pad & \key1[17]_pad  ;
  assign n73648 = ~n73646 & ~n73647 ;
  assign n73649 = decrypt_pad & \key3[2]_pad  ;
  assign n73650 = ~decrypt_pad & \key1[2]_pad  ;
  assign n73651 = ~n73649 & ~n73650 ;
  assign n73652 = decrypt_pad & \key1[10]_pad  ;
  assign n73653 = ~decrypt_pad & \key3[10]_pad  ;
  assign n73654 = ~n73652 & ~n73653 ;
  assign n73655 = decrypt_pad & \key3[3]_pad  ;
  assign n73656 = ~decrypt_pad & \key1[3]_pad  ;
  assign n73657 = ~n73655 & ~n73656 ;
  assign n73658 = decrypt_pad & \key1[37]_pad  ;
  assign n73659 = ~decrypt_pad & \key3[37]_pad  ;
  assign n73660 = ~n73658 & ~n73659 ;
  assign n73661 = decrypt_pad & \key1[40]_pad  ;
  assign n73662 = ~decrypt_pad & \key3[40]_pad  ;
  assign n73663 = ~n73661 & ~n73662 ;
  assign n73664 = decrypt_pad & \key3[33]_pad  ;
  assign n73665 = ~decrypt_pad & \key1[33]_pad  ;
  assign n73666 = ~n73664 & ~n73665 ;
  assign n73667 = decrypt_pad & \key1[6]_pad  ;
  assign n73668 = ~decrypt_pad & \key3[6]_pad  ;
  assign n73669 = ~n73667 & ~n73668 ;
  assign n73670 = decrypt_pad & \key1[53]_pad  ;
  assign n73671 = ~decrypt_pad & \key3[53]_pad  ;
  assign n73672 = ~n73670 & ~n73671 ;
  assign n73673 = decrypt_pad & \key3[24]_pad  ;
  assign n73674 = ~decrypt_pad & \key1[24]_pad  ;
  assign n73675 = ~n73673 & ~n73674 ;
  assign n73676 = decrypt_pad & \key1[34]_pad  ;
  assign n73677 = ~decrypt_pad & \key3[34]_pad  ;
  assign n73678 = ~n73676 & ~n73677 ;
  assign n73679 = decrypt_pad & \key3[49]_pad  ;
  assign n73680 = ~decrypt_pad & \key1[49]_pad  ;
  assign n73681 = ~n73679 & ~n73680 ;
  assign n73682 = decrypt_pad & \key1[14]_pad  ;
  assign n73683 = ~decrypt_pad & \key3[14]_pad  ;
  assign n73684 = ~n73682 & ~n73683 ;
  assign n73685 = decrypt_pad & \key1[29]_pad  ;
  assign n73686 = ~decrypt_pad & \key3[29]_pad  ;
  assign n73687 = ~n73685 & ~n73686 ;
  assign n73688 = decrypt_pad & \key1[21]_pad  ;
  assign n73689 = ~decrypt_pad & \key3[21]_pad  ;
  assign n73690 = ~n73688 & ~n73689 ;
  assign n73691 = decrypt_pad & \key3[4]_pad  ;
  assign n73692 = ~decrypt_pad & \key1[4]_pad  ;
  assign n73693 = ~n73691 & ~n73692 ;
  assign n73694 = decrypt_pad & \key3[37]_pad  ;
  assign n73695 = ~decrypt_pad & \key1[37]_pad  ;
  assign n73696 = ~n73694 & ~n73695 ;
  assign n73697 = decrypt_pad & \key3[53]_pad  ;
  assign n73698 = ~decrypt_pad & \key1[53]_pad  ;
  assign n73699 = ~n73697 & ~n73698 ;
  assign n73700 = decrypt_pad & \key3[31]_pad  ;
  assign n73701 = ~decrypt_pad & \key1[31]_pad  ;
  assign n73702 = ~n73700 & ~n73701 ;
  assign n73703 = decrypt_pad & \key1[42]_pad  ;
  assign n73704 = ~decrypt_pad & \key3[42]_pad  ;
  assign n73705 = ~n73703 & ~n73704 ;
  assign n73706 = decrypt_pad & \key3[43]_pad  ;
  assign n73707 = ~decrypt_pad & \key1[43]_pad  ;
  assign n73708 = ~n73706 & ~n73707 ;
  assign n73709 = decrypt_pad & \key1[55]_pad  ;
  assign n73710 = ~decrypt_pad & \key3[55]_pad  ;
  assign n73711 = ~n73709 & ~n73710 ;
  assign n73712 = decrypt_pad & \key3[20]_pad  ;
  assign n73713 = ~decrypt_pad & \key1[20]_pad  ;
  assign n73714 = ~n73712 & ~n73713 ;
  assign n73715 = decrypt_pad & \key3[36]_pad  ;
  assign n73716 = ~decrypt_pad & \key1[36]_pad  ;
  assign n73717 = ~n73715 & ~n73716 ;
  assign n73718 = decrypt_pad & \key1[22]_pad  ;
  assign n73719 = ~decrypt_pad & \key3[22]_pad  ;
  assign n73720 = ~n73718 & ~n73719 ;
  assign n73721 = decrypt_pad & \key3[55]_pad  ;
  assign n73722 = ~decrypt_pad & \key1[55]_pad  ;
  assign n73723 = ~n73721 & ~n73722 ;
  assign n73724 = decrypt_pad & \key3[15]_pad  ;
  assign n73725 = ~decrypt_pad & \key1[15]_pad  ;
  assign n73726 = ~n73724 & ~n73725 ;
  assign n73727 = decrypt_pad & \key3[40]_pad  ;
  assign n73728 = ~decrypt_pad & \key1[40]_pad  ;
  assign n73729 = ~n73727 & ~n73728 ;
  assign n73730 = decrypt_pad & \key3[8]_pad  ;
  assign n73731 = ~decrypt_pad & \key1[8]_pad  ;
  assign n73732 = ~n73730 & ~n73731 ;
  assign n73733 = decrypt_pad & \key1[16]_pad  ;
  assign n73734 = ~decrypt_pad & \key3[16]_pad  ;
  assign n73735 = ~n73733 & ~n73734 ;
  assign n73736 = decrypt_pad & \key3[22]_pad  ;
  assign n73737 = ~decrypt_pad & \key1[22]_pad  ;
  assign n73738 = ~n73736 & ~n73737 ;
  assign n73739 = decrypt_pad & \key3[27]_pad  ;
  assign n73740 = ~decrypt_pad & \key1[27]_pad  ;
  assign n73741 = ~n73739 & ~n73740 ;
  assign n73742 = decrypt_pad & \key1[31]_pad  ;
  assign n73743 = ~decrypt_pad & \key3[31]_pad  ;
  assign n73744 = ~n73742 & ~n73743 ;
  assign n73745 = decrypt_pad & \key1[46]_pad  ;
  assign n73746 = ~decrypt_pad & \key3[46]_pad  ;
  assign n73747 = ~n73745 & ~n73746 ;
  assign n73748 = decrypt_pad & \key3[26]_pad  ;
  assign n73749 = ~decrypt_pad & \key1[26]_pad  ;
  assign n73750 = ~n73748 & ~n73749 ;
  assign n73751 = decrypt_pad & \key1[24]_pad  ;
  assign n73752 = ~decrypt_pad & \key3[24]_pad  ;
  assign n73753 = ~n73751 & ~n73752 ;
  assign n73754 = decrypt_pad & \key3[35]_pad  ;
  assign n73755 = ~decrypt_pad & \key1[35]_pad  ;
  assign n73756 = ~n73754 & ~n73755 ;
  assign n73757 = decrypt_pad & \key3[28]_pad  ;
  assign n73758 = ~decrypt_pad & \key1[28]_pad  ;
  assign n73759 = ~n73757 & ~n73758 ;
  assign n73760 = decrypt_pad & \key3[48]_pad  ;
  assign n73761 = ~decrypt_pad & \key1[48]_pad  ;
  assign n73762 = ~n73760 & ~n73761 ;
  assign n73763 = decrypt_pad & \key1[15]_pad  ;
  assign n73764 = ~decrypt_pad & \key3[15]_pad  ;
  assign n73765 = ~n73763 & ~n73764 ;
  assign n73766 = decrypt_pad & \key3[38]_pad  ;
  assign n73767 = ~decrypt_pad & \key1[38]_pad  ;
  assign n73768 = ~n73766 & ~n73767 ;
  assign n73769 = decrypt_pad & \key3[45]_pad  ;
  assign n73770 = ~decrypt_pad & \key1[45]_pad  ;
  assign n73771 = ~n73769 & ~n73770 ;
  assign n73772 = decrypt_pad & \key1[50]_pad  ;
  assign n73773 = ~decrypt_pad & \key3[50]_pad  ;
  assign n73774 = ~n73772 & ~n73773 ;
  assign n73775 = decrypt_pad & \key1[26]_pad  ;
  assign n73776 = ~decrypt_pad & \key3[26]_pad  ;
  assign n73777 = ~n73775 & ~n73776 ;
  assign n73778 = decrypt_pad & \key3[9]_pad  ;
  assign n73779 = ~decrypt_pad & \key1[9]_pad  ;
  assign n73780 = ~n73778 & ~n73779 ;
  assign n73781 = decrypt_pad & \key1[39]_pad  ;
  assign n73782 = ~decrypt_pad & \key3[39]_pad  ;
  assign n73783 = ~n73781 & ~n73782 ;
  assign n73784 = decrypt_pad & \key3[54]_pad  ;
  assign n73785 = ~decrypt_pad & \key1[54]_pad  ;
  assign n73786 = ~n73784 & ~n73785 ;
  assign n73787 = decrypt_pad & \key3[25]_pad  ;
  assign n73788 = ~decrypt_pad & \key1[25]_pad  ;
  assign n73789 = ~n73787 & ~n73788 ;
  assign n73790 = decrypt_pad & \key1[8]_pad  ;
  assign n73791 = ~decrypt_pad & \key3[8]_pad  ;
  assign n73792 = ~n73790 & ~n73791 ;
  assign n73793 = decrypt_pad & \key1[0]_pad  ;
  assign n73794 = ~decrypt_pad & \key3[0]_pad  ;
  assign n73795 = ~n73793 & ~n73794 ;
  assign n73796 = decrypt_pad & \key1[20]_pad  ;
  assign n73797 = ~decrypt_pad & \key3[20]_pad  ;
  assign n73798 = ~n73796 & ~n73797 ;
  assign n73799 = decrypt_pad & \key3[46]_pad  ;
  assign n73800 = ~decrypt_pad & \key1[46]_pad  ;
  assign n73801 = ~n73799 & ~n73800 ;
  assign n73802 = decrypt_pad & \key1[25]_pad  ;
  assign n73803 = ~decrypt_pad & \key3[25]_pad  ;
  assign n73804 = ~n73802 & ~n73803 ;
  assign n73805 = decrypt_pad & \key1[44]_pad  ;
  assign n73806 = ~decrypt_pad & \key3[44]_pad  ;
  assign n73807 = ~n73805 & ~n73806 ;
  assign n73808 = decrypt_pad & \key1[51]_pad  ;
  assign n73809 = ~decrypt_pad & \key3[51]_pad  ;
  assign n73810 = ~n73808 & ~n73809 ;
  assign n73811 = decrypt_pad & \key3[50]_pad  ;
  assign n73812 = ~decrypt_pad & \key1[50]_pad  ;
  assign n73813 = ~n73811 & ~n73812 ;
  assign n73814 = decrypt_pad & \key3[32]_pad  ;
  assign n73815 = ~decrypt_pad & \key1[32]_pad  ;
  assign n73816 = ~n73814 & ~n73815 ;
  assign n73817 = decrypt_pad & \key1[43]_pad  ;
  assign n73818 = ~decrypt_pad & \key3[43]_pad  ;
  assign n73819 = ~n73817 & ~n73818 ;
  assign n73820 = decrypt_pad & \key1[3]_pad  ;
  assign n73821 = ~decrypt_pad & \key3[3]_pad  ;
  assign n73822 = ~n73820 & ~n73821 ;
  assign n73823 = decrypt_pad & \key3[7]_pad  ;
  assign n73824 = ~decrypt_pad & \key1[7]_pad  ;
  assign n73825 = ~n73823 & ~n73824 ;
  assign n73826 = decrypt_pad & \key3[44]_pad  ;
  assign n73827 = ~decrypt_pad & \key1[44]_pad  ;
  assign n73828 = ~n73826 & ~n73827 ;
  assign n73829 = decrypt_pad & \key1[54]_pad  ;
  assign n73830 = ~decrypt_pad & \key3[54]_pad  ;
  assign n73831 = ~n73829 & ~n73830 ;
  assign n73832 = decrypt_pad & \key1[30]_pad  ;
  assign n73833 = ~decrypt_pad & \key3[30]_pad  ;
  assign n73834 = ~n73832 & ~n73833 ;
  assign n73835 = decrypt_pad & \key3[1]_pad  ;
  assign n73836 = ~decrypt_pad & \key1[1]_pad  ;
  assign n73837 = ~n73835 & ~n73836 ;
  assign n73838 = decrypt_pad & \key1[18]_pad  ;
  assign n73839 = ~decrypt_pad & \key3[18]_pad  ;
  assign n73840 = ~n73838 & ~n73839 ;
  assign n73841 = decrypt_pad & \key1[28]_pad  ;
  assign n73842 = ~decrypt_pad & \key3[28]_pad  ;
  assign n73843 = ~n73841 & ~n73842 ;
  assign n73844 = decrypt_pad & \key3[39]_pad  ;
  assign n73845 = ~decrypt_pad & \key1[39]_pad  ;
  assign n73846 = ~n73844 & ~n73845 ;
  assign n73847 = decrypt_pad & \key1[17]_pad  ;
  assign n73848 = ~decrypt_pad & \key3[17]_pad  ;
  assign n73849 = ~n73847 & ~n73848 ;
  assign n73850 = decrypt_pad & \key1[1]_pad  ;
  assign n73851 = ~decrypt_pad & \key3[1]_pad  ;
  assign n73852 = ~n73850 & ~n73851 ;
  assign n73853 = decrypt_pad & \key3[13]_pad  ;
  assign n73854 = ~decrypt_pad & \key1[13]_pad  ;
  assign n73855 = ~n73853 & ~n73854 ;
  assign n73856 = decrypt_pad & \key1[19]_pad  ;
  assign n73857 = ~decrypt_pad & \key3[19]_pad  ;
  assign n73858 = ~n73856 & ~n73857 ;
  assign n73859 = decrypt_pad & \key3[6]_pad  ;
  assign n73860 = ~decrypt_pad & \key1[6]_pad  ;
  assign n73861 = ~n73859 & ~n73860 ;
  assign n73862 = decrypt_pad & \key1[47]_pad  ;
  assign n73863 = ~decrypt_pad & \key3[47]_pad  ;
  assign n73864 = ~n73862 & ~n73863 ;
  assign n73865 = decrypt_pad & \key1[23]_pad  ;
  assign n73866 = ~decrypt_pad & \key3[23]_pad  ;
  assign n73867 = ~n73865 & ~n73866 ;
  assign n73868 = decrypt_pad & \key1[12]_pad  ;
  assign n73869 = ~decrypt_pad & \key3[12]_pad  ;
  assign n73870 = ~n73868 & ~n73869 ;
  assign n73871 = decrypt_pad & \key3[52]_pad  ;
  assign n73872 = ~decrypt_pad & \key1[52]_pad  ;
  assign n73873 = ~n73871 & ~n73872 ;
  assign n73874 = decrypt_pad & \key1[5]_pad  ;
  assign n73875 = ~decrypt_pad & \key3[5]_pad  ;
  assign n73876 = ~n73874 & ~n73875 ;
  assign n73877 = decrypt_pad & \key1[9]_pad  ;
  assign n73878 = ~decrypt_pad & \key3[9]_pad  ;
  assign n73879 = ~n73877 & ~n73878 ;
  assign n73880 = decrypt_pad & \key3[0]_pad  ;
  assign n73881 = ~decrypt_pad & \key1[0]_pad  ;
  assign n73882 = ~n73880 & ~n73881 ;
  assign n73883 = decrypt_pad & \key1[4]_pad  ;
  assign n73884 = ~decrypt_pad & \key3[4]_pad  ;
  assign n73885 = ~n73883 & ~n73884 ;
  assign n73886 = decrypt_pad & \key3[11]_pad  ;
  assign n73887 = ~decrypt_pad & \key1[11]_pad  ;
  assign n73888 = ~n73886 & ~n73887 ;
  assign n73889 = decrypt_pad & \key1[52]_pad  ;
  assign n73890 = ~decrypt_pad & \key3[52]_pad  ;
  assign n73891 = ~n73889 & ~n73890 ;
  assign n73892 = decrypt_pad & \key3[18]_pad  ;
  assign n73893 = ~decrypt_pad & \key1[18]_pad  ;
  assign n73894 = ~n73892 & ~n73893 ;
  assign n73895 = decrypt_pad & \key1[36]_pad  ;
  assign n73896 = ~decrypt_pad & \key3[36]_pad  ;
  assign n73897 = ~n73895 & ~n73896 ;
  assign n73898 = decrypt_pad & \key3[5]_pad  ;
  assign n73899 = ~decrypt_pad & \key1[5]_pad  ;
  assign n73900 = ~n73898 & ~n73899 ;
  assign n73901 = decrypt_pad & \key3[42]_pad  ;
  assign n73902 = ~decrypt_pad & \key1[42]_pad  ;
  assign n73903 = ~n73901 & ~n73902 ;
  assign n73904 = decrypt_pad & \key1[2]_pad  ;
  assign n73905 = ~decrypt_pad & \key3[2]_pad  ;
  assign n73906 = ~n73904 & ~n73905 ;
  assign n73907 = decrypt_pad & \key1[48]_pad  ;
  assign n73908 = ~decrypt_pad & \key3[48]_pad  ;
  assign n73909 = ~n73907 & ~n73908 ;
  assign n73910 = decrypt_pad & \key3[34]_pad  ;
  assign n73911 = ~decrypt_pad & \key1[34]_pad  ;
  assign n73912 = ~n73910 & ~n73911 ;
  assign n73913 = decrypt_pad & \key3[21]_pad  ;
  assign n73914 = ~decrypt_pad & \key1[21]_pad  ;
  assign n73915 = ~n73913 & ~n73914 ;
  assign n73916 = decrypt_pad & \key1[49]_pad  ;
  assign n73917 = ~decrypt_pad & \key3[49]_pad  ;
  assign n73918 = ~n73916 & ~n73917 ;
  assign n73919 = decrypt_pad & \key3[47]_pad  ;
  assign n73920 = ~decrypt_pad & \key1[47]_pad  ;
  assign n73921 = ~n73919 & ~n73920 ;
  assign n73922 = decrypt_pad & \key3[29]_pad  ;
  assign n73923 = ~decrypt_pad & \key1[29]_pad  ;
  assign n73924 = ~n73922 & ~n73923 ;
  assign n73925 = decrypt_pad & \key1[13]_pad  ;
  assign n73926 = ~decrypt_pad & \key3[13]_pad  ;
  assign n73927 = ~n73925 & ~n73926 ;
  assign n73928 = decrypt_pad & \key1[41]_pad  ;
  assign n73929 = ~decrypt_pad & \key3[41]_pad  ;
  assign n73930 = ~n73928 & ~n73929 ;
  assign n73931 = decrypt_pad & \key3[41]_pad  ;
  assign n73932 = ~decrypt_pad & \key1[41]_pad  ;
  assign n73933 = ~n73931 & ~n73932 ;
  assign n73934 = decrypt_pad & \key3[16]_pad  ;
  assign n73935 = ~decrypt_pad & \key1[16]_pad  ;
  assign n73936 = ~n73934 & ~n73935 ;
  assign n73938 = n47023 & n47039 ;
  assign n73939 = n46984 & ~n47048 ;
  assign n73940 = ~n47233 & n73939 ;
  assign n73941 = ~n73938 & n73940 ;
  assign n73937 = ~n47023 & ~n47297 ;
  assign n73942 = ~n47224 & ~n73937 ;
  assign n73943 = n73941 & n73942 ;
  assign n73944 = ~n47023 & ~n47054 ;
  assign n73945 = ~n47208 & n73944 ;
  assign n73946 = n47023 & ~n47038 ;
  assign n73947 = ~n47279 & n73946 ;
  assign n73948 = ~n73945 & ~n73947 ;
  assign n73949 = ~n46984 & ~n47052 ;
  assign n73950 = ~n47027 & n73949 ;
  assign n73951 = ~n47056 & n73950 ;
  assign n73952 = ~n73948 & n73951 ;
  assign n73953 = ~n73943 & ~n73952 ;
  assign n73955 = ~n46996 & n47023 ;
  assign n73956 = ~n47277 & n73955 ;
  assign n73954 = ~n47023 & n47292 ;
  assign n73957 = ~n47049 & ~n73954 ;
  assign n73958 = ~n73956 & n73957 ;
  assign n73959 = ~n73953 & n73958 ;
  assign n73960 = ~\u1_L1_reg[20]/NET0131  & ~n73959 ;
  assign n73961 = \u1_L1_reg[20]/NET0131  & n73959 ;
  assign n73962 = ~n73960 & ~n73961 ;
  assign n73964 = ~n58296 & n58423 ;
  assign n73965 = n57468 & ~n73964 ;
  assign n73966 = ~n57524 & ~n58312 ;
  assign n73967 = ~n57468 & ~n73966 ;
  assign n73963 = n57474 & n58298 ;
  assign n73968 = ~n57474 & n58303 ;
  assign n73969 = ~n73963 & ~n73968 ;
  assign n73970 = ~n73967 & n73969 ;
  assign n73971 = ~n73965 & n73970 ;
  assign n73972 = ~n57495 & ~n73971 ;
  assign n73973 = ~n57481 & n58317 ;
  assign n73974 = ~n73968 & ~n73973 ;
  assign n73975 = ~n57468 & ~n73974 ;
  assign n73977 = n57474 & ~n57506 ;
  assign n73978 = ~n58298 & n73977 ;
  assign n73976 = n57475 & ~n73966 ;
  assign n73979 = ~n58316 & ~n73976 ;
  assign n73980 = ~n73978 & n73979 ;
  assign n73981 = n57495 & ~n73980 ;
  assign n73982 = ~n73975 & ~n73981 ;
  assign n73983 = ~n73972 & n73982 ;
  assign n73984 = ~\u0_L9_reg[9]/NET0131  & ~n73983 ;
  assign n73985 = \u0_L9_reg[9]/NET0131  & n73983 ;
  assign n73986 = ~n73984 & ~n73985 ;
  assign n74002 = ~n71092 & ~n71093 ;
  assign n74003 = n71038 & ~n74002 ;
  assign n73999 = n71055 & ~n71453 ;
  assign n74000 = ~n71054 & ~n73999 ;
  assign n74001 = ~n71038 & ~n74000 ;
  assign n74004 = n71444 & ~n74001 ;
  assign n74005 = ~n74003 & n74004 ;
  assign n74006 = n71067 & ~n74005 ;
  assign n73988 = ~n71106 & ~n71453 ;
  assign n73989 = n71031 & ~n73988 ;
  assign n73987 = n71039 & ~n71052 ;
  assign n73994 = ~n71094 & ~n73987 ;
  assign n73990 = ~n71031 & ~n71085 ;
  assign n73991 = n71785 & n73990 ;
  assign n73992 = n71031 & n71082 ;
  assign n73993 = ~n71105 & n73992 ;
  assign n73995 = ~n73991 & ~n73993 ;
  assign n73996 = n73994 & n73995 ;
  assign n73997 = ~n73989 & n73996 ;
  assign n73998 = ~n71067 & ~n73997 ;
  assign n74007 = ~n71096 & n71444 ;
  assign n74008 = ~n71038 & ~n74007 ;
  assign n74009 = ~n71086 & ~n71110 ;
  assign n74010 = ~n74008 & n74009 ;
  assign n74011 = ~n73998 & n74010 ;
  assign n74012 = ~n74006 & n74011 ;
  assign n74013 = \u0_L0_reg[10]/NET0131  & n74012 ;
  assign n74014 = ~\u0_L0_reg[10]/NET0131  & ~n74012 ;
  assign n74015 = ~n74013 & ~n74014 ;
  assign n74016 = ~n37946 & n37952 ;
  assign n74017 = n37948 & ~n74016 ;
  assign n74018 = ~n37962 & n38632 ;
  assign n74019 = ~n74017 & ~n74018 ;
  assign n74020 = ~n38507 & ~n74019 ;
  assign n74021 = n37976 & ~n74020 ;
  assign n74022 = ~n37939 & n38000 ;
  assign n74027 = ~n37993 & ~n74022 ;
  assign n74023 = ~n37945 & ~n38649 ;
  assign n74024 = n38638 & ~n74023 ;
  assign n74025 = ~n37953 & ~n38635 ;
  assign n74026 = n37959 & ~n74025 ;
  assign n74028 = ~n74024 & ~n74026 ;
  assign n74029 = n74027 & n74028 ;
  assign n74030 = n37964 & n74029 ;
  assign n74031 = ~n37976 & ~n74030 ;
  assign n74032 = ~n37951 & ~n38507 ;
  assign n74033 = ~n37920 & ~n74032 ;
  assign n74034 = ~n37961 & ~n37970 ;
  assign n74035 = ~n74033 & n74034 ;
  assign n74036 = ~n74031 & n74035 ;
  assign n74037 = ~n74021 & n74036 ;
  assign n74038 = \u1_L7_reg[10]/NET0131  & n74037 ;
  assign n74039 = ~\u1_L7_reg[10]/NET0131  & ~n74037 ;
  assign n74040 = ~n74038 & ~n74039 ;
  assign n74041 = ~n63624 & n63927 ;
  assign n74042 = ~n63599 & ~n63606 ;
  assign n74043 = ~n63627 & ~n74042 ;
  assign n74044 = ~n63583 & ~n74043 ;
  assign n74045 = ~n63616 & ~n64200 ;
  assign n74046 = ~n63615 & ~n74045 ;
  assign n74047 = ~n63577 & ~n74046 ;
  assign n74048 = ~n74044 & n74047 ;
  assign n74049 = ~n74041 & ~n74048 ;
  assign n74051 = n63583 & n63626 ;
  assign n74050 = n63634 & n63638 ;
  assign n74052 = ~n63577 & ~n74050 ;
  assign n74053 = ~n74051 & n74052 ;
  assign n74054 = ~n63636 & ~n74053 ;
  assign n74057 = ~n63608 & ~n64197 ;
  assign n74058 = n63583 & ~n74057 ;
  assign n74055 = ~n63639 & ~n64204 ;
  assign n74056 = n63590 & ~n74055 ;
  assign n74059 = n63615 & ~n74056 ;
  assign n74060 = ~n74058 & n74059 ;
  assign n74061 = ~n74054 & n74060 ;
  assign n74062 = ~n63607 & n63645 ;
  assign n74063 = ~n63615 & ~n63643 ;
  assign n74064 = n63625 & n74063 ;
  assign n74065 = ~n74062 & n74064 ;
  assign n74066 = ~n74061 & ~n74065 ;
  assign n74067 = ~n74049 & ~n74066 ;
  assign n74068 = ~\u0_L5_reg[26]/NET0131  & ~n74067 ;
  assign n74069 = \u0_L5_reg[26]/NET0131  & n74067 ;
  assign n74070 = ~n74068 & ~n74069 ;
  assign n74089 = ~n66783 & ~n66796 ;
  assign n74090 = ~n66822 & n74089 ;
  assign n74091 = n66803 & ~n67485 ;
  assign n74092 = ~n67226 & n74091 ;
  assign n74093 = ~n74090 & n74092 ;
  assign n74094 = ~n66790 & ~n66803 ;
  assign n74095 = ~n66818 & n74094 ;
  assign n74096 = ~n74093 & ~n74095 ;
  assign n74097 = ~n66807 & ~n67232 ;
  assign n74098 = ~n74096 & n74097 ;
  assign n74099 = n66770 & ~n74098 ;
  assign n74078 = ~n66804 & ~n66809 ;
  assign n74079 = n66776 & n66789 ;
  assign n74080 = ~n66803 & ~n74079 ;
  assign n74081 = ~n74078 & n74080 ;
  assign n74076 = ~n66796 & n66803 ;
  assign n74077 = n66783 & n74076 ;
  assign n74074 = n66842 & n67485 ;
  assign n74075 = n66809 & n66811 ;
  assign n74082 = ~n74074 & ~n74075 ;
  assign n74083 = ~n74077 & n74082 ;
  assign n74084 = ~n74081 & n74083 ;
  assign n74085 = ~n66770 & ~n74084 ;
  assign n74071 = n66805 & n66811 ;
  assign n74072 = n67233 & ~n74071 ;
  assign n74073 = n66803 & ~n74072 ;
  assign n74086 = ~n66803 & n66844 ;
  assign n74087 = ~n66807 & ~n74086 ;
  assign n74088 = n66789 & ~n74087 ;
  assign n74100 = ~n74073 & ~n74088 ;
  assign n74101 = ~n74085 & n74100 ;
  assign n74102 = ~n74099 & n74101 ;
  assign n74103 = \u0_L3_reg[25]/NET0131  & n74102 ;
  assign n74104 = ~\u0_L3_reg[25]/NET0131  & ~n74102 ;
  assign n74105 = ~n74103 & ~n74104 ;
  assign n74122 = ~n72537 & n73500 ;
  assign n74118 = ~n72557 & ~n72568 ;
  assign n74119 = ~n72562 & n74118 ;
  assign n74120 = n72543 & ~n73351 ;
  assign n74121 = n73376 & n74120 ;
  assign n74123 = ~n74119 & ~n74121 ;
  assign n74124 = ~n74122 & n74123 ;
  assign n74125 = ~n72569 & n74124 ;
  assign n74126 = n72524 & ~n74125 ;
  assign n74106 = ~n73358 & ~n73506 ;
  assign n74107 = n73498 & n74106 ;
  assign n74108 = n72557 & ~n74107 ;
  assign n74109 = n72559 & n72592 ;
  assign n74110 = ~n74108 & ~n74109 ;
  assign n74111 = ~n72524 & ~n74110 ;
  assign n74115 = n72594 & ~n73490 ;
  assign n74116 = ~n72524 & ~n72557 ;
  assign n74117 = ~n74115 & n74116 ;
  assign n74113 = n72537 & n72557 ;
  assign n74114 = n72566 & n74113 ;
  assign n74112 = n73352 & n73354 ;
  assign n74127 = ~n73501 & ~n74112 ;
  assign n74128 = ~n74114 & n74127 ;
  assign n74129 = ~n74117 & n74128 ;
  assign n74130 = ~n74111 & n74129 ;
  assign n74131 = ~n74126 & n74130 ;
  assign n74132 = \u0_desIn_r_reg[58]/NET0131  & n74131 ;
  assign n74133 = ~\u0_desIn_r_reg[58]/NET0131  & ~n74131 ;
  assign n74134 = ~n74132 & ~n74133 ;
  assign n74135 = ~n30875 & n30897 ;
  assign n74136 = n30785 & ~n74135 ;
  assign n74137 = n30792 & n74136 ;
  assign n74138 = n30794 & n30816 ;
  assign n74139 = ~n30785 & ~n31400 ;
  assign n74140 = ~n74138 & n74139 ;
  assign n74141 = ~n74137 & ~n74140 ;
  assign n74143 = n30785 & ~n30803 ;
  assign n74144 = ~n30880 & n74143 ;
  assign n74146 = ~n30793 & n74144 ;
  assign n74147 = n30771 & ~n74146 ;
  assign n74142 = ~n30785 & ~n30787 ;
  assign n74145 = ~n74142 & ~n74144 ;
  assign n74148 = n30785 & ~n30881 ;
  assign n74149 = n30818 & ~n74148 ;
  assign n74150 = ~n30816 & ~n74149 ;
  assign n74151 = ~n74145 & n74150 ;
  assign n74152 = ~n74147 & n74151 ;
  assign n74153 = ~n31400 & ~n31402 ;
  assign n74154 = n30785 & ~n74153 ;
  assign n74155 = ~n31407 & ~n74154 ;
  assign n74156 = ~n30805 & n30816 ;
  assign n74157 = ~n74155 & n74156 ;
  assign n74158 = ~n74152 & ~n74157 ;
  assign n74159 = ~n74141 & ~n74158 ;
  assign n74160 = \u1_L12_reg[5]/NET0131  & ~n74159 ;
  assign n74161 = ~\u1_L12_reg[5]/NET0131  & n74159 ;
  assign n74162 = ~n74160 & ~n74161 ;
  assign n74166 = n60746 & ~n60836 ;
  assign n74167 = ~n61252 & n74166 ;
  assign n74168 = ~n60746 & ~n61241 ;
  assign n74169 = ~n60846 & n74168 ;
  assign n74170 = ~n74167 & ~n74169 ;
  assign n74171 = ~n60718 & ~n60835 ;
  assign n74172 = ~n61242 & ~n61268 ;
  assign n74173 = n74171 & n74172 ;
  assign n74174 = ~n61253 & n74173 ;
  assign n74175 = ~n74170 & n74174 ;
  assign n74176 = ~n60746 & ~n60791 ;
  assign n74177 = n60763 & n60780 ;
  assign n74178 = n60718 & ~n74177 ;
  assign n74179 = n60762 & n74178 ;
  assign n74180 = ~n60837 & ~n60849 ;
  assign n74181 = n74179 & n74180 ;
  assign n74182 = ~n74176 & n74181 ;
  assign n74183 = ~n74175 & ~n74182 ;
  assign n74163 = ~n60846 & ~n60860 ;
  assign n74164 = n60780 & ~n74163 ;
  assign n74165 = ~n60746 & n60761 ;
  assign n74184 = ~n61256 & ~n74165 ;
  assign n74185 = ~n74164 & n74184 ;
  assign n74186 = ~n74183 & n74185 ;
  assign n74187 = ~\u0_L7_reg[20]/NET0131  & ~n74186 ;
  assign n74188 = \u0_L7_reg[20]/NET0131  & n74186 ;
  assign n74189 = ~n74187 & ~n74188 ;
  assign n74204 = n72953 & ~n73008 ;
  assign n74205 = n73044 & ~n74204 ;
  assign n74201 = ~n73011 & ~n73019 ;
  assign n74202 = n72947 & n72960 ;
  assign n74203 = ~n74201 & n74202 ;
  assign n74206 = ~n73053 & ~n73232 ;
  assign n74207 = ~n74203 & n74206 ;
  assign n74208 = ~n74205 & n74207 ;
  assign n74209 = ~n72985 & ~n74208 ;
  assign n74191 = n72941 & ~n72992 ;
  assign n74192 = ~n72954 & ~n72974 ;
  assign n74193 = ~n72941 & n72960 ;
  assign n74194 = ~n74192 & n74193 ;
  assign n74195 = ~n72968 & ~n74194 ;
  assign n74196 = ~n74191 & n74195 ;
  assign n74197 = n72985 & ~n74196 ;
  assign n74190 = ~n72941 & n72977 ;
  assign n74198 = n72947 & n72987 ;
  assign n74199 = ~n73237 & ~n74198 ;
  assign n74200 = n72941 & ~n74199 ;
  assign n74210 = ~n74190 & ~n74200 ;
  assign n74211 = ~n74197 & n74210 ;
  assign n74212 = ~n74209 & n74211 ;
  assign n74213 = \u0_desIn_r_reg[10]/NET0131  & n74212 ;
  assign n74214 = ~\u0_desIn_r_reg[10]/NET0131  & ~n74212 ;
  assign n74215 = ~n74213 & ~n74214 ;
  assign n74216 = n33823 & n33847 ;
  assign n74217 = n33831 & ~n74216 ;
  assign n74218 = ~n34308 & n74217 ;
  assign n74219 = n33868 & n74218 ;
  assign n74220 = n33842 & n33869 ;
  assign n74221 = ~n33831 & ~n34307 ;
  assign n74222 = ~n74220 & n74221 ;
  assign n74223 = ~n74219 & ~n74222 ;
  assign n74225 = ~n33807 & n33821 ;
  assign n74226 = ~n33801 & n33814 ;
  assign n74227 = ~n74225 & ~n74226 ;
  assign n74228 = n33831 & ~n34307 ;
  assign n74229 = ~n74227 & n74228 ;
  assign n74224 = ~n33831 & n34303 ;
  assign n74230 = n33842 & ~n33861 ;
  assign n74231 = ~n74224 & n74230 ;
  assign n74232 = ~n74229 & n74231 ;
  assign n74233 = ~n33824 & ~n33920 ;
  assign n74234 = n33831 & ~n74233 ;
  assign n74235 = ~n33917 & ~n34289 ;
  assign n74236 = n33814 & ~n74235 ;
  assign n74238 = ~n33850 & ~n33939 ;
  assign n74239 = ~n33808 & ~n33831 ;
  assign n74240 = ~n74238 & n74239 ;
  assign n74237 = n33807 & n33938 ;
  assign n74241 = ~n33842 & ~n74237 ;
  assign n74242 = ~n74240 & n74241 ;
  assign n74243 = ~n74236 & n74242 ;
  assign n74244 = ~n74234 & n74243 ;
  assign n74245 = ~n74232 & ~n74244 ;
  assign n74246 = ~n74223 & ~n74245 ;
  assign n74247 = \u1_L10_reg[5]/NET0131  & ~n74246 ;
  assign n74248 = ~\u1_L10_reg[5]/NET0131  & n74246 ;
  assign n74249 = ~n74247 & ~n74248 ;
  assign n74250 = n46550 & ~n46559 ;
  assign n74262 = ~n46528 & ~n46542 ;
  assign n74263 = n74250 & ~n74262 ;
  assign n74260 = n46522 & n46582 ;
  assign n74261 = ~n46550 & ~n46868 ;
  assign n74264 = ~n74260 & ~n74261 ;
  assign n74265 = ~n74263 & n74264 ;
  assign n74266 = ~n46516 & ~n74265 ;
  assign n74251 = ~n46550 & ~n46553 ;
  assign n74252 = ~n74250 & ~n74251 ;
  assign n74256 = ~n46564 & ~n74252 ;
  assign n74253 = ~n46542 & ~n46563 ;
  assign n74254 = ~n46522 & ~n74253 ;
  assign n74255 = n46522 & ~n46868 ;
  assign n74257 = ~n74254 & ~n74255 ;
  assign n74258 = n74256 & n74257 ;
  assign n74259 = n46516 & ~n74258 ;
  assign n74267 = ~n46554 & ~n46597 ;
  assign n74268 = n46551 & ~n74267 ;
  assign n74269 = ~n46590 & ~n74268 ;
  assign n74270 = ~n74259 & n74269 ;
  assign n74271 = ~n74266 & n74270 ;
  assign n74272 = ~\u1_L1_reg[19]/P0001  & ~n74271 ;
  assign n74273 = \u1_L1_reg[19]/P0001  & n74271 ;
  assign n74274 = ~n74272 & ~n74273 ;
  assign n74275 = n56245 & n56287 ;
  assign n74276 = n56258 & n56261 ;
  assign n74277 = ~n74275 & ~n74276 ;
  assign n74278 = ~n56219 & ~n74277 ;
  assign n74282 = n56247 & n56251 ;
  assign n74283 = n56274 & ~n74282 ;
  assign n74284 = ~n56265 & n74283 ;
  assign n74279 = ~n56219 & ~n56225 ;
  assign n74280 = n56238 & n56743 ;
  assign n74281 = ~n74279 & n74280 ;
  assign n74285 = ~n56754 & ~n74281 ;
  assign n74286 = n74284 & n74285 ;
  assign n74287 = ~n74278 & n74286 ;
  assign n74288 = n56262 & n56755 ;
  assign n74289 = ~n56267 & ~n56274 ;
  assign n74290 = ~n56284 & ~n56286 ;
  assign n74291 = n74289 & n74290 ;
  assign n74292 = ~n74288 & n74291 ;
  assign n74293 = ~n74287 & ~n74292 ;
  assign n74294 = ~n56238 & ~n56291 ;
  assign n74295 = ~n56288 & ~n74294 ;
  assign n74296 = ~n56245 & ~n74295 ;
  assign n74297 = ~n56254 & ~n56744 ;
  assign n74298 = ~n56274 & ~n74297 ;
  assign n74299 = ~n56219 & ~n74298 ;
  assign n74300 = ~n74296 & n74299 ;
  assign n74301 = n56219 & ~n56286 ;
  assign n74302 = ~n56268 & n74301 ;
  assign n74303 = ~n74300 & ~n74302 ;
  assign n74304 = ~n74293 & ~n74303 ;
  assign n74305 = ~\u0_L10_reg[26]/NET0131  & ~n74304 ;
  assign n74306 = \u0_L10_reg[26]/NET0131  & n74304 ;
  assign n74307 = ~n74305 & ~n74306 ;
  assign n74309 = ~n66274 & n67254 ;
  assign n74310 = ~n66268 & ~n74309 ;
  assign n74311 = n66288 & ~n74310 ;
  assign n74312 = ~n66288 & n66328 ;
  assign n74308 = n66313 & ~n66316 ;
  assign n74313 = n66255 & ~n74308 ;
  assign n74314 = ~n74312 & n74313 ;
  assign n74315 = ~n74311 & n74314 ;
  assign n74319 = ~n66298 & ~n66321 ;
  assign n74320 = n66290 & ~n74319 ;
  assign n74316 = ~n66267 & n67268 ;
  assign n74323 = ~n66255 & ~n74316 ;
  assign n74324 = ~n74320 & n74323 ;
  assign n74317 = ~n66317 & n67267 ;
  assign n74318 = ~n66288 & ~n74317 ;
  assign n74321 = n66291 & ~n67255 ;
  assign n74322 = n66322 & n74321 ;
  assign n74325 = ~n74318 & ~n74322 ;
  assign n74326 = n74324 & n74325 ;
  assign n74327 = ~n74315 & ~n74326 ;
  assign n74328 = \u0_L3_reg[12]/NET0131  & n74327 ;
  assign n74329 = ~\u0_L3_reg[12]/NET0131  & ~n74327 ;
  assign n74330 = ~n74328 & ~n74329 ;
  assign n74331 = ~n66350 & ~n66370 ;
  assign n74332 = ~n67193 & ~n74331 ;
  assign n74333 = n66377 & ~n74332 ;
  assign n74334 = n66420 & ~n74331 ;
  assign n74335 = n66400 & ~n66406 ;
  assign n74336 = ~n67208 & n74335 ;
  assign n74337 = ~n74334 & n74336 ;
  assign n74338 = ~n74333 & n74337 ;
  assign n74339 = n66357 & ~n66369 ;
  assign n74340 = n66363 & ~n74339 ;
  assign n74341 = ~n67592 & ~n74340 ;
  assign n74342 = ~n66377 & ~n74341 ;
  assign n74343 = ~n66369 & n66426 ;
  assign n74344 = ~n66385 & ~n74343 ;
  assign n74345 = n66363 & ~n74344 ;
  assign n74346 = n66377 & ~n67203 ;
  assign n74347 = ~n74345 & n74346 ;
  assign n74348 = ~n74342 & ~n74347 ;
  assign n74349 = ~n66400 & ~n66409 ;
  assign n74350 = ~n66427 & n74349 ;
  assign n74351 = ~n74348 & n74350 ;
  assign n74352 = ~n74338 & ~n74351 ;
  assign n74353 = \u0_L3_reg[17]/NET0131  & ~n74352 ;
  assign n74354 = ~\u0_L3_reg[17]/NET0131  & n74352 ;
  assign n74355 = ~n74353 & ~n74354 ;
  assign n74369 = n23141 & ~n23469 ;
  assign n74370 = ~n23473 & n74369 ;
  assign n74368 = ~n23102 & n23156 ;
  assign n74371 = ~n23464 & ~n23471 ;
  assign n74372 = ~n74368 & n74371 ;
  assign n74373 = ~n74370 & n74372 ;
  assign n74374 = n23134 & ~n74373 ;
  assign n74359 = ~n23151 & ~n23449 ;
  assign n74360 = n23134 & ~n74359 ;
  assign n74356 = ~n23118 & n23212 ;
  assign n74357 = n23134 & ~n23143 ;
  assign n74358 = n23219 & ~n74357 ;
  assign n74361 = ~n23473 & ~n74358 ;
  assign n74362 = ~n74356 & n74361 ;
  assign n74363 = ~n74360 & n74362 ;
  assign n74364 = ~n23141 & ~n74363 ;
  assign n74365 = n23111 & n23155 ;
  assign n74366 = ~n23166 & ~n74365 ;
  assign n74367 = n23141 & ~n74366 ;
  assign n74375 = ~n23474 & ~n74367 ;
  assign n74376 = ~n74364 & n74375 ;
  assign n74377 = ~n74374 & n74376 ;
  assign n74378 = \u2_L2_reg[5]/NET0131  & ~n74377 ;
  assign n74379 = ~\u2_L2_reg[5]/NET0131  & n74377 ;
  assign n74380 = ~n74378 & ~n74379 ;
  assign n74383 = ~n34695 & ~n35668 ;
  assign n74384 = n35954 & n74383 ;
  assign n74381 = n34695 & n35660 ;
  assign n74382 = n34701 & n35656 ;
  assign n74385 = ~n74381 & ~n74382 ;
  assign n74386 = ~n74384 & n74385 ;
  assign n74387 = ~n34747 & ~n74386 ;
  assign n74388 = ~n34701 & n34753 ;
  assign n74389 = ~n34750 & ~n74388 ;
  assign n74390 = n35652 & ~n74389 ;
  assign n74391 = ~n34708 & ~n34772 ;
  assign n74392 = ~n35680 & ~n74391 ;
  assign n74393 = n34695 & ~n74392 ;
  assign n74394 = ~n34695 & ~n34729 ;
  assign n74395 = ~n74391 & n74394 ;
  assign n74396 = ~n35672 & ~n35949 ;
  assign n74397 = ~n74395 & n74396 ;
  assign n74398 = ~n74393 & n74397 ;
  assign n74399 = n34747 & ~n74398 ;
  assign n74400 = ~n74390 & ~n74399 ;
  assign n74401 = ~n74387 & n74400 ;
  assign n74402 = \u1_L9_reg[17]/NET0131  & n74401 ;
  assign n74403 = ~\u1_L9_reg[17]/NET0131  & ~n74401 ;
  assign n74404 = ~n74402 & ~n74403 ;
  assign n74419 = n59579 & ~n59622 ;
  assign n74420 = ~n59617 & n74419 ;
  assign n74421 = ~n59636 & ~n59944 ;
  assign n74422 = n74420 & n74421 ;
  assign n74423 = ~n59579 & ~n59588 ;
  assign n74424 = ~n59935 & n74423 ;
  assign n74425 = ~n74422 & ~n74424 ;
  assign n74426 = n59552 & n59587 ;
  assign n74427 = ~n59938 & ~n74426 ;
  assign n74428 = ~n74425 & n74427 ;
  assign n74429 = n59604 & ~n74428 ;
  assign n74408 = ~n59565 & n59620 ;
  assign n74409 = ~n59597 & ~n74408 ;
  assign n74410 = ~n59552 & n59579 ;
  assign n74411 = ~n74409 & ~n74410 ;
  assign n74413 = ~n59559 & n59579 ;
  assign n74412 = ~n59579 & ~n59622 ;
  assign n74414 = ~n59572 & ~n74412 ;
  assign n74415 = ~n74413 & n74414 ;
  assign n74416 = ~n74411 & ~n74415 ;
  assign n74417 = ~n59604 & ~n74416 ;
  assign n74405 = ~n59558 & n60024 ;
  assign n74406 = n59939 & ~n74405 ;
  assign n74407 = n59579 & ~n74406 ;
  assign n74418 = n59596 & n59607 ;
  assign n74430 = ~n59618 & ~n74418 ;
  assign n74431 = ~n74407 & n74430 ;
  assign n74432 = ~n74417 & n74431 ;
  assign n74433 = ~n74429 & n74432 ;
  assign n74434 = \u0_L8_reg[25]/NET0131  & n74433 ;
  assign n74435 = ~\u0_L8_reg[25]/NET0131  & ~n74433 ;
  assign n74436 = ~n74434 & ~n74435 ;
  assign n74439 = n37322 & n37466 ;
  assign n74438 = ~n37386 & ~n37485 ;
  assign n74440 = ~n37388 & n74438 ;
  assign n74441 = ~n74439 & n74440 ;
  assign n74442 = ~n37341 & ~n74441 ;
  assign n74443 = ~n37341 & n37381 ;
  assign n74444 = ~n37373 & ~n74443 ;
  assign n74445 = ~n37322 & ~n74444 ;
  assign n74446 = ~n37377 & ~n74445 ;
  assign n74447 = ~n74442 & n74446 ;
  assign n74448 = n37362 & ~n74447 ;
  assign n74452 = ~n37342 & n74438 ;
  assign n74453 = n37322 & ~n37349 ;
  assign n74454 = ~n74452 & ~n74453 ;
  assign n74455 = ~n37348 & ~n37484 ;
  assign n74456 = n37322 & ~n37335 ;
  assign n74457 = ~n37485 & n74456 ;
  assign n74458 = ~n74455 & n74457 ;
  assign n74459 = ~n74454 & ~n74458 ;
  assign n74460 = ~n37362 & ~n74459 ;
  assign n74437 = ~n37322 & n37467 ;
  assign n74449 = ~n37348 & n37373 ;
  assign n74450 = ~n37379 & ~n74449 ;
  assign n74451 = n37322 & ~n74450 ;
  assign n74461 = ~n74437 & ~n74451 ;
  assign n74462 = ~n74460 & n74461 ;
  assign n74463 = ~n74448 & n74462 ;
  assign n74464 = ~\u1_L8_reg[16]/NET0131  & ~n74463 ;
  assign n74465 = \u1_L8_reg[16]/NET0131  & n74463 ;
  assign n74466 = ~n74464 & ~n74465 ;
  assign n74479 = ~n43834 & ~n44404 ;
  assign n74480 = ~n43849 & ~n74479 ;
  assign n74481 = n43799 & n44414 ;
  assign n74482 = ~n43872 & ~n74481 ;
  assign n74483 = ~n43812 & ~n74482 ;
  assign n74484 = ~n74480 & ~n74483 ;
  assign n74485 = ~n43806 & ~n74484 ;
  assign n74473 = n43806 & n43835 ;
  assign n74467 = ~n43812 & n43827 ;
  assign n74474 = ~n44396 & ~n74467 ;
  assign n74475 = ~n74473 & n74474 ;
  assign n74468 = ~n43853 & ~n43856 ;
  assign n74469 = n43812 & ~n74468 ;
  assign n74470 = n43831 & n43852 ;
  assign n74471 = ~n43858 & ~n74470 ;
  assign n74472 = ~n43806 & ~n74471 ;
  assign n74476 = ~n74469 & ~n74472 ;
  assign n74477 = n74475 & n74476 ;
  assign n74478 = n43849 & ~n74477 ;
  assign n74486 = ~n43854 & ~n44147 ;
  assign n74487 = n43806 & ~n74486 ;
  assign n74488 = n43799 & n43838 ;
  assign n74489 = ~n43852 & n74488 ;
  assign n74490 = ~n44146 & ~n74489 ;
  assign n74491 = n43855 & n74490 ;
  assign n74492 = ~n43849 & ~n74491 ;
  assign n74493 = ~n74487 & ~n74492 ;
  assign n74494 = ~n74478 & n74493 ;
  assign n74495 = ~n74485 & n74494 ;
  assign n74496 = ~\u1_L3_reg[26]/NET0131  & ~n74495 ;
  assign n74497 = \u1_L3_reg[26]/NET0131  & n74495 ;
  assign n74498 = ~n74496 & ~n74497 ;
  assign n74499 = n44059 & ~n44078 ;
  assign n74500 = ~n44568 & ~n74499 ;
  assign n74501 = n44046 & ~n74500 ;
  assign n74504 = ~n44086 & ~n44576 ;
  assign n74505 = ~n44101 & n74504 ;
  assign n74502 = n44078 & ~n44087 ;
  assign n74503 = n44554 & n74502 ;
  assign n74506 = ~n44119 & ~n74503 ;
  assign n74507 = n74505 & n74506 ;
  assign n74508 = ~n74501 & n74507 ;
  assign n74509 = ~n44071 & ~n44078 ;
  assign n74510 = ~n44317 & n74509 ;
  assign n74511 = ~n44066 & n44078 ;
  assign n74512 = ~n44094 & ~n44553 ;
  assign n74513 = n74511 & n74512 ;
  assign n74514 = ~n74510 & ~n74513 ;
  assign n74515 = n44046 & ~n44099 ;
  assign n74516 = n44569 & n74515 ;
  assign n74517 = n44086 & ~n44298 ;
  assign n74518 = ~n74516 & n74517 ;
  assign n74519 = ~n74514 & n74518 ;
  assign n74520 = ~n74508 & ~n74519 ;
  assign n74521 = n44078 & n44088 ;
  assign n74522 = n44086 & ~n44575 ;
  assign n74523 = ~n44046 & ~n44313 ;
  assign n74524 = n44577 & n74523 ;
  assign n74525 = ~n74522 & n74524 ;
  assign n74526 = ~n74521 & ~n74525 ;
  assign n74527 = ~n74520 & n74526 ;
  assign n74528 = ~\u1_L3_reg[21]/NET0131  & ~n74527 ;
  assign n74529 = \u1_L3_reg[21]/NET0131  & n74527 ;
  assign n74530 = ~n74528 & ~n74529 ;
  assign n74544 = n54819 & ~n54841 ;
  assign n74545 = ~n54835 & ~n74544 ;
  assign n74546 = ~n54840 & ~n74545 ;
  assign n74547 = ~n54806 & ~n74546 ;
  assign n74543 = n54858 & ~n54910 ;
  assign n74548 = ~n54948 & ~n74543 ;
  assign n74549 = ~n74547 & n74548 ;
  assign n74550 = ~n54850 & ~n74549 ;
  assign n74531 = n54872 & n54928 ;
  assign n74535 = ~n54857 & ~n74531 ;
  assign n74532 = n54842 & n54862 ;
  assign n74533 = n54876 & ~n54927 ;
  assign n74534 = ~n54872 & n74533 ;
  assign n74536 = ~n74532 & ~n74534 ;
  assign n74537 = n74535 & n74536 ;
  assign n74538 = n54850 & ~n74537 ;
  assign n74540 = ~n54838 & ~n54875 ;
  assign n74539 = ~n54837 & ~n54882 ;
  assign n74541 = ~n54812 & ~n74539 ;
  assign n74542 = ~n74540 & n74541 ;
  assign n74551 = ~n74538 & ~n74542 ;
  assign n74552 = ~n74550 & n74551 ;
  assign n74553 = ~\u0_L11_reg[26]/NET0131  & ~n74552 ;
  assign n74554 = \u0_L11_reg[26]/NET0131  & n74552 ;
  assign n74555 = ~n74553 & ~n74554 ;
  assign n74556 = ~n6226 & n6252 ;
  assign n74557 = ~n6229 & ~n6250 ;
  assign n74558 = ~n74556 & n74557 ;
  assign n74559 = n6198 & ~n74558 ;
  assign n74560 = ~n6210 & n6570 ;
  assign n74561 = ~n74559 & ~n74560 ;
  assign n74562 = ~n6244 & ~n74561 ;
  assign n74573 = n6564 & n6587 ;
  assign n74565 = n6227 & n6268 ;
  assign n74574 = ~n6563 & ~n74565 ;
  assign n74575 = ~n74573 & n74574 ;
  assign n74572 = n6198 & n6247 ;
  assign n74576 = ~n6569 & ~n74572 ;
  assign n74577 = n74575 & n74576 ;
  assign n74578 = n6244 & ~n74577 ;
  assign n74563 = ~n6236 & ~n6564 ;
  assign n74564 = ~n6268 & ~n74563 ;
  assign n74566 = ~n6198 & ~n74565 ;
  assign n74567 = ~n6248 & n74566 ;
  assign n74568 = ~n74564 & n74567 ;
  assign n74569 = n6198 & ~n6237 ;
  assign n74570 = ~n6577 & n74569 ;
  assign n74571 = ~n74568 & ~n74570 ;
  assign n74579 = ~n6198 & ~n6210 ;
  assign n74580 = n6217 & ~n6244 ;
  assign n74581 = n74579 & n74580 ;
  assign n74582 = ~n74571 & ~n74581 ;
  assign n74583 = ~n74578 & n74582 ;
  assign n74584 = ~n74562 & n74583 ;
  assign n74585 = \u2_L13_reg[15]/NET0131  & n74584 ;
  assign n74586 = ~\u2_L13_reg[15]/NET0131  & ~n74584 ;
  assign n74587 = ~n74585 & ~n74586 ;
  assign n74597 = ~n31782 & ~n31796 ;
  assign n74598 = ~n32641 & ~n74597 ;
  assign n74599 = n31768 & ~n74598 ;
  assign n74600 = n31829 & ~n74597 ;
  assign n74601 = ~n31844 & ~n33094 ;
  assign n74602 = ~n74600 & n74601 ;
  assign n74603 = ~n74599 & n74602 ;
  assign n74604 = n31813 & ~n74603 ;
  assign n74589 = ~n31823 & ~n32635 ;
  assign n74590 = ~n31768 & ~n74589 ;
  assign n74588 = n31827 & n32629 ;
  assign n74591 = n31832 & ~n33077 ;
  assign n74592 = ~n74588 & ~n74591 ;
  assign n74593 = ~n74590 & n74592 ;
  assign n74594 = ~n31813 & ~n74593 ;
  assign n74595 = ~n31834 & ~n33080 ;
  assign n74596 = n31820 & ~n74595 ;
  assign n74605 = ~n74594 & ~n74596 ;
  assign n74606 = ~n74604 & n74605 ;
  assign n74607 = ~\u1_L11_reg[17]/NET0131  & ~n74606 ;
  assign n74608 = \u1_L11_reg[17]/NET0131  & n74606 ;
  assign n74609 = ~n74607 & ~n74608 ;
  assign n74615 = ~n36783 & ~n36796 ;
  assign n74624 = n36768 & ~n74615 ;
  assign n74625 = n36774 & ~n74624 ;
  assign n74626 = ~n37226 & ~n74625 ;
  assign n74627 = n36790 & ~n74626 ;
  assign n74612 = n36768 & ~n36790 ;
  assign n74623 = n36783 & n74612 ;
  assign n74628 = n36783 & ~n36798 ;
  assign n74629 = ~n36768 & ~n36808 ;
  assign n74630 = ~n74628 & n74629 ;
  assign n74631 = ~n74623 & ~n74630 ;
  assign n74632 = ~n74627 & n74631 ;
  assign n74633 = n36819 & ~n74632 ;
  assign n74616 = ~n37214 & ~n74615 ;
  assign n74617 = ~n36776 & ~n36790 ;
  assign n74618 = ~n74616 & n74617 ;
  assign n74610 = ~n36808 & ~n37235 ;
  assign n74611 = n36768 & ~n74610 ;
  assign n74613 = n36774 & n36826 ;
  assign n74614 = ~n74612 & n74613 ;
  assign n74619 = ~n37225 & ~n74614 ;
  assign n74620 = ~n74611 & n74619 ;
  assign n74621 = ~n74618 & n74620 ;
  assign n74622 = ~n36819 & ~n74621 ;
  assign n74635 = ~n36776 & ~n36798 ;
  assign n74636 = ~n36824 & ~n37213 ;
  assign n74637 = ~n74635 & n74636 ;
  assign n74638 = ~n37218 & ~n74637 ;
  assign n74639 = ~n36790 & ~n74638 ;
  assign n74634 = n37213 & n37561 ;
  assign n74640 = ~n37228 & ~n74634 ;
  assign n74641 = ~n74639 & n74640 ;
  assign n74642 = ~n74622 & n74641 ;
  assign n74643 = ~n74633 & n74642 ;
  assign n74644 = ~\u1_L8_reg[31]/NET0131  & ~n74643 ;
  assign n74645 = \u1_L8_reg[31]/NET0131  & n74643 ;
  assign n74646 = ~n74644 & ~n74645 ;
  assign n74648 = n39917 & ~n39931 ;
  assign n74649 = n39972 & ~n74648 ;
  assign n74650 = n39940 & ~n39981 ;
  assign n74651 = ~n40506 & n74650 ;
  assign n74652 = ~n74649 & ~n74651 ;
  assign n74653 = n39947 & ~n40523 ;
  assign n74654 = n40040 & n74653 ;
  assign n74655 = ~n74652 & n74654 ;
  assign n74657 = ~n39910 & ~n39948 ;
  assign n74656 = n39916 & ~n39955 ;
  assign n74658 = ~n39961 & ~n74656 ;
  assign n74659 = ~n74657 & n74658 ;
  assign n74660 = ~n39982 & n40031 ;
  assign n74661 = ~n74659 & n74660 ;
  assign n74662 = ~n74655 & ~n74661 ;
  assign n74647 = n39931 & n40057 ;
  assign n74663 = ~n39933 & ~n74647 ;
  assign n74664 = ~n74662 & n74663 ;
  assign n74668 = ~n39916 & n39951 ;
  assign n74665 = ~n39932 & ~n39962 ;
  assign n74666 = ~n40505 & n74665 ;
  assign n74667 = ~n39981 & n74666 ;
  assign n74669 = n39940 & ~n39947 ;
  assign n74670 = ~n74667 & n74669 ;
  assign n74671 = ~n74668 & n74670 ;
  assign n74672 = ~n74664 & ~n74671 ;
  assign n74673 = ~\u1_L6_reg[13]/NET0131  & ~n74672 ;
  assign n74674 = \u1_L6_reg[13]/NET0131  & n74672 ;
  assign n74675 = ~n74673 & ~n74674 ;
  assign n74678 = n6310 & n6329 ;
  assign n74679 = ~n6301 & n74678 ;
  assign n74677 = ~n6304 & n6342 ;
  assign n74680 = n6324 & ~n74677 ;
  assign n74681 = ~n74679 & n74680 ;
  assign n74682 = ~n6619 & n74681 ;
  assign n74683 = n6304 & ~n6310 ;
  assign n74684 = ~n6324 & ~n6328 ;
  assign n74685 = ~n74683 & n74684 ;
  assign n74686 = ~n74682 & ~n74685 ;
  assign n74687 = n6310 & n6354 ;
  assign n74688 = n6289 & ~n6328 ;
  assign n74676 = n6326 & n6356 ;
  assign n74689 = ~n6543 & ~n74676 ;
  assign n74690 = n74688 & n74689 ;
  assign n74691 = ~n74687 & n74690 ;
  assign n74692 = ~n74686 & n74691 ;
  assign n74693 = ~n6603 & ~n74678 ;
  assign n74694 = n74684 & n74693 ;
  assign n74695 = ~n6346 & ~n6602 ;
  assign n74696 = n6301 & ~n74695 ;
  assign n74697 = ~n6353 & ~n74696 ;
  assign n74698 = n74681 & n74697 ;
  assign n74699 = ~n74694 & ~n74698 ;
  assign n74700 = ~n6289 & ~n6628 ;
  assign n74701 = n6363 & n74700 ;
  assign n74702 = ~n74699 & n74701 ;
  assign n74703 = ~n74692 & ~n74702 ;
  assign n74704 = ~\u2_L13_reg[20]/NET0131  & n74703 ;
  assign n74705 = \u2_L13_reg[20]/NET0131  & ~n74703 ;
  assign n74706 = ~n74704 & ~n74705 ;
  assign n74721 = ~n51073 & n51104 ;
  assign n74723 = n51092 & n74721 ;
  assign n74718 = ~n51079 & n51092 ;
  assign n74722 = ~n74718 & ~n74721 ;
  assign n74724 = n51086 & ~n74722 ;
  assign n74725 = ~n74723 & n74724 ;
  assign n74708 = ~n51086 & ~n51104 ;
  assign n74719 = ~n51106 & n74708 ;
  assign n74720 = ~n74718 & n74719 ;
  assign n74726 = ~n51067 & ~n74720 ;
  assign n74727 = ~n74725 & n74726 ;
  assign n74728 = ~n51079 & n51121 ;
  assign n74729 = ~n51104 & ~n51107 ;
  assign n74730 = ~n74728 & n74729 ;
  assign n74731 = ~n51116 & ~n74718 ;
  assign n74732 = ~n51073 & ~n74731 ;
  assign n74733 = n51086 & n51106 ;
  assign n74734 = ~n51079 & ~n51086 ;
  assign n74735 = n51104 & ~n74734 ;
  assign n74736 = ~n74733 & n74735 ;
  assign n74737 = ~n74732 & n74736 ;
  assign n74738 = ~n74730 & ~n74737 ;
  assign n74712 = n51092 & n51095 ;
  assign n74707 = n51073 & n51121 ;
  assign n74739 = n51067 & ~n74707 ;
  assign n74740 = ~n74712 & n74739 ;
  assign n74741 = ~n74738 & n74740 ;
  assign n74742 = ~n74727 & ~n74741 ;
  assign n74709 = n51092 & n74708 ;
  assign n74710 = ~n74707 & ~n74709 ;
  assign n74711 = n51079 & ~n74710 ;
  assign n74713 = n51092 & n51124 ;
  assign n74714 = ~n74712 & ~n74713 ;
  assign n74715 = n51096 & n51116 ;
  assign n74716 = n74714 & ~n74715 ;
  assign n74717 = n51104 & ~n74716 ;
  assign n74743 = ~n74711 & ~n74717 ;
  assign n74744 = ~n74742 & n74743 ;
  assign n74745 = \u0_L14_reg[25]/P0001  & n74744 ;
  assign n74746 = ~\u0_L14_reg[25]/P0001  & ~n74744 ;
  assign n74747 = ~n74745 & ~n74746 ;
  assign n74800 = decrypt_pad & ~\u0_uk_K_r14_reg[40]/NET0131  ;
  assign n74801 = ~decrypt_pad & ~\u0_uk_K_r14_reg[33]/NET0131  ;
  assign n74802 = ~n74800 & ~n74801 ;
  assign n74803 = \u0_R14_reg[16]/NET0131  & ~n74802 ;
  assign n74804 = ~\u0_R14_reg[16]/NET0131  & n74802 ;
  assign n74805 = ~n74803 & ~n74804 ;
  assign n74748 = decrypt_pad & ~\u0_uk_K_r14_reg[4]/NET0131  ;
  assign n74749 = ~decrypt_pad & ~\u0_uk_K_r14_reg[54]/NET0131  ;
  assign n74750 = ~n74748 & ~n74749 ;
  assign n74751 = \u0_R14_reg[12]/NET0131  & ~n74750 ;
  assign n74752 = ~\u0_R14_reg[12]/NET0131  & n74750 ;
  assign n74753 = ~n74751 & ~n74752 ;
  assign n74782 = decrypt_pad & ~\u0_uk_K_r14_reg[32]/NET0131  ;
  assign n74783 = ~decrypt_pad & ~\u0_uk_K_r14_reg[25]/NET0131  ;
  assign n74784 = ~n74782 & ~n74783 ;
  assign n74785 = \u0_R14_reg[15]/NET0131  & ~n74784 ;
  assign n74786 = ~\u0_R14_reg[15]/NET0131  & n74784 ;
  assign n74787 = ~n74785 & ~n74786 ;
  assign n74761 = decrypt_pad & ~\u0_uk_K_r14_reg[24]/NET0131  ;
  assign n74762 = ~decrypt_pad & ~\u0_uk_K_r14_reg[17]/NET0131  ;
  assign n74763 = ~n74761 & ~n74762 ;
  assign n74764 = \u0_R14_reg[14]/NET0131  & ~n74763 ;
  assign n74765 = ~\u0_R14_reg[14]/NET0131  & n74763 ;
  assign n74766 = ~n74764 & ~n74765 ;
  assign n74768 = decrypt_pad & ~\u0_uk_K_r14_reg[55]/NET0131  ;
  assign n74769 = ~decrypt_pad & ~\u0_uk_K_r14_reg[48]/NET0131  ;
  assign n74770 = ~n74768 & ~n74769 ;
  assign n74771 = \u0_R14_reg[13]/NET0131  & ~n74770 ;
  assign n74772 = ~\u0_R14_reg[13]/NET0131  & n74770 ;
  assign n74773 = ~n74771 & ~n74772 ;
  assign n74775 = n74766 & ~n74773 ;
  assign n74754 = decrypt_pad & ~\u0_uk_K_r14_reg[20]/NET0131  ;
  assign n74755 = ~decrypt_pad & ~\u0_uk_K_r14_reg[13]/NET0131  ;
  assign n74756 = ~n74754 & ~n74755 ;
  assign n74757 = \u0_R14_reg[17]/NET0131  & ~n74756 ;
  assign n74758 = ~\u0_R14_reg[17]/NET0131  & n74756 ;
  assign n74759 = ~n74757 & ~n74758 ;
  assign n74811 = ~n74759 & ~n74773 ;
  assign n74812 = ~n74775 & ~n74811 ;
  assign n74813 = n74787 & ~n74812 ;
  assign n74779 = ~n74766 & n74773 ;
  assign n74814 = ~n74766 & ~n74787 ;
  assign n74815 = n74759 & n74814 ;
  assign n74816 = ~n74779 & ~n74815 ;
  assign n74817 = ~n74813 & n74816 ;
  assign n74818 = n74753 & ~n74817 ;
  assign n74792 = ~n74753 & ~n74759 ;
  assign n74793 = n74773 & n74792 ;
  assign n74807 = n74766 & n74793 ;
  assign n74808 = ~n74766 & n74792 ;
  assign n74809 = ~n74773 & n74808 ;
  assign n74810 = ~n74807 & ~n74809 ;
  assign n74819 = ~n74773 & n74792 ;
  assign n74820 = ~n74787 & n74819 ;
  assign n74788 = ~n74753 & n74759 ;
  assign n74821 = n74787 & n74788 ;
  assign n74822 = ~n74766 & n74821 ;
  assign n74823 = ~n74820 & ~n74822 ;
  assign n74824 = n74810 & n74823 ;
  assign n74825 = ~n74818 & n74824 ;
  assign n74826 = ~n74805 & ~n74825 ;
  assign n74760 = n74753 & n74759 ;
  assign n74767 = n74760 & n74766 ;
  assign n74774 = n74767 & n74773 ;
  assign n74776 = ~n74753 & n74775 ;
  assign n74777 = n74759 & n74776 ;
  assign n74778 = ~n74774 & ~n74777 ;
  assign n74780 = n74753 & ~n74759 ;
  assign n74781 = ~n74779 & n74780 ;
  assign n74789 = n74779 & n74788 ;
  assign n74790 = ~n74787 & ~n74789 ;
  assign n74791 = ~n74781 & n74790 ;
  assign n74794 = n74760 & ~n74773 ;
  assign n74795 = ~n74766 & n74794 ;
  assign n74796 = n74787 & ~n74793 ;
  assign n74797 = ~n74795 & n74796 ;
  assign n74798 = ~n74791 & ~n74797 ;
  assign n74799 = n74778 & ~n74798 ;
  assign n74806 = ~n74799 & n74805 ;
  assign n74830 = n74778 & ~n74809 ;
  assign n74831 = ~n74787 & ~n74830 ;
  assign n74827 = n74773 & n74787 ;
  assign n74828 = n74766 & n74827 ;
  assign n74829 = ~n74753 & n74828 ;
  assign n74832 = n74780 & n74827 ;
  assign n74833 = ~n74766 & n74832 ;
  assign n74834 = ~n74829 & ~n74833 ;
  assign n74835 = ~n74831 & n74834 ;
  assign n74836 = ~n74806 & n74835 ;
  assign n74837 = ~n74826 & n74836 ;
  assign n74838 = \u0_L14_reg[10]/P0001  & n74837 ;
  assign n74839 = ~\u0_L14_reg[10]/P0001  & ~n74837 ;
  assign n74840 = ~n74838 & ~n74839 ;
  assign n74843 = ~n51227 & ~n51239 ;
  assign n74844 = ~n51215 & ~n74843 ;
  assign n74845 = ~n51223 & ~n51238 ;
  assign n74846 = ~n51188 & n51219 ;
  assign n74847 = n74845 & n74846 ;
  assign n74848 = ~n51181 & ~n51187 ;
  assign n74849 = ~n51194 & ~n51201 ;
  assign n74850 = n74848 & n74849 ;
  assign n74841 = n51194 & n51201 ;
  assign n74842 = ~n51244 & n74841 ;
  assign n74851 = n51208 & ~n74842 ;
  assign n74852 = ~n74850 & n74851 ;
  assign n74853 = ~n74847 & n74852 ;
  assign n74854 = ~n74844 & n74853 ;
  assign n74856 = n51215 & ~n74845 ;
  assign n74857 = ~n51235 & ~n74856 ;
  assign n74858 = ~n51201 & ~n74857 ;
  assign n74855 = n51201 & n51217 ;
  assign n74864 = ~n51208 & ~n74855 ;
  assign n74859 = ~n51215 & ~n51236 ;
  assign n74860 = n51187 & ~n51201 ;
  assign n74861 = n51218 & n74860 ;
  assign n74862 = n51195 & n51215 ;
  assign n74863 = ~n74861 & ~n74862 ;
  assign n74865 = ~n74859 & n74863 ;
  assign n74866 = n74864 & n74865 ;
  assign n74867 = ~n74858 & n74866 ;
  assign n74868 = ~n74854 & ~n74867 ;
  assign n74869 = n51188 & n51218 ;
  assign n74870 = ~n51201 & ~n74869 ;
  assign n74871 = ~n74862 & n74870 ;
  assign n74872 = n51194 & n51240 ;
  assign n74873 = n51201 & ~n74872 ;
  assign n74874 = ~n51246 & n74873 ;
  assign n74875 = ~n74871 & ~n74874 ;
  assign n74876 = ~n74868 & ~n74875 ;
  assign n74877 = \u0_L14_reg[2]/P0001  & n74876 ;
  assign n74878 = ~\u0_L14_reg[2]/P0001  & ~n74876 ;
  assign n74879 = ~n74877 & ~n74878 ;
  assign n74880 = decrypt_pad & ~\u0_uk_K_r14_reg[9]/NET0131  ;
  assign n74881 = ~decrypt_pad & ~\u0_uk_K_r14_reg[2]/NET0131  ;
  assign n74882 = ~n74880 & ~n74881 ;
  assign n74883 = \u0_R14_reg[23]/NET0131  & ~n74882 ;
  assign n74884 = ~\u0_R14_reg[23]/NET0131  & n74882 ;
  assign n74885 = ~n74883 & ~n74884 ;
  assign n74899 = decrypt_pad & ~\u0_uk_K_r14_reg[29]/NET0131  ;
  assign n74900 = ~decrypt_pad & ~\u0_uk_K_r14_reg[22]/NET0131  ;
  assign n74901 = ~n74899 & ~n74900 ;
  assign n74902 = \u0_R14_reg[21]/NET0131  & ~n74901 ;
  assign n74903 = ~\u0_R14_reg[21]/NET0131  & n74901 ;
  assign n74904 = ~n74902 & ~n74903 ;
  assign n74886 = decrypt_pad & ~\u0_uk_K_r14_reg[14]/NET0131  ;
  assign n74887 = ~decrypt_pad & ~\u0_uk_K_r14_reg[7]/NET0131  ;
  assign n74888 = ~n74886 & ~n74887 ;
  assign n74889 = \u0_R14_reg[20]/NET0131  & ~n74888 ;
  assign n74890 = ~\u0_R14_reg[20]/NET0131  & n74888 ;
  assign n74891 = ~n74889 & ~n74890 ;
  assign n74892 = decrypt_pad & ~\u0_uk_K_r14_reg[30]/NET0131  ;
  assign n74893 = ~decrypt_pad & ~\u0_uk_K_r14_reg[23]/NET0131  ;
  assign n74894 = ~n74892 & ~n74893 ;
  assign n74895 = \u0_R14_reg[25]/NET0131  & ~n74894 ;
  assign n74896 = ~\u0_R14_reg[25]/NET0131  & n74894 ;
  assign n74897 = ~n74895 & ~n74896 ;
  assign n74916 = ~n74891 & ~n74897 ;
  assign n74922 = n74904 & n74916 ;
  assign n74905 = decrypt_pad & ~\u0_uk_K_r14_reg[51]/NET0131  ;
  assign n74906 = ~decrypt_pad & ~\u0_uk_K_r14_reg[44]/NET0131  ;
  assign n74907 = ~n74905 & ~n74906 ;
  assign n74908 = \u0_R14_reg[22]/P0001  & ~n74907 ;
  assign n74909 = ~\u0_R14_reg[22]/P0001  & n74907 ;
  assign n74910 = ~n74908 & ~n74909 ;
  assign n74923 = n74904 & ~n74910 ;
  assign n74924 = n74891 & ~n74923 ;
  assign n74925 = ~n74922 & ~n74924 ;
  assign n74926 = n74885 & ~n74925 ;
  assign n74917 = ~n74904 & n74916 ;
  assign n74918 = ~n74891 & n74897 ;
  assign n74919 = n74904 & n74918 ;
  assign n74920 = ~n74917 & ~n74919 ;
  assign n74921 = ~n74885 & ~n74920 ;
  assign n74898 = n74891 & n74897 ;
  assign n74914 = n74898 & n74904 ;
  assign n74915 = n74910 & n74914 ;
  assign n74927 = decrypt_pad & ~\u0_uk_K_r14_reg[35]/P0001  ;
  assign n74928 = ~decrypt_pad & ~\u0_uk_K_r14_reg[28]/NET0131  ;
  assign n74929 = ~n74927 & ~n74928 ;
  assign n74930 = \u0_R14_reg[24]/NET0131  & ~n74929 ;
  assign n74931 = ~\u0_R14_reg[24]/NET0131  & n74929 ;
  assign n74932 = ~n74930 & ~n74931 ;
  assign n74933 = ~n74915 & ~n74932 ;
  assign n74934 = ~n74921 & n74933 ;
  assign n74935 = ~n74926 & n74934 ;
  assign n74937 = ~n74904 & n74918 ;
  assign n74940 = n74891 & n74923 ;
  assign n74941 = ~n74937 & ~n74940 ;
  assign n74942 = n74885 & ~n74941 ;
  assign n74936 = n74910 & n74917 ;
  assign n74938 = ~n74910 & n74937 ;
  assign n74939 = ~n74936 & ~n74938 ;
  assign n74943 = ~n74897 & n74923 ;
  assign n74949 = n74932 & ~n74943 ;
  assign n74944 = n74891 & ~n74904 ;
  assign n74945 = ~n74885 & n74944 ;
  assign n74946 = n74897 & n74904 ;
  assign n74947 = ~n74891 & n74910 ;
  assign n74948 = n74946 & n74947 ;
  assign n74950 = ~n74945 & ~n74948 ;
  assign n74951 = n74949 & n74950 ;
  assign n74952 = n74939 & n74951 ;
  assign n74953 = ~n74942 & n74952 ;
  assign n74954 = ~n74935 & ~n74953 ;
  assign n74911 = ~n74904 & ~n74910 ;
  assign n74912 = n74898 & n74911 ;
  assign n74913 = ~n74885 & n74912 ;
  assign n74955 = n74885 & n74937 ;
  assign n74956 = ~n74910 & n74955 ;
  assign n74957 = ~n74885 & ~n74910 ;
  assign n74958 = n74891 & ~n74897 ;
  assign n74959 = n74904 & n74958 ;
  assign n74960 = n74957 & n74959 ;
  assign n74961 = ~n74956 & ~n74960 ;
  assign n74962 = ~n74913 & n74961 ;
  assign n74963 = ~n74954 & n74962 ;
  assign n74964 = \u0_L14_reg[19]/P0001  & n74963 ;
  assign n74965 = ~\u0_L14_reg[19]/P0001  & ~n74963 ;
  assign n74966 = ~n74964 & ~n74965 ;
  assign n74968 = ~n74910 & ~n74946 ;
  assign n74967 = n74904 & n74947 ;
  assign n74969 = ~n74898 & ~n74967 ;
  assign n74970 = ~n74968 & n74969 ;
  assign n74971 = ~n74885 & ~n74912 ;
  assign n74972 = ~n74970 & n74971 ;
  assign n74973 = ~n74904 & n74958 ;
  assign n74974 = ~n74910 & n74973 ;
  assign n74975 = n74885 & ~n74914 ;
  assign n74976 = ~n74967 & n74975 ;
  assign n74977 = ~n74974 & n74976 ;
  assign n74978 = ~n74972 & ~n74977 ;
  assign n74979 = n74932 & ~n74978 ;
  assign n74980 = n74891 & n74943 ;
  assign n74990 = ~n74932 & ~n74955 ;
  assign n74991 = ~n74980 & n74990 ;
  assign n74982 = n74910 & n74944 ;
  assign n74987 = ~n74891 & ~n74910 ;
  assign n74988 = ~n74982 & ~n74987 ;
  assign n74989 = n74885 & ~n74988 ;
  assign n74981 = n74957 & n74958 ;
  assign n74983 = n74897 & n74982 ;
  assign n74984 = ~n74981 & ~n74983 ;
  assign n74985 = ~n74940 & ~n74967 ;
  assign n74986 = ~n74885 & ~n74985 ;
  assign n74992 = n74984 & ~n74986 ;
  assign n74993 = ~n74989 & n74992 ;
  assign n74994 = n74991 & n74993 ;
  assign n74995 = ~n74979 & ~n74994 ;
  assign n74997 = n74898 & n74910 ;
  assign n74998 = ~n74891 & n74943 ;
  assign n74999 = ~n74997 & ~n74998 ;
  assign n75000 = n74885 & ~n74999 ;
  assign n74996 = n74917 & n74957 ;
  assign n75001 = n74961 & ~n74996 ;
  assign n75002 = ~n75000 & n75001 ;
  assign n75003 = ~n74995 & n75002 ;
  assign n75004 = ~\u0_L14_reg[11]/P0001  & n75003 ;
  assign n75005 = \u0_L14_reg[11]/P0001  & ~n75003 ;
  assign n75006 = ~n75004 & ~n75005 ;
  assign n75008 = ~n51215 & n74848 ;
  assign n75009 = ~n51195 & ~n75008 ;
  assign n75007 = ~n51201 & ~n51245 ;
  assign n75010 = ~n51225 & n75007 ;
  assign n75011 = n75009 & n75010 ;
  assign n75012 = n51215 & n51250 ;
  assign n75013 = n51201 & n74843 ;
  assign n75014 = ~n75012 & n75013 ;
  assign n75015 = ~n75011 & ~n75014 ;
  assign n75018 = n51188 & n51215 ;
  assign n75019 = ~n51194 & n75018 ;
  assign n75016 = ~n51194 & n51241 ;
  assign n75017 = n51201 & n51240 ;
  assign n75020 = n51208 & ~n75017 ;
  assign n75021 = ~n75016 & n75020 ;
  assign n75022 = ~n75019 & n75021 ;
  assign n75023 = ~n75015 & n75022 ;
  assign n75024 = n51201 & n75009 ;
  assign n75025 = ~n51215 & n51238 ;
  assign n75026 = ~n51223 & ~n51235 ;
  assign n75027 = ~n75025 & n75026 ;
  assign n75028 = n75007 & n75027 ;
  assign n75029 = ~n75024 & ~n75028 ;
  assign n75030 = ~n51188 & ~n51194 ;
  assign n75031 = n51215 & ~n51238 ;
  assign n75032 = n75030 & n75031 ;
  assign n75033 = ~n51208 & ~n51225 ;
  assign n75034 = ~n75032 & n75033 ;
  assign n75035 = ~n75029 & n75034 ;
  assign n75036 = ~n75023 & ~n75035 ;
  assign n75037 = \u0_L14_reg[28]/P0001  & ~n75036 ;
  assign n75038 = ~\u0_L14_reg[28]/P0001  & n75036 ;
  assign n75039 = ~n75037 & ~n75038 ;
  assign n75048 = ~n74805 & ~n74829 ;
  assign n75040 = n74787 & n74819 ;
  assign n75045 = ~n74766 & ~n74773 ;
  assign n75046 = ~n74827 & ~n75045 ;
  assign n75047 = n74760 & ~n75046 ;
  assign n75049 = ~n75040 & ~n75047 ;
  assign n75050 = n75048 & n75049 ;
  assign n75041 = n74759 & ~n74773 ;
  assign n75042 = n74766 & n74780 ;
  assign n75043 = ~n75041 & ~n75042 ;
  assign n75044 = ~n74787 & ~n75043 ;
  assign n75051 = n74810 & ~n75044 ;
  assign n75052 = n75050 & n75051 ;
  assign n75060 = ~n74774 & n74805 ;
  assign n75054 = ~n74773 & n74821 ;
  assign n75055 = ~n74789 & ~n74832 ;
  assign n75061 = ~n75054 & n75055 ;
  assign n75062 = n75060 & n75061 ;
  assign n75053 = n74766 & n74820 ;
  assign n75056 = ~n74753 & n74779 ;
  assign n75057 = n74753 & n75045 ;
  assign n75058 = ~n75056 & ~n75057 ;
  assign n75059 = ~n74787 & ~n75058 ;
  assign n75063 = ~n75053 & ~n75059 ;
  assign n75064 = n75062 & n75063 ;
  assign n75065 = ~n75052 & ~n75064 ;
  assign n75066 = n74775 & n74780 ;
  assign n75067 = n74787 & ~n75066 ;
  assign n75068 = ~n74809 & n75067 ;
  assign n75069 = ~n74790 & ~n75068 ;
  assign n75070 = ~n74833 & ~n75069 ;
  assign n75071 = ~n75065 & n75070 ;
  assign n75072 = ~\u0_L14_reg[20]/P0001  & ~n75071 ;
  assign n75073 = \u0_L14_reg[20]/P0001  & n75071 ;
  assign n75074 = ~n75072 & ~n75073 ;
  assign n75090 = decrypt_pad & ~\u0_uk_K_r14_reg[2]/NET0131  ;
  assign n75091 = ~decrypt_pad & ~\u0_uk_K_r14_reg[50]/NET0131  ;
  assign n75092 = ~n75090 & ~n75091 ;
  assign n75093 = \u0_R14_reg[24]/NET0131  & ~n75092 ;
  assign n75094 = ~\u0_R14_reg[24]/NET0131  & n75092 ;
  assign n75095 = ~n75093 & ~n75094 ;
  assign n75096 = decrypt_pad & ~\u0_uk_K_r14_reg[37]/NET0131  ;
  assign n75097 = ~decrypt_pad & ~\u0_uk_K_r14_reg[30]/NET0131  ;
  assign n75098 = ~n75096 & ~n75097 ;
  assign n75099 = \u0_R14_reg[25]/NET0131  & ~n75098 ;
  assign n75100 = ~\u0_R14_reg[25]/NET0131  & n75098 ;
  assign n75101 = ~n75099 & ~n75100 ;
  assign n75102 = ~n75095 & ~n75101 ;
  assign n75103 = n75095 & n75101 ;
  assign n75104 = ~n75102 & ~n75103 ;
  assign n75081 = decrypt_pad & ~\u0_uk_K_r14_reg[22]/NET0131  ;
  assign n75082 = ~decrypt_pad & ~\u0_uk_K_r14_reg[15]/NET0131  ;
  assign n75083 = ~n75081 & ~n75082 ;
  assign n75084 = \u0_R14_reg[26]/P0001  & ~n75083 ;
  assign n75085 = ~\u0_R14_reg[26]/P0001  & n75083 ;
  assign n75086 = ~n75084 & ~n75085 ;
  assign n75121 = n75086 & ~n75095 ;
  assign n75107 = decrypt_pad & ~\u0_uk_K_r14_reg[0]/NET0131  ;
  assign n75108 = ~decrypt_pad & ~\u0_uk_K_r14_reg[52]/NET0131  ;
  assign n75109 = ~n75107 & ~n75108 ;
  assign n75110 = \u0_R14_reg[27]/P0001  & ~n75109 ;
  assign n75111 = ~\u0_R14_reg[27]/P0001  & n75109 ;
  assign n75112 = ~n75110 & ~n75111 ;
  assign n75075 = decrypt_pad & ~\u0_uk_K_r14_reg[38]/NET0131  ;
  assign n75076 = ~decrypt_pad & ~\u0_uk_K_r14_reg[31]/NET0131  ;
  assign n75077 = ~n75075 & ~n75076 ;
  assign n75078 = \u0_R14_reg[29]/NET0131  & ~n75077 ;
  assign n75079 = ~\u0_R14_reg[29]/NET0131  & n75077 ;
  assign n75080 = ~n75078 & ~n75079 ;
  assign n75120 = n75080 & ~n75095 ;
  assign n75122 = n75112 & ~n75120 ;
  assign n75123 = ~n75121 & n75122 ;
  assign n75124 = ~n75104 & n75123 ;
  assign n75087 = n75080 & n75086 ;
  assign n75106 = n75087 & n75102 ;
  assign n75113 = n75106 & ~n75112 ;
  assign n75088 = ~n75080 & ~n75086 ;
  assign n75089 = ~n75087 & ~n75088 ;
  assign n75105 = n75089 & n75104 ;
  assign n75114 = decrypt_pad & ~\u0_uk_K_r14_reg[42]/P0001  ;
  assign n75115 = ~decrypt_pad & ~\u0_uk_K_r14_reg[35]/P0001  ;
  assign n75116 = ~n75114 & ~n75115 ;
  assign n75117 = \u0_R14_reg[28]/NET0131  & ~n75116 ;
  assign n75118 = ~\u0_R14_reg[28]/NET0131  & n75116 ;
  assign n75119 = ~n75117 & ~n75118 ;
  assign n75125 = ~n75105 & n75119 ;
  assign n75126 = ~n75113 & n75125 ;
  assign n75127 = ~n75124 & n75126 ;
  assign n75140 = n75086 & ~n75112 ;
  assign n75141 = ~n75089 & ~n75101 ;
  assign n75142 = ~n75140 & ~n75141 ;
  assign n75143 = n75095 & ~n75142 ;
  assign n75128 = n75086 & n75101 ;
  assign n75129 = ~n75101 & n75112 ;
  assign n75130 = ~n75128 & ~n75129 ;
  assign n75131 = n75120 & ~n75130 ;
  assign n75144 = ~n75119 & ~n75131 ;
  assign n75132 = ~n75080 & ~n75101 ;
  assign n75133 = n75080 & n75101 ;
  assign n75134 = ~n75132 & ~n75133 ;
  assign n75135 = ~n75112 & ~n75134 ;
  assign n75136 = ~n75080 & ~n75095 ;
  assign n75137 = ~n75086 & ~n75101 ;
  assign n75138 = ~n75128 & ~n75137 ;
  assign n75139 = n75136 & n75138 ;
  assign n75145 = ~n75135 & ~n75139 ;
  assign n75146 = n75144 & n75145 ;
  assign n75147 = ~n75143 & n75146 ;
  assign n75148 = ~n75127 & ~n75147 ;
  assign n75149 = \u0_L14_reg[12]/P0001  & n75148 ;
  assign n75150 = ~\u0_L14_reg[12]/P0001  & ~n75148 ;
  assign n75151 = ~n75149 & ~n75150 ;
  assign n75152 = ~n50917 & ~n50942 ;
  assign n75155 = ~n50978 & ~n75152 ;
  assign n75156 = n50904 & ~n75155 ;
  assign n75153 = ~n50904 & ~n50951 ;
  assign n75154 = ~n75152 & n75153 ;
  assign n75157 = ~n50955 & ~n75154 ;
  assign n75158 = n51168 & n75157 ;
  assign n75159 = ~n75156 & n75158 ;
  assign n75161 = ~n50924 & n50958 ;
  assign n75162 = ~n50904 & ~n75161 ;
  assign n75163 = ~n51155 & n75162 ;
  assign n75164 = ~n50932 & n50937 ;
  assign n75165 = ~n50973 & ~n75164 ;
  assign n75166 = ~n50917 & ~n75165 ;
  assign n75167 = n50904 & ~n51165 ;
  assign n75168 = ~n75166 & n75167 ;
  assign n75169 = ~n75163 & ~n75168 ;
  assign n75160 = ~n50910 & n50934 ;
  assign n75170 = ~n50898 & ~n50974 ;
  assign n75171 = ~n75160 & n75170 ;
  assign n75172 = ~n75169 & n75171 ;
  assign n75173 = ~n75159 & ~n75172 ;
  assign n75174 = \u0_L14_reg[17]/P0001  & ~n75173 ;
  assign n75175 = ~\u0_L14_reg[17]/P0001  & n75173 ;
  assign n75176 = ~n75174 & ~n75175 ;
  assign n75195 = ~n74943 & ~n74987 ;
  assign n75196 = ~n74885 & ~n75195 ;
  assign n75193 = n74885 & ~n74910 ;
  assign n75194 = n74898 & n75193 ;
  assign n75197 = n74932 & ~n75194 ;
  assign n75198 = ~n74998 & n75197 ;
  assign n75199 = ~n75196 & n75198 ;
  assign n75200 = n74897 & ~n74988 ;
  assign n75201 = ~n74959 & ~n75200 ;
  assign n75202 = n74885 & ~n75201 ;
  assign n75203 = ~n74932 & ~n74974 ;
  assign n75204 = ~n75202 & n75203 ;
  assign n75205 = ~n75199 & ~n75204 ;
  assign n75178 = n74910 & n74937 ;
  assign n75177 = n74898 & ~n74910 ;
  assign n75179 = ~n74922 & ~n75177 ;
  assign n75180 = ~n75178 & n75179 ;
  assign n75181 = ~n74932 & ~n75180 ;
  assign n75182 = ~n74910 & n74916 ;
  assign n75183 = ~n75181 & ~n75182 ;
  assign n75184 = ~n74885 & ~n75183 ;
  assign n75187 = n74920 & ~n74959 ;
  assign n75188 = n74885 & ~n75187 ;
  assign n75185 = ~n74914 & ~n74973 ;
  assign n75186 = ~n74885 & ~n75185 ;
  assign n75189 = n74932 & n74946 ;
  assign n75190 = ~n75186 & ~n75189 ;
  assign n75191 = ~n75188 & n75190 ;
  assign n75192 = n74910 & ~n75191 ;
  assign n75206 = ~n75184 & ~n75192 ;
  assign n75207 = ~n75205 & n75206 ;
  assign n75208 = \u0_L14_reg[4]/P0001  & n75207 ;
  assign n75209 = ~\u0_L14_reg[4]/P0001  & ~n75207 ;
  assign n75210 = ~n75208 & ~n75209 ;
  assign n75217 = n74910 & n74958 ;
  assign n75218 = ~n74987 & ~n75217 ;
  assign n75219 = n74904 & ~n75218 ;
  assign n75220 = ~n74919 & ~n75219 ;
  assign n75221 = n74885 & ~n75220 ;
  assign n75222 = n74916 & ~n74923 ;
  assign n75223 = ~n74997 & ~n75222 ;
  assign n75224 = ~n74885 & ~n75223 ;
  assign n75225 = n74939 & n74984 ;
  assign n75226 = ~n75224 & n75225 ;
  assign n75227 = ~n75221 & n75226 ;
  assign n75228 = n74932 & ~n75227 ;
  assign n75211 = ~n74911 & ~n74967 ;
  assign n75212 = ~n74897 & ~n75211 ;
  assign n75213 = n75185 & ~n75212 ;
  assign n75214 = n74885 & ~n75213 ;
  assign n75215 = ~n75178 & ~n75214 ;
  assign n75216 = ~n74932 & ~n75215 ;
  assign n75230 = ~n75177 & ~n75219 ;
  assign n75231 = ~n74885 & ~n74932 ;
  assign n75232 = ~n75230 & n75231 ;
  assign n75229 = n74946 & n75193 ;
  assign n75233 = ~n74974 & ~n75229 ;
  assign n75234 = ~n75232 & n75233 ;
  assign n75235 = ~n75216 & n75234 ;
  assign n75236 = ~n75228 & n75235 ;
  assign n75237 = ~\u0_L14_reg[29]/P0001  & n75236 ;
  assign n75238 = \u0_L14_reg[29]/P0001  & ~n75236 ;
  assign n75239 = ~n75237 & ~n75238 ;
  assign n75245 = n50809 & n50869 ;
  assign n75246 = ~n51029 & ~n51031 ;
  assign n75247 = ~n75245 & n75246 ;
  assign n75248 = n50848 & ~n75247 ;
  assign n75241 = ~n50990 & ~n51005 ;
  assign n75242 = ~n50848 & ~n75241 ;
  assign n75243 = ~n50876 & ~n50993 ;
  assign n75244 = n50856 & ~n75243 ;
  assign n75240 = n50815 & n50877 ;
  assign n75249 = n50866 & ~n75240 ;
  assign n75250 = ~n75244 & n75249 ;
  assign n75251 = ~n75242 & n75250 ;
  assign n75252 = ~n75248 & n75251 ;
  assign n75257 = ~n50867 & ~n50993 ;
  assign n75258 = n50815 & ~n50829 ;
  assign n75259 = ~n75257 & n75258 ;
  assign n75260 = ~n50866 & ~n50885 ;
  assign n75253 = n50816 & n50999 ;
  assign n75261 = ~n51047 & ~n75253 ;
  assign n75262 = n75260 & n75261 ;
  assign n75263 = ~n75259 & n75262 ;
  assign n75254 = ~n50815 & ~n50878 ;
  assign n75255 = ~n50841 & ~n51030 ;
  assign n75256 = n50848 & ~n75255 ;
  assign n75264 = ~n75254 & ~n75256 ;
  assign n75265 = n75263 & n75264 ;
  assign n75266 = ~n75252 & ~n75265 ;
  assign n75267 = n50848 & n50877 ;
  assign n75268 = n50855 & n50868 ;
  assign n75269 = ~n75267 & ~n75268 ;
  assign n75270 = ~n75266 & n75269 ;
  assign n75271 = \u0_L14_reg[21]/P0001  & n75270 ;
  assign n75272 = ~\u0_L14_reg[21]/P0001  & ~n75270 ;
  assign n75273 = ~n75271 & ~n75272 ;
  assign n75274 = n51194 & n51241 ;
  assign n75275 = ~n51225 & ~n75274 ;
  assign n75276 = n51218 & n51238 ;
  assign n75277 = ~n51250 & ~n75276 ;
  assign n75278 = ~n75019 & n75277 ;
  assign n75279 = ~n51208 & ~n75278 ;
  assign n75280 = n75275 & ~n75279 ;
  assign n75281 = ~n51201 & ~n75280 ;
  assign n75282 = ~n75025 & n75030 ;
  assign n75283 = ~n51216 & ~n75282 ;
  assign n75284 = n51201 & ~n75283 ;
  assign n75286 = n51188 & ~n51215 ;
  assign n75287 = ~n74849 & n75286 ;
  assign n75285 = n74841 & n75025 ;
  assign n75288 = ~n51208 & ~n75285 ;
  assign n75289 = ~n75287 & n75288 ;
  assign n75290 = ~n75284 & n75289 ;
  assign n75293 = ~n51219 & ~n74860 ;
  assign n75294 = n75030 & ~n75293 ;
  assign n75295 = n51208 & ~n51251 ;
  assign n75296 = ~n75294 & n75295 ;
  assign n75291 = ~n51226 & ~n75018 ;
  assign n75292 = n51201 & ~n75291 ;
  assign n75297 = n74863 & n75275 ;
  assign n75298 = ~n75292 & n75297 ;
  assign n75299 = n75296 & n75298 ;
  assign n75300 = ~n75290 & ~n75299 ;
  assign n75301 = ~n75281 & ~n75300 ;
  assign n75302 = ~\u0_L14_reg[13]/P0001  & n75301 ;
  assign n75303 = \u0_L14_reg[13]/P0001  & ~n75301 ;
  assign n75304 = ~n75302 & ~n75303 ;
  assign n75309 = n75136 & n75140 ;
  assign n75310 = n75095 & n75112 ;
  assign n75311 = ~n75086 & n75310 ;
  assign n75312 = ~n75309 & ~n75311 ;
  assign n75313 = ~n75101 & ~n75312 ;
  assign n75305 = ~n75086 & n75095 ;
  assign n75306 = ~n75121 & ~n75305 ;
  assign n75317 = n75080 & ~n75129 ;
  assign n75318 = n75306 & n75317 ;
  assign n75314 = ~n75088 & ~n75128 ;
  assign n75315 = n75095 & ~n75112 ;
  assign n75316 = ~n75314 & n75315 ;
  assign n75319 = ~n75119 & ~n75316 ;
  assign n75320 = ~n75318 & n75319 ;
  assign n75321 = ~n75313 & n75320 ;
  assign n75322 = ~n75089 & n75102 ;
  assign n75330 = n75119 & ~n75322 ;
  assign n75323 = ~n75095 & n75101 ;
  assign n75324 = ~n75305 & ~n75323 ;
  assign n75325 = n75080 & ~n75112 ;
  assign n75326 = ~n75103 & n75325 ;
  assign n75327 = ~n75324 & n75326 ;
  assign n75328 = ~n75137 & n75310 ;
  assign n75329 = n75314 & n75328 ;
  assign n75331 = ~n75327 & ~n75329 ;
  assign n75332 = n75330 & n75331 ;
  assign n75333 = ~n75321 & ~n75332 ;
  assign n75337 = n75095 & n75132 ;
  assign n75335 = ~n75080 & n75086 ;
  assign n75336 = n75323 & n75335 ;
  assign n75338 = ~n75106 & ~n75336 ;
  assign n75339 = ~n75337 & n75338 ;
  assign n75340 = n75112 & ~n75339 ;
  assign n75307 = n75101 & ~n75112 ;
  assign n75308 = n75306 & n75307 ;
  assign n75334 = n75088 & n75129 ;
  assign n75341 = ~n75308 & ~n75334 ;
  assign n75342 = ~n75340 & n75341 ;
  assign n75343 = ~n75333 & n75342 ;
  assign n75344 = ~\u0_L14_reg[22]/P0001  & ~n75343 ;
  assign n75345 = \u0_L14_reg[22]/P0001  & n75343 ;
  assign n75346 = ~n75344 & ~n75345 ;
  assign n75368 = n51096 & ~n51121 ;
  assign n75369 = ~n51095 & ~n51135 ;
  assign n75370 = ~n75368 & n75369 ;
  assign n75371 = n51104 & ~n75370 ;
  assign n75363 = ~n51104 & n51124 ;
  assign n75364 = ~n51107 & ~n51132 ;
  assign n75365 = ~n75363 & n75364 ;
  assign n75366 = ~n51092 & ~n75365 ;
  assign n75355 = n51092 & n51106 ;
  assign n75367 = n51131 & n75355 ;
  assign n75372 = ~n51122 & ~n51130 ;
  assign n75373 = ~n75367 & n75372 ;
  assign n75374 = ~n75366 & n75373 ;
  assign n75375 = ~n75371 & n75374 ;
  assign n75376 = n51067 & ~n75375 ;
  assign n75348 = ~n51073 & n51092 ;
  assign n75349 = ~n51135 & ~n75348 ;
  assign n75350 = n51086 & ~n75349 ;
  assign n75351 = ~n51086 & n51096 ;
  assign n75352 = ~n51117 & ~n75351 ;
  assign n75353 = ~n75350 & n75352 ;
  assign n75354 = ~n51104 & ~n75353 ;
  assign n75356 = ~n51124 & ~n74728 ;
  assign n75357 = ~n75355 & n75356 ;
  assign n75358 = n51104 & ~n75357 ;
  assign n75347 = ~n51092 & n51133 ;
  assign n75359 = ~n51123 & ~n75347 ;
  assign n75360 = ~n75358 & n75359 ;
  assign n75361 = ~n75354 & n75360 ;
  assign n75362 = ~n51067 & ~n75361 ;
  assign n75377 = ~n51133 & ~n75351 ;
  assign n75378 = n51092 & ~n75377 ;
  assign n75379 = ~n51104 & n75378 ;
  assign n75380 = ~n51122 & ~n74713 ;
  assign n75381 = n51104 & ~n75380 ;
  assign n75382 = ~n75379 & ~n75381 ;
  assign n75383 = ~n75362 & n75382 ;
  assign n75384 = ~n75376 & n75383 ;
  assign n75385 = \u0_L14_reg[14]/P0001  & n75384 ;
  assign n75386 = ~\u0_L14_reg[14]/P0001  & ~n75384 ;
  assign n75387 = ~n75385 & ~n75386 ;
  assign n75401 = ~n51315 & ~n51318 ;
  assign n75402 = ~n51324 & ~n75401 ;
  assign n75403 = ~n51357 & ~n51402 ;
  assign n75404 = ~n75402 & n75403 ;
  assign n75400 = ~n51278 & n51407 ;
  assign n75405 = n51369 & ~n75400 ;
  assign n75406 = n75404 & n75405 ;
  assign n75407 = ~n51292 & ~n75406 ;
  assign n75388 = n51265 & ~n51271 ;
  assign n75389 = n51363 & ~n75388 ;
  assign n75390 = n51292 & ~n75389 ;
  assign n75391 = n51284 & n75388 ;
  assign n75392 = ~n51397 & ~n75391 ;
  assign n75393 = ~n75390 & n75392 ;
  assign n75394 = n51278 & ~n75393 ;
  assign n75395 = n51310 & n51335 ;
  assign n75396 = ~n51298 & ~n51318 ;
  assign n75397 = n51292 & ~n75388 ;
  assign n75398 = n51327 & n75397 ;
  assign n75399 = ~n75396 & n75398 ;
  assign n75408 = ~n75395 & ~n75399 ;
  assign n75409 = ~n75394 & n75408 ;
  assign n75410 = ~n75407 & n75409 ;
  assign n75411 = \u0_L14_reg[6]/P0001  & n75410 ;
  assign n75412 = ~\u0_L14_reg[6]/P0001  & ~n75410 ;
  assign n75413 = ~n75411 & ~n75412 ;
  assign n75434 = ~n50934 & ~n75161 ;
  assign n75435 = n50910 & ~n75162 ;
  assign n75436 = ~n75434 & n75435 ;
  assign n75432 = ~n50974 & ~n51148 ;
  assign n75433 = n50904 & ~n75432 ;
  assign n75437 = ~n50978 & ~n75433 ;
  assign n75438 = ~n75436 & n75437 ;
  assign n75439 = ~n50898 & ~n75438 ;
  assign n75425 = ~n50957 & n50958 ;
  assign n75426 = ~n50967 & ~n75425 ;
  assign n75427 = ~n50898 & ~n75426 ;
  assign n75428 = ~n50953 & ~n50956 ;
  assign n75429 = ~n75160 & n75428 ;
  assign n75430 = ~n75427 & n75429 ;
  assign n75431 = ~n50904 & ~n75430 ;
  assign n75417 = ~n50957 & ~n50971 ;
  assign n75418 = n50904 & ~n75417 ;
  assign n75415 = ~n50911 & ~n50943 ;
  assign n75416 = n50917 & ~n75415 ;
  assign n75414 = ~n50910 & n50933 ;
  assign n75419 = n50910 & ~n50948 ;
  assign n75420 = n51153 & ~n75419 ;
  assign n75421 = ~n75414 & ~n75420 ;
  assign n75422 = ~n75416 & n75421 ;
  assign n75423 = ~n75418 & n75422 ;
  assign n75424 = n50898 & ~n75423 ;
  assign n75440 = ~n50952 & ~n50972 ;
  assign n75441 = ~n75424 & n75440 ;
  assign n75442 = ~n75431 & n75441 ;
  assign n75443 = ~n75439 & n75442 ;
  assign n75444 = \u0_L14_reg[31]/P0001  & n75443 ;
  assign n75445 = ~\u0_L14_reg[31]/P0001  & ~n75443 ;
  assign n75446 = ~n75444 & ~n75445 ;
  assign n75459 = ~n75095 & ~n75133 ;
  assign n75460 = n75138 & n75459 ;
  assign n75457 = ~n75080 & ~n75137 ;
  assign n75458 = n75095 & ~n75457 ;
  assign n75461 = ~n75112 & ~n75458 ;
  assign n75462 = ~n75460 & n75461 ;
  assign n75447 = n75080 & n75095 ;
  assign n75448 = ~n75136 & ~n75447 ;
  assign n75449 = n75128 & n75448 ;
  assign n75450 = ~n75101 & n75447 ;
  assign n75451 = n75086 & n75450 ;
  assign n75452 = ~n75449 & ~n75451 ;
  assign n75454 = ~n75086 & ~n75448 ;
  assign n75455 = ~n75132 & n75454 ;
  assign n75456 = n75112 & n75455 ;
  assign n75463 = n75452 & ~n75456 ;
  assign n75464 = ~n75462 & n75463 ;
  assign n75465 = n75119 & ~n75464 ;
  assign n75466 = ~n75112 & n75119 ;
  assign n75467 = ~n75112 & n75455 ;
  assign n75468 = n75121 & n75132 ;
  assign n75469 = ~n75467 & ~n75468 ;
  assign n75470 = ~n75466 & ~n75469 ;
  assign n75453 = ~n75112 & ~n75452 ;
  assign n75471 = n75112 & ~n75119 ;
  assign n75472 = ~n75450 & n75471 ;
  assign n75473 = ~n75449 & n75472 ;
  assign n75474 = ~n75454 & n75473 ;
  assign n75475 = ~n75453 & ~n75474 ;
  assign n75476 = ~n75470 & n75475 ;
  assign n75477 = ~n75465 & n75476 ;
  assign n75478 = \u0_L14_reg[7]/P0001  & n75477 ;
  assign n75479 = ~\u0_L14_reg[7]/P0001  & ~n75477 ;
  assign n75480 = ~n75478 & ~n75479 ;
  assign n75486 = n75137 & n75448 ;
  assign n75487 = n75104 & ~n75137 ;
  assign n75488 = n75134 & n75487 ;
  assign n75489 = ~n75486 & ~n75488 ;
  assign n75490 = ~n75112 & ~n75489 ;
  assign n75481 = n75103 & n75335 ;
  assign n75482 = ~n75086 & n75133 ;
  assign n75483 = ~n75080 & n75324 ;
  assign n75484 = ~n75482 & ~n75483 ;
  assign n75485 = n75112 & ~n75484 ;
  assign n75491 = ~n75481 & ~n75485 ;
  assign n75492 = ~n75490 & n75491 ;
  assign n75493 = n75119 & ~n75492 ;
  assign n75498 = n75088 & n75095 ;
  assign n75500 = ~n75450 & ~n75498 ;
  assign n75501 = n75112 & ~n75500 ;
  assign n75499 = n75135 & ~n75498 ;
  assign n75497 = ~n75089 & n75103 ;
  assign n75502 = ~n75336 & ~n75497 ;
  assign n75503 = ~n75499 & n75502 ;
  assign n75504 = ~n75501 & n75503 ;
  assign n75505 = ~n75119 & ~n75504 ;
  assign n75494 = n75106 & ~n75466 ;
  assign n75495 = ~n75088 & n75307 ;
  assign n75496 = ~n75306 & n75495 ;
  assign n75506 = ~n75494 & ~n75496 ;
  assign n75507 = ~n75505 & n75506 ;
  assign n75508 = ~n75493 & n75507 ;
  assign n75509 = \u0_L14_reg[32]/P0001  & n75508 ;
  assign n75510 = ~\u0_L14_reg[32]/P0001  & ~n75508 ;
  assign n75511 = ~n75509 & ~n75510 ;
  assign n75518 = ~n51093 & n51096 ;
  assign n75519 = n74729 & ~n75518 ;
  assign n75520 = n51118 & ~n74733 ;
  assign n75521 = ~n75519 & ~n75520 ;
  assign n75522 = n74714 & ~n74728 ;
  assign n75523 = ~n75521 & n75522 ;
  assign n75524 = ~n51067 & ~n75523 ;
  assign n75512 = ~n51107 & ~n51125 ;
  assign n75513 = n51104 & ~n75512 ;
  assign n75514 = ~n51104 & n51134 ;
  assign n75515 = ~n75378 & ~n75514 ;
  assign n75516 = ~n75513 & n75515 ;
  assign n75517 = n51067 & ~n75516 ;
  assign n75525 = ~n51104 & n51130 ;
  assign n75526 = ~n51097 & ~n75348 ;
  assign n75527 = n51086 & ~n75526 ;
  assign n75528 = ~n51119 & ~n75527 ;
  assign n75529 = n51104 & ~n75528 ;
  assign n75530 = ~n75525 & ~n75529 ;
  assign n75531 = ~n75517 & n75530 ;
  assign n75532 = ~n75524 & n75531 ;
  assign n75533 = \u0_L14_reg[8]/P0001  & n75532 ;
  assign n75534 = ~\u0_L14_reg[8]/P0001  & ~n75532 ;
  assign n75535 = ~n75533 & ~n75534 ;
  assign n75536 = ~n74808 & n75067 ;
  assign n75537 = ~n74766 & n74780 ;
  assign n75538 = ~n74787 & ~n74794 ;
  assign n75539 = ~n75537 & n75538 ;
  assign n75540 = ~n75536 & ~n75539 ;
  assign n75541 = ~n74760 & ~n74792 ;
  assign n75542 = n74779 & n75541 ;
  assign n75543 = ~n74774 & ~n74805 ;
  assign n75544 = ~n75542 & n75543 ;
  assign n75545 = ~n75540 & n75544 ;
  assign n75549 = n74773 & n74788 ;
  assign n75548 = n74779 & ~n74780 ;
  assign n75550 = ~n74787 & ~n75548 ;
  assign n75551 = ~n75549 & n75550 ;
  assign n75552 = n74787 & ~n75041 ;
  assign n75553 = ~n75057 & n75552 ;
  assign n75554 = ~n75551 & ~n75553 ;
  assign n75546 = n74773 & n75042 ;
  assign n75547 = n74805 & ~n75546 ;
  assign n75555 = ~n74776 & n75547 ;
  assign n75556 = ~n75554 & n75555 ;
  assign n75557 = ~n75545 & ~n75556 ;
  assign n75558 = ~n74787 & ~n75546 ;
  assign n75559 = n74787 & ~n74807 ;
  assign n75560 = n74778 & n75559 ;
  assign n75561 = ~n75558 & ~n75560 ;
  assign n75562 = ~n75053 & ~n75561 ;
  assign n75563 = ~n75557 & n75562 ;
  assign n75564 = \u0_L14_reg[1]/P0001  & n75563 ;
  assign n75565 = ~\u0_L14_reg[1]/P0001  & ~n75563 ;
  assign n75566 = ~n75564 & ~n75565 ;
  assign n75572 = n74779 & n74792 ;
  assign n75573 = ~n75040 & ~n75572 ;
  assign n75574 = n75547 & n75573 ;
  assign n75567 = n74788 & n75045 ;
  assign n75568 = ~n74767 & ~n75567 ;
  assign n75569 = ~n74787 & ~n75568 ;
  assign n75570 = ~n74821 & ~n75549 ;
  assign n75571 = n74766 & ~n75570 ;
  assign n75575 = ~n75569 & ~n75571 ;
  assign n75576 = n75574 & n75575 ;
  assign n75577 = ~n74776 & ~n74811 ;
  assign n75578 = ~n74787 & ~n75577 ;
  assign n75579 = ~n74788 & n74828 ;
  assign n75580 = ~n74805 & ~n75057 ;
  assign n75581 = n75055 & n75580 ;
  assign n75582 = ~n75579 & n75581 ;
  assign n75583 = ~n75578 & n75582 ;
  assign n75584 = ~n75576 & ~n75583 ;
  assign n75586 = n74773 & n75541 ;
  assign n75585 = ~n74773 & ~n74780 ;
  assign n75587 = n74814 & ~n75585 ;
  assign n75588 = ~n75586 & n75587 ;
  assign n75589 = n74759 & n74787 ;
  assign n75590 = ~n75058 & n75589 ;
  assign n75591 = ~n75588 & ~n75590 ;
  assign n75592 = ~n75584 & n75591 ;
  assign n75593 = \u0_L14_reg[26]/P0001  & n75592 ;
  assign n75594 = ~\u0_L14_reg[26]/P0001  & ~n75592 ;
  assign n75595 = ~n75593 & ~n75594 ;
  assign n75609 = decrypt_pad & ~\u1_uk_K_r14_reg[51]/NET0131  ;
  assign n75610 = ~decrypt_pad & ~\u1_uk_K_r14_reg[31]/NET0131  ;
  assign n75611 = ~n75609 & ~n75610 ;
  assign n75612 = \u1_R14_reg[17]/NET0131  & ~n75611 ;
  assign n75613 = ~\u1_R14_reg[17]/NET0131  & n75611 ;
  assign n75614 = ~n75612 & ~n75613 ;
  assign n75596 = decrypt_pad & ~\u1_uk_K_r14_reg[45]/NET0131  ;
  assign n75597 = ~decrypt_pad & ~\u1_uk_K_r14_reg[52]/NET0131  ;
  assign n75598 = ~n75596 & ~n75597 ;
  assign n75599 = \u1_R14_reg[21]/NET0131  & ~n75598 ;
  assign n75600 = ~\u1_R14_reg[21]/NET0131  & n75598 ;
  assign n75601 = ~n75599 & ~n75600 ;
  assign n75616 = decrypt_pad & ~\u1_uk_K_r14_reg[29]/NET0131  ;
  assign n75617 = ~decrypt_pad & ~\u1_uk_K_r14_reg[36]/NET0131  ;
  assign n75618 = ~n75616 & ~n75617 ;
  assign n75619 = \u1_R14_reg[16]/NET0131  & ~n75618 ;
  assign n75620 = ~\u1_R14_reg[16]/NET0131  & n75618 ;
  assign n75621 = ~n75619 & ~n75620 ;
  assign n75633 = n75601 & n75621 ;
  assign n75634 = ~n75614 & n75633 ;
  assign n75625 = decrypt_pad & ~\u1_uk_K_r14_reg[1]/NET0131  ;
  assign n75626 = ~decrypt_pad & ~\u1_uk_K_r14_reg[8]/P0001  ;
  assign n75627 = ~n75625 & ~n75626 ;
  assign n75628 = \u1_R14_reg[19]/P0001  & ~n75627 ;
  assign n75629 = ~\u1_R14_reg[19]/P0001  & n75627 ;
  assign n75630 = ~n75628 & ~n75629 ;
  assign n75602 = decrypt_pad & ~\u1_uk_K_r14_reg[14]/NET0131  ;
  assign n75603 = ~decrypt_pad & ~\u1_uk_K_r14_reg[21]/NET0131  ;
  assign n75604 = ~n75602 & ~n75603 ;
  assign n75605 = \u1_R14_reg[18]/NET0131  & ~n75604 ;
  assign n75606 = ~\u1_R14_reg[18]/NET0131  & n75604 ;
  assign n75607 = ~n75605 & ~n75606 ;
  assign n75631 = n75614 & ~n75621 ;
  assign n75632 = ~n75607 & n75631 ;
  assign n75635 = ~n75630 & ~n75632 ;
  assign n75636 = ~n75634 & n75635 ;
  assign n75638 = n75614 & n75633 ;
  assign n75637 = ~n75614 & ~n75621 ;
  assign n75643 = n75630 & ~n75637 ;
  assign n75644 = ~n75638 & n75643 ;
  assign n75639 = ~n75601 & ~n75614 ;
  assign n75640 = ~n75607 & n75639 ;
  assign n75641 = ~n75601 & ~n75621 ;
  assign n75642 = n75607 & n75641 ;
  assign n75645 = ~n75640 & ~n75642 ;
  assign n75646 = n75644 & n75645 ;
  assign n75647 = ~n75636 & ~n75646 ;
  assign n75608 = n75601 & ~n75607 ;
  assign n75615 = n75608 & n75614 ;
  assign n75622 = ~n75601 & n75621 ;
  assign n75623 = n75614 & n75622 ;
  assign n75624 = n75607 & n75623 ;
  assign n75648 = ~n75615 & ~n75624 ;
  assign n75649 = ~n75647 & n75648 ;
  assign n75650 = decrypt_pad & ~\u1_uk_K_r14_reg[16]/NET0131  ;
  assign n75651 = ~decrypt_pad & ~\u1_uk_K_r14_reg[23]/NET0131  ;
  assign n75652 = ~n75650 & ~n75651 ;
  assign n75653 = \u1_R14_reg[20]/NET0131  & ~n75652 ;
  assign n75654 = ~\u1_R14_reg[20]/NET0131  & n75652 ;
  assign n75655 = ~n75653 & ~n75654 ;
  assign n75656 = ~n75649 & n75655 ;
  assign n75671 = ~n75614 & n75642 ;
  assign n75672 = ~n75624 & ~n75671 ;
  assign n75673 = n75601 & n75637 ;
  assign n75674 = ~n75607 & n75673 ;
  assign n75675 = n75672 & ~n75674 ;
  assign n75676 = n75630 & ~n75675 ;
  assign n75659 = ~n75601 & n75630 ;
  assign n75660 = n75607 & n75631 ;
  assign n75661 = ~n75614 & n75622 ;
  assign n75662 = ~n75660 & ~n75661 ;
  assign n75663 = ~n75659 & ~n75662 ;
  assign n75665 = ~n75601 & n75614 ;
  assign n75666 = n75630 & ~n75665 ;
  assign n75664 = ~n75630 & ~n75637 ;
  assign n75667 = ~n75607 & ~n75664 ;
  assign n75668 = ~n75666 & n75667 ;
  assign n75669 = ~n75663 & ~n75668 ;
  assign n75670 = ~n75655 & ~n75669 ;
  assign n75657 = n75608 & n75621 ;
  assign n75658 = n75614 & n75657 ;
  assign n75677 = ~n75614 & n75621 ;
  assign n75678 = n75607 & ~n75630 ;
  assign n75679 = n75677 & n75678 ;
  assign n75680 = ~n75658 & ~n75679 ;
  assign n75681 = ~n75670 & n75680 ;
  assign n75682 = ~n75676 & n75681 ;
  assign n75683 = ~n75656 & n75682 ;
  assign n75684 = \u1_L14_reg[25]/P0001  & n75683 ;
  assign n75685 = ~\u1_L14_reg[25]/P0001  & ~n75683 ;
  assign n75686 = ~n75684 & ~n75685 ;
  assign n75687 = decrypt_pad & ~\u1_uk_K_r14_reg[33]/NET0131  ;
  assign n75688 = ~decrypt_pad & ~\u1_uk_K_r14_reg[40]/NET0131  ;
  assign n75689 = ~n75687 & ~n75688 ;
  assign n75690 = \u1_R14_reg[16]/NET0131  & ~n75689 ;
  assign n75691 = ~\u1_R14_reg[16]/NET0131  & n75689 ;
  assign n75692 = ~n75690 & ~n75691 ;
  assign n75699 = decrypt_pad & ~\u1_uk_K_r14_reg[54]/NET0131  ;
  assign n75700 = ~decrypt_pad & ~\u1_uk_K_r14_reg[4]/NET0131  ;
  assign n75701 = ~n75699 & ~n75700 ;
  assign n75702 = \u1_R14_reg[12]/NET0131  & ~n75701 ;
  assign n75703 = ~\u1_R14_reg[12]/NET0131  & n75701 ;
  assign n75704 = ~n75702 & ~n75703 ;
  assign n75730 = decrypt_pad & ~\u1_uk_K_r14_reg[25]/NET0131  ;
  assign n75731 = ~decrypt_pad & ~\u1_uk_K_r14_reg[32]/NET0131  ;
  assign n75732 = ~n75730 & ~n75731 ;
  assign n75733 = \u1_R14_reg[15]/NET0131  & ~n75732 ;
  assign n75734 = ~\u1_R14_reg[15]/NET0131  & n75732 ;
  assign n75735 = ~n75733 & ~n75734 ;
  assign n75706 = decrypt_pad & ~\u1_uk_K_r14_reg[17]/NET0131  ;
  assign n75707 = ~decrypt_pad & ~\u1_uk_K_r14_reg[24]/NET0131  ;
  assign n75708 = ~n75706 & ~n75707 ;
  assign n75709 = \u1_R14_reg[14]/NET0131  & ~n75708 ;
  assign n75710 = ~\u1_R14_reg[14]/NET0131  & n75708 ;
  assign n75711 = ~n75709 & ~n75710 ;
  assign n75713 = decrypt_pad & ~\u1_uk_K_r14_reg[48]/NET0131  ;
  assign n75714 = ~decrypt_pad & ~\u1_uk_K_r14_reg[55]/NET0131  ;
  assign n75715 = ~n75713 & ~n75714 ;
  assign n75716 = \u1_R14_reg[13]/NET0131  & ~n75715 ;
  assign n75717 = ~\u1_R14_reg[13]/NET0131  & n75715 ;
  assign n75718 = ~n75716 & ~n75717 ;
  assign n75720 = n75711 & ~n75718 ;
  assign n75693 = decrypt_pad & ~\u1_uk_K_r14_reg[13]/NET0131  ;
  assign n75694 = ~decrypt_pad & ~\u1_uk_K_r14_reg[20]/NET0131  ;
  assign n75695 = ~n75693 & ~n75694 ;
  assign n75696 = \u1_R14_reg[17]/NET0131  & ~n75695 ;
  assign n75697 = ~\u1_R14_reg[17]/NET0131  & n75695 ;
  assign n75698 = ~n75696 & ~n75697 ;
  assign n75747 = ~n75698 & ~n75718 ;
  assign n75751 = ~n75720 & ~n75747 ;
  assign n75752 = n75735 & ~n75751 ;
  assign n75724 = ~n75711 & n75718 ;
  assign n75753 = ~n75711 & ~n75735 ;
  assign n75754 = n75698 & n75753 ;
  assign n75755 = ~n75724 & ~n75754 ;
  assign n75756 = ~n75752 & n75755 ;
  assign n75757 = n75704 & ~n75756 ;
  assign n75737 = ~n75704 & n75718 ;
  assign n75738 = ~n75698 & n75737 ;
  assign n75746 = n75711 & n75738 ;
  assign n75748 = ~n75704 & ~n75711 ;
  assign n75749 = n75747 & n75748 ;
  assign n75750 = ~n75746 & ~n75749 ;
  assign n75758 = ~n75704 & n75747 ;
  assign n75759 = ~n75735 & n75758 ;
  assign n75727 = n75698 & ~n75704 ;
  assign n75760 = n75727 & n75735 ;
  assign n75761 = ~n75711 & n75760 ;
  assign n75762 = ~n75759 & ~n75761 ;
  assign n75763 = n75750 & n75762 ;
  assign n75764 = ~n75757 & n75763 ;
  assign n75765 = ~n75692 & ~n75764 ;
  assign n75705 = n75698 & n75704 ;
  assign n75739 = n75705 & ~n75718 ;
  assign n75740 = ~n75711 & n75739 ;
  assign n75741 = ~n75738 & ~n75740 ;
  assign n75742 = n75735 & ~n75741 ;
  assign n75712 = n75705 & n75711 ;
  assign n75719 = n75712 & n75718 ;
  assign n75721 = ~n75704 & n75720 ;
  assign n75722 = n75698 & n75721 ;
  assign n75723 = ~n75719 & ~n75722 ;
  assign n75725 = ~n75698 & n75704 ;
  assign n75726 = ~n75724 & n75725 ;
  assign n75728 = n75724 & n75727 ;
  assign n75729 = ~n75726 & ~n75728 ;
  assign n75736 = ~n75729 & ~n75735 ;
  assign n75743 = n75723 & ~n75736 ;
  assign n75744 = ~n75742 & n75743 ;
  assign n75745 = n75692 & ~n75744 ;
  assign n75769 = n75723 & ~n75749 ;
  assign n75770 = ~n75735 & ~n75769 ;
  assign n75766 = n75718 & n75735 ;
  assign n75767 = n75711 & n75766 ;
  assign n75768 = ~n75704 & n75767 ;
  assign n75771 = n75725 & n75766 ;
  assign n75772 = ~n75711 & n75771 ;
  assign n75773 = ~n75768 & ~n75772 ;
  assign n75774 = ~n75770 & n75773 ;
  assign n75775 = ~n75745 & n75774 ;
  assign n75776 = ~n75765 & n75775 ;
  assign n75777 = \u1_L14_reg[10]/P0001  & n75776 ;
  assign n75778 = ~\u1_L14_reg[10]/P0001  & ~n75776 ;
  assign n75779 = ~n75777 & ~n75778 ;
  assign n75780 = n28728 & n28753 ;
  assign n75781 = ~n28728 & ~n28753 ;
  assign n75782 = ~n75780 & ~n75781 ;
  assign n75783 = n28728 & ~n28747 ;
  assign n75784 = ~n28722 & ~n75783 ;
  assign n75785 = n75782 & n75784 ;
  assign n75792 = n28722 & n28753 ;
  assign n75793 = n28766 & n75792 ;
  assign n75794 = ~n28716 & ~n75793 ;
  assign n75795 = ~n75785 & n75794 ;
  assign n75786 = ~n28747 & n28755 ;
  assign n75787 = ~n28728 & n28748 ;
  assign n75788 = n28740 & n75787 ;
  assign n75789 = ~n28722 & ~n28747 ;
  assign n75790 = n28753 & n75789 ;
  assign n75791 = ~n75788 & ~n75790 ;
  assign n75796 = ~n75786 & n75791 ;
  assign n75797 = n75795 & n75796 ;
  assign n75803 = ~n28752 & ~n28763 ;
  assign n75801 = ~n28734 & n28747 ;
  assign n75802 = n28740 & ~n75801 ;
  assign n75804 = n75784 & ~n75802 ;
  assign n75805 = ~n75803 & n75804 ;
  assign n75798 = n28728 & n28754 ;
  assign n75799 = ~n28747 & n75798 ;
  assign n75800 = ~n28758 & n28771 ;
  assign n75806 = n28716 & ~n75800 ;
  assign n75807 = ~n75799 & n75806 ;
  assign n75808 = ~n75805 & n75807 ;
  assign n75809 = ~n75797 & ~n75808 ;
  assign n75810 = n28734 & ~n28770 ;
  assign n75811 = n28773 & n75810 ;
  assign n75812 = ~n28722 & ~n75811 ;
  assign n75813 = n28728 & n28764 ;
  assign n75814 = n28722 & ~n28759 ;
  assign n75815 = ~n75813 & n75814 ;
  assign n75816 = ~n75812 & ~n75815 ;
  assign n75817 = ~n75809 & ~n75816 ;
  assign n75818 = \u1_L14_reg[2]/P0001  & n75817 ;
  assign n75819 = ~\u1_L14_reg[2]/P0001  & ~n75817 ;
  assign n75820 = ~n75818 & ~n75819 ;
  assign n75823 = ~n28441 & ~n28508 ;
  assign n75824 = n28453 & n28460 ;
  assign n75825 = ~n28494 & ~n75824 ;
  assign n75826 = n28447 & n75825 ;
  assign n75827 = n75823 & ~n75826 ;
  assign n75821 = ~n28453 & n28469 ;
  assign n75828 = n28447 & ~n75821 ;
  assign n75829 = ~n75825 & n75828 ;
  assign n75830 = n28441 & ~n75829 ;
  assign n75831 = ~n75827 & ~n75830 ;
  assign n75833 = n28490 & n75821 ;
  assign n75832 = n28454 & ~n28469 ;
  assign n75834 = n28482 & ~n75832 ;
  assign n75835 = ~n75833 & n75834 ;
  assign n75836 = ~n28514 & n75835 ;
  assign n75837 = ~n75831 & n75836 ;
  assign n75842 = ~n28441 & n75824 ;
  assign n75843 = ~n28461 & ~n75842 ;
  assign n75844 = n28469 & ~n75843 ;
  assign n75839 = n28441 & ~n28470 ;
  assign n75838 = n28453 & ~n28488 ;
  assign n75840 = ~n28486 & ~n75838 ;
  assign n75841 = n75839 & n75840 ;
  assign n75845 = ~n28441 & ~n28460 ;
  assign n75846 = n28463 & n75845 ;
  assign n75847 = ~n28482 & ~n75846 ;
  assign n75848 = ~n75841 & n75847 ;
  assign n75849 = ~n75844 & n75848 ;
  assign n75850 = ~n75837 & ~n75849 ;
  assign n75851 = n28460 & n75832 ;
  assign n75852 = ~n28487 & ~n75851 ;
  assign n75853 = ~n28441 & ~n75852 ;
  assign n75822 = n28493 & n75821 ;
  assign n75854 = n28460 & n28470 ;
  assign n75855 = ~n28441 & n75854 ;
  assign n75856 = ~n75822 & ~n75855 ;
  assign n75857 = ~n75853 & n75856 ;
  assign n75858 = ~n75850 & n75857 ;
  assign n75859 = \u1_L14_reg[27]/P0001  & n75858 ;
  assign n75860 = ~\u1_L14_reg[27]/P0001  & ~n75858 ;
  assign n75861 = ~n75859 & ~n75860 ;
  assign n75862 = decrypt_pad & ~\u1_uk_K_r14_reg[7]/NET0131  ;
  assign n75863 = ~decrypt_pad & ~\u1_uk_K_r14_reg[14]/NET0131  ;
  assign n75864 = ~n75862 & ~n75863 ;
  assign n75865 = \u1_R14_reg[20]/NET0131  & ~n75864 ;
  assign n75866 = ~\u1_R14_reg[20]/NET0131  & n75864 ;
  assign n75867 = ~n75865 & ~n75866 ;
  assign n75868 = decrypt_pad & ~\u1_uk_K_r14_reg[22]/NET0131  ;
  assign n75869 = ~decrypt_pad & ~\u1_uk_K_r14_reg[29]/NET0131  ;
  assign n75870 = ~n75868 & ~n75869 ;
  assign n75871 = \u1_R14_reg[21]/NET0131  & ~n75870 ;
  assign n75872 = ~\u1_R14_reg[21]/NET0131  & n75870 ;
  assign n75873 = ~n75871 & ~n75872 ;
  assign n75882 = decrypt_pad & ~\u1_uk_K_r14_reg[44]/NET0131  ;
  assign n75883 = ~decrypt_pad & ~\u1_uk_K_r14_reg[51]/NET0131  ;
  assign n75884 = ~n75882 & ~n75883 ;
  assign n75885 = \u1_R14_reg[22]/P0001  & ~n75884 ;
  assign n75886 = ~\u1_R14_reg[22]/P0001  & n75884 ;
  assign n75887 = ~n75885 & ~n75886 ;
  assign n75888 = n75873 & ~n75887 ;
  assign n75902 = n75867 & n75888 ;
  assign n75874 = decrypt_pad & ~\u1_uk_K_r14_reg[2]/NET0131  ;
  assign n75875 = ~decrypt_pad & ~\u1_uk_K_r14_reg[9]/NET0131  ;
  assign n75876 = ~n75874 & ~n75875 ;
  assign n75877 = \u1_R14_reg[23]/P0001  & ~n75876 ;
  assign n75878 = ~\u1_R14_reg[23]/P0001  & n75876 ;
  assign n75879 = ~n75877 & ~n75878 ;
  assign n75889 = decrypt_pad & ~\u1_uk_K_r14_reg[23]/NET0131  ;
  assign n75890 = ~decrypt_pad & ~\u1_uk_K_r14_reg[30]/NET0131  ;
  assign n75891 = ~n75889 & ~n75890 ;
  assign n75892 = \u1_R14_reg[25]/NET0131  & ~n75891 ;
  assign n75893 = ~\u1_R14_reg[25]/NET0131  & n75891 ;
  assign n75894 = ~n75892 & ~n75893 ;
  assign n75903 = ~n75867 & n75894 ;
  assign n75904 = ~n75873 & n75903 ;
  assign n75905 = n75879 & ~n75904 ;
  assign n75906 = ~n75902 & n75905 ;
  assign n75907 = n75867 & n75894 ;
  assign n75908 = ~n75873 & ~n75887 ;
  assign n75909 = n75907 & n75908 ;
  assign n75910 = ~n75879 & ~n75909 ;
  assign n75911 = ~n75906 & ~n75910 ;
  assign n75912 = ~n75867 & ~n75894 ;
  assign n75913 = n75887 & n75912 ;
  assign n75914 = ~n75887 & n75903 ;
  assign n75915 = ~n75913 & ~n75914 ;
  assign n75916 = ~n75873 & ~n75915 ;
  assign n75917 = ~n75867 & n75873 ;
  assign n75918 = n75887 & n75917 ;
  assign n75919 = n75894 & n75918 ;
  assign n75895 = n75888 & ~n75894 ;
  assign n75880 = n75867 & ~n75873 ;
  assign n75881 = ~n75879 & n75880 ;
  assign n75896 = decrypt_pad & ~\u1_uk_K_r14_reg[28]/NET0131  ;
  assign n75897 = ~decrypt_pad & ~\u1_uk_K_r14_reg[35]/P0001  ;
  assign n75898 = ~n75896 & ~n75897 ;
  assign n75899 = \u1_R14_reg[24]/NET0131  & ~n75898 ;
  assign n75900 = ~\u1_R14_reg[24]/NET0131  & n75898 ;
  assign n75901 = ~n75899 & ~n75900 ;
  assign n75920 = ~n75881 & n75901 ;
  assign n75921 = ~n75895 & n75920 ;
  assign n75922 = ~n75919 & n75921 ;
  assign n75923 = ~n75916 & n75922 ;
  assign n75924 = ~n75911 & n75923 ;
  assign n75927 = ~n75873 & n75912 ;
  assign n75928 = n75873 & n75894 ;
  assign n75929 = ~n75867 & n75928 ;
  assign n75930 = ~n75927 & ~n75929 ;
  assign n75931 = n75910 & n75930 ;
  assign n75933 = ~n75894 & n75917 ;
  assign n75932 = n75867 & ~n75888 ;
  assign n75934 = n75879 & ~n75932 ;
  assign n75935 = ~n75933 & n75934 ;
  assign n75936 = ~n75931 & ~n75935 ;
  assign n75925 = n75873 & n75907 ;
  assign n75926 = n75887 & n75925 ;
  assign n75937 = ~n75901 & ~n75926 ;
  assign n75938 = ~n75936 & n75937 ;
  assign n75939 = ~n75924 & ~n75938 ;
  assign n75940 = n75879 & ~n75887 ;
  assign n75941 = n75904 & n75940 ;
  assign n75942 = ~n75879 & ~n75887 ;
  assign n75943 = n75867 & ~n75894 ;
  assign n75944 = n75873 & n75943 ;
  assign n75945 = n75942 & n75944 ;
  assign n75946 = ~n75941 & ~n75945 ;
  assign n75947 = ~n75939 & n75946 ;
  assign n75948 = \u1_L14_reg[19]/P0001  & n75947 ;
  assign n75949 = ~\u1_L14_reg[19]/P0001  & ~n75947 ;
  assign n75950 = ~n75948 & ~n75949 ;
  assign n75973 = ~n75887 & ~n75928 ;
  assign n75974 = ~n75907 & ~n75918 ;
  assign n75975 = ~n75973 & n75974 ;
  assign n75976 = n75910 & ~n75975 ;
  assign n75968 = ~n75873 & n75943 ;
  assign n75969 = ~n75887 & n75968 ;
  assign n75970 = n75879 & ~n75918 ;
  assign n75971 = ~n75925 & n75970 ;
  assign n75972 = ~n75969 & n75971 ;
  assign n75977 = n75901 & ~n75972 ;
  assign n75978 = ~n75976 & n75977 ;
  assign n75960 = ~n75867 & ~n75887 ;
  assign n75961 = n75905 & ~n75960 ;
  assign n75962 = ~n75879 & ~n75902 ;
  assign n75963 = ~n75918 & n75962 ;
  assign n75964 = ~n75961 & ~n75963 ;
  assign n75952 = n75942 & n75943 ;
  assign n75953 = n75887 & n75907 ;
  assign n75954 = ~n75873 & n75953 ;
  assign n75955 = ~n75952 & ~n75954 ;
  assign n75956 = n75879 & n75887 ;
  assign n75957 = ~n75873 & n75956 ;
  assign n75958 = ~n75895 & ~n75957 ;
  assign n75959 = n75867 & ~n75958 ;
  assign n75965 = n75955 & ~n75959 ;
  assign n75966 = ~n75964 & n75965 ;
  assign n75967 = ~n75901 & ~n75966 ;
  assign n75979 = n75888 & n75912 ;
  assign n75980 = ~n75953 & ~n75979 ;
  assign n75981 = n75879 & ~n75980 ;
  assign n75951 = n75927 & n75942 ;
  assign n75982 = n75946 & ~n75951 ;
  assign n75983 = ~n75981 & n75982 ;
  assign n75984 = ~n75967 & n75983 ;
  assign n75985 = ~n75978 & n75984 ;
  assign n75986 = ~\u1_L14_reg[11]/P0001  & n75985 ;
  assign n75987 = \u1_L14_reg[11]/P0001  & ~n75985 ;
  assign n75988 = ~n75986 & ~n75987 ;
  assign n75989 = n75607 & n75673 ;
  assign n75990 = n75630 & ~n75989 ;
  assign n75991 = n75621 & n75640 ;
  assign n75992 = n75990 & ~n75991 ;
  assign n75993 = ~n75621 & n75640 ;
  assign n75996 = ~n75630 & ~n75993 ;
  assign n75994 = ~n75607 & n75623 ;
  assign n75995 = n75607 & n75634 ;
  assign n75997 = ~n75994 & ~n75995 ;
  assign n75998 = n75996 & n75997 ;
  assign n75999 = ~n75992 & ~n75998 ;
  assign n76000 = n75607 & ~n75614 ;
  assign n76001 = n75608 & ~n75677 ;
  assign n76002 = ~n75630 & ~n76001 ;
  assign n76003 = ~n76000 & ~n76002 ;
  assign n76004 = ~n75622 & ~n76003 ;
  assign n76005 = n75608 & ~n75621 ;
  assign n76006 = ~n75623 & ~n76005 ;
  assign n76007 = n75630 & ~n76006 ;
  assign n76008 = ~n75655 & ~n76007 ;
  assign n76009 = ~n76004 & n76008 ;
  assign n76012 = ~n75621 & n75665 ;
  assign n76013 = ~n75657 & ~n76012 ;
  assign n76014 = n75630 & ~n76013 ;
  assign n76015 = n75601 & n75631 ;
  assign n76016 = ~n75630 & n76015 ;
  assign n76010 = n75622 & n76000 ;
  assign n76011 = n75655 & ~n76010 ;
  assign n76017 = ~n75658 & n76011 ;
  assign n76018 = ~n76016 & n76017 ;
  assign n76019 = ~n76014 & n76018 ;
  assign n76020 = ~n76009 & ~n76019 ;
  assign n76021 = ~n75999 & ~n76020 ;
  assign n76022 = \u1_L14_reg[3]/P0001  & n76021 ;
  assign n76023 = ~\u1_L14_reg[3]/P0001  & ~n76021 ;
  assign n76024 = ~n76022 & ~n76023 ;
  assign n76025 = n28753 & n28758 ;
  assign n76026 = ~n75783 & ~n76025 ;
  assign n76027 = n28741 & n28758 ;
  assign n76028 = n28722 & ~n76027 ;
  assign n76029 = ~n75798 & n76028 ;
  assign n76030 = n76026 & n76029 ;
  assign n76034 = n28753 & ~n76026 ;
  assign n76031 = ~n28740 & n28758 ;
  assign n76032 = ~n28722 & ~n28776 ;
  assign n76033 = ~n76031 & n76032 ;
  assign n76035 = n75781 & ~n75801 ;
  assign n76036 = n76033 & ~n76035 ;
  assign n76037 = ~n76034 & n76036 ;
  assign n76038 = ~n76030 & ~n76037 ;
  assign n76039 = n28716 & ~n76038 ;
  assign n76040 = n28722 & ~n76035 ;
  assign n76041 = ~n28740 & n75801 ;
  assign n76042 = n75782 & ~n76041 ;
  assign n76043 = n76033 & ~n76042 ;
  assign n76044 = ~n76040 & ~n76043 ;
  assign n76045 = n28728 & n28741 ;
  assign n76046 = ~n28740 & ~n75803 ;
  assign n76047 = ~n76045 & ~n76046 ;
  assign n76048 = n28747 & ~n76047 ;
  assign n76049 = ~n28716 & ~n76048 ;
  assign n76050 = ~n76044 & n76049 ;
  assign n76051 = ~n76039 & ~n76050 ;
  assign n76052 = \u1_L14_reg[28]/P0001  & ~n76051 ;
  assign n76053 = ~\u1_L14_reg[28]/P0001  & n76051 ;
  assign n76054 = ~n76052 & ~n76053 ;
  assign n76060 = ~n75718 & n75760 ;
  assign n76055 = n75704 & ~n75718 ;
  assign n76056 = ~n75737 & ~n76055 ;
  assign n76057 = n75753 & ~n76056 ;
  assign n76059 = ~n75728 & ~n75771 ;
  assign n76062 = ~n76057 & n76059 ;
  assign n76063 = ~n76060 & n76062 ;
  assign n76058 = n75711 & n75759 ;
  assign n76061 = n75692 & ~n75719 ;
  assign n76064 = ~n76058 & n76061 ;
  assign n76065 = n76063 & n76064 ;
  assign n76073 = ~n75692 & ~n75740 ;
  assign n76066 = n75698 & ~n75718 ;
  assign n76067 = n75735 & ~n76066 ;
  assign n76068 = ~n75725 & ~n75737 ;
  assign n76069 = n76067 & n76068 ;
  assign n76074 = ~n75768 & ~n76069 ;
  assign n76075 = n76073 & n76074 ;
  assign n76070 = n75711 & n75725 ;
  assign n76071 = ~n76066 & ~n76070 ;
  assign n76072 = ~n75735 & ~n76071 ;
  assign n76076 = n75750 & ~n76072 ;
  assign n76077 = n76075 & n76076 ;
  assign n76078 = ~n76065 & ~n76077 ;
  assign n76079 = ~n75728 & ~n75735 ;
  assign n76080 = n75720 & n75725 ;
  assign n76081 = n75735 & ~n76080 ;
  assign n76082 = ~n75749 & n76081 ;
  assign n76083 = ~n76079 & ~n76082 ;
  assign n76084 = ~n75772 & ~n76083 ;
  assign n76085 = ~n76078 & n76084 ;
  assign n76086 = ~\u1_L14_reg[20]/P0001  & ~n76085 ;
  assign n76087 = \u1_L14_reg[20]/P0001  & n76085 ;
  assign n76088 = ~n76086 & ~n76087 ;
  assign n76102 = decrypt_pad & ~\u1_uk_K_r14_reg[15]/NET0131  ;
  assign n76103 = ~decrypt_pad & ~\u1_uk_K_r14_reg[22]/NET0131  ;
  assign n76104 = ~n76102 & ~n76103 ;
  assign n76105 = \u1_R14_reg[26]/NET0131  & ~n76104 ;
  assign n76106 = ~\u1_R14_reg[26]/NET0131  & n76104 ;
  assign n76107 = ~n76105 & ~n76106 ;
  assign n76108 = decrypt_pad & ~\u1_uk_K_r14_reg[50]/NET0131  ;
  assign n76109 = ~decrypt_pad & ~\u1_uk_K_r14_reg[2]/NET0131  ;
  assign n76110 = ~n76108 & ~n76109 ;
  assign n76111 = \u1_R14_reg[24]/NET0131  & ~n76110 ;
  assign n76112 = ~\u1_R14_reg[24]/NET0131  & n76110 ;
  assign n76113 = ~n76111 & ~n76112 ;
  assign n76089 = decrypt_pad & ~\u1_uk_K_r14_reg[30]/NET0131  ;
  assign n76090 = ~decrypt_pad & ~\u1_uk_K_r14_reg[37]/NET0131  ;
  assign n76091 = ~n76089 & ~n76090 ;
  assign n76092 = \u1_R14_reg[25]/NET0131  & ~n76091 ;
  assign n76093 = ~\u1_R14_reg[25]/NET0131  & n76091 ;
  assign n76094 = ~n76092 & ~n76093 ;
  assign n76095 = decrypt_pad & ~\u1_uk_K_r14_reg[31]/NET0131  ;
  assign n76096 = ~decrypt_pad & ~\u1_uk_K_r14_reg[38]/NET0131  ;
  assign n76097 = ~n76095 & ~n76096 ;
  assign n76098 = \u1_R14_reg[29]/NET0131  & ~n76097 ;
  assign n76099 = ~\u1_R14_reg[29]/NET0131  & n76097 ;
  assign n76100 = ~n76098 & ~n76099 ;
  assign n76129 = n76094 & ~n76100 ;
  assign n76130 = ~n76113 & n76129 ;
  assign n76131 = ~n76094 & ~n76100 ;
  assign n76132 = n76113 & n76131 ;
  assign n76133 = ~n76130 & ~n76132 ;
  assign n76134 = n76107 & n76133 ;
  assign n76101 = ~n76094 & n76100 ;
  assign n76135 = n76101 & n76113 ;
  assign n76136 = n76094 & n76100 ;
  assign n76137 = ~n76113 & n76136 ;
  assign n76138 = ~n76135 & ~n76137 ;
  assign n76139 = ~n76107 & n76138 ;
  assign n76140 = ~n76134 & ~n76139 ;
  assign n76142 = ~n76107 & ~n76113 ;
  assign n76143 = ~n76094 & ~n76142 ;
  assign n76116 = decrypt_pad & ~\u1_uk_K_r14_reg[52]/NET0131  ;
  assign n76117 = ~decrypt_pad & ~\u1_uk_K_r14_reg[0]/P0001  ;
  assign n76118 = ~n76116 & ~n76117 ;
  assign n76119 = \u1_R14_reg[27]/P0001  & ~n76118 ;
  assign n76120 = ~\u1_R14_reg[27]/P0001  & n76118 ;
  assign n76121 = ~n76119 & ~n76120 ;
  assign n76141 = ~n76113 & ~n76131 ;
  assign n76144 = n76121 & ~n76141 ;
  assign n76145 = ~n76143 & n76144 ;
  assign n76114 = n76107 & ~n76113 ;
  assign n76115 = n76101 & n76114 ;
  assign n76122 = n76115 & ~n76121 ;
  assign n76123 = decrypt_pad & ~\u1_uk_K_r14_reg[35]/P0001  ;
  assign n76124 = ~decrypt_pad & ~\u1_uk_K_r14_reg[42]/P0001  ;
  assign n76125 = ~n76123 & ~n76124 ;
  assign n76126 = \u1_R14_reg[28]/NET0131  & ~n76125 ;
  assign n76127 = ~\u1_R14_reg[28]/NET0131  & n76125 ;
  assign n76128 = ~n76126 & ~n76127 ;
  assign n76146 = ~n76122 & n76128 ;
  assign n76147 = ~n76145 & n76146 ;
  assign n76148 = ~n76140 & n76147 ;
  assign n76155 = ~n76107 & ~n76133 ;
  assign n76153 = n76107 & n76113 ;
  assign n76154 = ~n76121 & n76153 ;
  assign n76150 = n76100 & ~n76113 ;
  assign n76151 = ~n76094 & n76121 ;
  assign n76152 = n76150 & n76151 ;
  assign n76159 = ~n76128 & ~n76152 ;
  assign n76160 = ~n76154 & n76159 ;
  assign n76149 = n76107 & n76135 ;
  assign n76156 = ~n76131 & ~n76136 ;
  assign n76157 = ~n76114 & n76121 ;
  assign n76158 = ~n76156 & ~n76157 ;
  assign n76161 = ~n76149 & ~n76158 ;
  assign n76162 = n76160 & n76161 ;
  assign n76163 = ~n76155 & n76162 ;
  assign n76164 = ~n76148 & ~n76163 ;
  assign n76165 = \u1_L14_reg[12]/P0001  & n76164 ;
  assign n76166 = ~\u1_L14_reg[12]/P0001  & ~n76164 ;
  assign n76167 = ~n76165 & ~n76166 ;
  assign n76168 = ~n28557 & ~n28579 ;
  assign n76169 = ~n28601 & ~n76168 ;
  assign n76170 = n28531 & ~n76169 ;
  assign n76173 = n28576 & ~n28586 ;
  assign n76171 = ~n28531 & ~n28557 ;
  assign n76172 = n28579 & n76171 ;
  assign n76174 = ~n28591 & ~n76172 ;
  assign n76175 = n76173 & n76174 ;
  assign n76176 = ~n28558 & n76175 ;
  assign n76177 = ~n76170 & n76176 ;
  assign n76182 = n28550 & n28560 ;
  assign n76183 = ~n28563 & ~n76182 ;
  assign n76181 = ~n28537 & n28604 ;
  assign n76180 = n28559 & n28565 ;
  assign n76184 = n28531 & ~n76180 ;
  assign n76185 = ~n76181 & n76184 ;
  assign n76186 = n76183 & n76185 ;
  assign n76187 = ~n28560 & ~n28565 ;
  assign n76188 = ~n28550 & ~n76187 ;
  assign n76189 = n28544 & ~n28557 ;
  assign n76190 = ~n28531 & ~n76189 ;
  assign n76191 = ~n76188 & n76190 ;
  assign n76192 = ~n76186 & ~n76191 ;
  assign n76178 = ~n28550 & n28587 ;
  assign n76179 = n28543 & n76178 ;
  assign n76193 = ~n28576 & ~n28603 ;
  assign n76194 = ~n76179 & n76193 ;
  assign n76195 = ~n76192 & n76194 ;
  assign n76196 = ~n76177 & ~n76195 ;
  assign n76197 = \u1_L14_reg[17]/P0001  & ~n76196 ;
  assign n76198 = ~\u1_L14_reg[17]/P0001  & n76196 ;
  assign n76199 = ~n76197 & ~n76198 ;
  assign n76219 = n75887 & n75904 ;
  assign n76200 = ~n75887 & n75907 ;
  assign n76220 = ~n75933 & ~n76200 ;
  assign n76221 = ~n76219 & n76220 ;
  assign n76222 = ~n75879 & ~n76221 ;
  assign n76216 = ~n75914 & ~n75944 ;
  assign n76217 = ~n75954 & n76216 ;
  assign n76218 = n75879 & ~n76217 ;
  assign n76223 = ~n75969 & ~n76218 ;
  assign n76224 = ~n76222 & n76223 ;
  assign n76225 = ~n75901 & ~n76224 ;
  assign n76202 = ~n75895 & ~n75960 ;
  assign n76203 = ~n75879 & ~n76202 ;
  assign n76201 = n75879 & n76200 ;
  assign n76204 = n75887 & n75928 ;
  assign n76205 = ~n75979 & ~n76204 ;
  assign n76206 = ~n76201 & n76205 ;
  assign n76207 = ~n76203 & n76206 ;
  assign n76208 = n75901 & ~n76207 ;
  assign n76209 = n75930 & ~n75944 ;
  assign n76210 = n75956 & ~n76209 ;
  assign n76211 = ~n75925 & ~n75968 ;
  assign n76212 = n75887 & n76211 ;
  assign n76213 = ~n75887 & ~n75912 ;
  assign n76214 = ~n75879 & ~n76213 ;
  assign n76215 = ~n76212 & n76214 ;
  assign n76226 = ~n76210 & ~n76215 ;
  assign n76227 = ~n76208 & n76226 ;
  assign n76228 = ~n76225 & n76227 ;
  assign n76229 = \u1_L14_reg[4]/P0001  & n76228 ;
  assign n76230 = ~\u1_L14_reg[4]/P0001  & ~n76228 ;
  assign n76231 = ~n76229 & ~n76230 ;
  assign n76239 = n75887 & n75943 ;
  assign n76240 = ~n75960 & ~n76239 ;
  assign n76241 = n75873 & ~n76240 ;
  assign n76245 = ~n75929 & ~n76241 ;
  assign n76246 = n75879 & ~n76245 ;
  assign n76247 = ~n75888 & n75912 ;
  assign n76248 = ~n75953 & ~n76247 ;
  assign n76249 = ~n75879 & ~n76248 ;
  assign n76250 = ~n75916 & n75955 ;
  assign n76251 = ~n76249 & n76250 ;
  assign n76252 = ~n76246 & n76251 ;
  assign n76253 = n75901 & ~n76252 ;
  assign n76232 = ~n75908 & ~n75918 ;
  assign n76233 = ~n75894 & ~n76232 ;
  assign n76234 = n76211 & ~n76233 ;
  assign n76235 = n75879 & ~n76234 ;
  assign n76236 = ~n76219 & ~n76235 ;
  assign n76237 = ~n75901 & ~n76236 ;
  assign n76242 = ~n76200 & ~n76241 ;
  assign n76243 = ~n75879 & ~n75901 ;
  assign n76244 = ~n76242 & n76243 ;
  assign n76238 = n75928 & n75940 ;
  assign n76254 = ~n75969 & ~n76238 ;
  assign n76255 = ~n76244 & n76254 ;
  assign n76256 = ~n76237 & n76255 ;
  assign n76257 = ~n76253 & n76256 ;
  assign n76258 = ~\u1_L14_reg[29]/P0001  & n76257 ;
  assign n76259 = \u1_L14_reg[29]/P0001  & ~n76257 ;
  assign n76260 = ~n76258 & ~n76259 ;
  assign n76267 = ~n28469 & ~n28493 ;
  assign n76268 = n75824 & n76267 ;
  assign n76271 = ~n28509 & n75847 ;
  assign n76272 = ~n76268 & n76271 ;
  assign n76264 = ~n28453 & n28462 ;
  assign n76265 = ~n28491 & ~n76264 ;
  assign n76266 = n28441 & ~n76265 ;
  assign n76263 = n28496 & n28504 ;
  assign n76269 = ~n28486 & ~n75833 ;
  assign n76270 = ~n76263 & n76269 ;
  assign n76273 = ~n76266 & n76270 ;
  assign n76274 = n76272 & n76273 ;
  assign n76277 = ~n28441 & ~n28475 ;
  assign n76278 = ~n28492 & n76277 ;
  assign n76280 = n28441 & ~n28505 ;
  assign n76279 = n28462 & n28469 ;
  assign n76281 = ~n75832 & ~n76279 ;
  assign n76282 = n76280 & n76281 ;
  assign n76283 = ~n76278 & ~n76282 ;
  assign n76275 = ~n28462 & ~n28507 ;
  assign n76276 = n75821 & ~n76275 ;
  assign n76284 = n28482 & ~n28515 ;
  assign n76285 = ~n76276 & n76284 ;
  assign n76286 = ~n76283 & n76285 ;
  assign n76287 = ~n76274 & ~n76286 ;
  assign n76261 = n28488 & n75842 ;
  assign n76262 = n28441 & n28508 ;
  assign n76288 = ~n76261 & ~n76262 ;
  assign n76289 = ~n76287 & n76288 ;
  assign n76290 = \u1_L14_reg[21]/P0001  & n76289 ;
  assign n76291 = ~\u1_L14_reg[21]/P0001  & ~n76289 ;
  assign n76292 = ~n76290 & ~n76291 ;
  assign n76295 = ~n28716 & ~n28722 ;
  assign n76296 = ~n76025 & n76295 ;
  assign n76293 = n28757 & n75783 ;
  assign n76294 = ~n28748 & n28782 ;
  assign n76297 = ~n76293 & ~n76294 ;
  assign n76298 = n76296 & n76297 ;
  assign n76299 = n28722 & ~n28775 ;
  assign n76300 = ~n75787 & n76299 ;
  assign n76301 = ~n28722 & ~n75780 ;
  assign n76302 = ~n76041 & n76301 ;
  assign n76303 = ~n76300 & ~n76302 ;
  assign n76304 = n28716 & ~n28765 ;
  assign n76305 = n75791 & n76304 ;
  assign n76306 = ~n76303 & n76305 ;
  assign n76307 = ~n76298 & ~n76306 ;
  assign n76308 = n28734 & n75813 ;
  assign n76309 = ~n28776 & ~n76308 ;
  assign n76310 = ~n76307 & n76309 ;
  assign n76311 = ~n28747 & ~n28757 ;
  assign n76312 = n75803 & n76311 ;
  assign n76313 = ~n28741 & n28766 ;
  assign n76314 = ~n28716 & n28722 ;
  assign n76315 = ~n76313 & n76314 ;
  assign n76316 = ~n76046 & n76315 ;
  assign n76317 = ~n76312 & n76316 ;
  assign n76318 = ~n76310 & ~n76317 ;
  assign n76319 = ~\u1_L14_reg[13]/P0001  & ~n76318 ;
  assign n76320 = \u1_L14_reg[13]/P0001  & n76318 ;
  assign n76321 = ~n76319 & ~n76320 ;
  assign n76334 = ~n28482 & ~n75855 ;
  assign n76335 = ~n28463 & ~n28474 ;
  assign n76336 = ~n75854 & ~n76335 ;
  assign n76337 = n28441 & ~n76336 ;
  assign n76338 = ~n28491 & n75823 ;
  assign n76339 = ~n75854 & n76338 ;
  assign n76340 = ~n76337 & ~n76339 ;
  assign n76341 = ~n28514 & ~n76340 ;
  assign n76342 = ~n76334 & ~n76341 ;
  assign n76323 = ~n28461 & ~n75833 ;
  assign n76324 = n28441 & ~n76323 ;
  assign n76327 = ~n28453 & ~n28485 ;
  assign n76328 = ~n28441 & ~n28454 ;
  assign n76329 = ~n76327 & n76328 ;
  assign n76322 = n28453 & n76279 ;
  assign n76325 = n28441 & ~n28463 ;
  assign n76326 = n28474 & ~n76325 ;
  assign n76330 = ~n76322 & ~n76326 ;
  assign n76331 = ~n76329 & n76330 ;
  assign n76332 = ~n76324 & n76331 ;
  assign n76333 = ~n28482 & ~n76332 ;
  assign n76343 = n28461 & n28469 ;
  assign n76344 = ~n28509 & ~n76343 ;
  assign n76345 = n75852 & n76344 ;
  assign n76346 = n28441 & ~n76345 ;
  assign n76347 = ~n76333 & ~n76346 ;
  assign n76348 = ~n76342 & n76347 ;
  assign n76349 = ~\u1_L14_reg[5]/P0001  & n76348 ;
  assign n76350 = \u1_L14_reg[5]/P0001  & ~n76348 ;
  assign n76351 = ~n76349 & ~n76350 ;
  assign n76370 = ~n76121 & ~n76132 ;
  assign n76368 = ~n76100 & n76113 ;
  assign n76369 = ~n76107 & ~n76368 ;
  assign n76371 = ~n76141 & ~n76369 ;
  assign n76372 = n76370 & n76371 ;
  assign n76376 = ~n76107 & n76150 ;
  assign n76377 = ~n76151 & n76376 ;
  assign n76355 = ~n76094 & ~n76107 ;
  assign n76354 = n76113 & n76121 ;
  assign n76373 = ~n76354 & ~n76368 ;
  assign n76374 = n76355 & ~n76373 ;
  assign n76375 = n76136 & n76153 ;
  assign n76378 = ~n76374 & ~n76375 ;
  assign n76379 = ~n76377 & n76378 ;
  assign n76380 = ~n76372 & n76379 ;
  assign n76381 = ~n76128 & ~n76380 ;
  assign n76361 = n76107 & ~n76137 ;
  assign n76362 = ~n76121 & ~n76138 ;
  assign n76363 = ~n76361 & n76362 ;
  assign n76356 = n76094 & n76107 ;
  assign n76357 = ~n76355 & ~n76356 ;
  assign n76352 = ~n76100 & ~n76107 ;
  assign n76358 = ~n76352 & n76354 ;
  assign n76359 = n76357 & n76358 ;
  assign n76360 = n76131 & n76142 ;
  assign n76364 = ~n76115 & ~n76360 ;
  assign n76365 = ~n76359 & n76364 ;
  assign n76366 = ~n76363 & n76365 ;
  assign n76367 = n76128 & ~n76366 ;
  assign n76382 = n76114 & n76156 ;
  assign n76383 = ~n76132 & ~n76382 ;
  assign n76384 = n76121 & ~n76383 ;
  assign n76353 = n76151 & n76352 ;
  assign n76385 = ~n76142 & ~n76153 ;
  assign n76386 = n76094 & ~n76121 ;
  assign n76387 = ~n76385 & n76386 ;
  assign n76388 = ~n76353 & ~n76387 ;
  assign n76389 = ~n76384 & n76388 ;
  assign n76390 = ~n76367 & n76389 ;
  assign n76391 = ~n76381 & n76390 ;
  assign n76392 = ~\u1_L14_reg[22]/P0001  & ~n76391 ;
  assign n76393 = \u1_L14_reg[22]/P0001  & n76391 ;
  assign n76394 = ~n76392 & ~n76393 ;
  assign n76395 = ~n75614 & n75641 ;
  assign n76396 = n75607 & n75633 ;
  assign n76397 = n75630 & ~n75632 ;
  assign n76398 = ~n76396 & n76397 ;
  assign n76399 = ~n76395 & n76398 ;
  assign n76400 = n75607 & n75665 ;
  assign n76401 = ~n75630 & ~n75673 ;
  assign n76402 = ~n76400 & n76401 ;
  assign n76403 = ~n75658 & ~n75991 ;
  assign n76404 = n76402 & n76403 ;
  assign n76405 = ~n76399 & ~n76404 ;
  assign n76406 = ~n75607 & n76012 ;
  assign n76407 = ~n75655 & ~n75995 ;
  assign n76408 = ~n76406 & n76407 ;
  assign n76409 = ~n76405 & n76408 ;
  assign n76415 = ~n75639 & ~n75641 ;
  assign n76416 = n76398 & n76415 ;
  assign n76412 = ~n76015 & ~n76395 ;
  assign n76413 = ~n75607 & ~n75630 ;
  assign n76414 = ~n76412 & n76413 ;
  assign n76417 = ~n75994 & n76011 ;
  assign n76410 = ~n75614 & n75657 ;
  assign n76411 = n75638 & n75678 ;
  assign n76418 = ~n76410 & ~n76411 ;
  assign n76419 = n76417 & n76418 ;
  assign n76420 = ~n76414 & n76419 ;
  assign n76421 = ~n76416 & n76420 ;
  assign n76422 = ~n76409 & ~n76421 ;
  assign n76423 = ~n75673 & ~n76012 ;
  assign n76424 = n75607 & ~n76423 ;
  assign n76425 = ~n75630 & n76424 ;
  assign n76426 = ~n75671 & ~n75994 ;
  assign n76427 = n75630 & ~n76426 ;
  assign n76428 = ~n76425 & ~n76427 ;
  assign n76429 = ~n76422 & n76428 ;
  assign n76430 = \u1_L14_reg[14]/P0001  & n76429 ;
  assign n76431 = ~\u1_L14_reg[14]/P0001  & ~n76429 ;
  assign n76432 = ~n76430 & ~n76431 ;
  assign n76441 = n28668 & n28669 ;
  assign n76436 = ~n28639 & n28665 ;
  assign n76440 = n28683 & n76436 ;
  assign n76442 = ~n28627 & ~n76440 ;
  assign n76443 = ~n76441 & n76442 ;
  assign n76439 = n28688 & n28698 ;
  assign n76433 = ~n28633 & n28653 ;
  assign n76434 = ~n28683 & ~n76433 ;
  assign n76435 = ~n28681 & ~n76434 ;
  assign n76437 = n28678 & ~n76436 ;
  assign n76438 = n28681 & n76437 ;
  assign n76444 = ~n76435 & ~n76438 ;
  assign n76445 = ~n76439 & n76444 ;
  assign n76446 = n76443 & n76445 ;
  assign n76448 = ~n28639 & ~n28683 ;
  assign n76449 = ~n28665 & ~n28669 ;
  assign n76450 = ~n28675 & n76449 ;
  assign n76451 = ~n76448 & n76450 ;
  assign n76447 = n28657 & n28669 ;
  assign n76452 = n28627 & ~n76447 ;
  assign n76453 = ~n76451 & n76452 ;
  assign n76454 = ~n76446 & ~n76453 ;
  assign n76457 = ~n28657 & ~n28669 ;
  assign n76458 = ~n28680 & ~n76457 ;
  assign n76459 = ~n28675 & ~n76458 ;
  assign n76460 = n28627 & ~n76459 ;
  assign n76455 = ~n28653 & n28680 ;
  assign n76456 = ~n28633 & n76455 ;
  assign n76461 = ~n28676 & ~n76456 ;
  assign n76462 = ~n76460 & n76461 ;
  assign n76463 = n28665 & ~n76462 ;
  assign n76464 = ~n76454 & ~n76463 ;
  assign n76465 = \u1_L14_reg[6]/P0001  & n76464 ;
  assign n76466 = ~\u1_L14_reg[6]/P0001  & ~n76464 ;
  assign n76467 = ~n76465 & ~n76466 ;
  assign n76485 = n28531 & ~n28600 ;
  assign n76486 = ~n28603 & n76485 ;
  assign n76487 = ~n28537 & ~n28557 ;
  assign n76488 = ~n28567 & n76487 ;
  assign n76489 = ~n28531 & ~n76488 ;
  assign n76490 = ~n28564 & n76489 ;
  assign n76491 = ~n76486 & ~n76490 ;
  assign n76482 = n28543 & n28588 ;
  assign n76483 = ~n76189 & ~n76482 ;
  assign n76484 = n28550 & ~n76483 ;
  assign n76492 = ~n28601 & ~n76484 ;
  assign n76493 = ~n76491 & n76492 ;
  assign n76494 = ~n28576 & ~n76493 ;
  assign n76472 = ~n28543 & n28587 ;
  assign n76473 = ~n28567 & ~n76472 ;
  assign n76474 = n28531 & ~n76473 ;
  assign n76469 = n28557 & ~n28592 ;
  assign n76468 = n28550 & ~n28614 ;
  assign n76470 = ~n28565 & ~n76468 ;
  assign n76471 = ~n76469 & n76470 ;
  assign n76475 = ~n28594 & ~n76178 ;
  assign n76476 = ~n76471 & n76475 ;
  assign n76477 = ~n76474 & n76476 ;
  assign n76478 = n28576 & ~n76477 ;
  assign n76479 = ~n28551 & ~n28561 ;
  assign n76480 = ~n76179 & n76479 ;
  assign n76481 = ~n28531 & ~n76480 ;
  assign n76495 = ~n28607 & ~n28613 ;
  assign n76496 = ~n76481 & n76495 ;
  assign n76497 = ~n76478 & n76496 ;
  assign n76498 = ~n76494 & n76497 ;
  assign n76499 = \u1_L14_reg[31]/P0001  & n76498 ;
  assign n76500 = ~\u1_L14_reg[31]/P0001  & ~n76498 ;
  assign n76501 = ~n76499 & ~n76500 ;
  assign n76513 = n28568 & ~n28602 ;
  assign n76514 = n28531 & ~n76513 ;
  assign n76509 = ~n28537 & ~n76182 ;
  assign n76510 = n28537 & ~n76188 ;
  assign n76511 = ~n76509 & ~n76510 ;
  assign n76504 = ~n28562 & ~n28604 ;
  assign n76512 = ~n28531 & ~n76504 ;
  assign n76515 = ~n76511 & ~n76512 ;
  assign n76516 = ~n76514 & n76515 ;
  assign n76517 = ~n28576 & ~n76516 ;
  assign n76502 = ~n28569 & n76183 ;
  assign n76503 = n28537 & ~n76502 ;
  assign n76505 = n28614 & ~n76504 ;
  assign n76506 = ~n28558 & ~n76505 ;
  assign n76507 = ~n76503 & n76506 ;
  assign n76508 = n28576 & ~n76507 ;
  assign n76518 = n28537 & ~n28604 ;
  assign n76519 = ~n28531 & ~n76509 ;
  assign n76520 = ~n76518 & n76519 ;
  assign n76521 = ~n76508 & ~n76520 ;
  assign n76522 = ~n76517 & n76521 ;
  assign n76523 = \u1_L14_reg[9]/P0001  & n76522 ;
  assign n76524 = ~\u1_L14_reg[9]/P0001  & ~n76522 ;
  assign n76525 = ~n76523 & ~n76524 ;
  assign n76527 = ~n76150 & ~n76368 ;
  assign n76528 = ~n76356 & ~n76527 ;
  assign n76529 = ~n76107 & ~n76131 ;
  assign n76530 = n76527 & ~n76529 ;
  assign n76531 = ~n76528 & ~n76530 ;
  assign n76526 = n76121 & ~n76128 ;
  assign n76532 = ~n76121 & n76128 ;
  assign n76533 = ~n76526 & ~n76532 ;
  assign n76534 = ~n76135 & n76533 ;
  assign n76535 = ~n76531 & n76534 ;
  assign n76536 = ~n76128 & ~n76375 ;
  assign n76537 = ~n76100 & n76114 ;
  assign n76538 = n76121 & ~n76537 ;
  assign n76539 = ~n76528 & n76538 ;
  assign n76540 = n76536 & n76539 ;
  assign n76541 = ~n76535 & ~n76540 ;
  assign n76542 = ~n76113 & n76131 ;
  assign n76543 = n76107 & n76542 ;
  assign n76544 = ~n76541 & ~n76543 ;
  assign n76547 = ~n76113 & ~n76357 ;
  assign n76546 = n76094 & ~n76527 ;
  assign n76545 = ~n76136 & n76153 ;
  assign n76548 = n76532 & ~n76545 ;
  assign n76549 = ~n76546 & n76548 ;
  assign n76550 = ~n76547 & n76549 ;
  assign n76551 = ~n76544 & ~n76550 ;
  assign n76552 = \u1_L14_reg[7]/P0001  & ~n76551 ;
  assign n76553 = ~\u1_L14_reg[7]/P0001  & n76551 ;
  assign n76554 = ~n76552 & ~n76553 ;
  assign n76559 = n76355 & ~n76527 ;
  assign n76560 = ~n76121 & ~n76130 ;
  assign n76561 = ~n76149 & n76560 ;
  assign n76562 = ~n76559 & n76561 ;
  assign n76563 = n76107 & ~n76368 ;
  assign n76564 = ~n76101 & ~n76352 ;
  assign n76565 = ~n76563 & n76564 ;
  assign n76566 = n76121 & ~n76542 ;
  assign n76567 = ~n76565 & n76566 ;
  assign n76568 = ~n76562 & ~n76567 ;
  assign n76558 = n76356 & n76368 ;
  assign n76569 = n76128 & ~n76558 ;
  assign n76570 = ~n76568 & n76569 ;
  assign n76571 = n76113 & n76352 ;
  assign n76574 = ~n76121 & ~n76156 ;
  assign n76575 = ~n76571 & n76574 ;
  assign n76576 = ~n76382 & n76536 ;
  assign n76572 = n76094 & n76571 ;
  assign n76573 = n76354 & ~n76564 ;
  assign n76577 = ~n76572 & ~n76573 ;
  assign n76578 = n76576 & n76577 ;
  assign n76579 = ~n76575 & n76578 ;
  assign n76580 = ~n76570 & ~n76579 ;
  assign n76555 = n76115 & n76121 ;
  assign n76556 = ~n76352 & n76386 ;
  assign n76557 = n76385 & n76556 ;
  assign n76581 = ~n76555 & ~n76557 ;
  assign n76582 = ~n76580 & n76581 ;
  assign n76583 = \u1_L14_reg[32]/P0001  & n76582 ;
  assign n76584 = ~\u1_L14_reg[32]/P0001  & ~n76582 ;
  assign n76585 = ~n76583 & ~n76584 ;
  assign n76604 = ~n28633 & n28668 ;
  assign n76605 = ~n28670 & ~n76604 ;
  assign n76606 = n28659 & n76605 ;
  assign n76607 = n28665 & ~n76606 ;
  assign n76608 = n28647 & n28653 ;
  assign n76609 = ~n76607 & ~n76608 ;
  assign n76610 = ~n28627 & ~n76609 ;
  assign n76588 = ~n28682 & ~n76458 ;
  assign n76589 = ~n28665 & ~n76588 ;
  assign n76590 = ~n28627 & ~n76589 ;
  assign n76599 = n28627 & ~n76438 ;
  assign n76597 = ~n28665 & ~n28678 ;
  assign n76598 = ~n28681 & n76597 ;
  assign n76591 = ~n28653 & n28665 ;
  assign n76592 = ~n28633 & ~n28655 ;
  assign n76593 = n76591 & n76592 ;
  assign n76594 = n28665 & ~n28680 ;
  assign n76595 = ~n28640 & n28653 ;
  assign n76596 = n76594 & n76595 ;
  assign n76600 = ~n76593 & ~n76596 ;
  assign n76601 = ~n76598 & n76600 ;
  assign n76602 = n76599 & n76601 ;
  assign n76603 = ~n76590 & ~n76602 ;
  assign n76586 = n28633 & n28679 ;
  assign n76587 = n28698 & n76586 ;
  assign n76611 = ~n28647 & ~n28688 ;
  assign n76612 = n76591 & ~n76611 ;
  assign n76613 = ~n76587 & ~n76612 ;
  assign n76614 = ~n76603 & n76613 ;
  assign n76615 = ~n76610 & n76614 ;
  assign n76616 = \u1_L14_reg[24]/P0001  & n76615 ;
  assign n76617 = ~\u1_L14_reg[24]/P0001  & ~n76615 ;
  assign n76618 = ~n76616 & ~n76617 ;
  assign n76619 = n28653 & ~n28688 ;
  assign n76620 = ~n28700 & ~n76592 ;
  assign n76621 = n28669 & n76436 ;
  assign n76622 = ~n28647 & ~n28653 ;
  assign n76623 = ~n76621 & n76622 ;
  assign n76624 = ~n76620 & n76623 ;
  assign n76625 = ~n76619 & ~n76624 ;
  assign n76626 = ~n28657 & ~n28689 ;
  assign n76627 = ~n28646 & ~n28665 ;
  assign n76628 = ~n76626 & n76627 ;
  assign n76629 = ~n76625 & ~n76628 ;
  assign n76630 = n28627 & ~n76629 ;
  assign n76635 = ~n76455 & ~n76620 ;
  assign n76636 = ~n28665 & ~n76635 ;
  assign n76637 = ~n28633 & ~n28679 ;
  assign n76638 = ~n76586 & n76594 ;
  assign n76639 = ~n76637 & n76638 ;
  assign n76640 = ~n76456 & ~n76639 ;
  assign n76641 = ~n76636 & n76640 ;
  assign n76642 = ~n28627 & ~n76641 ;
  assign n76631 = n28680 & n76433 ;
  assign n76632 = ~n76441 & ~n76631 ;
  assign n76633 = n28665 & ~n76632 ;
  assign n76634 = n28640 & n28698 ;
  assign n76643 = ~n76633 & ~n76634 ;
  assign n76644 = ~n76642 & n76643 ;
  assign n76645 = ~n76630 & n76644 ;
  assign n76646 = \u1_L14_reg[16]/P0001  & n76645 ;
  assign n76647 = ~\u1_L14_reg[16]/P0001  & ~n76645 ;
  assign n76648 = ~n76646 & ~n76647 ;
  assign n76662 = ~n75634 & ~n76005 ;
  assign n76663 = ~n76015 & n76662 ;
  assign n76664 = ~n75630 & ~n76663 ;
  assign n76660 = ~n75638 & ~n75991 ;
  assign n76661 = n75630 & ~n76660 ;
  assign n76665 = ~n75632 & n75672 ;
  assign n76666 = ~n76661 & n76665 ;
  assign n76667 = ~n76664 & n76666 ;
  assign n76668 = ~n75655 & ~n76667 ;
  assign n76649 = ~n75634 & ~n75993 ;
  assign n76650 = n75630 & ~n76649 ;
  assign n76651 = n75621 & n76413 ;
  assign n76652 = ~n76424 & ~n76651 ;
  assign n76653 = ~n76650 & n76652 ;
  assign n76654 = n75655 & ~n76653 ;
  assign n76655 = ~n75630 & ~n76010 ;
  assign n76656 = n75601 & n75632 ;
  assign n76657 = ~n76400 & ~n76656 ;
  assign n76658 = n75990 & n76657 ;
  assign n76659 = ~n76655 & ~n76658 ;
  assign n76669 = ~n76654 & ~n76659 ;
  assign n76670 = ~n76668 & n76669 ;
  assign n76671 = \u1_L14_reg[8]/P0001  & n76670 ;
  assign n76672 = ~\u1_L14_reg[8]/P0001  & ~n76670 ;
  assign n76673 = ~n76671 & ~n76672 ;
  assign n76678 = ~n75698 & n75748 ;
  assign n76679 = n76081 & ~n76678 ;
  assign n76680 = ~n75711 & n75725 ;
  assign n76681 = ~n75735 & ~n75739 ;
  assign n76682 = ~n76680 & n76681 ;
  assign n76683 = ~n76679 & ~n76682 ;
  assign n76684 = n75724 & n75725 ;
  assign n76685 = ~n75692 & ~n75728 ;
  assign n76686 = ~n76684 & n76685 ;
  assign n76687 = ~n75719 & n76686 ;
  assign n76688 = ~n76683 & n76687 ;
  assign n76690 = ~n75711 & n76055 ;
  assign n76691 = n76067 & ~n76690 ;
  assign n76693 = n75718 & n75727 ;
  assign n76692 = n75724 & ~n75725 ;
  assign n76694 = ~n75735 & ~n76692 ;
  assign n76695 = ~n76693 & n76694 ;
  assign n76696 = ~n76691 & ~n76695 ;
  assign n76674 = n75718 & n76070 ;
  assign n76689 = n75692 & ~n76674 ;
  assign n76697 = ~n75721 & n76689 ;
  assign n76698 = ~n76696 & n76697 ;
  assign n76699 = ~n76688 & ~n76698 ;
  assign n76676 = n75723 & ~n75746 ;
  assign n76677 = n75735 & ~n76676 ;
  assign n76675 = ~n75735 & n76674 ;
  assign n76700 = ~n76058 & ~n76675 ;
  assign n76701 = ~n76677 & n76700 ;
  assign n76702 = ~n76699 & n76701 ;
  assign n76703 = \u1_L14_reg[1]/P0001  & n76702 ;
  assign n76704 = ~\u1_L14_reg[1]/P0001  & ~n76702 ;
  assign n76705 = ~n76703 & ~n76704 ;
  assign n76709 = ~n75698 & ~n76056 ;
  assign n76708 = n75705 & n75718 ;
  assign n76710 = ~n75735 & ~n76708 ;
  assign n76711 = ~n76709 & n76710 ;
  assign n76706 = n75698 & ~n76056 ;
  assign n76707 = n75735 & ~n76706 ;
  assign n76712 = ~n75711 & ~n76707 ;
  assign n76713 = ~n76711 & n76712 ;
  assign n76714 = ~n75711 & n75738 ;
  assign n76720 = n75735 & n75758 ;
  assign n76721 = ~n76714 & ~n76720 ;
  assign n76722 = n76689 & n76721 ;
  assign n76715 = n75748 & n76066 ;
  assign n76716 = ~n75712 & ~n76715 ;
  assign n76717 = ~n75735 & ~n76716 ;
  assign n76718 = ~n75760 & ~n76693 ;
  assign n76719 = n75711 & ~n76718 ;
  assign n76723 = ~n76717 & ~n76719 ;
  assign n76724 = n76722 & n76723 ;
  assign n76725 = ~n75721 & ~n75747 ;
  assign n76726 = ~n75735 & ~n76725 ;
  assign n76727 = ~n75727 & n75767 ;
  assign n76728 = ~n75692 & ~n76690 ;
  assign n76729 = n76059 & n76728 ;
  assign n76730 = ~n76727 & n76729 ;
  assign n76731 = ~n76726 & n76730 ;
  assign n76732 = ~n76724 & ~n76731 ;
  assign n76733 = ~n76713 & ~n76732 ;
  assign n76734 = \u1_L14_reg[26]/P0001  & n76733 ;
  assign n76735 = ~\u1_L14_reg[26]/P0001  & ~n76733 ;
  assign n76736 = ~n76734 & ~n76735 ;
  assign n76774 = decrypt_pad & ~\u2_uk_K_r14_reg[23]/NET0131  ;
  assign n76775 = ~decrypt_pad & ~\u2_uk_K_r14_reg[16]/NET0131  ;
  assign n76776 = ~n76774 & ~n76775 ;
  assign n76777 = \u2_R14_reg[20]/NET0131  & ~n76776 ;
  assign n76778 = ~\u2_R14_reg[20]/NET0131  & n76776 ;
  assign n76779 = ~n76777 & ~n76778 ;
  assign n76767 = decrypt_pad & ~\u2_uk_K_r14_reg[8]/NET0131  ;
  assign n76768 = ~decrypt_pad & ~\u2_uk_K_r14_reg[1]/NET0131  ;
  assign n76769 = ~n76767 & ~n76768 ;
  assign n76770 = \u2_R14_reg[19]/P0001  & ~n76769 ;
  assign n76771 = ~\u2_R14_reg[19]/P0001  & n76769 ;
  assign n76772 = ~n76770 & ~n76771 ;
  assign n76737 = decrypt_pad & ~\u2_uk_K_r14_reg[31]/NET0131  ;
  assign n76738 = ~decrypt_pad & ~\u2_uk_K_r14_reg[51]/NET0131  ;
  assign n76739 = ~n76737 & ~n76738 ;
  assign n76740 = \u2_R14_reg[17]/NET0131  & ~n76739 ;
  assign n76741 = ~\u2_R14_reg[17]/NET0131  & n76739 ;
  assign n76742 = ~n76740 & ~n76741 ;
  assign n76743 = decrypt_pad & ~\u2_uk_K_r14_reg[36]/NET0131  ;
  assign n76744 = ~decrypt_pad & ~\u2_uk_K_r14_reg[29]/NET0131  ;
  assign n76745 = ~n76743 & ~n76744 ;
  assign n76746 = \u2_R14_reg[16]/NET0131  & ~n76745 ;
  assign n76747 = ~\u2_R14_reg[16]/NET0131  & n76745 ;
  assign n76748 = ~n76746 & ~n76747 ;
  assign n76750 = decrypt_pad & ~\u2_uk_K_r14_reg[52]/NET0131  ;
  assign n76751 = ~decrypt_pad & ~\u2_uk_K_r14_reg[45]/NET0131  ;
  assign n76752 = ~n76750 & ~n76751 ;
  assign n76753 = \u2_R14_reg[21]/NET0131  & ~n76752 ;
  assign n76754 = ~\u2_R14_reg[21]/NET0131  & n76752 ;
  assign n76755 = ~n76753 & ~n76754 ;
  assign n76780 = n76748 & n76755 ;
  assign n76781 = ~n76742 & n76780 ;
  assign n76782 = ~n76772 & ~n76781 ;
  assign n76760 = decrypt_pad & ~\u2_uk_K_r14_reg[21]/NET0131  ;
  assign n76761 = ~decrypt_pad & ~\u2_uk_K_r14_reg[14]/NET0131  ;
  assign n76762 = ~n76760 & ~n76761 ;
  assign n76763 = \u2_R14_reg[18]/NET0131  & ~n76762 ;
  assign n76764 = ~\u2_R14_reg[18]/NET0131  & n76762 ;
  assign n76765 = ~n76763 & ~n76764 ;
  assign n76783 = n76742 & ~n76765 ;
  assign n76784 = ~n76748 & n76783 ;
  assign n76785 = n76782 & ~n76784 ;
  assign n76788 = n76748 & n76765 ;
  assign n76789 = ~n76755 & ~n76783 ;
  assign n76790 = ~n76788 & n76789 ;
  assign n76749 = ~n76742 & ~n76748 ;
  assign n76786 = n76742 & n76780 ;
  assign n76787 = n76772 & ~n76786 ;
  assign n76791 = ~n76749 & n76787 ;
  assign n76792 = ~n76790 & n76791 ;
  assign n76793 = ~n76785 & ~n76792 ;
  assign n76757 = n76748 & ~n76755 ;
  assign n76795 = n76755 & ~n76765 ;
  assign n76796 = ~n76757 & ~n76795 ;
  assign n76794 = ~n76755 & ~n76765 ;
  assign n76797 = n76742 & ~n76794 ;
  assign n76798 = ~n76796 & n76797 ;
  assign n76799 = ~n76793 & ~n76798 ;
  assign n76800 = n76779 & ~n76799 ;
  assign n76801 = ~n76755 & n76772 ;
  assign n76802 = ~n76748 & n76765 ;
  assign n76803 = ~n76801 & n76802 ;
  assign n76804 = n76772 & n76794 ;
  assign n76805 = ~n76803 & ~n76804 ;
  assign n76806 = ~n76779 & ~n76805 ;
  assign n76807 = ~n76765 & n76780 ;
  assign n76808 = ~n76806 & ~n76807 ;
  assign n76809 = n76742 & ~n76808 ;
  assign n76756 = n76749 & ~n76755 ;
  assign n76758 = n76742 & n76757 ;
  assign n76759 = ~n76756 & ~n76758 ;
  assign n76766 = ~n76759 & n76765 ;
  assign n76773 = n76766 & n76772 ;
  assign n76813 = ~n76765 & ~n76779 ;
  assign n76814 = ~n76780 & n76813 ;
  assign n76815 = ~n76772 & ~n76788 ;
  assign n76816 = ~n76814 & n76815 ;
  assign n76810 = ~n76748 & n76755 ;
  assign n76811 = ~n76765 & n76810 ;
  assign n76812 = n76772 & ~n76811 ;
  assign n76817 = ~n76742 & ~n76812 ;
  assign n76818 = ~n76816 & n76817 ;
  assign n76819 = ~n76773 & ~n76818 ;
  assign n76820 = ~n76809 & n76819 ;
  assign n76821 = ~n76800 & n76820 ;
  assign n76822 = \u2_L14_reg[25]/P0001  & n76821 ;
  assign n76823 = ~\u2_L14_reg[25]/P0001  & ~n76821 ;
  assign n76824 = ~n76822 & ~n76823 ;
  assign n76852 = decrypt_pad & ~\u2_uk_K_r14_reg[39]/P0001  ;
  assign n76853 = ~decrypt_pad & ~\u2_uk_K_r14_reg[32]/NET0131  ;
  assign n76854 = ~n76852 & ~n76853 ;
  assign n76855 = \u2_R14_reg[8]/NET0131  & ~n76854 ;
  assign n76856 = ~\u2_R14_reg[8]/NET0131  & n76854 ;
  assign n76857 = ~n76855 & ~n76856 ;
  assign n76838 = decrypt_pad & ~\u2_uk_K_r14_reg[48]/NET0131  ;
  assign n76839 = ~decrypt_pad & ~\u2_uk_K_r14_reg[41]/NET0131  ;
  assign n76840 = ~n76838 & ~n76839 ;
  assign n76841 = \u2_R14_reg[7]/P0001  & ~n76840 ;
  assign n76842 = ~\u2_R14_reg[7]/P0001  & n76840 ;
  assign n76843 = ~n76841 & ~n76842 ;
  assign n76844 = decrypt_pad & ~\u2_uk_K_r14_reg[6]/NET0131  ;
  assign n76845 = ~decrypt_pad & ~\u2_uk_K_r14_reg[24]/NET0131  ;
  assign n76846 = ~n76844 & ~n76845 ;
  assign n76847 = \u2_R14_reg[5]/NET0131  & ~n76846 ;
  assign n76848 = ~\u2_R14_reg[5]/NET0131  & n76846 ;
  assign n76849 = ~n76847 & ~n76848 ;
  assign n76825 = decrypt_pad & ~\u2_uk_K_r14_reg[19]/NET0131  ;
  assign n76826 = ~decrypt_pad & ~\u2_uk_K_r14_reg[12]/NET0131  ;
  assign n76827 = ~n76825 & ~n76826 ;
  assign n76828 = \u2_R14_reg[9]/NET0131  & ~n76827 ;
  assign n76829 = ~\u2_R14_reg[9]/NET0131  & n76827 ;
  assign n76830 = ~n76828 & ~n76829 ;
  assign n76831 = decrypt_pad & ~\u2_uk_K_r14_reg[27]/NET0131  ;
  assign n76832 = ~decrypt_pad & ~\u2_uk_K_r14_reg[20]/NET0131  ;
  assign n76833 = ~n76831 & ~n76832 ;
  assign n76834 = \u2_R14_reg[4]/NET0131  & ~n76833 ;
  assign n76835 = ~\u2_R14_reg[4]/NET0131  & n76833 ;
  assign n76836 = ~n76834 & ~n76835 ;
  assign n76862 = ~n76830 & n76836 ;
  assign n76863 = ~n76849 & n76862 ;
  assign n76864 = n76830 & n76836 ;
  assign n76865 = decrypt_pad & ~\u2_uk_K_r14_reg[54]/NET0131  ;
  assign n76866 = ~decrypt_pad & ~\u2_uk_K_r14_reg[47]/NET0131  ;
  assign n76867 = ~n76865 & ~n76866 ;
  assign n76868 = \u2_R14_reg[6]/NET0131  & ~n76867 ;
  assign n76869 = ~\u2_R14_reg[6]/NET0131  & n76867 ;
  assign n76870 = ~n76868 & ~n76869 ;
  assign n76871 = n76864 & ~n76870 ;
  assign n76872 = ~n76863 & ~n76871 ;
  assign n76873 = ~n76843 & ~n76872 ;
  assign n76858 = ~n76830 & n76849 ;
  assign n76837 = n76830 & ~n76836 ;
  assign n76859 = n76837 & ~n76849 ;
  assign n76860 = ~n76858 & ~n76859 ;
  assign n76861 = n76843 & ~n76860 ;
  assign n76874 = ~n76849 & n76870 ;
  assign n76875 = ~n76836 & n76874 ;
  assign n76876 = ~n76830 & n76875 ;
  assign n76877 = ~n76861 & ~n76876 ;
  assign n76878 = ~n76873 & n76877 ;
  assign n76879 = n76857 & ~n76878 ;
  assign n76887 = ~n76843 & n76870 ;
  assign n76888 = n76849 & ~n76887 ;
  assign n76889 = ~n76836 & ~n76874 ;
  assign n76890 = ~n76888 & n76889 ;
  assign n76880 = ~n76849 & ~n76870 ;
  assign n76850 = ~n76843 & n76849 ;
  assign n76885 = ~n76850 & n76864 ;
  assign n76886 = ~n76880 & n76885 ;
  assign n76881 = ~n76830 & n76880 ;
  assign n76882 = n76836 & n76849 ;
  assign n76883 = ~n76830 & n76870 ;
  assign n76884 = n76882 & n76883 ;
  assign n76891 = ~n76881 & ~n76884 ;
  assign n76892 = ~n76886 & n76891 ;
  assign n76893 = ~n76890 & n76892 ;
  assign n76894 = ~n76857 & ~n76893 ;
  assign n76851 = n76837 & n76850 ;
  assign n76895 = ~n76830 & ~n76836 ;
  assign n76896 = n76849 & n76895 ;
  assign n76897 = ~n76870 & n76896 ;
  assign n76898 = n76864 & n76870 ;
  assign n76899 = ~n76897 & ~n76898 ;
  assign n76900 = n76843 & ~n76899 ;
  assign n76901 = ~n76851 & ~n76900 ;
  assign n76902 = ~n76894 & n76901 ;
  assign n76903 = ~n76879 & n76902 ;
  assign n76904 = \u2_L14_reg[18]/P0001  & n76903 ;
  assign n76905 = ~\u2_L14_reg[18]/P0001  & ~n76903 ;
  assign n76906 = ~n76904 & ~n76905 ;
  assign n76934 = decrypt_pad & ~\u2_uk_K_r14_reg[40]/NET0131  ;
  assign n76935 = ~decrypt_pad & ~\u2_uk_K_r14_reg[33]/NET0131  ;
  assign n76936 = ~n76934 & ~n76935 ;
  assign n76937 = \u2_R14_reg[16]/NET0131  & ~n76936 ;
  assign n76938 = ~\u2_R14_reg[16]/NET0131  & n76936 ;
  assign n76939 = ~n76937 & ~n76938 ;
  assign n76907 = decrypt_pad & ~\u2_uk_K_r14_reg[32]/NET0131  ;
  assign n76908 = ~decrypt_pad & ~\u2_uk_K_r14_reg[25]/NET0131  ;
  assign n76909 = ~n76907 & ~n76908 ;
  assign n76910 = \u2_R14_reg[15]/NET0131  & ~n76909 ;
  assign n76911 = ~\u2_R14_reg[15]/NET0131  & n76909 ;
  assign n76912 = ~n76910 & ~n76911 ;
  assign n76913 = decrypt_pad & ~\u2_uk_K_r14_reg[24]/NET0131  ;
  assign n76914 = ~decrypt_pad & ~\u2_uk_K_r14_reg[17]/NET0131  ;
  assign n76915 = ~n76913 & ~n76914 ;
  assign n76916 = \u2_R14_reg[14]/NET0131  & ~n76915 ;
  assign n76917 = ~\u2_R14_reg[14]/NET0131  & n76915 ;
  assign n76918 = ~n76916 & ~n76917 ;
  assign n76920 = decrypt_pad & ~\u2_uk_K_r14_reg[55]/NET0131  ;
  assign n76921 = ~decrypt_pad & ~\u2_uk_K_r14_reg[48]/NET0131  ;
  assign n76922 = ~n76920 & ~n76921 ;
  assign n76923 = \u2_R14_reg[13]/NET0131  & ~n76922 ;
  assign n76924 = ~\u2_R14_reg[13]/NET0131  & n76922 ;
  assign n76925 = ~n76923 & ~n76924 ;
  assign n76960 = ~n76918 & n76925 ;
  assign n76927 = decrypt_pad & ~\u2_uk_K_r14_reg[4]/NET0131  ;
  assign n76928 = ~decrypt_pad & ~\u2_uk_K_r14_reg[54]/NET0131  ;
  assign n76929 = ~n76927 & ~n76928 ;
  assign n76930 = \u2_R14_reg[12]/NET0131  & ~n76929 ;
  assign n76931 = ~\u2_R14_reg[12]/NET0131  & n76929 ;
  assign n76932 = ~n76930 & ~n76931 ;
  assign n76940 = decrypt_pad & ~\u2_uk_K_r14_reg[20]/NET0131  ;
  assign n76941 = ~decrypt_pad & ~\u2_uk_K_r14_reg[13]/NET0131  ;
  assign n76942 = ~n76940 & ~n76941 ;
  assign n76943 = \u2_R14_reg[17]/NET0131  & ~n76942 ;
  assign n76944 = ~\u2_R14_reg[17]/NET0131  & n76942 ;
  assign n76945 = ~n76943 & ~n76944 ;
  assign n76961 = n76932 & ~n76945 ;
  assign n76962 = ~n76960 & n76961 ;
  assign n76963 = ~n76932 & n76945 ;
  assign n76964 = n76925 & n76963 ;
  assign n76965 = ~n76918 & n76964 ;
  assign n76966 = ~n76962 & ~n76965 ;
  assign n76967 = ~n76912 & ~n76966 ;
  assign n76946 = n76932 & n76945 ;
  assign n76947 = n76925 & n76946 ;
  assign n76948 = n76918 & n76947 ;
  assign n76949 = n76918 & ~n76925 ;
  assign n76950 = ~n76932 & n76949 ;
  assign n76951 = n76945 & n76950 ;
  assign n76952 = ~n76948 & ~n76951 ;
  assign n76953 = n76925 & ~n76932 ;
  assign n76954 = ~n76945 & n76953 ;
  assign n76955 = ~n76925 & n76932 ;
  assign n76956 = ~n76918 & n76955 ;
  assign n76957 = n76945 & n76956 ;
  assign n76958 = ~n76954 & ~n76957 ;
  assign n76959 = n76912 & ~n76958 ;
  assign n76968 = n76952 & ~n76959 ;
  assign n76969 = ~n76967 & n76968 ;
  assign n76970 = n76939 & ~n76969 ;
  assign n76971 = ~n76925 & ~n76945 ;
  assign n76972 = ~n76949 & ~n76971 ;
  assign n76973 = n76912 & ~n76972 ;
  assign n76974 = ~n76912 & ~n76918 ;
  assign n76975 = n76945 & n76974 ;
  assign n76976 = ~n76960 & ~n76975 ;
  assign n76977 = ~n76973 & n76976 ;
  assign n76978 = n76932 & ~n76977 ;
  assign n76979 = n76918 & n76954 ;
  assign n76919 = n76912 & n76918 ;
  assign n76980 = ~n76932 & n76971 ;
  assign n76981 = n76912 & n76963 ;
  assign n76982 = ~n76980 & ~n76981 ;
  assign n76983 = ~n76919 & ~n76982 ;
  assign n76984 = ~n76979 & ~n76983 ;
  assign n76985 = ~n76978 & n76984 ;
  assign n76986 = ~n76939 & ~n76985 ;
  assign n76987 = ~n76918 & n76980 ;
  assign n76988 = n76952 & ~n76987 ;
  assign n76989 = ~n76912 & ~n76988 ;
  assign n76926 = n76919 & n76925 ;
  assign n76933 = n76926 & ~n76932 ;
  assign n76990 = n76912 & n76925 ;
  assign n76991 = n76961 & n76990 ;
  assign n76992 = ~n76918 & n76991 ;
  assign n76993 = ~n76933 & ~n76992 ;
  assign n76994 = ~n76989 & n76993 ;
  assign n76995 = ~n76986 & n76994 ;
  assign n76996 = ~n76970 & n76995 ;
  assign n76997 = \u2_L14_reg[10]/P0001  & n76996 ;
  assign n76998 = ~\u2_L14_reg[10]/P0001  & ~n76996 ;
  assign n76999 = ~n76997 & ~n76998 ;
  assign n77001 = n76837 & n76870 ;
  assign n77002 = n76849 & n77001 ;
  assign n77000 = n76837 & n76880 ;
  assign n77003 = ~n76843 & ~n77000 ;
  assign n77004 = ~n77002 & n77003 ;
  assign n77005 = ~n76870 & n76882 ;
  assign n77006 = n76843 & ~n77005 ;
  assign n77007 = ~n76876 & n77006 ;
  assign n77008 = ~n77004 & ~n77007 ;
  assign n77009 = n76830 & ~n76849 ;
  assign n77010 = n76836 & n76870 ;
  assign n77011 = ~n77009 & n77010 ;
  assign n77012 = ~n76859 & ~n77011 ;
  assign n77013 = ~n76843 & ~n77012 ;
  assign n77014 = n76836 & n76843 ;
  assign n77015 = n76830 & n76874 ;
  assign n77016 = n77014 & n77015 ;
  assign n77021 = ~n76857 & ~n77016 ;
  assign n77022 = ~n77013 & n77021 ;
  assign n77017 = ~n76860 & ~n76870 ;
  assign n77018 = n76830 & ~n76843 ;
  assign n77019 = n76880 & n77018 ;
  assign n77020 = ~n77002 & ~n77019 ;
  assign n77023 = ~n77017 & n77020 ;
  assign n77024 = n77022 & n77023 ;
  assign n77034 = ~n76843 & ~n76849 ;
  assign n77035 = n76895 & n77034 ;
  assign n77031 = ~n76836 & n76870 ;
  assign n77032 = n76843 & n76849 ;
  assign n77033 = ~n77031 & n77032 ;
  assign n77036 = n76857 & ~n77033 ;
  assign n77037 = ~n77035 & n77036 ;
  assign n77028 = ~n76837 & ~n76862 ;
  assign n77029 = ~n76882 & n76887 ;
  assign n77030 = n77028 & n77029 ;
  assign n77025 = n76849 & n76871 ;
  assign n77026 = n76862 & ~n76870 ;
  assign n77027 = ~n76849 & n77026 ;
  assign n77038 = ~n77025 & ~n77027 ;
  assign n77039 = ~n77030 & n77038 ;
  assign n77040 = n77037 & n77039 ;
  assign n77041 = ~n77024 & ~n77040 ;
  assign n77042 = ~n77008 & ~n77041 ;
  assign n77043 = \u2_L14_reg[2]/P0001  & n77042 ;
  assign n77044 = ~\u2_L14_reg[2]/P0001  & ~n77042 ;
  assign n77045 = ~n77043 & ~n77044 ;
  assign n77046 = decrypt_pad & ~\u2_uk_K_r14_reg[7]/NET0131  ;
  assign n77047 = ~decrypt_pad & ~\u2_uk_K_r14_reg[0]/NET0131  ;
  assign n77048 = ~n77046 & ~n77047 ;
  assign n77049 = \u2_R14_reg[32]/NET0131  & ~n77048 ;
  assign n77050 = ~\u2_R14_reg[32]/NET0131  & n77048 ;
  assign n77051 = ~n77049 & ~n77050 ;
  assign n77082 = decrypt_pad & ~\u2_uk_K_r14_reg[1]/NET0131  ;
  assign n77083 = ~decrypt_pad & ~\u2_uk_K_r14_reg[49]/P0001  ;
  assign n77084 = ~n77082 & ~n77083 ;
  assign n77085 = \u2_R14_reg[31]/P0001  & ~n77084 ;
  assign n77086 = ~\u2_R14_reg[31]/P0001  & n77084 ;
  assign n77087 = ~n77085 & ~n77086 ;
  assign n77073 = decrypt_pad & ~\u2_uk_K_r14_reg[16]/NET0131  ;
  assign n77074 = ~decrypt_pad & ~\u2_uk_K_r14_reg[9]/NET0131  ;
  assign n77075 = ~n77073 & ~n77074 ;
  assign n77076 = \u2_R14_reg[28]/NET0131  & ~n77075 ;
  assign n77077 = ~\u2_R14_reg[28]/NET0131  & n77075 ;
  assign n77078 = ~n77076 & ~n77077 ;
  assign n77058 = decrypt_pad & ~\u2_uk_K_r14_reg[44]/NET0131  ;
  assign n77059 = ~decrypt_pad & ~\u2_uk_K_r14_reg[37]/NET0131  ;
  assign n77060 = ~n77058 & ~n77059 ;
  assign n77061 = \u2_R14_reg[30]/NET0131  & ~n77060 ;
  assign n77062 = ~\u2_R14_reg[30]/NET0131  & n77060 ;
  assign n77063 = ~n77061 & ~n77062 ;
  assign n77065 = decrypt_pad & ~\u2_uk_K_r14_reg[43]/NET0131  ;
  assign n77066 = ~decrypt_pad & ~\u2_uk_K_r14_reg[36]/NET0131  ;
  assign n77067 = ~n77065 & ~n77066 ;
  assign n77068 = \u2_R14_reg[29]/NET0131  & ~n77067 ;
  assign n77069 = ~\u2_R14_reg[29]/NET0131  & n77067 ;
  assign n77070 = ~n77068 & ~n77069 ;
  assign n77108 = ~n77063 & ~n77070 ;
  assign n77127 = ~n77078 & n77108 ;
  assign n77052 = decrypt_pad & ~\u2_uk_K_r14_reg[28]/NET0131  ;
  assign n77053 = ~decrypt_pad & ~\u2_uk_K_r14_reg[21]/NET0131  ;
  assign n77054 = ~n77052 & ~n77053 ;
  assign n77055 = \u2_R14_reg[1]/NET0131  & ~n77054 ;
  assign n77056 = ~\u2_R14_reg[1]/NET0131  & n77054 ;
  assign n77057 = ~n77055 & ~n77056 ;
  assign n77091 = n77057 & ~n77078 ;
  assign n77120 = n77070 & n77091 ;
  assign n77094 = ~n77057 & n77070 ;
  assign n77126 = n77078 & n77094 ;
  assign n77128 = ~n77120 & ~n77126 ;
  assign n77129 = ~n77127 & n77128 ;
  assign n77130 = ~n77087 & ~n77129 ;
  assign n77064 = ~n77057 & ~n77063 ;
  assign n77116 = ~n77064 & ~n77078 ;
  assign n77117 = n77070 & ~n77116 ;
  assign n77115 = ~n77057 & n77078 ;
  assign n77118 = n77087 & ~n77115 ;
  assign n77119 = n77117 & n77118 ;
  assign n77123 = ~n77070 & n77078 ;
  assign n77124 = n77063 & n77123 ;
  assign n77125 = ~n77057 & n77124 ;
  assign n77121 = n77063 & n77120 ;
  assign n77122 = n77057 & n77108 ;
  assign n77131 = ~n77121 & ~n77122 ;
  assign n77132 = ~n77125 & n77131 ;
  assign n77133 = ~n77119 & n77132 ;
  assign n77134 = ~n77130 & n77133 ;
  assign n77135 = n77051 & ~n77134 ;
  assign n77071 = n77064 & n77070 ;
  assign n77088 = ~n77071 & n77087 ;
  assign n77072 = n77063 & n77070 ;
  assign n77079 = n77072 & ~n77078 ;
  assign n77080 = ~n77063 & n77070 ;
  assign n77081 = n77057 & ~n77080 ;
  assign n77089 = ~n77079 & ~n77081 ;
  assign n77090 = n77088 & n77089 ;
  assign n77092 = ~n77070 & n77091 ;
  assign n77093 = n77063 & n77092 ;
  assign n77095 = ~n77078 & ~n77087 ;
  assign n77096 = n77094 & n77095 ;
  assign n77097 = n77063 & ~n77087 ;
  assign n77098 = n77057 & n77078 ;
  assign n77099 = n77097 & n77098 ;
  assign n77100 = ~n77096 & ~n77099 ;
  assign n77101 = ~n77093 & n77100 ;
  assign n77102 = ~n77090 & n77101 ;
  assign n77103 = ~n77051 & ~n77102 ;
  assign n77107 = ~n77057 & n77079 ;
  assign n77109 = n77098 & n77108 ;
  assign n77110 = ~n77107 & ~n77109 ;
  assign n77111 = ~n77087 & ~n77110 ;
  assign n77104 = ~n77057 & ~n77070 ;
  assign n77105 = n77063 & n77087 ;
  assign n77106 = n77104 & n77105 ;
  assign n77112 = ~n77063 & n77078 ;
  assign n77113 = ~n77087 & n77112 ;
  assign n77114 = n77094 & n77113 ;
  assign n77136 = ~n77106 & ~n77114 ;
  assign n77137 = ~n77111 & n77136 ;
  assign n77138 = ~n77103 & n77137 ;
  assign n77139 = ~n77135 & n77138 ;
  assign n77140 = \u2_L14_reg[27]/P0001  & n77139 ;
  assign n77141 = ~\u2_L14_reg[27]/P0001  & ~n77139 ;
  assign n77142 = ~n77140 & ~n77141 ;
  assign n77169 = decrypt_pad & ~\u2_uk_K_r14_reg[9]/NET0131  ;
  assign n77170 = ~decrypt_pad & ~\u2_uk_K_r14_reg[2]/NET0131  ;
  assign n77171 = ~n77169 & ~n77170 ;
  assign n77172 = \u2_R14_reg[23]/P0001  & ~n77171 ;
  assign n77173 = ~\u2_R14_reg[23]/P0001  & n77171 ;
  assign n77174 = ~n77172 & ~n77173 ;
  assign n77162 = decrypt_pad & ~\u2_uk_K_r14_reg[14]/NET0131  ;
  assign n77163 = ~decrypt_pad & ~\u2_uk_K_r14_reg[7]/NET0131  ;
  assign n77164 = ~n77162 & ~n77163 ;
  assign n77165 = \u2_R14_reg[20]/NET0131  & ~n77164 ;
  assign n77166 = ~\u2_R14_reg[20]/NET0131  & n77164 ;
  assign n77167 = ~n77165 & ~n77166 ;
  assign n77149 = decrypt_pad & ~\u2_uk_K_r14_reg[51]/NET0131  ;
  assign n77150 = ~decrypt_pad & ~\u2_uk_K_r14_reg[44]/NET0131  ;
  assign n77151 = ~n77149 & ~n77150 ;
  assign n77152 = \u2_R14_reg[22]/P0001  & ~n77151 ;
  assign n77153 = ~\u2_R14_reg[22]/P0001  & n77151 ;
  assign n77154 = ~n77152 & ~n77153 ;
  assign n77175 = decrypt_pad & ~\u2_uk_K_r14_reg[29]/NET0131  ;
  assign n77176 = ~decrypt_pad & ~\u2_uk_K_r14_reg[22]/NET0131  ;
  assign n77177 = ~n77175 & ~n77176 ;
  assign n77178 = \u2_R14_reg[21]/NET0131  & ~n77177 ;
  assign n77179 = ~\u2_R14_reg[21]/NET0131  & n77177 ;
  assign n77180 = ~n77178 & ~n77179 ;
  assign n77183 = ~n77154 & n77180 ;
  assign n77184 = n77167 & n77183 ;
  assign n77155 = decrypt_pad & ~\u2_uk_K_r14_reg[30]/NET0131  ;
  assign n77156 = ~decrypt_pad & ~\u2_uk_K_r14_reg[23]/NET0131  ;
  assign n77157 = ~n77155 & ~n77156 ;
  assign n77158 = \u2_R14_reg[25]/NET0131  & ~n77157 ;
  assign n77159 = ~\u2_R14_reg[25]/NET0131  & n77157 ;
  assign n77160 = ~n77158 & ~n77159 ;
  assign n77185 = n77160 & ~n77167 ;
  assign n77186 = ~n77180 & n77185 ;
  assign n77187 = ~n77184 & ~n77186 ;
  assign n77188 = n77174 & ~n77187 ;
  assign n77161 = ~n77154 & n77160 ;
  assign n77168 = ~n77161 & ~n77167 ;
  assign n77181 = ~n77174 & ~n77180 ;
  assign n77182 = ~n77168 & n77181 ;
  assign n77143 = decrypt_pad & ~\u2_uk_K_r14_reg[35]/P0001  ;
  assign n77144 = ~decrypt_pad & ~\u2_uk_K_r14_reg[28]/NET0131  ;
  assign n77145 = ~n77143 & ~n77144 ;
  assign n77146 = \u2_R14_reg[24]/NET0131  & ~n77145 ;
  assign n77147 = ~\u2_R14_reg[24]/NET0131  & n77145 ;
  assign n77148 = ~n77146 & ~n77147 ;
  assign n77189 = ~n77154 & ~n77160 ;
  assign n77190 = n77180 & n77189 ;
  assign n77191 = n77148 & ~n77190 ;
  assign n77192 = ~n77182 & n77191 ;
  assign n77193 = ~n77188 & n77192 ;
  assign n77197 = ~n77167 & ~n77180 ;
  assign n77198 = n77174 & ~n77185 ;
  assign n77199 = ~n77197 & n77198 ;
  assign n77200 = ~n77184 & n77199 ;
  assign n77194 = n77160 & n77167 ;
  assign n77195 = n77180 & n77194 ;
  assign n77196 = n77154 & n77195 ;
  assign n77201 = ~n77148 & ~n77196 ;
  assign n77202 = ~n77200 & n77201 ;
  assign n77203 = ~n77193 & ~n77202 ;
  assign n77216 = ~n77160 & n77167 ;
  assign n77217 = n77180 & n77216 ;
  assign n77218 = ~n77174 & ~n77217 ;
  assign n77215 = n77174 & ~n77186 ;
  assign n77219 = ~n77154 & ~n77215 ;
  assign n77220 = ~n77218 & n77219 ;
  assign n77204 = ~n77160 & n77197 ;
  assign n77205 = n77160 & n77180 ;
  assign n77206 = ~n77167 & n77205 ;
  assign n77207 = ~n77204 & ~n77206 ;
  assign n77208 = ~n77148 & ~n77174 ;
  assign n77209 = n77148 & n77154 ;
  assign n77210 = ~n77208 & ~n77209 ;
  assign n77211 = ~n77207 & ~n77210 ;
  assign n77212 = ~n77154 & ~n77174 ;
  assign n77213 = n77194 & n77212 ;
  assign n77214 = ~n77180 & n77213 ;
  assign n77221 = ~n77211 & ~n77214 ;
  assign n77222 = ~n77220 & n77221 ;
  assign n77223 = ~n77203 & n77222 ;
  assign n77224 = \u2_L14_reg[19]/P0001  & n77223 ;
  assign n77225 = ~\u2_L14_reg[19]/P0001  & ~n77223 ;
  assign n77226 = ~n77224 & ~n77225 ;
  assign n77227 = ~n77167 & n77180 ;
  assign n77231 = n77154 & ~n77227 ;
  assign n77232 = ~n77194 & n77231 ;
  assign n77228 = n77167 & ~n77180 ;
  assign n77229 = ~n77227 & ~n77228 ;
  assign n77230 = n77161 & ~n77229 ;
  assign n77233 = ~n77174 & ~n77230 ;
  assign n77234 = ~n77232 & n77233 ;
  assign n77237 = n77174 & ~n77195 ;
  assign n77235 = n77154 & n77227 ;
  assign n77236 = n77189 & n77228 ;
  assign n77238 = ~n77235 & ~n77236 ;
  assign n77239 = n77237 & n77238 ;
  assign n77240 = ~n77234 & ~n77239 ;
  assign n77241 = n77148 & ~n77240 ;
  assign n77242 = n77154 & n77228 ;
  assign n77246 = ~n77154 & ~n77167 ;
  assign n77247 = ~n77242 & ~n77246 ;
  assign n77248 = n77215 & n77247 ;
  assign n77249 = ~n77174 & ~n77184 ;
  assign n77250 = ~n77235 & n77249 ;
  assign n77251 = ~n77248 & ~n77250 ;
  assign n77244 = ~n77183 & ~n77212 ;
  assign n77245 = n77216 & ~n77244 ;
  assign n77243 = n77160 & n77242 ;
  assign n77252 = ~n77148 & ~n77243 ;
  assign n77253 = ~n77245 & n77252 ;
  assign n77254 = ~n77251 & n77253 ;
  assign n77255 = ~n77241 & ~n77254 ;
  assign n77256 = n77154 & n77194 ;
  assign n77257 = ~n77160 & n77227 ;
  assign n77258 = ~n77154 & n77257 ;
  assign n77259 = ~n77256 & ~n77258 ;
  assign n77260 = n77174 & ~n77259 ;
  assign n77261 = n77204 & n77212 ;
  assign n77262 = ~n77220 & ~n77261 ;
  assign n77263 = ~n77260 & n77262 ;
  assign n77264 = ~n77255 & n77263 ;
  assign n77265 = ~\u2_L14_reg[11]/P0001  & n77264 ;
  assign n77266 = \u2_L14_reg[11]/P0001  & ~n77264 ;
  assign n77267 = ~n77265 & ~n77266 ;
  assign n77271 = n76742 & n76810 ;
  assign n77272 = ~n76759 & ~n76765 ;
  assign n77269 = ~n76742 & n76765 ;
  assign n77273 = n76780 & n77269 ;
  assign n77274 = ~n76772 & ~n77273 ;
  assign n77275 = ~n77272 & n77274 ;
  assign n77276 = ~n77271 & n77275 ;
  assign n77277 = ~n76742 & n76757 ;
  assign n77278 = ~n76765 & n77277 ;
  assign n77279 = n76749 & n76755 ;
  assign n77280 = n76765 & n77279 ;
  assign n77281 = ~n77278 & ~n77280 ;
  assign n77282 = n76742 & ~n76755 ;
  assign n77283 = ~n76748 & n77282 ;
  assign n77284 = n76772 & ~n76807 ;
  assign n77285 = ~n77283 & n77284 ;
  assign n77286 = n77281 & n77285 ;
  assign n77287 = ~n77276 & ~n77286 ;
  assign n77268 = n76780 & n76783 ;
  assign n77270 = n76757 & n77269 ;
  assign n77288 = ~n77268 & ~n77270 ;
  assign n77289 = ~n77287 & n77288 ;
  assign n77290 = n76779 & ~n77289 ;
  assign n77291 = ~n76757 & n77269 ;
  assign n77292 = ~n76781 & ~n76796 ;
  assign n77293 = n77275 & n77292 ;
  assign n77294 = ~n76758 & n76812 ;
  assign n77295 = n77281 & n77294 ;
  assign n77296 = ~n77293 & ~n77295 ;
  assign n77297 = ~n77291 & ~n77296 ;
  assign n77298 = ~n76779 & ~n77297 ;
  assign n77299 = ~n77290 & ~n77298 ;
  assign n77300 = \u2_L14_reg[3]/P0001  & ~n77299 ;
  assign n77301 = ~\u2_L14_reg[3]/P0001  & n77299 ;
  assign n77302 = ~n77300 & ~n77301 ;
  assign n77306 = ~n76836 & ~n76883 ;
  assign n77307 = n76849 & ~n76862 ;
  assign n77308 = ~n77306 & n77307 ;
  assign n77309 = n76843 & ~n76863 ;
  assign n77310 = ~n77308 & n77309 ;
  assign n77312 = ~n77009 & n77306 ;
  assign n77311 = ~n76843 & ~n76875 ;
  assign n77313 = ~n76884 & n77311 ;
  assign n77314 = ~n77312 & n77313 ;
  assign n77315 = ~n77310 & ~n77314 ;
  assign n77303 = n76864 & n76880 ;
  assign n77316 = n76857 & ~n77303 ;
  assign n77304 = ~n76870 & n77014 ;
  assign n77305 = n76837 & n76874 ;
  assign n77317 = ~n77304 & ~n77305 ;
  assign n77318 = n77316 & n77317 ;
  assign n77319 = ~n77315 & n77318 ;
  assign n77320 = n76843 & ~n77312 ;
  assign n77321 = ~n76859 & ~n76882 ;
  assign n77322 = ~n77026 & n77321 ;
  assign n77323 = n77311 & n77322 ;
  assign n77324 = ~n77320 & ~n77323 ;
  assign n77325 = n76874 & n77028 ;
  assign n77326 = ~n76857 & ~n76884 ;
  assign n77327 = ~n77325 & n77326 ;
  assign n77328 = ~n77324 & n77327 ;
  assign n77329 = ~n77319 & ~n77328 ;
  assign n77330 = \u2_L14_reg[28]/P0001  & ~n77329 ;
  assign n77331 = ~\u2_L14_reg[28]/P0001  & n77329 ;
  assign n77332 = ~n77330 & ~n77331 ;
  assign n77343 = ~n76948 & ~n76965 ;
  assign n77338 = ~n76953 & ~n76955 ;
  assign n77339 = n76974 & ~n77338 ;
  assign n77344 = n76939 & ~n76991 ;
  assign n77345 = ~n77339 & n77344 ;
  assign n77340 = ~n76925 & n76981 ;
  assign n77341 = ~n76912 & n76918 ;
  assign n77342 = n76980 & n77341 ;
  assign n77346 = ~n77340 & ~n77342 ;
  assign n77347 = n77345 & n77346 ;
  assign n77348 = n77343 & n77347 ;
  assign n77357 = ~n76957 & ~n76979 ;
  assign n77349 = ~n76925 & n76945 ;
  assign n77350 = n76912 & ~n77349 ;
  assign n77351 = ~n76953 & ~n76961 ;
  assign n77352 = n77350 & n77351 ;
  assign n77358 = ~n76987 & ~n77352 ;
  assign n77359 = n77357 & n77358 ;
  assign n77353 = n76918 & n76961 ;
  assign n77354 = ~n77349 & ~n77353 ;
  assign n77355 = ~n76912 & ~n77354 ;
  assign n77356 = ~n76933 & ~n76939 ;
  assign n77360 = ~n77355 & n77356 ;
  assign n77361 = n77359 & n77360 ;
  assign n77362 = ~n77348 & ~n77361 ;
  assign n77333 = n76960 & n76961 ;
  assign n77334 = n76949 & n76961 ;
  assign n77335 = ~n77333 & ~n77334 ;
  assign n77336 = ~n76987 & n77335 ;
  assign n77337 = n76912 & ~n77336 ;
  assign n77363 = n76953 & n76975 ;
  assign n77364 = ~n77337 & ~n77363 ;
  assign n77365 = ~n77362 & n77364 ;
  assign n77366 = ~\u2_L14_reg[20]/P0001  & ~n77365 ;
  assign n77367 = \u2_L14_reg[20]/P0001  & n77365 ;
  assign n77368 = ~n77366 & ~n77367 ;
  assign n77369 = decrypt_pad & ~\u2_uk_K_r14_reg[2]/NET0131  ;
  assign n77370 = ~decrypt_pad & ~\u2_uk_K_r14_reg[50]/NET0131  ;
  assign n77371 = ~n77369 & ~n77370 ;
  assign n77372 = \u2_R14_reg[24]/NET0131  & ~n77371 ;
  assign n77373 = ~\u2_R14_reg[24]/NET0131  & n77371 ;
  assign n77374 = ~n77372 & ~n77373 ;
  assign n77375 = decrypt_pad & ~\u2_uk_K_r14_reg[37]/NET0131  ;
  assign n77376 = ~decrypt_pad & ~\u2_uk_K_r14_reg[30]/NET0131  ;
  assign n77377 = ~n77375 & ~n77376 ;
  assign n77378 = \u2_R14_reg[25]/NET0131  & ~n77377 ;
  assign n77379 = ~\u2_R14_reg[25]/NET0131  & n77377 ;
  assign n77380 = ~n77378 & ~n77379 ;
  assign n77381 = n77374 & n77380 ;
  assign n77384 = decrypt_pad & ~\u2_uk_K_r14_reg[22]/NET0131  ;
  assign n77385 = ~decrypt_pad & ~\u2_uk_K_r14_reg[15]/NET0131  ;
  assign n77386 = ~n77384 & ~n77385 ;
  assign n77387 = \u2_R14_reg[26]/P0001  & ~n77386 ;
  assign n77388 = ~\u2_R14_reg[26]/P0001  & n77386 ;
  assign n77389 = ~n77387 & ~n77388 ;
  assign n77408 = ~n77380 & ~n77389 ;
  assign n77390 = decrypt_pad & ~\u2_uk_K_r14_reg[38]/NET0131  ;
  assign n77391 = ~decrypt_pad & ~\u2_uk_K_r14_reg[31]/NET0131  ;
  assign n77392 = ~n77390 & ~n77391 ;
  assign n77393 = \u2_R14_reg[29]/NET0131  & ~n77392 ;
  assign n77394 = ~\u2_R14_reg[29]/NET0131  & n77392 ;
  assign n77395 = ~n77393 & ~n77394 ;
  assign n77410 = ~n77374 & ~n77395 ;
  assign n77411 = n77408 & n77410 ;
  assign n77412 = ~n77381 & ~n77411 ;
  assign n77413 = decrypt_pad & ~\u2_uk_K_r14_reg[0]/NET0131  ;
  assign n77414 = ~decrypt_pad & ~\u2_uk_K_r14_reg[52]/NET0131  ;
  assign n77415 = ~n77413 & ~n77414 ;
  assign n77416 = \u2_R14_reg[27]/P0001  & ~n77415 ;
  assign n77417 = ~\u2_R14_reg[27]/P0001  & n77415 ;
  assign n77418 = ~n77416 & ~n77417 ;
  assign n77419 = ~n77412 & n77418 ;
  assign n77382 = ~n77374 & ~n77380 ;
  assign n77383 = ~n77381 & ~n77382 ;
  assign n77396 = n77389 & ~n77395 ;
  assign n77397 = n77383 & n77396 ;
  assign n77398 = decrypt_pad & ~\u2_uk_K_r14_reg[42]/P0001  ;
  assign n77399 = ~decrypt_pad & ~\u2_uk_K_r14_reg[35]/P0001  ;
  assign n77400 = ~n77398 & ~n77399 ;
  assign n77401 = \u2_R14_reg[28]/NET0131  & ~n77400 ;
  assign n77402 = ~\u2_R14_reg[28]/NET0131  & n77400 ;
  assign n77403 = ~n77401 & ~n77402 ;
  assign n77407 = n77374 & n77395 ;
  assign n77409 = n77407 & n77408 ;
  assign n77423 = n77403 & ~n77409 ;
  assign n77424 = ~n77397 & n77423 ;
  assign n77404 = n77380 & n77395 ;
  assign n77405 = ~n77374 & n77404 ;
  assign n77406 = ~n77389 & n77405 ;
  assign n77420 = n77389 & n77395 ;
  assign n77421 = n77382 & n77420 ;
  assign n77422 = ~n77418 & n77421 ;
  assign n77425 = ~n77406 & ~n77422 ;
  assign n77426 = n77424 & n77425 ;
  assign n77427 = ~n77419 & n77426 ;
  assign n77431 = n77383 & n77420 ;
  assign n77428 = n77380 & n77389 ;
  assign n77429 = ~n77408 & ~n77428 ;
  assign n77430 = n77410 & n77429 ;
  assign n77444 = ~n77403 & ~n77430 ;
  assign n77445 = ~n77431 & n77444 ;
  assign n77432 = n77374 & n77389 ;
  assign n77433 = ~n77380 & ~n77395 ;
  assign n77434 = ~n77404 & ~n77433 ;
  assign n77435 = ~n77432 & n77434 ;
  assign n77436 = ~n77418 & ~n77435 ;
  assign n77438 = n77374 & ~n77389 ;
  assign n77439 = ~n77395 & n77438 ;
  assign n77440 = ~n77418 & ~n77439 ;
  assign n77437 = ~n77407 & ~n77410 ;
  assign n77441 = ~n77380 & ~n77432 ;
  assign n77442 = n77437 & n77441 ;
  assign n77443 = ~n77440 & n77442 ;
  assign n77446 = ~n77436 & ~n77443 ;
  assign n77447 = n77445 & n77446 ;
  assign n77448 = ~n77427 & ~n77447 ;
  assign n77449 = \u2_L14_reg[12]/P0001  & n77448 ;
  assign n77450 = ~\u2_L14_reg[12]/P0001  & ~n77448 ;
  assign n77451 = ~n77449 & ~n77450 ;
  assign n77471 = decrypt_pad & ~\u2_uk_K_r14_reg[11]/NET0131  ;
  assign n77472 = ~decrypt_pad & ~\u2_uk_K_r14_reg[4]/NET0131  ;
  assign n77473 = ~n77471 & ~n77472 ;
  assign n77474 = \u2_R14_reg[1]/NET0131  & ~n77473 ;
  assign n77475 = ~\u2_R14_reg[1]/NET0131  & n77473 ;
  assign n77476 = ~n77474 & ~n77475 ;
  assign n77458 = decrypt_pad & ~\u2_uk_K_r14_reg[41]/NET0131  ;
  assign n77459 = ~decrypt_pad & ~\u2_uk_K_r14_reg[34]/NET0131  ;
  assign n77460 = ~n77458 & ~n77459 ;
  assign n77461 = \u2_R14_reg[5]/NET0131  & ~n77460 ;
  assign n77462 = ~\u2_R14_reg[5]/NET0131  & n77460 ;
  assign n77463 = ~n77461 & ~n77462 ;
  assign n77464 = decrypt_pad & ~\u2_uk_K_r14_reg[47]/NET0131  ;
  assign n77465 = ~decrypt_pad & ~\u2_uk_K_r14_reg[40]/NET0131  ;
  assign n77466 = ~n77464 & ~n77465 ;
  assign n77467 = \u2_R14_reg[32]/NET0131  & ~n77466 ;
  assign n77468 = ~\u2_R14_reg[32]/NET0131  & n77466 ;
  assign n77469 = ~n77467 & ~n77468 ;
  assign n77477 = decrypt_pad & ~\u2_uk_K_r14_reg[26]/NET0131  ;
  assign n77478 = ~decrypt_pad & ~\u2_uk_K_r14_reg[19]/NET0131  ;
  assign n77479 = ~n77477 & ~n77478 ;
  assign n77480 = \u2_R14_reg[2]/NET0131  & ~n77479 ;
  assign n77481 = ~\u2_R14_reg[2]/NET0131  & n77479 ;
  assign n77482 = ~n77480 & ~n77481 ;
  assign n77485 = ~n77469 & n77482 ;
  assign n77494 = ~n77463 & n77485 ;
  assign n77495 = n77463 & ~n77469 ;
  assign n77496 = ~n77482 & n77495 ;
  assign n77497 = ~n77494 & ~n77496 ;
  assign n77498 = n77476 & ~n77497 ;
  assign n77489 = ~n77463 & ~n77476 ;
  assign n77490 = n77469 & n77489 ;
  assign n77491 = n77469 & n77476 ;
  assign n77492 = n77463 & n77491 ;
  assign n77493 = ~n77490 & ~n77492 ;
  assign n77499 = decrypt_pad & ~\u2_uk_K_r14_reg[3]/NET0131  ;
  assign n77500 = ~decrypt_pad & ~\u2_uk_K_r14_reg[53]/NET0131  ;
  assign n77501 = ~n77499 & ~n77500 ;
  assign n77502 = \u2_R14_reg[3]/NET0131  & ~n77501 ;
  assign n77503 = ~\u2_R14_reg[3]/NET0131  & n77501 ;
  assign n77504 = ~n77502 & ~n77503 ;
  assign n77505 = n77493 & n77504 ;
  assign n77506 = ~n77498 & n77505 ;
  assign n77470 = ~n77463 & ~n77469 ;
  assign n77507 = n77463 & n77469 ;
  assign n77508 = ~n77470 & ~n77507 ;
  assign n77509 = ~n77476 & ~n77508 ;
  assign n77510 = ~n77469 & ~n77482 ;
  assign n77511 = ~n77463 & n77510 ;
  assign n77512 = ~n77504 & ~n77511 ;
  assign n77513 = ~n77509 & n77512 ;
  assign n77514 = ~n77506 & ~n77513 ;
  assign n77452 = decrypt_pad & ~\u2_uk_K_r14_reg[13]/NET0131  ;
  assign n77453 = ~decrypt_pad & ~\u2_uk_K_r14_reg[6]/NET0131  ;
  assign n77454 = ~n77452 & ~n77453 ;
  assign n77455 = \u2_R14_reg[4]/NET0131  & ~n77454 ;
  assign n77456 = ~\u2_R14_reg[4]/NET0131  & n77454 ;
  assign n77457 = ~n77455 & ~n77456 ;
  assign n77483 = n77476 & n77482 ;
  assign n77484 = ~n77463 & n77483 ;
  assign n77486 = ~n77476 & n77485 ;
  assign n77487 = ~n77484 & ~n77486 ;
  assign n77488 = ~n77470 & ~n77487 ;
  assign n77515 = ~n77457 & ~n77488 ;
  assign n77516 = ~n77514 & n77515 ;
  assign n77518 = ~n77476 & n77510 ;
  assign n77517 = n77469 & n77482 ;
  assign n77519 = ~n77504 & ~n77517 ;
  assign n77520 = ~n77518 & n77519 ;
  assign n77521 = ~n77476 & ~n77482 ;
  assign n77523 = n77469 & n77521 ;
  assign n77524 = n77463 & n77523 ;
  assign n77522 = ~n77469 & ~n77521 ;
  assign n77525 = n77504 & ~n77522 ;
  assign n77526 = ~n77524 & n77525 ;
  assign n77527 = ~n77520 & ~n77526 ;
  assign n77528 = ~n77463 & n77491 ;
  assign n77529 = ~n77482 & n77528 ;
  assign n77530 = n77463 & n77483 ;
  assign n77531 = n77457 & ~n77530 ;
  assign n77532 = ~n77529 & n77531 ;
  assign n77533 = ~n77527 & n77532 ;
  assign n77534 = ~n77516 & ~n77533 ;
  assign n77535 = ~\u2_L14_reg[17]/P0001  & n77534 ;
  assign n77536 = \u2_L14_reg[17]/P0001  & ~n77534 ;
  assign n77537 = ~n77535 & ~n77536 ;
  assign n77538 = n77174 & ~n77217 ;
  assign n77539 = n77160 & ~n77247 ;
  assign n77540 = n77538 & ~n77539 ;
  assign n77541 = n77154 & n77186 ;
  assign n77542 = ~n77174 & ~n77257 ;
  assign n77543 = ~n77541 & n77542 ;
  assign n77544 = ~n77540 & ~n77543 ;
  assign n77545 = ~n77213 & ~n77236 ;
  assign n77546 = ~n77544 & n77545 ;
  assign n77547 = ~n77148 & ~n77546 ;
  assign n77559 = ~n77190 & ~n77246 ;
  assign n77560 = ~n77174 & ~n77559 ;
  assign n77556 = n77154 & n77205 ;
  assign n77557 = ~n77154 & n77174 ;
  assign n77558 = n77194 & n77557 ;
  assign n77561 = ~n77556 & ~n77558 ;
  assign n77562 = ~n77258 & n77561 ;
  assign n77563 = ~n77560 & n77562 ;
  assign n77564 = n77148 & ~n77563 ;
  assign n77551 = n77207 & n77538 ;
  assign n77548 = ~n77180 & n77216 ;
  assign n77549 = ~n77195 & ~n77548 ;
  assign n77550 = ~n77174 & n77549 ;
  assign n77552 = n77154 & ~n77550 ;
  assign n77553 = ~n77551 & n77552 ;
  assign n77554 = ~n77167 & ~n77174 ;
  assign n77555 = n77189 & n77554 ;
  assign n77565 = ~n77553 & ~n77555 ;
  assign n77566 = ~n77564 & n77565 ;
  assign n77567 = ~n77547 & n77566 ;
  assign n77568 = \u2_L14_reg[4]/P0001  & n77567 ;
  assign n77569 = ~\u2_L14_reg[4]/P0001  & ~n77567 ;
  assign n77570 = ~n77568 & ~n77569 ;
  assign n77583 = ~n77180 & ~n77189 ;
  assign n77584 = n77174 & ~n77583 ;
  assign n77572 = ~n77154 & ~n77197 ;
  assign n77573 = ~n77216 & n77572 ;
  assign n77581 = ~n77185 & ~n77216 ;
  assign n77582 = n77154 & ~n77581 ;
  assign n77585 = ~n77573 & ~n77582 ;
  assign n77586 = ~n77584 & n77585 ;
  assign n77571 = n77154 & n77217 ;
  assign n77577 = n77154 & ~n77160 ;
  assign n77578 = n77227 & ~n77577 ;
  assign n77579 = ~n77571 & ~n77578 ;
  assign n77580 = n77174 & ~n77579 ;
  assign n77587 = n77148 & ~n77580 ;
  assign n77588 = ~n77586 & n77587 ;
  assign n77589 = ~n77160 & ~n77183 ;
  assign n77590 = ~n77231 & n77589 ;
  assign n77591 = n77549 & ~n77590 ;
  assign n77592 = n77174 & ~n77591 ;
  assign n77593 = ~n77148 & ~n77541 ;
  assign n77594 = ~n77592 & n77593 ;
  assign n77595 = ~n77588 & ~n77594 ;
  assign n77574 = ~n77571 & ~n77573 ;
  assign n77575 = n77208 & ~n77574 ;
  assign n77576 = n77205 & n77557 ;
  assign n77596 = ~n77236 & ~n77576 ;
  assign n77597 = ~n77575 & n77596 ;
  assign n77598 = ~n77595 & n77597 ;
  assign n77599 = ~\u2_L14_reg[29]/P0001  & n77598 ;
  assign n77600 = \u2_L14_reg[29]/P0001  & ~n77598 ;
  assign n77601 = ~n77599 & ~n77600 ;
  assign n77609 = n77057 & n77124 ;
  assign n77610 = ~n77064 & ~n77087 ;
  assign n77611 = ~n77095 & ~n77610 ;
  assign n77612 = ~n77609 & ~n77611 ;
  assign n77614 = n77087 & ~n77120 ;
  assign n77613 = n77072 & n77078 ;
  assign n77615 = ~n77122 & ~n77613 ;
  assign n77616 = n77614 & n77615 ;
  assign n77617 = ~n77612 & ~n77616 ;
  assign n77606 = ~n77078 & n77104 ;
  assign n77607 = ~n77126 & ~n77606 ;
  assign n77608 = n77063 & ~n77607 ;
  assign n77605 = ~n77063 & n77092 ;
  assign n77618 = n77051 & ~n77605 ;
  assign n77619 = ~n77608 & n77618 ;
  assign n77620 = ~n77617 & n77619 ;
  assign n77626 = ~n77051 & ~n77079 ;
  assign n77629 = ~n77125 & n77626 ;
  assign n77602 = n77057 & n77113 ;
  assign n77625 = ~n77063 & n77606 ;
  assign n77630 = ~n77602 & ~n77625 ;
  assign n77631 = n77629 & n77630 ;
  assign n77621 = ~n77124 & ~n77126 ;
  assign n77622 = n77087 & ~n77621 ;
  assign n77624 = n77080 & n77098 ;
  assign n77623 = n77091 & n77097 ;
  assign n77627 = ~n77096 & ~n77623 ;
  assign n77628 = ~n77624 & n77627 ;
  assign n77632 = ~n77622 & n77628 ;
  assign n77633 = n77631 & n77632 ;
  assign n77634 = ~n77620 & ~n77633 ;
  assign n77603 = n77070 & n77602 ;
  assign n77604 = n77087 & n77127 ;
  assign n77635 = ~n77603 & ~n77604 ;
  assign n77636 = ~n77634 & n77635 ;
  assign n77637 = \u2_L14_reg[21]/P0001  & n77636 ;
  assign n77638 = ~\u2_L14_reg[21]/P0001  & ~n77636 ;
  assign n77639 = ~n77637 & ~n77638 ;
  assign n77640 = ~n76884 & ~n77025 ;
  assign n77641 = ~n76896 & ~n77305 ;
  assign n77642 = ~n77027 & n77641 ;
  assign n77643 = ~n76857 & ~n77642 ;
  assign n77644 = n77640 & ~n77643 ;
  assign n77645 = ~n76843 & ~n77644 ;
  assign n77646 = ~n76837 & ~n76849 ;
  assign n77647 = ~n77026 & n77646 ;
  assign n77648 = ~n76898 & ~n77647 ;
  assign n77649 = n76843 & ~n77648 ;
  assign n77651 = n76837 & ~n76870 ;
  assign n77652 = ~n77034 & n77651 ;
  assign n77650 = n76858 & n77304 ;
  assign n77653 = ~n76857 & ~n77650 ;
  assign n77654 = ~n77652 & n77653 ;
  assign n77655 = ~n77649 & n77654 ;
  assign n77658 = ~n76864 & ~n76883 ;
  assign n77659 = n77034 & ~n77658 ;
  assign n77660 = n76857 & ~n76897 ;
  assign n77661 = ~n77659 & n77660 ;
  assign n77656 = ~n76881 & ~n77001 ;
  assign n77657 = n76843 & ~n77656 ;
  assign n77662 = n77020 & n77640 ;
  assign n77663 = ~n77657 & n77662 ;
  assign n77664 = n77661 & n77663 ;
  assign n77665 = ~n77655 & ~n77664 ;
  assign n77666 = ~n77645 & ~n77665 ;
  assign n77667 = \u2_L14_reg[13]/P0001  & ~n77666 ;
  assign n77668 = ~\u2_L14_reg[13]/P0001  & n77666 ;
  assign n77669 = ~n77667 & ~n77668 ;
  assign n77675 = ~n77092 & ~n77125 ;
  assign n77676 = n77087 & ~n77675 ;
  assign n77671 = n77057 & ~n77070 ;
  assign n77672 = n77610 & ~n77671 ;
  assign n77673 = ~n77613 & ~n77672 ;
  assign n77674 = ~n77115 & ~n77673 ;
  assign n77670 = n77094 & n77112 ;
  assign n77677 = ~n77113 & ~n77670 ;
  assign n77678 = ~n77674 & n77677 ;
  assign n77679 = ~n77676 & n77678 ;
  assign n77680 = ~n77051 & ~n77679 ;
  assign n77685 = ~n77094 & ~n77112 ;
  assign n77686 = ~n77670 & ~n77685 ;
  assign n77687 = n77087 & ~n77686 ;
  assign n77688 = ~n77087 & ~n77124 ;
  assign n77689 = ~n77127 & n77688 ;
  assign n77690 = ~n77687 & ~n77689 ;
  assign n77691 = ~n77121 & ~n77690 ;
  assign n77692 = n77051 & ~n77691 ;
  assign n77681 = ~n77107 & ~n77625 ;
  assign n77682 = ~n77093 & ~n77109 ;
  assign n77683 = n77681 & n77682 ;
  assign n77684 = n77087 & ~n77683 ;
  assign n77693 = ~n77114 & ~n77684 ;
  assign n77694 = ~n77692 & n77693 ;
  assign n77695 = ~n77680 & n77694 ;
  assign n77696 = ~\u2_L14_reg[5]/P0001  & n77695 ;
  assign n77697 = \u2_L14_reg[5]/P0001  & ~n77695 ;
  assign n77698 = ~n77696 & ~n77697 ;
  assign n77699 = decrypt_pad & ~\u2_uk_K_r14_reg[17]/NET0131  ;
  assign n77700 = ~decrypt_pad & ~\u2_uk_K_r14_reg[10]/P0001  ;
  assign n77701 = ~n77699 & ~n77700 ;
  assign n77702 = \u2_R14_reg[12]/NET0131  & ~n77701 ;
  assign n77703 = ~\u2_R14_reg[12]/NET0131  & n77701 ;
  assign n77704 = ~n77702 & ~n77703 ;
  assign n77712 = decrypt_pad & ~\u2_uk_K_r14_reg[53]/NET0131  ;
  assign n77713 = ~decrypt_pad & ~\u2_uk_K_r14_reg[46]/NET0131  ;
  assign n77714 = ~n77712 & ~n77713 ;
  assign n77715 = \u2_R14_reg[8]/NET0131  & ~n77714 ;
  assign n77716 = ~\u2_R14_reg[8]/NET0131  & n77714 ;
  assign n77717 = ~n77715 & ~n77716 ;
  assign n77725 = decrypt_pad & ~\u2_uk_K_r14_reg[33]/NET0131  ;
  assign n77726 = ~decrypt_pad & ~\u2_uk_K_r14_reg[26]/NET0131  ;
  assign n77727 = ~n77725 & ~n77726 ;
  assign n77728 = \u2_R14_reg[10]/P0001  & ~n77727 ;
  assign n77729 = ~\u2_R14_reg[10]/P0001  & n77727 ;
  assign n77730 = ~n77728 & ~n77729 ;
  assign n77746 = n77717 & n77730 ;
  assign n77718 = decrypt_pad & ~\u2_uk_K_r14_reg[5]/NET0131  ;
  assign n77719 = ~decrypt_pad & ~\u2_uk_K_r14_reg[55]/NET0131  ;
  assign n77720 = ~n77718 & ~n77719 ;
  assign n77721 = \u2_R14_reg[13]/NET0131  & ~n77720 ;
  assign n77722 = ~\u2_R14_reg[13]/NET0131  & n77720 ;
  assign n77723 = ~n77721 & ~n77722 ;
  assign n77735 = decrypt_pad & ~\u2_uk_K_r14_reg[25]/NET0131  ;
  assign n77736 = ~decrypt_pad & ~\u2_uk_K_r14_reg[18]/NET0131  ;
  assign n77737 = ~n77735 & ~n77736 ;
  assign n77738 = \u2_R14_reg[9]/NET0131  & ~n77737 ;
  assign n77739 = ~\u2_R14_reg[9]/NET0131  & n77737 ;
  assign n77740 = ~n77738 & ~n77739 ;
  assign n77758 = n77723 & ~n77740 ;
  assign n77759 = n77730 & n77758 ;
  assign n77705 = decrypt_pad & ~\u2_uk_K_r14_reg[34]/NET0131  ;
  assign n77706 = ~decrypt_pad & ~\u2_uk_K_r14_reg[27]/NET0131  ;
  assign n77707 = ~n77705 & ~n77706 ;
  assign n77708 = \u2_R14_reg[11]/P0001  & ~n77707 ;
  assign n77709 = ~\u2_R14_reg[11]/P0001  & n77707 ;
  assign n77710 = ~n77708 & ~n77709 ;
  assign n77755 = ~n77723 & n77740 ;
  assign n77764 = ~n77717 & ~n77740 ;
  assign n77765 = ~n77755 & ~n77764 ;
  assign n77766 = ~n77710 & n77765 ;
  assign n77767 = ~n77759 & ~n77766 ;
  assign n77768 = ~n77746 & ~n77767 ;
  assign n77742 = n77717 & ~n77723 ;
  assign n77724 = ~n77717 & n77723 ;
  assign n77741 = ~n77730 & ~n77740 ;
  assign n77762 = ~n77724 & n77741 ;
  assign n77763 = ~n77742 & n77762 ;
  assign n77769 = n77746 & ~n77755 ;
  assign n77770 = ~n77730 & n77740 ;
  assign n77771 = ~n77723 & n77770 ;
  assign n77772 = ~n77769 & ~n77771 ;
  assign n77773 = n77710 & ~n77772 ;
  assign n77774 = ~n77763 & ~n77773 ;
  assign n77775 = ~n77768 & n77774 ;
  assign n77776 = ~n77704 & ~n77775 ;
  assign n77711 = n77704 & n77710 ;
  assign n77731 = n77724 & ~n77730 ;
  assign n77732 = ~n77717 & ~n77723 ;
  assign n77733 = n77730 & n77732 ;
  assign n77734 = ~n77731 & ~n77733 ;
  assign n77743 = n77741 & n77742 ;
  assign n77744 = n77734 & ~n77743 ;
  assign n77745 = n77711 & ~n77744 ;
  assign n77747 = n77732 & n77740 ;
  assign n77748 = ~n77746 & ~n77747 ;
  assign n77749 = n77704 & ~n77710 ;
  assign n77750 = ~n77748 & n77749 ;
  assign n77760 = n77710 & n77717 ;
  assign n77761 = n77759 & n77760 ;
  assign n77751 = n77717 & n77723 ;
  assign n77752 = n77730 & n77740 ;
  assign n77753 = n77704 & n77752 ;
  assign n77754 = ~n77751 & n77753 ;
  assign n77756 = ~n77710 & n77730 ;
  assign n77757 = n77755 & n77756 ;
  assign n77777 = ~n77754 & ~n77757 ;
  assign n77778 = ~n77761 & n77777 ;
  assign n77779 = ~n77750 & n77778 ;
  assign n77780 = ~n77745 & n77779 ;
  assign n77781 = ~n77776 & n77780 ;
  assign n77782 = ~\u2_L14_reg[30]/P0001  & n77781 ;
  assign n77783 = \u2_L14_reg[30]/P0001  & ~n77781 ;
  assign n77784 = ~n77782 & ~n77783 ;
  assign n77808 = ~n77380 & n77410 ;
  assign n77809 = n77389 & n77808 ;
  assign n77806 = n77432 & ~n77433 ;
  assign n77807 = ~n77389 & n77437 ;
  assign n77810 = ~n77806 & ~n77807 ;
  assign n77811 = ~n77809 & n77810 ;
  assign n77812 = ~n77418 & ~n77811 ;
  assign n77813 = n77374 & ~n77380 ;
  assign n77814 = n77418 & n77813 ;
  assign n77815 = ~n77405 & ~n77814 ;
  assign n77816 = ~n77389 & ~n77815 ;
  assign n77817 = n77381 & n77420 ;
  assign n77818 = ~n77816 & ~n77817 ;
  assign n77819 = ~n77812 & n77818 ;
  assign n77820 = ~n77403 & ~n77819 ;
  assign n77798 = n77404 & n77438 ;
  assign n77799 = ~n77380 & n77432 ;
  assign n77800 = ~n77798 & ~n77799 ;
  assign n77801 = n77418 & ~n77800 ;
  assign n77796 = ~n77405 & ~n77409 ;
  assign n77797 = ~n77418 & ~n77796 ;
  assign n77802 = ~n77411 & ~n77421 ;
  assign n77803 = ~n77797 & n77802 ;
  assign n77804 = ~n77801 & n77803 ;
  assign n77805 = n77403 & ~n77804 ;
  assign n77785 = n77410 & n77428 ;
  assign n77786 = ~n77421 & ~n77785 ;
  assign n77787 = n77374 & n77433 ;
  assign n77788 = n77786 & ~n77787 ;
  assign n77789 = n77418 & ~n77788 ;
  assign n77790 = ~n77389 & n77418 ;
  assign n77791 = n77433 & n77790 ;
  assign n77792 = ~n77374 & ~n77389 ;
  assign n77793 = ~n77432 & ~n77792 ;
  assign n77794 = n77380 & ~n77418 ;
  assign n77795 = ~n77793 & n77794 ;
  assign n77821 = ~n77791 & ~n77795 ;
  assign n77822 = ~n77789 & n77821 ;
  assign n77823 = ~n77805 & n77822 ;
  assign n77824 = ~n77820 & n77823 ;
  assign n77825 = ~\u2_L14_reg[22]/P0001  & ~n77824 ;
  assign n77826 = \u2_L14_reg[22]/P0001  & n77824 ;
  assign n77827 = ~n77825 & ~n77826 ;
  assign n77844 = ~n76756 & n76772 ;
  assign n77843 = n76755 & n76788 ;
  assign n77845 = ~n76784 & ~n77843 ;
  assign n77846 = n77844 & n77845 ;
  assign n77848 = ~n76772 & ~n77268 ;
  assign n77847 = n76765 & n77282 ;
  assign n77849 = ~n77279 & ~n77847 ;
  assign n77850 = n77848 & n77849 ;
  assign n77851 = ~n77278 & n77850 ;
  assign n77852 = ~n77846 & ~n77851 ;
  assign n77853 = ~n76755 & n76784 ;
  assign n77854 = ~n77273 & ~n77853 ;
  assign n77855 = ~n77852 & n77854 ;
  assign n77856 = ~n76779 & ~n77855 ;
  assign n77829 = ~n76756 & ~n77271 ;
  assign n77830 = ~n76772 & ~n77829 ;
  assign n77828 = ~n76758 & ~n76765 ;
  assign n77831 = ~n76781 & n77828 ;
  assign n77832 = ~n77830 & n77831 ;
  assign n77833 = ~n76772 & n76786 ;
  assign n77834 = n76765 & ~n77277 ;
  assign n77835 = ~n77833 & n77834 ;
  assign n77836 = ~n77832 & ~n77835 ;
  assign n77837 = ~n76783 & n76810 ;
  assign n77838 = ~n76758 & ~n76807 ;
  assign n77839 = ~n77837 & n77838 ;
  assign n77840 = n76772 & ~n77839 ;
  assign n77841 = ~n77836 & ~n77840 ;
  assign n77842 = n76779 & ~n77841 ;
  assign n77857 = ~n76756 & n76765 ;
  assign n77858 = ~n77828 & ~n77857 ;
  assign n77859 = n76772 & ~n77858 ;
  assign n77860 = ~n77280 & ~n77847 ;
  assign n77861 = ~n76748 & ~n77860 ;
  assign n77862 = ~n76772 & ~n77861 ;
  assign n77863 = ~n77859 & ~n77862 ;
  assign n77864 = ~n77842 & ~n77863 ;
  assign n77865 = ~n77856 & n77864 ;
  assign n77866 = \u2_L14_reg[14]/P0001  & n77865 ;
  assign n77867 = ~\u2_L14_reg[14]/P0001  & ~n77865 ;
  assign n77868 = ~n77866 & ~n77867 ;
  assign n77883 = ~n77724 & ~n77742 ;
  assign n77888 = ~n77741 & n77883 ;
  assign n77889 = ~n77752 & n77888 ;
  assign n77886 = n77724 & n77752 ;
  assign n77887 = ~n77710 & n77886 ;
  assign n77882 = n77710 & ~n77717 ;
  assign n77884 = n77741 & ~n77882 ;
  assign n77885 = ~n77883 & n77884 ;
  assign n77890 = n77770 & n77882 ;
  assign n77891 = n77746 & n77755 ;
  assign n77892 = ~n77890 & ~n77891 ;
  assign n77893 = ~n77885 & n77892 ;
  assign n77894 = ~n77887 & n77893 ;
  assign n77895 = ~n77889 & n77894 ;
  assign n77896 = ~n77704 & ~n77895 ;
  assign n77875 = ~n77730 & n77732 ;
  assign n77876 = ~n77740 & n77875 ;
  assign n77877 = ~n77759 & ~n77876 ;
  assign n77878 = n77710 & ~n77877 ;
  assign n77869 = n77724 & n77730 ;
  assign n77870 = ~n77755 & ~n77758 ;
  assign n77871 = ~n77732 & ~n77870 ;
  assign n77872 = ~n77869 & ~n77871 ;
  assign n77873 = n77711 & ~n77872 ;
  assign n77874 = n77732 & n77753 ;
  assign n77879 = ~n77717 & ~n77770 ;
  assign n77880 = n77749 & n77870 ;
  assign n77881 = ~n77879 & n77880 ;
  assign n77897 = ~n77874 & ~n77881 ;
  assign n77898 = ~n77873 & n77897 ;
  assign n77899 = ~n77878 & n77898 ;
  assign n77900 = ~n77896 & n77899 ;
  assign n77901 = \u2_L14_reg[6]/P0001  & n77900 ;
  assign n77902 = ~\u2_L14_reg[6]/P0001  & ~n77900 ;
  assign n77903 = ~n77901 & ~n77902 ;
  assign n77915 = ~n77482 & n77504 ;
  assign n77916 = n77476 & ~n77915 ;
  assign n77917 = n77463 & ~n77916 ;
  assign n77918 = ~n77523 & ~n77917 ;
  assign n77919 = ~n77507 & ~n77918 ;
  assign n77912 = n77463 & ~n77476 ;
  assign n77913 = ~n77494 & ~n77912 ;
  assign n77914 = n77504 & ~n77913 ;
  assign n77920 = n77491 & ~n77504 ;
  assign n77921 = n77457 & ~n77486 ;
  assign n77922 = ~n77920 & n77921 ;
  assign n77923 = ~n77914 & n77922 ;
  assign n77924 = ~n77919 & n77923 ;
  assign n77934 = ~n77521 & ~n77915 ;
  assign n77935 = n77507 & ~n77934 ;
  assign n77929 = n77482 & n77504 ;
  assign n77930 = n77528 & n77929 ;
  assign n77936 = ~n77457 & ~n77930 ;
  assign n77937 = ~n77935 & n77936 ;
  assign n77925 = n77510 & ~n77912 ;
  assign n77926 = n77489 & n77517 ;
  assign n77927 = ~n77925 & ~n77926 ;
  assign n77928 = ~n77504 & ~n77927 ;
  assign n77931 = n77495 & n77929 ;
  assign n77932 = ~n77511 & ~n77931 ;
  assign n77933 = n77476 & ~n77932 ;
  assign n77938 = ~n77928 & ~n77933 ;
  assign n77939 = n77937 & n77938 ;
  assign n77940 = ~n77924 & ~n77939 ;
  assign n77904 = n77504 & ~n77523 ;
  assign n77905 = n77463 & ~n77485 ;
  assign n77906 = ~n77483 & ~n77489 ;
  assign n77907 = ~n77905 & n77906 ;
  assign n77908 = n77483 & n77507 ;
  assign n77909 = ~n77504 & ~n77908 ;
  assign n77910 = ~n77907 & n77909 ;
  assign n77911 = ~n77904 & ~n77910 ;
  assign n77941 = n77470 & ~n77476 ;
  assign n77942 = n77929 & n77941 ;
  assign n77943 = ~n77911 & ~n77942 ;
  assign n77944 = ~n77940 & n77943 ;
  assign n77945 = \u2_L14_reg[31]/P0001  & n77944 ;
  assign n77946 = ~\u2_L14_reg[31]/P0001  & ~n77944 ;
  assign n77947 = ~n77945 & ~n77946 ;
  assign n77955 = n77470 & n77476 ;
  assign n77956 = ~n77912 & ~n77955 ;
  assign n77964 = ~n77469 & ~n77956 ;
  assign n77965 = n77493 & ~n77964 ;
  assign n77966 = n77482 & ~n77965 ;
  assign n77952 = n77476 & n77495 ;
  assign n77953 = ~n77489 & ~n77952 ;
  assign n77967 = n77915 & ~n77953 ;
  assign n77968 = ~n77529 & ~n77967 ;
  assign n77969 = ~n77966 & n77968 ;
  assign n77970 = n77457 & ~n77969 ;
  assign n77948 = ~n77482 & n77492 ;
  assign n77949 = ~n77469 & n77530 ;
  assign n77950 = ~n77948 & ~n77949 ;
  assign n77951 = ~n77504 & ~n77950 ;
  assign n77957 = ~n77484 & n77956 ;
  assign n77958 = n77504 & ~n77957 ;
  assign n77959 = n77482 & n77509 ;
  assign n77954 = ~n77504 & ~n77953 ;
  assign n77960 = ~n77948 & ~n77954 ;
  assign n77961 = ~n77959 & n77960 ;
  assign n77962 = ~n77958 & n77961 ;
  assign n77963 = ~n77457 & ~n77962 ;
  assign n77971 = ~n77951 & ~n77963 ;
  assign n77972 = ~n77970 & n77971 ;
  assign n77973 = \u2_L14_reg[9]/P0001  & n77972 ;
  assign n77974 = ~\u2_L14_reg[9]/P0001  & ~n77972 ;
  assign n77975 = ~n77973 & ~n77974 ;
  assign n77976 = ~n77482 & n77955 ;
  assign n77977 = n77904 & ~n77976 ;
  assign n77981 = n77457 & n77964 ;
  assign n77978 = ~n77457 & ~n77492 ;
  assign n77979 = n77482 & ~n77493 ;
  assign n77980 = ~n77978 & n77979 ;
  assign n77982 = n77463 & n77518 ;
  assign n77983 = ~n77504 & ~n77529 ;
  assign n77984 = ~n77982 & n77983 ;
  assign n77985 = ~n77980 & n77984 ;
  assign n77986 = ~n77981 & n77985 ;
  assign n77987 = ~n77977 & ~n77986 ;
  assign n77989 = ~n77504 & n77517 ;
  assign n77990 = ~n77483 & ~n77989 ;
  assign n77991 = n77463 & ~n77990 ;
  assign n77992 = n77504 & n77955 ;
  assign n77993 = ~n77457 & ~n77920 ;
  assign n77988 = ~n77482 & n77489 ;
  assign n77994 = ~n77931 & ~n77988 ;
  assign n77995 = n77993 & n77994 ;
  assign n77996 = ~n77992 & n77995 ;
  assign n77997 = ~n77991 & n77996 ;
  assign n77999 = n77457 & ~n77524 ;
  assign n77998 = n77504 & n77952 ;
  assign n78000 = ~n77930 & ~n77942 ;
  assign n78001 = ~n77998 & n78000 ;
  assign n78002 = n77999 & n78001 ;
  assign n78003 = ~n77997 & ~n78002 ;
  assign n78004 = ~n77987 & ~n78003 ;
  assign n78005 = ~\u2_L14_reg[23]/P0001  & n78004 ;
  assign n78006 = \u2_L14_reg[23]/P0001  & ~n78004 ;
  assign n78007 = ~n78005 & ~n78006 ;
  assign n78009 = ~n77092 & ~n77117 ;
  assign n78010 = n77087 & ~n78009 ;
  assign n78008 = n77104 & n77112 ;
  assign n78011 = ~n77051 & ~n78008 ;
  assign n78012 = ~n78010 & n78011 ;
  assign n78015 = n77097 & n77671 ;
  assign n78014 = n77070 & n77112 ;
  assign n78016 = n77051 & ~n78014 ;
  assign n78017 = ~n78015 & n78016 ;
  assign n78013 = n77087 & n77606 ;
  assign n78018 = ~n77107 & ~n77609 ;
  assign n78019 = ~n78013 & n78018 ;
  assign n78020 = n78017 & n78019 ;
  assign n78021 = ~n78012 & ~n78020 ;
  assign n78022 = n77080 & n77091 ;
  assign n78023 = ~n77051 & n77123 ;
  assign n78024 = ~n78022 & ~n78023 ;
  assign n78025 = n77688 & n78024 ;
  assign n78026 = n77681 & n78025 ;
  assign n78027 = n77087 & ~n77121 ;
  assign n78028 = ~n77605 & n78027 ;
  assign n78029 = ~n78026 & ~n78028 ;
  assign n78030 = ~n78021 & ~n78029 ;
  assign n78031 = \u2_L14_reg[15]/P0001  & n78030 ;
  assign n78032 = ~\u2_L14_reg[15]/P0001  & ~n78030 ;
  assign n78033 = ~n78031 & ~n78032 ;
  assign n78036 = ~n77389 & ~n77437 ;
  assign n78037 = ~n77382 & n78036 ;
  assign n78038 = n77428 & n77437 ;
  assign n78034 = n77403 & ~n77418 ;
  assign n78035 = ~n77403 & n77418 ;
  assign n78039 = ~n78034 & ~n78035 ;
  assign n78040 = ~n77809 & n78039 ;
  assign n78041 = ~n78038 & n78040 ;
  assign n78042 = ~n78037 & n78041 ;
  assign n78044 = n77437 & ~n77441 ;
  assign n78043 = ~n77374 & ~n77429 ;
  assign n78045 = n78034 & ~n78043 ;
  assign n78046 = ~n78044 & n78045 ;
  assign n78047 = ~n78042 & ~n78046 ;
  assign n78048 = n77395 & n77799 ;
  assign n78049 = ~n78047 & ~n78048 ;
  assign n78050 = n77395 & n77813 ;
  assign n78051 = ~n78036 & ~n78050 ;
  assign n78052 = ~n78038 & n78051 ;
  assign n78053 = ~n77809 & n78035 ;
  assign n78054 = ~n78052 & n78053 ;
  assign n78055 = ~n78049 & ~n78054 ;
  assign n78056 = \u2_L14_reg[7]/P0001  & ~n78055 ;
  assign n78057 = ~\u2_L14_reg[7]/P0001  & n78055 ;
  assign n78058 = ~n78056 & ~n78057 ;
  assign n78060 = ~n77380 & n77807 ;
  assign n78061 = ~n77381 & n77434 ;
  assign n78062 = ~n77441 & n78061 ;
  assign n78063 = ~n78060 & ~n78062 ;
  assign n78064 = ~n77418 & ~n78063 ;
  assign n78059 = n77381 & n77396 ;
  assign n78065 = ~n77404 & ~n77432 ;
  assign n78066 = ~n77808 & n78065 ;
  assign n78067 = n77418 & ~n77420 ;
  assign n78068 = ~n78066 & n78067 ;
  assign n78069 = ~n78059 & ~n78068 ;
  assign n78070 = ~n78064 & n78069 ;
  assign n78071 = n77403 & ~n78070 ;
  assign n78072 = n77380 & n77439 ;
  assign n78076 = n77786 & ~n77817 ;
  assign n78077 = ~n78072 & n78076 ;
  assign n78073 = ~n77439 & ~n78050 ;
  assign n78074 = n77418 & ~n78073 ;
  assign n78075 = ~n77434 & n77440 ;
  assign n78078 = ~n78074 & ~n78075 ;
  assign n78079 = n78077 & n78078 ;
  assign n78080 = ~n77403 & ~n78079 ;
  assign n78081 = n77418 & n77421 ;
  assign n78082 = ~n77374 & n77428 ;
  assign n78083 = ~n77798 & ~n78082 ;
  assign n78084 = ~n77418 & ~n78083 ;
  assign n78085 = ~n78081 & ~n78084 ;
  assign n78086 = ~n78080 & n78085 ;
  assign n78087 = ~n78071 & n78086 ;
  assign n78088 = \u2_L14_reg[32]/P0001  & n78087 ;
  assign n78089 = ~\u2_L14_reg[32]/P0001  & ~n78087 ;
  assign n78090 = ~n78088 & ~n78089 ;
  assign n78096 = ~n77730 & ~n77755 ;
  assign n78097 = ~n77883 & ~n78096 ;
  assign n78098 = ~n77710 & ~n77763 ;
  assign n78099 = ~n78097 & n78098 ;
  assign n78100 = n77710 & ~n77747 ;
  assign n78101 = ~n77740 & n77746 ;
  assign n78102 = n77734 & ~n78101 ;
  assign n78103 = n78100 & n78102 ;
  assign n78104 = ~n78099 & ~n78103 ;
  assign n78105 = ~n77704 & ~n78104 ;
  assign n78106 = ~n77710 & ~n77888 ;
  assign n78108 = n77710 & ~n77762 ;
  assign n78107 = n77717 & n77752 ;
  assign n78109 = ~n77869 & ~n78107 ;
  assign n78110 = n78108 & n78109 ;
  assign n78111 = ~n78106 & ~n78110 ;
  assign n78112 = n77704 & ~n77885 ;
  assign n78113 = ~n78111 & n78112 ;
  assign n78114 = ~n78105 & ~n78113 ;
  assign n78091 = n77740 & n77751 ;
  assign n78092 = n77756 & n78091 ;
  assign n78093 = n77710 & ~n77730 ;
  assign n78094 = ~n77751 & n78093 ;
  assign n78095 = n77765 & n78094 ;
  assign n78115 = ~n78092 & ~n78095 ;
  assign n78116 = ~n78114 & n78115 ;
  assign n78117 = \u2_L14_reg[24]/P0001  & n78116 ;
  assign n78118 = ~\u2_L14_reg[24]/P0001  & ~n78116 ;
  assign n78119 = ~n78117 & ~n78118 ;
  assign n78123 = ~n77740 & ~n77751 ;
  assign n78124 = ~n78091 & ~n78123 ;
  assign n78125 = ~n77732 & ~n78124 ;
  assign n78126 = n77710 & n77747 ;
  assign n78127 = ~n78125 & ~n78126 ;
  assign n78128 = ~n77730 & ~n78127 ;
  assign n78120 = ~n77730 & n77742 ;
  assign n78121 = ~n77733 & ~n78120 ;
  assign n78122 = ~n77710 & ~n78121 ;
  assign n78129 = ~n77886 & ~n78122 ;
  assign n78130 = ~n78128 & n78129 ;
  assign n78131 = n77704 & ~n78130 ;
  assign n78132 = n78100 & n78124 ;
  assign n78133 = n77710 & ~n77876 ;
  assign n78134 = n77723 & n77764 ;
  assign n78135 = ~n77875 & ~n78091 ;
  assign n78136 = ~n78134 & n78135 ;
  assign n78137 = ~n78133 & ~n78136 ;
  assign n78138 = ~n78132 & ~n78137 ;
  assign n78139 = ~n77704 & ~n78138 ;
  assign n78140 = n77733 & ~n77740 ;
  assign n78141 = ~n77891 & ~n78140 ;
  assign n78142 = n77710 & ~n78141 ;
  assign n78143 = ~n77710 & n78101 ;
  assign n78144 = ~n78142 & ~n78143 ;
  assign n78145 = ~n78139 & n78144 ;
  assign n78146 = ~n78131 & n78145 ;
  assign n78147 = \u2_L14_reg[16]/P0001  & n78146 ;
  assign n78148 = ~\u2_L14_reg[16]/P0001  & ~n78146 ;
  assign n78149 = ~n78147 & ~n78148 ;
  assign n78157 = n76756 & ~n76765 ;
  assign n78158 = ~n76781 & ~n78157 ;
  assign n78159 = n76772 & ~n78158 ;
  assign n78160 = n76748 & ~n76765 ;
  assign n78161 = ~n76772 & n78160 ;
  assign n78162 = ~n77861 & ~n78161 ;
  assign n78163 = ~n78159 & n78162 ;
  assign n78164 = n76779 & ~n78163 ;
  assign n78150 = n76810 & ~n77269 ;
  assign n78151 = n76782 & ~n78150 ;
  assign n78152 = n76787 & ~n77278 ;
  assign n78153 = ~n78151 & ~n78152 ;
  assign n78154 = ~n76766 & ~n76784 ;
  assign n78155 = ~n78153 & n78154 ;
  assign n78156 = ~n76779 & ~n78155 ;
  assign n78165 = ~n76772 & n77270 ;
  assign n78166 = n76755 & n76784 ;
  assign n78167 = n77860 & ~n78166 ;
  assign n78168 = n76772 & ~n78167 ;
  assign n78169 = ~n78165 & ~n78168 ;
  assign n78170 = ~n78156 & n78169 ;
  assign n78171 = ~n78164 & n78170 ;
  assign n78172 = \u2_L14_reg[8]/P0001  & n78171 ;
  assign n78173 = ~\u2_L14_reg[8]/P0001  & ~n78171 ;
  assign n78174 = ~n78172 & ~n78173 ;
  assign n78179 = ~n76918 & ~n76945 ;
  assign n78180 = ~n77349 & ~n78179 ;
  assign n78181 = n76932 & ~n78180 ;
  assign n78182 = ~n76912 & ~n78181 ;
  assign n78183 = ~n76932 & n78179 ;
  assign n78184 = n76912 & ~n77334 ;
  assign n78185 = ~n78183 & n78184 ;
  assign n78186 = ~n78182 & ~n78185 ;
  assign n78187 = ~n76939 & ~n77333 ;
  assign n78188 = n77343 & n78187 ;
  assign n78189 = ~n78186 & n78188 ;
  assign n78190 = ~n76956 & n77350 ;
  assign n78191 = n76960 & ~n76961 ;
  assign n78192 = ~n76912 & ~n76964 ;
  assign n78193 = ~n78191 & n78192 ;
  assign n78194 = ~n78190 & ~n78193 ;
  assign n78175 = n76925 & n77353 ;
  assign n78195 = n76939 & ~n76950 ;
  assign n78196 = ~n78175 & n78195 ;
  assign n78197 = ~n78194 & n78196 ;
  assign n78198 = ~n78189 & ~n78197 ;
  assign n78177 = n76952 & ~n76979 ;
  assign n78178 = n76912 & ~n78177 ;
  assign n78176 = ~n76912 & n78175 ;
  assign n78199 = ~n77342 & ~n78176 ;
  assign n78200 = ~n78178 & n78199 ;
  assign n78201 = ~n78198 & n78200 ;
  assign n78202 = \u2_L14_reg[1]/P0001  & n78201 ;
  assign n78203 = ~\u2_L14_reg[1]/P0001  & ~n78201 ;
  assign n78204 = ~n78202 & ~n78203 ;
  assign n78206 = ~n76918 & n77349 ;
  assign n78207 = ~n76946 & ~n78206 ;
  assign n78208 = ~n76912 & ~n78207 ;
  assign n78209 = ~n76964 & ~n76981 ;
  assign n78210 = ~n78208 & n78209 ;
  assign n78211 = n76918 & ~n78210 ;
  assign n78212 = ~n76932 & n78208 ;
  assign n78213 = n76912 & n76980 ;
  assign n78205 = ~n76918 & n76954 ;
  assign n78214 = ~n78175 & ~n78205 ;
  assign n78215 = ~n78213 & n78214 ;
  assign n78216 = ~n78212 & n78215 ;
  assign n78217 = ~n78211 & n78216 ;
  assign n78218 = n76939 & ~n78217 ;
  assign n78219 = n76926 & ~n76963 ;
  assign n78220 = ~n76956 & ~n76991 ;
  assign n78221 = ~n76965 & n78220 ;
  assign n78222 = ~n78219 & n78221 ;
  assign n78223 = ~n76939 & ~n78222 ;
  assign n78224 = ~n76945 & ~n77338 ;
  assign n78225 = ~n76947 & ~n78224 ;
  assign n78226 = ~n76918 & ~n78225 ;
  assign n78227 = ~n76950 & ~n76971 ;
  assign n78228 = ~n76939 & ~n78227 ;
  assign n78229 = ~n76912 & ~n78228 ;
  assign n78230 = ~n78226 & n78229 ;
  assign n78231 = n76912 & ~n76957 ;
  assign n78232 = ~n76965 & n78231 ;
  assign n78233 = ~n78230 & ~n78232 ;
  assign n78234 = ~n78223 & ~n78233 ;
  assign n78235 = ~n78218 & n78234 ;
  assign n78236 = \u2_L14_reg[26]/P0001  & n78235 ;
  assign n78237 = ~\u2_L14_reg[26]/P0001  & ~n78235 ;
  assign n78238 = ~n78236 & ~n78237 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g16/_0_  = ~n5910 ;
  assign \g191647/_3_  = ~n6000 ;
  assign \g191648/_3_  = ~n6094 ;
  assign \g191819/_3_  = ~n6192 ;
  assign \g191821/_0_  = ~n6283 ;
  assign \g191940/_3_  = ~n6374 ;
  assign \g191941/_0_  = n6400 ;
  assign \g191942/_0_  = ~n6500 ;
  assign \g191944/_0_  = ~n6529 ;
  assign \g191945/_0_  = ~n6560 ;
  assign \g191946/_0_  = ~n6601 ;
  assign \g191947/_3_  = ~n6635 ;
  assign \g191948/_0_  = ~n6672 ;
  assign \g191949/_0_  = ~n6711 ;
  assign \g191950/_0_  = ~n6790 ;
  assign \g191951/_3_  = ~n6835 ;
  assign \g191952/_0_  = ~n6867 ;
  assign \g192015/_3_  = ~n6896 ;
  assign \g192016/_3_  = ~n6920 ;
  assign \g192017/_3_  = ~n6952 ;
  assign \g192018/_3_  = ~n6981 ;
  assign \g192019/_3_  = ~n7015 ;
  assign \g192020/_0_  = ~n7106 ;
  assign \g192021/_3_  = ~n7130 ;
  assign \g192022/_0_  = ~n7158 ;
  assign \g192047/_0_  = ~n7193 ;
  assign \g192048/_0_  = ~n7227 ;
  assign \g192049/_0_  = ~n7254 ;
  assign \g192050/_0_  = ~n7283 ;
  assign \g192051/_0_  = ~n7308 ;
  assign \g192081/_0_  = ~n7335 ;
  assign \g193428/_3_  = ~n7431 ;
  assign \g193720/_0_  = ~n7529 ;
  assign \g193721/_0_  = ~n7621 ;
  assign \g193877/_0_  = ~n7716 ;
  assign \g193878/_0_  = ~n7746 ;
  assign \g193879/_0_  = ~n7785 ;
  assign \g193880/_3_  = ~n7878 ;
  assign \g193881/_0_  = ~n7976 ;
  assign \g193882/_0_  = ~n8008 ;
  assign \g193998/_0_  = ~n8042 ;
  assign \g193999/_0_  = n8074 ;
  assign \g194000/_3_  = ~n8112 ;
  assign \g194001/_0_  = ~n8146 ;
  assign \g194002/_0_  = ~n8247 ;
  assign \g194003/_0_  = ~n8271 ;
  assign \g194004/_0_  = ~n8306 ;
  assign \g194005/_0_  = ~n8342 ;
  assign \g194006/_0_  = ~n8377 ;
  assign \g194007/_0_  = ~n8418 ;
  assign \g194008/_0_  = ~n8449 ;
  assign \g194009/_0_  = ~n8477 ;
  assign \g194010/_0_  = ~n8504 ;
  assign \g194055/_3_  = ~n8534 ;
  assign \g194056/_3_  = ~n8563 ;
  assign \g194057/_0_  = ~n8589 ;
  assign \g194058/_0_  = ~n8676 ;
  assign \g194059/_0_  = ~n8701 ;
  assign \g194060/_0_  = ~n8724 ;
  assign \g194090/_0_  = ~n8760 ;
  assign \g194091/_0_  = ~n8786 ;
  assign \g194092/_0_  = ~n8819 ;
  assign \g194093/_0_  = ~n8848 ;
  assign \g195671/_0_  = ~n8938 ;
  assign \g195672/_3_  = ~n9035 ;
  assign \g195868/_0_  = ~n9132 ;
  assign \g195869/_0_  = ~n9230 ;
  assign \g195870/_0_  = ~n9323 ;
  assign \g196010/_0_  = ~n9355 ;
  assign \g196011/_0_  = n9388 ;
  assign \g196012/_0_  = ~n9488 ;
  assign \g196013/_0_  = ~n9522 ;
  assign \g196014/_0_  = ~n9553 ;
  assign \g196015/_0_  = ~n9585 ;
  assign \g196016/_0_  = ~n9623 ;
  assign \g196017/_0_  = ~n9702 ;
  assign \g196018/_0_  = ~n9738 ;
  assign \g196019/_3_  = ~n9783 ;
  assign \g196020/_0_  = ~n9816 ;
  assign \g196021/_0_  = ~n9857 ;
  assign \g196022/_0_  = ~n9890 ;
  assign \g196096/_3_  = ~n9919 ;
  assign \g196097/_0_  = ~n9944 ;
  assign \g196098/_0_  = ~n9977 ;
  assign \g196099/_0_  = ~n10006 ;
  assign \g196100/_3_  = ~n10041 ;
  assign \g196101/_0_  = ~n10128 ;
  assign \g196102/_0_  = ~n10150 ;
  assign \g196103/_0_  = ~n10177 ;
  assign \g196136/_0_  = ~n10213 ;
  assign \g196137/_0_  = ~n10246 ;
  assign \g196138/_0_  = ~n10275 ;
  assign \g196139/_0_  = ~n10304 ;
  assign \g196140/_0_  = ~n10330 ;
  assign \g196170/_0_  = ~n10357 ;
  assign \g197520/_3_  = ~n10453 ;
  assign \g197821/_0_  = ~n10549 ;
  assign \g197923/_0_  = ~n10646 ;
  assign \g197996/_0_  = ~n10744 ;
  assign \g197997/_3_  = ~n10835 ;
  assign \g197998/_0_  = ~n10872 ;
  assign \g197999/_0_  = ~n10969 ;
  assign \g198000/_0_  = ~n11001 ;
  assign \g198071/_0_  = ~n11031 ;
  assign \g198123/_0_  = ~n11054 ;
  assign \g198124/_0_  = ~n11090 ;
  assign \g198125/_0_  = ~n11130 ;
  assign \g198126/_0_  = ~n11165 ;
  assign \g198127/_0_  = ~n11257 ;
  assign \g198128/_0_  = ~n11290 ;
  assign \g198129/_0_  = ~n11328 ;
  assign \g198130/_0_  = ~n11365 ;
  assign \g198131/_0_  = ~n11392 ;
  assign \g198132/_0_  = n11422 ;
  assign \g198133/_0_  = ~n11460 ;
  assign \g198134/_3_  = ~n11494 ;
  assign \g198135/_0_  = ~n11527 ;
  assign \g198182/_0_  = ~n11554 ;
  assign \g198183/_3_  = ~n11588 ;
  assign \g198184/_0_  = ~n11615 ;
  assign \g198185/_0_  = ~n11698 ;
  assign \g198186/_0_  = ~n11727 ;
  assign \g198187/_0_  = ~n11750 ;
  assign \g198219/_0_  = ~n11776 ;
  assign \g198220/_0_  = ~n11815 ;
  assign \g198221/_0_  = ~n11846 ;
  assign \g198222/_0_  = ~n11876 ;
  assign \g199794/_0_  = ~n11967 ;
  assign \g199795/_3_  = ~n12064 ;
  assign \g200006/_0_  = ~n12159 ;
  assign \g200007/_0_  = ~n12252 ;
  assign \g200008/_0_  = ~n12349 ;
  assign \g200139/_0_  = ~n12382 ;
  assign \g200140/_0_  = n12414 ;
  assign \g200141/_0_  = ~n12511 ;
  assign \g200142/_0_  = ~n12543 ;
  assign \g200143/_0_  = ~n12574 ;
  assign \g200144/_0_  = ~n12609 ;
  assign \g200145/_0_  = ~n12647 ;
  assign \g200146/_0_  = ~n12685 ;
  assign \g200147/_0_  = ~n12764 ;
  assign \g200148/_0_  = ~n12798 ;
  assign \g200149/_0_  = ~n12831 ;
  assign \g200150/_3_  = ~n12876 ;
  assign \g200151/_0_  = ~n12911 ;
  assign \g200228/_3_  = ~n12940 ;
  assign \g200229/_0_  = ~n12965 ;
  assign \g200230/_0_  = ~n12998 ;
  assign \g200231/_0_  = ~n13027 ;
  assign \g200232/_3_  = ~n13059 ;
  assign \g200233/_0_  = ~n13146 ;
  assign \g200234/_0_  = ~n13176 ;
  assign \g200235/_0_  = ~n13203 ;
  assign \g200268/_0_  = ~n13239 ;
  assign \g200269/_0_  = ~n13272 ;
  assign \g200270/_0_  = ~n13301 ;
  assign \g200271/_0_  = ~n13330 ;
  assign \g200272/_0_  = ~n13356 ;
  assign \g200299/_0_  = ~n13383 ;
  assign \g201655/_3_  = ~n13474 ;
  assign \g201960/_0_  = ~n13569 ;
  assign \g201961/_0_  = ~n13659 ;
  assign \g202131/_0_  = ~n13692 ;
  assign \g202132/_0_  = ~n13789 ;
  assign \g202133/_3_  = ~n13881 ;
  assign \g202134/_0_  = ~n13915 ;
  assign \g202135/_0_  = ~n13950 ;
  assign \g202136/_0_  = ~n14041 ;
  assign \g202257/_0_  = ~n14072 ;
  assign \g202258/_0_  = n14106 ;
  assign \g202259/_3_  = ~n14144 ;
  assign \g202260/_0_  = ~n14246 ;
  assign \g202261/_0_  = ~n14282 ;
  assign \g202262/_0_  = ~n14314 ;
  assign \g202263/_0_  = ~n14339 ;
  assign \g202264/_0_  = ~n14375 ;
  assign \g202265/_0_  = ~n14409 ;
  assign \g202266/_0_  = ~n14447 ;
  assign \g202267/_0_  = ~n14479 ;
  assign \g202268/_0_  = ~n14505 ;
  assign \g202269/_0_  = ~n14530 ;
  assign \g202317/_0_  = ~n14558 ;
  assign \g202318/_3_  = ~n14592 ;
  assign \g202319/_0_  = ~n14617 ;
  assign \g202320/_0_  = ~n14701 ;
  assign \g202321/_0_  = ~n14724 ;
  assign \g202322/_0_  = ~n14746 ;
  assign \g202354/_0_  = ~n14780 ;
  assign \g202355/_0_  = ~n14807 ;
  assign \g202356/_0_  = ~n14841 ;
  assign \g202357/_0_  = ~n14870 ;
  assign \g203927/_0_  = ~n14957 ;
  assign \g203928/_3_  = ~n15050 ;
  assign \g204142/_0_  = ~n15147 ;
  assign \g204143/_0_  = ~n15240 ;
  assign \g204144/_0_  = ~n15333 ;
  assign \g204275/_0_  = ~n15368 ;
  assign \g204276/_0_  = n15399 ;
  assign \g204277/_0_  = ~n15432 ;
  assign \g204278/_0_  = ~n15464 ;
  assign \g204279/_0_  = ~n15563 ;
  assign \g204280/_0_  = ~n15591 ;
  assign \g204281/_0_  = ~n15630 ;
  assign \g204282/_0_  = ~n15669 ;
  assign \g204283/_0_  = ~n15700 ;
  assign \g204284/_0_  = ~n15786 ;
  assign \g204285/_0_  = ~n15821 ;
  assign \g204286/_3_  = ~n15863 ;
  assign \g204287/_0_  = ~n15896 ;
  assign \g204363/_3_  = ~n15928 ;
  assign \g204364/_0_  = ~n15952 ;
  assign \g204365/_0_  = ~n15983 ;
  assign \g204366/_0_  = ~n16013 ;
  assign \g204367/_3_  = ~n16051 ;
  assign \g204368/_0_  = ~n16142 ;
  assign \g204369/_0_  = ~n16171 ;
  assign \g204370/_0_  = ~n16197 ;
  assign \g204403/_0_  = ~n16232 ;
  assign \g204404/_0_  = ~n16266 ;
  assign \g204405/_0_  = ~n16293 ;
  assign \g204406/_0_  = ~n16323 ;
  assign \g204407/_0_  = ~n16347 ;
  assign \g204434/_0_  = ~n16372 ;
  assign \g205833/_3_  = ~n16467 ;
  assign \g206103/_0_  = ~n16565 ;
  assign \g206104/_0_  = ~n16650 ;
  assign \g206266/_0_  = ~n16683 ;
  assign \g206267/_0_  = ~n16782 ;
  assign \g206268/_0_  = ~n16821 ;
  assign \g206269/_3_  = ~n16911 ;
  assign \g206270/_0_  = ~n16943 ;
  assign \g206271/_0_  = ~n17028 ;
  assign \g206387/_0_  = ~n17060 ;
  assign \g206388/_0_  = n17092 ;
  assign \g206389/_3_  = ~n17129 ;
  assign \g206390/_0_  = ~n17231 ;
  assign \g206391/_0_  = ~n17268 ;
  assign \g206392/_0_  = ~n17292 ;
  assign \g206393/_0_  = ~n17323 ;
  assign \g206394/_0_  = ~n17359 ;
  assign \g206395/_0_  = ~n17393 ;
  assign \g206396/_0_  = ~n17431 ;
  assign \g206397/_0_  = ~n17464 ;
  assign \g206398/_0_  = ~n17495 ;
  assign \g206399/_0_  = ~n17520 ;
  assign \g206446/_0_  = ~n17550 ;
  assign \g206447/_3_  = ~n17581 ;
  assign \g206448/_0_  = ~n17606 ;
  assign \g206449/_0_  = ~n17690 ;
  assign \g206450/_0_  = ~n17711 ;
  assign \g206451/_0_  = ~n17736 ;
  assign \g206483/_0_  = ~n17770 ;
  assign \g206484/_0_  = ~n17795 ;
  assign \g206485/_0_  = ~n17829 ;
  assign \g206486/_0_  = ~n17858 ;
  assign \g208069/_0_  = ~n17952 ;
  assign \g208070/_3_  = ~n18047 ;
  assign \g208253/_0_  = ~n18142 ;
  assign \g208254/_0_  = ~n18236 ;
  assign \g208255/_0_  = ~n18323 ;
  assign \g208406/_0_  = ~n18355 ;
  assign \g208407/_0_  = n18387 ;
  assign \g208408/_0_  = ~n18486 ;
  assign \g208409/_0_  = ~n18522 ;
  assign \g208410/_0_  = ~n18556 ;
  assign \g208411/_0_  = ~n18589 ;
  assign \g208412/_0_  = ~n18629 ;
  assign \g208413/_0_  = ~n18668 ;
  assign \g208414/_0_  = ~n18699 ;
  assign \g208415/_3_  = ~n18790 ;
  assign \g208416/_0_  = ~n18824 ;
  assign \g208417/_0_  = ~n18859 ;
  assign \g208418/_0_  = ~n18894 ;
  assign \g208493/_3_  = ~n18926 ;
  assign \g208494/_0_  = ~n18951 ;
  assign \g208495/_0_  = ~n18983 ;
  assign \g208496/_0_  = ~n19010 ;
  assign \g208497/_3_  = ~n19043 ;
  assign \g208498/_0_  = ~n19130 ;
  assign \g208499/_0_  = ~n19155 ;
  assign \g208500/_0_  = ~n19181 ;
  assign \g208533/_0_  = ~n19217 ;
  assign \g208534/_0_  = ~n19250 ;
  assign \g208535/_0_  = ~n19279 ;
  assign \g208536/_0_  = ~n19309 ;
  assign \g208537/_0_  = ~n19334 ;
  assign \g208564/_0_  = ~n19358 ;
  assign \g209938/_3_  = ~n19454 ;
  assign \g210205/_0_  = ~n19549 ;
  assign \g210206/_0_  = ~n19635 ;
  assign \g210380/_0_  = ~n19668 ;
  assign \g210381/_0_  = ~n19765 ;
  assign \g210382/_0_  = ~n19799 ;
  assign \g210383/_3_  = ~n19889 ;
  assign \g210384/_0_  = ~n19924 ;
  assign \g210385/_0_  = ~n20012 ;
  assign \g210499/_0_  = ~n20044 ;
  assign \g210500/_0_  = n20075 ;
  assign \g210501/_3_  = ~n20112 ;
  assign \g210502/_0_  = ~n20147 ;
  assign \g210503/_0_  = ~n20250 ;
  assign \g210504/_0_  = ~n20275 ;
  assign \g210505/_0_  = ~n20307 ;
  assign \g210506/_0_  = ~n20344 ;
  assign \g210507/_0_  = ~n20378 ;
  assign \g210508/_0_  = ~n20410 ;
  assign \g210509/_0_  = ~n20445 ;
  assign \g210510/_0_  = ~n20476 ;
  assign \g210511/_0_  = ~n20501 ;
  assign \g210558/_0_  = ~n20530 ;
  assign \g210559/_3_  = ~n20566 ;
  assign \g210560/_0_  = ~n20592 ;
  assign \g210561/_0_  = ~n20678 ;
  assign \g210562/_0_  = ~n20702 ;
  assign \g210563/_0_  = ~n20727 ;
  assign \g210595/_0_  = ~n20762 ;
  assign \g210596/_0_  = ~n20787 ;
  assign \g210597/_0_  = ~n20822 ;
  assign \g210598/_0_  = ~n20852 ;
  assign \g212159/_0_  = ~n20944 ;
  assign \g212160/_3_  = ~n21042 ;
  assign \g212384/_0_  = ~n21137 ;
  assign \g212385/_0_  = ~n21234 ;
  assign \g212386/_0_  = ~n21328 ;
  assign \g212536/_0_  = ~n21359 ;
  assign \g212537/_0_  = n21390 ;
  assign \g212538/_0_  = ~n21489 ;
  assign \g212539/_0_  = ~n21520 ;
  assign \g212540/_0_  = ~n21554 ;
  assign \g212541/_0_  = ~n21586 ;
  assign \g212542/_0_  = ~n21625 ;
  assign \g212543/_0_  = ~n21658 ;
  assign \g212544/_0_  = ~n21692 ;
  assign \g212545/_0_  = ~n21731 ;
  assign \g212546/_3_  = ~n21821 ;
  assign \g212547/_0_  = ~n21856 ;
  assign \g212623/_3_  = ~n21893 ;
  assign \g212624/_0_  = ~n21918 ;
  assign \g212625/_0_  = ~n21952 ;
  assign \g212626/_0_  = ~n21982 ;
  assign \g212627/_0_  = ~n22013 ;
  assign \g212628/_3_  = ~n22048 ;
  assign \g212629/_0_  = ~n22135 ;
  assign \g212630/_0_  = ~n22159 ;
  assign \g212631/_0_  = ~n22185 ;
  assign \g212667/_0_  = ~n22221 ;
  assign \g212668/_0_  = ~n22254 ;
  assign \g212669/_0_  = ~n22283 ;
  assign \g212670/_0_  = ~n22313 ;
  assign \g212671/_0_  = ~n22338 ;
  assign \g212699/_0_  = ~n22363 ;
  assign \g214033/_3_  = ~n22456 ;
  assign \g214309/_3_  = ~n22551 ;
  assign \g214310/_0_  = ~n22640 ;
  assign \g214494/_0_  = ~n22673 ;
  assign \g214495/_0_  = ~n22769 ;
  assign \g214496/_0_  = ~n22803 ;
  assign \g214497/_3_  = ~n22893 ;
  assign \g214632/_0_  = ~n22923 ;
  assign \g214633/_0_  = n22958 ;
  assign \g214634/_3_  = ~n22995 ;
  assign \g214635/_0_  = ~n23096 ;
  assign \g214636/_0_  = ~n23174 ;
  assign \g214637/_0_  = ~n23208 ;
  assign \g214638/_0_  = ~n23254 ;
  assign \g214639/_0_  = ~n23287 ;
  assign \g214640/_0_  = ~n23321 ;
  assign \g214641/_0_  = ~n23352 ;
  assign \g214642/_0_  = ~n23383 ;
  assign \g214643/_0_  = ~n23418 ;
  assign \g214691/_0_  = ~n23443 ;
  assign \g214692/_0_  = ~n23481 ;
  assign \g214693/_3_  = ~n23512 ;
  assign \g214694/_0_  = ~n23596 ;
  assign \g214695/_0_  = ~n23624 ;
  assign \g214696/_0_  = ~n23654 ;
  assign \g214697/_0_  = ~n23678 ;
  assign \g214729/_0_  = ~n23712 ;
  assign \g214730/_0_  = ~n23737 ;
  assign \g214731/_0_  = ~n23771 ;
  assign \g214732/_0_  = ~n23800 ;
  assign \g214733/_0_  = ~n23827 ;
  assign \g216157/_0_  = ~n23914 ;
  assign \g216158/_3_  = ~n24012 ;
  assign \g216492/_0_  = ~n24107 ;
  assign \g216493/_0_  = ~n24195 ;
  assign \g216671/_0_  = n24226 ;
  assign \g216672/_0_  = ~n24257 ;
  assign \g216673/_0_  = ~n24353 ;
  assign \g216674/_0_  = ~n24436 ;
  assign \g216675/_0_  = ~n24472 ;
  assign \g216676/_3_  = ~n24517 ;
  assign \g216677/_0_  = ~n24550 ;
  assign \g216735/_0_  = ~n24583 ;
  assign \g216736/_3_  = ~n24619 ;
  assign \g216737/_0_  = ~n24654 ;
  assign \g216738/_0_  = ~n24754 ;
  assign \g216739/_0_  = ~n24779 ;
  assign \g216740/_0_  = ~n24816 ;
  assign \g216741/_0_  = ~n24851 ;
  assign \g216742/_0_  = ~n24885 ;
  assign \g216743/_0_  = ~n24922 ;
  assign \g216744/_0_  = ~n24951 ;
  assign \g216745/_0_  = ~n24980 ;
  assign \g216746/_3_  = ~n25018 ;
  assign \g216747/_0_  = ~n25105 ;
  assign \g216748/_0_  = ~n25134 ;
  assign \g216749/_0_  = ~n25160 ;
  assign \g216788/_0_  = ~n25196 ;
  assign \g216789/_0_  = ~n25229 ;
  assign \g216790/_0_  = ~n25258 ;
  assign \g216791/_0_  = ~n25285 ;
  assign \g216792/_0_  = ~n25310 ;
  assign \g216829/_0_  = ~n25335 ;
  assign \g218407/_3_  = ~n25433 ;
  assign \g218408/_0_  = ~n25520 ;
  assign \g218423/_3_  = ~n25618 ;
  assign \g218601/_0_  = ~n25715 ;
  assign \g218602/_0_  = ~n25754 ;
  assign \g218603/_0_  = ~n25786 ;
  assign \g218604/_0_  = ~n25874 ;
  assign \g218724/_0_  = ~n25904 ;
  assign \g218725/_0_  = n25937 ;
  assign \g218726/_0_  = ~n26039 ;
  assign \g218727/_0_  = ~n26070 ;
  assign \g218728/_0_  = ~n26094 ;
  assign \g218729/_0_  = ~n26129 ;
  assign \g218730/_0_  = ~n26164 ;
  assign \g218731/_0_  = ~n26201 ;
  assign \g218732/_0_  = ~n26236 ;
  assign \g218733/_0_  = ~n26267 ;
  assign \g218734/_0_  = ~n26353 ;
  assign \g218735/_3_  = ~n26395 ;
  assign \g218736/_0_  = ~n26423 ;
  assign \g218808/_3_  = ~n26455 ;
  assign \g218809/_0_  = ~n26489 ;
  assign \g218810/_0_  = ~n26518 ;
  assign \g218811/_3_  = ~n26554 ;
  assign \g218812/_0_  = ~n26580 ;
  assign \g218813/_0_  = ~n26667 ;
  assign \g218814/_0_  = ~n26696 ;
  assign \g218846/_0_  = ~n26733 ;
  assign \g218847/_0_  = ~n26765 ;
  assign \g218848/_0_  = ~n26793 ;
  assign \g218849/_0_  = ~n26818 ;
  assign \g218877/_0_  = ~n26843 ;
  assign \g22/_0_  = ~n26931 ;
  assign \g220545/_0_  = ~n27018 ;
  assign \g220546/_3_  = ~n27114 ;
  assign \g220725/_3_  = ~n27208 ;
  assign \g220726/_0_  = ~n27304 ;
  assign \g220793/_0_  = ~n27337 ;
  assign \g220794/_0_  = n27372 ;
  assign \g220795/_0_  = ~n27475 ;
  assign \g220796/_0_  = ~n27558 ;
  assign \g220797/_0_  = ~n27587 ;
  assign \g220798/_0_  = ~n27619 ;
  assign \g220799/_0_  = ~n27654 ;
  assign \g220800/_0_  = ~n27701 ;
  assign \g220801/_0_  = ~n27730 ;
  assign \g220802/_0_  = ~n27816 ;
  assign \g220803/_0_  = ~n27852 ;
  assign \g220804/_3_  = ~n27894 ;
  assign \g220805/_0_  = ~n27930 ;
  assign \g220806/_0_  = ~n27959 ;
  assign \g220807/_0_  = ~n27994 ;
  assign \g220872/_3_  = ~n28026 ;
  assign \g220873/_0_  = ~n28059 ;
  assign \g220874/_3_  = ~n28093 ;
  assign \g220875/_0_  = ~n28180 ;
  assign \g220876/_0_  = ~n28210 ;
  assign \g220877/_0_  = ~n28237 ;
  assign \g220921/_0_  = ~n28273 ;
  assign \g220922/_0_  = ~n28306 ;
  assign \g220923/_0_  = ~n28332 ;
  assign \g220924/_0_  = ~n28361 ;
  assign \g220925/_0_  = ~n28386 ;
  assign \g220926/_0_  = ~n28410 ;
  assign \g220969/_0_  = ~n28435 ;
  assign \g221011/_3_  = ~n28525 ;
  assign \g221039/_3_  = ~n28621 ;
  assign \g221086/_3_  = ~n28710 ;
  assign \g221131/_0_  = ~n28790 ;
  assign \g224010/_3_  = ~n28882 ;
  assign \g224368/_3_  = ~n28972 ;
  assign \g224369/_3_  = ~n29066 ;
  assign \g224532/_0_  = ~n29108 ;
  assign \g224533/_0_  = ~n29142 ;
  assign \g224534/_0_  = ~n29238 ;
  assign \g224535/_3_  = ~n29326 ;
  assign \g224536/_0_  = ~n29353 ;
  assign \g224537/_0_  = ~n29453 ;
  assign \g224640/_3_  = ~n29492 ;
  assign \g224641/_0_  = ~n29592 ;
  assign \g224642/_0_  = ~n29630 ;
  assign \g224643/_3_  = ~n29660 ;
  assign \g224644/_0_  = n29694 ;
  assign \g224645/_0_  = ~n29723 ;
  assign \g224646/_3_  = ~n29745 ;
  assign \g224647/_0_  = ~n29777 ;
  assign \g224648/_3_  = ~n29812 ;
  assign \g224649/_0_  = ~n29852 ;
  assign \g224650/_0_  = ~n29884 ;
  assign \g224651/_0_  = ~n29916 ;
  assign \g224652/_0_  = ~n29942 ;
  assign \g224690/_0_  = ~n29968 ;
  assign \g224691/_3_  = ~n29998 ;
  assign \g224692/_3_  = ~n30029 ;
  assign \g224693/_0_  = ~n30057 ;
  assign \g224694/_0_  = ~n30135 ;
  assign \g224695/_3_  = ~n30165 ;
  assign \g224723/_0_  = ~n30207 ;
  assign \g224724/_0_  = ~n30241 ;
  assign \g224725/_0_  = ~n30267 ;
  assign \g224726/_0_  = ~n30299 ;
  assign \g226372/_0_  = ~n30397 ;
  assign \g226373/_3_  = ~n30490 ;
  assign \g226549/_3_  = ~n30586 ;
  assign \g226550/_0_  = ~n30683 ;
  assign \g226616/_0_  = ~n30720 ;
  assign \g226635/_0_  = n30751 ;
  assign \g226636/_0_  = ~n30838 ;
  assign \g226637/_0_  = ~n30872 ;
  assign \g226638/_0_  = ~n30912 ;
  assign \g226639/_0_  = ~n30942 ;
  assign \g226640/_0_  = ~n30978 ;
  assign \g226641/_3_  = ~n31068 ;
  assign \g226642/_0_  = ~n31103 ;
  assign \g226643/_0_  = ~n31135 ;
  assign \g226644/_0_  = ~n31162 ;
  assign \g226645/_0_  = ~n31258 ;
  assign \g226646/_0_  = ~n31299 ;
  assign \g226692/_3_  = ~n31332 ;
  assign \g226693/_0_  = ~n31354 ;
  assign \g226694/_3_  = ~n31387 ;
  assign \g226695/_3_  = ~n31420 ;
  assign \g226696/_3_  = ~n31453 ;
  assign \g226697/_0_  = ~n31536 ;
  assign \g226698/_0_  = ~n31565 ;
  assign \g226699/_0_  = ~n31595 ;
  assign \g226728/_0_  = ~n31631 ;
  assign \g226729/_0_  = ~n31663 ;
  assign \g226730/_0_  = ~n31690 ;
  assign \g226731/_0_  = ~n31714 ;
  assign \g226732/_0_  = ~n31739 ;
  assign \g226759/_0_  = ~n31762 ;
  assign \g228250/_0_  = ~n31858 ;
  assign \g228396/_0_  = ~n31955 ;
  assign \g228397/_0_  = ~n32042 ;
  assign \g228566/_0_  = ~n32138 ;
  assign \g228567/_0_  = ~n32175 ;
  assign \g228568/_0_  = ~n32267 ;
  assign \g228609/_0_  = ~n32296 ;
  assign \g228610/_3_  = ~n32390 ;
  assign \g228688/_0_  = ~n32422 ;
  assign \g228689/_0_  = n32453 ;
  assign \g228690/_3_  = ~n32492 ;
  assign \g228691/_0_  = ~n32526 ;
  assign \g228692/_0_  = ~n32548 ;
  assign \g228693/_0_  = ~n32587 ;
  assign \g228694/_0_  = ~n32618 ;
  assign \g228695/_0_  = ~n32654 ;
  assign \g228696/_0_  = ~n32743 ;
  assign \g228697/_0_  = n32773 ;
  assign \g228698/_0_  = ~n32822 ;
  assign \g228699/_0_  = ~n32853 ;
  assign \g228700/_0_  = ~n32879 ;
  assign \g228748/_0_  = ~n32910 ;
  assign \g228749/_3_  = ~n32942 ;
  assign \g228750/_0_  = ~n32969 ;
  assign \g228751/_0_  = ~n33047 ;
  assign \g228752/_0_  = ~n33075 ;
  assign \g228753/_0_  = ~n33102 ;
  assign \g228784/_0_  = ~n33140 ;
  assign \g228785/_0_  = ~n33175 ;
  assign \g228786/_0_  = ~n33202 ;
  assign \g228787/_3_  = ~n33226 ;
  assign \g230339/_0_  = ~n33318 ;
  assign \g230340/_0_  = ~n33414 ;
  assign \g230546/_0_  = ~n33512 ;
  assign \g230580/_0_  = ~n33605 ;
  assign \g230679/_0_  = ~n33636 ;
  assign \g230680/_0_  = n33666 ;
  assign \g230681/_0_  = ~n33767 ;
  assign \g230682/_0_  = ~n33795 ;
  assign \g230683/_0_  = ~n33880 ;
  assign \g230684/_0_  = ~n33915 ;
  assign \g230685/_0_  = ~n33959 ;
  assign \g230686/_0_  = ~n33999 ;
  assign \g230687/_0_  = ~n34085 ;
  assign \g230688/_0_  = ~n34119 ;
  assign \g230689/_3_  = ~n34163 ;
  assign \g230690/_0_  = ~n34194 ;
  assign \g230710/_0_  = ~n34226 ;
  assign \g230766/_0_  = ~n34249 ;
  assign \g230767/_0_  = ~n34283 ;
  assign \g230768/_0_  = ~n34318 ;
  assign \g230769/_3_  = ~n34351 ;
  assign \g230770/_0_  = ~n34431 ;
  assign \g230771/_0_  = ~n34462 ;
  assign \g230772/_0_  = ~n34489 ;
  assign \g230773/_3_  = ~n34521 ;
  assign \g230810/_0_  = ~n34557 ;
  assign \g230811/_0_  = ~n34590 ;
  assign \g230812/_0_  = ~n34617 ;
  assign \g230813/_0_  = ~n34643 ;
  assign \g230814/_0_  = ~n34664 ;
  assign \g230840/_3_  = ~n34689 ;
  assign \g232196/_3_  = ~n34781 ;
  assign \g232469/_0_  = ~n34875 ;
  assign \g232470/_0_  = ~n34967 ;
  assign \g232633/_0_  = ~n35060 ;
  assign \g232635/_3_  = ~n35155 ;
  assign \g232636/_0_  = ~n35190 ;
  assign \g232637/_0_  = ~n35222 ;
  assign \g232691/_0_  = ~n35319 ;
  assign \g232747/_0_  = ~n35351 ;
  assign \g232748/_0_  = n35381 ;
  assign \g232749/_3_  = ~n35419 ;
  assign \g232750/_0_  = ~n35522 ;
  assign \g232751/_0_  = ~n35557 ;
  assign \g232752/_0_  = ~n35587 ;
  assign \g232753/_0_  = ~n35613 ;
  assign \g232754/_0_  = ~n35651 ;
  assign \g232755/_0_  = ~n35692 ;
  assign \g232756/_0_  = ~n35729 ;
  assign \g232757/_0_  = ~n35759 ;
  assign \g232758/_0_  = ~n35786 ;
  assign \g232759/_0_  = ~n35812 ;
  assign \g232804/_0_  = ~n35840 ;
  assign \g232805/_0_  = ~n35866 ;
  assign \g232806/_0_  = ~n35945 ;
  assign \g232807/_0_  = ~n35969 ;
  assign \g232808/_3_  = ~n36002 ;
  assign \g232809/_0_  = ~n36033 ;
  assign \g232841/_0_  = ~n36075 ;
  assign \g232842/_3_  = ~n36100 ;
  assign \g232843/_0_  = ~n36134 ;
  assign \g232844/_0_  = ~n36162 ;
  assign \g234520/_0_  = ~n36248 ;
  assign \g234687/_0_  = ~n36342 ;
  assign \g234688/_0_  = ~n36437 ;
  assign \g234689/_0_  = ~n36525 ;
  assign \g234764/_0_  = ~n36561 ;
  assign \g234765/_0_  = n36596 ;
  assign \g234766/_0_  = ~n36694 ;
  assign \g234767/_3_  = ~n36731 ;
  assign \g234768/_0_  = ~n36762 ;
  assign \g234769/_0_  = n36840 ;
  assign \g234770/_0_  = ~n36879 ;
  assign \g234771/_0_  = ~n36919 ;
  assign \g234772/_0_  = ~n36951 ;
  assign \g234773/_0_  = ~n36992 ;
  assign \g234774/_3_  = ~n37086 ;
  assign \g234775/_0_  = ~n37123 ;
  assign \g234776/_0_  = ~n37155 ;
  assign \g234824/_3_  = ~n37188 ;
  assign \g234825/_0_  = ~n37211 ;
  assign \g234826/_0_  = ~n37253 ;
  assign \g234827/_0_  = ~n37282 ;
  assign \g234828/_3_  = ~n37316 ;
  assign \g234829/_0_  = ~n37403 ;
  assign \g234830/_0_  = ~n37431 ;
  assign \g234831/_0_  = ~n37453 ;
  assign \g234867/_0_  = ~n37492 ;
  assign \g234868/_0_  = ~n37521 ;
  assign \g234869/_0_  = ~n37546 ;
  assign \g234870/_0_  = ~n37572 ;
  assign \g234896/_0_  = ~n37597 ;
  assign \g236294/_3_  = ~n37689 ;
  assign \g236541/_0_  = ~n37789 ;
  assign \g236542/_0_  = ~n37881 ;
  assign \g236724/_0_  = ~n37914 ;
  assign \g236725/_0_  = ~n38012 ;
  assign \g236726/_0_  = ~n38050 ;
  assign \g236727/_3_  = ~n38140 ;
  assign \g236728/_0_  = ~n38170 ;
  assign \g236729/_0_  = ~n38258 ;
  assign \g236821/_0_  = n38288 ;
  assign \g236822/_3_  = ~n38330 ;
  assign \g236823/_0_  = ~n38432 ;
  assign \g236824/_3_  = ~n38469 ;
  assign \g236825/_0_  = ~n38493 ;
  assign \g236826/_0_  = ~n38525 ;
  assign \g236827/_0_  = ~n38558 ;
  assign \g236828/_0_  = ~n38591 ;
  assign \g236829/_0_  = ~n38631 ;
  assign \g236830/_0_  = ~n38665 ;
  assign \g236831/_0_  = ~n38695 ;
  assign \g236832/_0_  = ~n38720 ;
  assign \g236877/_0_  = ~n38753 ;
  assign \g236878/_3_  = ~n38786 ;
  assign \g236879/_0_  = ~n38814 ;
  assign \g236880/_0_  = ~n38893 ;
  assign \g236881/_0_  = ~n38924 ;
  assign \g236882/_0_  = ~n38945 ;
  assign \g236914/_0_  = ~n38983 ;
  assign \g236915/_0_  = ~n39009 ;
  assign \g236916/_0_  = ~n39047 ;
  assign \g236917/_0_  = ~n39075 ;
  assign \g238530/_0_  = ~n39167 ;
  assign \g238531/_3_  = ~n39261 ;
  assign \g238723/_0_  = ~n39358 ;
  assign \g238724/_0_  = ~n39451 ;
  assign \g238725/_0_  = ~n39543 ;
  assign \g238840/_0_  = ~n39575 ;
  assign \g238841/_0_  = n39605 ;
  assign \g238842/_0_  = ~n39694 ;
  assign \g238843/_3_  = ~n39730 ;
  assign \g238844/_0_  = ~n39765 ;
  assign \g238845/_0_  = ~n39795 ;
  assign \g238846/_0_  = ~n39832 ;
  assign \g238847/_0_  = ~n39874 ;
  assign \g238848/_0_  = ~n39904 ;
  assign \g238849/_0_  = ~n39991 ;
  assign \g238850/_0_  = ~n40028 ;
  assign \g238851/_3_  = ~n40065 ;
  assign \g238852/_0_  = ~n40094 ;
  assign \g238924/_0_  = ~n40116 ;
  assign \g238925/_0_  = ~n40147 ;
  assign \g238926/_0_  = ~n40176 ;
  assign \g238927/_3_  = ~n40209 ;
  assign \g238928/_0_  = ~n40287 ;
  assign \g238929/_0_  = ~n40318 ;
  assign \g238930/_0_  = ~n40345 ;
  assign \g238965/_0_  = ~n40382 ;
  assign \g238966/_0_  = ~n40421 ;
  assign \g238967/_0_  = ~n40450 ;
  assign \g238968/_0_  = ~n40479 ;
  assign \g238969/_0_  = ~n40503 ;
  assign \g238996/_0_  = ~n40531 ;
  assign \g240353/_3_  = ~n40622 ;
  assign \g240640/_0_  = ~n40719 ;
  assign \g240641/_0_  = ~n40811 ;
  assign \g240813/_0_  = ~n40849 ;
  assign \g240814/_0_  = ~n40947 ;
  assign \g240815/_3_  = ~n41040 ;
  assign \g240816/_0_  = ~n41076 ;
  assign \g240817/_0_  = ~n41165 ;
  assign \g240818/_0_  = ~n41196 ;
  assign \g240925/_0_  = ~n41229 ;
  assign \g240926/_0_  = n41259 ;
  assign \g240927/_3_  = ~n41297 ;
  assign \g240928/_0_  = ~n41398 ;
  assign \g240929/_3_  = ~n41433 ;
  assign \g240930/_0_  = ~n41458 ;
  assign \g240931/_0_  = ~n41489 ;
  assign \g240932/_0_  = ~n41527 ;
  assign \g240933/_0_  = ~n41559 ;
  assign \g240934/_0_  = ~n41598 ;
  assign \g240935/_0_  = ~n41632 ;
  assign \g240936/_0_  = ~n41660 ;
  assign \g240937/_0_  = ~n41685 ;
  assign \g240984/_0_  = ~n41717 ;
  assign \g240985/_3_  = ~n41750 ;
  assign \g240986/_0_  = ~n41777 ;
  assign \g240987/_0_  = ~n41860 ;
  assign \g240988/_0_  = ~n41891 ;
  assign \g240989/_0_  = ~n41915 ;
  assign \g241021/_0_  = ~n41951 ;
  assign \g241022/_0_  = ~n41977 ;
  assign \g241023/_0_  = ~n42012 ;
  assign \g241024/_0_  = ~n42043 ;
  assign \g242616/_0_  = ~n42134 ;
  assign \g242617/_3_  = ~n42228 ;
  assign \g242815/_0_  = ~n42325 ;
  assign \g242816/_0_  = ~n42423 ;
  assign \g242817/_0_  = ~n42518 ;
  assign \g242955/_0_  = ~n42548 ;
  assign \g242956/_0_  = n42582 ;
  assign \g242957/_0_  = ~n42681 ;
  assign \g242958/_3_  = ~n42713 ;
  assign \g242959/_0_  = ~n42745 ;
  assign \g242960/_0_  = ~n42780 ;
  assign \g242961/_0_  = ~n42814 ;
  assign \g242962/_0_  = ~n42854 ;
  assign \g242963/_3_  = ~n42944 ;
  assign \g242964/_0_  = ~n42975 ;
  assign \g242965/_0_  = ~n43012 ;
  assign \g242966/_0_  = ~n43049 ;
  assign \g242967/_0_  = ~n43080 ;
  assign \g243037/_3_  = ~n43116 ;
  assign \g243038/_0_  = ~n43140 ;
  assign \g243039/_0_  = ~n43175 ;
  assign \g243040/_0_  = ~n43205 ;
  assign \g243041/_3_  = ~n43236 ;
  assign \g243042/_0_  = ~n43323 ;
  assign \g243043/_0_  = ~n43351 ;
  assign \g243044/_0_  = ~n43378 ;
  assign \g243078/_0_  = ~n43412 ;
  assign \g243079/_0_  = ~n43447 ;
  assign \g243080/_0_  = ~n43478 ;
  assign \g243081/_0_  = ~n43507 ;
  assign \g243082/_0_  = ~n43531 ;
  assign \g243109/_0_  = ~n43555 ;
  assign \g244465/_3_  = ~n43598 ;
  assign \g244753/_3_  = ~n43695 ;
  assign \g244754/_0_  = ~n43787 ;
  assign \g244924/_0_  = ~n43883 ;
  assign \g244925/_0_  = ~n43917 ;
  assign \g244926/_3_  = ~n44007 ;
  assign \g244927/_0_  = ~n44040 ;
  assign \g244928/_0_  = ~n44131 ;
  assign \g245035/_0_  = ~n44164 ;
  assign \g245036/_0_  = n44194 ;
  assign \g245037/_0_  = ~n44294 ;
  assign \g245038/_3_  = ~n44328 ;
  assign \g245039/_3_  = ~n44370 ;
  assign \g245040/_0_  = ~n44393 ;
  assign \g245041/_0_  = ~n44426 ;
  assign \g245043/_0_  = ~n44460 ;
  assign \g245045/_0_  = ~n44490 ;
  assign \g245046/_0_  = ~n44529 ;
  assign \g245047/_0_  = ~n44552 ;
  assign \g245092/_0_  = ~n44590 ;
  assign \g245093/_3_  = ~n44623 ;
  assign \g245094/_0_  = ~n44649 ;
  assign \g245095/_0_  = ~n44680 ;
  assign \g245096/_0_  = ~n44757 ;
  assign \g245097/_0_  = ~n44782 ;
  assign \g245129/_0_  = ~n44823 ;
  assign \g245130/_0_  = ~n44849 ;
  assign \g245131/_0_  = ~n44885 ;
  assign \g245132/_0_  = ~n44915 ;
  assign \g246715/_0_  = ~n45007 ;
  assign \g246716/_3_  = ~n45100 ;
  assign \g246911/_0_  = ~n45197 ;
  assign \g246912/_0_  = ~n45293 ;
  assign \g246913/_0_  = ~n45384 ;
  assign \g247057/_0_  = ~n45416 ;
  assign \g247058/_0_  = n45446 ;
  assign \g247059/_0_  = ~n45545 ;
  assign \g247060/_0_  = ~n45577 ;
  assign \g247061/_0_  = ~n45608 ;
  assign \g247062/_3_  = ~n45646 ;
  assign \g247063/_0_  = ~n45680 ;
  assign \g247064/_0_  = ~n45720 ;
  assign \g247065/_0_  = ~n45751 ;
  assign \g247066/_0_  = ~n45788 ;
  assign \g247067/_3_  = ~n45878 ;
  assign \g247068/_0_  = ~n45915 ;
  assign \g247069/_0_  = ~n45944 ;
  assign \g247137/_3_  = ~n45980 ;
  assign \g247138/_0_  = ~n46002 ;
  assign \g247139/_0_  = ~n46035 ;
  assign \g247140/_0_  = ~n46063 ;
  assign \g247141/_3_  = ~n46096 ;
  assign \g247142/_0_  = ~n46180 ;
  assign \g247143/_0_  = ~n46211 ;
  assign \g247144/_0_  = ~n46238 ;
  assign \g247179/_0_  = ~n46274 ;
  assign \g247180/_0_  = ~n46309 ;
  assign \g247181/_0_  = ~n46338 ;
  assign \g247182/_0_  = ~n46367 ;
  assign \g247183/_0_  = ~n46393 ;
  assign \g247210/_0_  = ~n46417 ;
  assign \g248581/_3_  = ~n46510 ;
  assign \g248828/_0_  = ~n46606 ;
  assign \g248829/_0_  = ~n46697 ;
  assign \g249033/_0_  = ~n46729 ;
  assign \g249035/_0_  = ~n46768 ;
  assign \g249036/_3_  = ~n46857 ;
  assign \g249037/_0_  = ~n46887 ;
  assign \g249038/_0_  = ~n46978 ;
  assign \g249147/_0_  = ~n47072 ;
  assign \g249148/_0_  = n47106 ;
  assign \g249149/_3_  = ~n47149 ;
  assign \g249150/_0_  = ~n47199 ;
  assign \g249152/_0_  = ~n47239 ;
  assign \g249153/_0_  = ~n47272 ;
  assign \g249155/_0_  = ~n47306 ;
  assign \g249156/_0_  = ~n47336 ;
  assign \g249157/_0_  = ~n47363 ;
  assign \g249200/_3_  = ~n47398 ;
  assign \g249201/_0_  = ~n47434 ;
  assign \g249202/_0_  = ~n47465 ;
  assign \g249203/_3_  = ~n47496 ;
  assign \g249204/_0_  = ~n47525 ;
  assign \g249205/_0_  = ~n47612 ;
  assign \g249206/_0_  = ~n47640 ;
  assign \g249207/_0_  = ~n47666 ;
  assign \g249239/_0_  = ~n47700 ;
  assign \g249240/_0_  = ~n47726 ;
  assign \g249241/_0_  = ~n47761 ;
  assign \g249242/_0_  = ~n47792 ;
  assign \g250815/_0_  = ~n47886 ;
  assign \g251006/_0_  = ~n47986 ;
  assign \g251007/_0_  = ~n48080 ;
  assign \g251008/_0_  = ~n48171 ;
  assign \g251009/_3_  = ~n48262 ;
  assign \g251160/_0_  = ~n48293 ;
  assign \g251161/_0_  = n48324 ;
  assign \g251162/_0_  = ~n48429 ;
  assign \g251163/_3_  = ~n48467 ;
  assign \g251164/_0_  = ~n48505 ;
  assign \g251165/_0_  = ~n48532 ;
  assign \g251166/_0_  = ~n48566 ;
  assign \g251167/_0_  = ~n48600 ;
  assign \g251168/_0_  = ~n48683 ;
  assign \g251169/_0_  = ~n48721 ;
  assign \g251170/_3_  = ~n48764 ;
  assign \g251171/_0_  = ~n48794 ;
  assign \g251245/_3_  = ~n48825 ;
  assign \g251246/_0_  = ~n48864 ;
  assign \g251247/_0_  = ~n48888 ;
  assign \g251248/_0_  = ~n48916 ;
  assign \g251249/_3_  = ~n48949 ;
  assign \g251250/_0_  = ~n49028 ;
  assign \g251251/_0_  = ~n49057 ;
  assign \g251252/_0_  = ~n49084 ;
  assign \g251286/_0_  = ~n49125 ;
  assign \g251287/_0_  = ~n49157 ;
  assign \g251288/_0_  = ~n49193 ;
  assign \g251289/_0_  = ~n49224 ;
  assign \g251290/_0_  = ~n49251 ;
  assign \g251291/_0_  = ~n49275 ;
  assign \g251318/_0_  = ~n49300 ;
  assign \g252698/_3_  = ~n49393 ;
  assign \g252942/_0_  = ~n49486 ;
  assign \g252943/_0_  = ~n49576 ;
  assign \g253118/_0_  = ~n49608 ;
  assign \g253119/_0_  = ~n49636 ;
  assign \g253120/_0_  = ~n49734 ;
  assign \g253121/_0_  = ~n49770 ;
  assign \g253122/_3_  = ~n49860 ;
  assign \g253123/_0_  = ~n49890 ;
  assign \g253236/_0_  = n49925 ;
  assign \g253237/_3_  = ~n49967 ;
  assign \g253238/_3_  = ~n50058 ;
  assign \g253239/_0_  = ~n50160 ;
  assign \g253240/_0_  = ~n50197 ;
  assign \g253241/_0_  = ~n50237 ;
  assign \g253242/_0_  = ~n50270 ;
  assign \g253243/_0_  = ~n50310 ;
  assign \g253244/_0_  = ~n50340 ;
  assign \g253245/_0_  = ~n50372 ;
  assign \g253246/_0_  = ~n50399 ;
  assign \g253247/_0_  = ~n50425 ;
  assign \g253248/_0_  = ~n50452 ;
  assign \g253306/_0_  = ~n50482 ;
  assign \g253307/_3_  = ~n50513 ;
  assign \g253308/_0_  = ~n50539 ;
  assign \g253309/_0_  = ~n50630 ;
  assign \g253310/_0_  = ~n50659 ;
  assign \g253311/_0_  = ~n50685 ;
  assign \g253356/_0_  = ~n50718 ;
  assign \g253357/_0_  = ~n50744 ;
  assign \g253358/_0_  = ~n50775 ;
  assign \g253359/_0_  = ~n50803 ;
  assign \g253436/_3_  = ~n50892 ;
  assign \g253437/_0_  = ~n50989 ;
  assign \g253438/_0_  = ~n51024 ;
  assign \g253469/_3_  = ~n51061 ;
  assign \g253470/_3_  = ~n51147 ;
  assign \g253471/_3_  = ~n51175 ;
  assign \g253521/_0_  = ~n51259 ;
  assign \g253522/_0_  = ~n51346 ;
  assign \g253523/_0_  = ~n51389 ;
  assign \g253524/_3_  = ~n51422 ;
  assign \g256730/_3_  = ~n51513 ;
  assign \g256731/_3_  = ~n51607 ;
  assign \g256927/_0_  = ~n51697 ;
  assign \g256928/_0_  = ~n51792 ;
  assign \g256929/_3_  = ~n51890 ;
  assign \g257049/_0_  = ~n51924 ;
  assign \g257050/_0_  = ~n51956 ;
  assign \g257051/_3_  = ~n51990 ;
  assign \g257052/_0_  = ~n52028 ;
  assign \g257053/_0_  = n52051 ;
  assign \g257054/_0_  = ~n52141 ;
  assign \g257055/_3_  = ~n52175 ;
  assign \g257056/_0_  = ~n52261 ;
  assign \g257057/_0_  = ~n52299 ;
  assign \g257058/_3_  = ~n52341 ;
  assign \g257059/_0_  = ~n52384 ;
  assign \g257060/_0_  = ~n52415 ;
  assign \g257082/_0_  = ~n52446 ;
  assign \g257125/_3_  = ~n52481 ;
  assign \g257126/_0_  = ~n52504 ;
  assign \g257127/_0_  = ~n52536 ;
  assign \g257128/_3_  = ~n52567 ;
  assign \g257129/_3_  = ~n52605 ;
  assign \g257130/_0_  = ~n52688 ;
  assign \g257131/_0_  = ~n52712 ;
  assign \g257132/_0_  = ~n52741 ;
  assign \g257163/_0_  = ~n52779 ;
  assign \g257164/_0_  = ~n52811 ;
  assign \g257165/_0_  = ~n52839 ;
  assign \g257166/_0_  = ~n52864 ;
  assign \g257167/_0_  = ~n52892 ;
  assign \g257194/_0_  = ~n52916 ;
  assign \g258552/_0_  = ~n53010 ;
  assign \g258850/_0_  = ~n53102 ;
  assign \g258851/_3_  = ~n53196 ;
  assign \g258993/_0_  = ~n53231 ;
  assign \g258994/_0_  = ~n53327 ;
  assign \g258995/_0_  = ~n53361 ;
  assign \g258996/_0_  = ~n53451 ;
  assign \g259026/_3_  = ~n53541 ;
  assign \g259027/_0_  = ~n53573 ;
  assign \g259105/_0_  = n53602 ;
  assign \g259106/_0_  = ~n53637 ;
  assign \g259107/_3_  = ~n53679 ;
  assign \g259108/_0_  = ~n53780 ;
  assign \g259109/_3_  = ~n53814 ;
  assign \g259110/_0_  = ~n53848 ;
  assign \g259111/_0_  = ~n53886 ;
  assign \g259112/_0_  = ~n53925 ;
  assign \g259113/_0_  = ~n53955 ;
  assign \g259114/_0_  = ~n53984 ;
  assign \g259115/_0_  = ~n54016 ;
  assign \g259116/_0_  = ~n54042 ;
  assign \g259117/_0_  = ~n54072 ;
  assign \g259163/_3_  = ~n54103 ;
  assign \g259164/_3_  = ~n54135 ;
  assign \g259165/_0_  = ~n54158 ;
  assign \g259166/_0_  = ~n54239 ;
  assign \g259167/_0_  = ~n54263 ;
  assign \g259168/_0_  = ~n54292 ;
  assign \g259197/_0_  = ~n54331 ;
  assign \g259198/_0_  = ~n54367 ;
  assign \g259199/_0_  = ~n54395 ;
  assign \g259200/_0_  = ~n54421 ;
  assign \g260774/_0_  = ~n54513 ;
  assign \g260792/_3_  = ~n54607 ;
  assign \g260991/_0_  = ~n54702 ;
  assign \g261013/_0_  = ~n54800 ;
  assign \g261070/_0_  = ~n54894 ;
  assign \g261125/_0_  = ~n54926 ;
  assign \g261126/_0_  = ~n54959 ;
  assign \g261128/_0_  = ~n55042 ;
  assign \g261129/_0_  = ~n55083 ;
  assign \g261130/_0_  = n55112 ;
  assign \g261131/_0_  = ~n55148 ;
  assign \g261132/_0_  = ~n55238 ;
  assign \g261133/_0_  = ~n55272 ;
  assign \g261134/_3_  = ~n55311 ;
  assign \g261135/_0_  = ~n55354 ;
  assign \g261136/_0_  = ~n55386 ;
  assign \g261158/_3_  = ~n55415 ;
  assign \g261206/_0_  = ~n55445 ;
  assign \g261207/_0_  = ~n55474 ;
  assign \g261208/_0_  = ~n55498 ;
  assign \g261209/_0_  = ~n55531 ;
  assign \g261210/_3_  = ~n55567 ;
  assign \g261211/_0_  = ~n55646 ;
  assign \g261212/_3_  = ~n55681 ;
  assign \g261213/_0_  = ~n55705 ;
  assign \g261248/_0_  = ~n55746 ;
  assign \g261249/_0_  = ~n55778 ;
  assign \g261250/_0_  = ~n55806 ;
  assign \g261251/_0_  = ~n55830 ;
  assign \g261252/_0_  = ~n55864 ;
  assign \g261279/_0_  = ~n55891 ;
  assign \g262658/_3_  = ~n55986 ;
  assign \g262949/_0_  = ~n56080 ;
  assign \g263008/_3_  = ~n56179 ;
  assign \g263092/_0_  = ~n56213 ;
  assign \g263093/_0_  = ~n56308 ;
  assign \g263099/_0_  = ~n56344 ;
  assign \g263100/_0_  = ~n56433 ;
  assign \g263101/_0_  = ~n56464 ;
  assign \g263159/_3_  = ~n56554 ;
  assign \g263204/_3_  = ~n56589 ;
  assign \g263205/_0_  = ~n56627 ;
  assign \g263206/_0_  = ~n56716 ;
  assign \g263208/_0_  = ~n56742 ;
  assign \g263209/_0_  = ~n56778 ;
  assign \g263210/_0_  = ~n56808 ;
  assign \g263211/_0_  = ~n56844 ;
  assign \g263212/_0_  = ~n56881 ;
  assign \g263213/_0_  = n56911 ;
  assign \g263214/_0_  = ~n56940 ;
  assign \g263215/_3_  = ~n56974 ;
  assign \g263216/_0_  = ~n57015 ;
  assign \g263260/_0_  = ~n57041 ;
  assign \g263261/_0_  = ~n57073 ;
  assign \g263262/_3_  = ~n57105 ;
  assign \g263263/_0_  = ~n57192 ;
  assign \g263264/_0_  = ~n57220 ;
  assign \g263265/_0_  = ~n57249 ;
  assign \g263297/_0_  = ~n57274 ;
  assign \g263298/_0_  = ~n57308 ;
  assign \g263299/_0_  = ~n57343 ;
  assign \g263300/_0_  = ~n57374 ;
  assign \g264930/_0_  = ~n57462 ;
  assign \g264946/_3_  = ~n57553 ;
  assign \g265143/_0_  = ~n57653 ;
  assign \g265144/_0_  = ~n57751 ;
  assign \g265152/_0_  = ~n57846 ;
  assign \g265222/_0_  = ~n57882 ;
  assign \g265223/_0_  = ~n57965 ;
  assign \g265224/_0_  = ~n57998 ;
  assign \g265225/_0_  = ~n58027 ;
  assign \g265226/_0_  = ~n58128 ;
  assign \g265227/_3_  = ~n58160 ;
  assign \g265228/_0_  = n58192 ;
  assign \g265229/_0_  = ~n58220 ;
  assign \g265230/_0_  = ~n58254 ;
  assign \g265231/_0_  = ~n58294 ;
  assign \g265232/_0_  = ~n58333 ;
  assign \g265233/_3_  = ~n58376 ;
  assign \g265234/_0_  = ~n58406 ;
  assign \g265306/_0_  = ~n58438 ;
  assign \g265307/_0_  = ~n58468 ;
  assign \g265308/_3_  = ~n58500 ;
  assign \g265309/_3_  = ~n58534 ;
  assign \g265310/_0_  = ~n58617 ;
  assign \g265311/_0_  = ~n58642 ;
  assign \g265312/_0_  = ~n58669 ;
  assign \g265313/_0_  = ~n58691 ;
  assign \g265348/_0_  = ~n58727 ;
  assign \g265349/_0_  = ~n58762 ;
  assign \g265350/_0_  = ~n58790 ;
  assign \g265351/_0_  = ~n58816 ;
  assign \g265379/_0_  = ~n58842 ;
  assign \g266965/_3_  = ~n58937 ;
  assign \g267049/_3_  = ~n59033 ;
  assign \g267050/_0_  = ~n59123 ;
  assign \g267215/_0_  = ~n59157 ;
  assign \g267216/_0_  = ~n59252 ;
  assign \g267263/_0_  = ~n59286 ;
  assign \g267264/_3_  = ~n59380 ;
  assign \g267265/_0_  = ~n59413 ;
  assign \g267266/_0_  = ~n59504 ;
  assign \g267314/_3_  = ~n59546 ;
  assign \g267315/_0_  = ~n59648 ;
  assign \g267316/_0_  = ~n59688 ;
  assign \g267317/_0_  = ~n59715 ;
  assign \g267318/_0_  = n59743 ;
  assign \g267319/_0_  = ~n59787 ;
  assign \g267320/_3_  = ~n59818 ;
  assign \g267321/_0_  = ~n59842 ;
  assign \g267322/_0_  = ~n59872 ;
  assign \g267324/_0_  = ~n59902 ;
  assign \g267325/_0_  = ~n59931 ;
  assign \g267326/_0_  = ~n59962 ;
  assign \g267372/_0_  = ~n59991 ;
  assign \g267373/_3_  = ~n60023 ;
  assign \g267374/_0_  = ~n60051 ;
  assign \g267375/_0_  = ~n60138 ;
  assign \g267376/_0_  = ~n60162 ;
  assign \g267377/_0_  = ~n60188 ;
  assign \g267409/_0_  = ~n60222 ;
  assign \g267410/_0_  = ~n60257 ;
  assign \g267411/_0_  = ~n60288 ;
  assign \g267412/_0_  = ~n60312 ;
  assign \g269004/_0_  = ~n60398 ;
  assign \g269099/_3_  = ~n60492 ;
  assign \g269202/_0_  = ~n60591 ;
  assign \g269226/_0_  = ~n60678 ;
  assign \g269333/_3_  = ~n60712 ;
  assign \g269334/_0_  = ~n60799 ;
  assign \g269335/_0_  = ~n60833 ;
  assign \g269355/_0_  = ~n60876 ;
  assign \g269356/_0_  = ~n60910 ;
  assign \g269357/_3_  = ~n61000 ;
  assign \g269358/_0_  = ~n61038 ;
  assign \g269359/_0_  = ~n61070 ;
  assign \g269360/_0_  = ~n61171 ;
  assign \g269361/_0_  = ~n61207 ;
  assign \g269362/_0_  = n61240 ;
  assign \g269363/_0_  = ~n61275 ;
  assign \g269364/_0_  = ~n61315 ;
  assign \g269414/_0_  = ~n61338 ;
  assign \g269415/_0_  = ~n61367 ;
  assign \g269416/_0_  = ~n61399 ;
  assign \g269417/_0_  = ~n61426 ;
  assign \g269418/_3_  = ~n61458 ;
  assign \g269419/_0_  = ~n61491 ;
  assign \g269420/_3_  = ~n61525 ;
  assign \g269421/_0_  = ~n61603 ;
  assign \g269456/_0_  = ~n61648 ;
  assign \g269457/_0_  = ~n61671 ;
  assign \g269458/_0_  = ~n61702 ;
  assign \g269459/_0_  = ~n61728 ;
  assign \g269460/_0_  = ~n61759 ;
  assign \g269487/_0_  = ~n61784 ;
  assign \g271006/_3_  = ~n61878 ;
  assign \g271186/_3_  = ~n61973 ;
  assign \g271187/_0_  = ~n62062 ;
  assign \g271299/_0_  = ~n62161 ;
  assign \g271300/_0_  = ~n62251 ;
  assign \g271301/_3_  = ~n62341 ;
  assign \g271302/_0_  = ~n62377 ;
  assign \g271303/_0_  = ~n62412 ;
  assign \g271352/_0_  = ~n62445 ;
  assign \g271410/_0_  = n62480 ;
  assign \g271411/_0_  = ~n62504 ;
  assign \g271412/_0_  = ~n62593 ;
  assign \g271413/_0_  = ~n62632 ;
  assign \g271414/_0_  = ~n62666 ;
  assign \g271415/_0_  = ~n62702 ;
  assign \g271416/_0_  = ~n62746 ;
  assign \g271417/_3_  = ~n62782 ;
  assign \g271418/_3_  = ~n62816 ;
  assign \g271419/_0_  = ~n62847 ;
  assign \g271420/_0_  = ~n62880 ;
  assign \g271421/_0_  = ~n62913 ;
  assign \g271422/_0_  = ~n62944 ;
  assign \g271468/_3_  = ~n62975 ;
  assign \g271469/_0_  = ~n63003 ;
  assign \g271470/_0_  = ~n63087 ;
  assign \g271471/_0_  = ~n63113 ;
  assign \g271472/_0_  = ~n63137 ;
  assign \g271473/_0_  = ~n63159 ;
  assign \g271505/_0_  = ~n63184 ;
  assign \g271506/_0_  = ~n63219 ;
  assign \g271507/_0_  = ~n63254 ;
  assign \g271508/_0_  = ~n63282 ;
  assign \g273135/_0_  = ~n63379 ;
  assign \g273136/_3_  = ~n63472 ;
  assign \g273362/_0_  = ~n63571 ;
  assign \g273373/_0_  = ~n63666 ;
  assign \g273374/_0_  = ~n63761 ;
  assign \g273431/_0_  = ~n63795 ;
  assign \g273432/_0_  = ~n63832 ;
  assign \g273433/_3_  = ~n63926 ;
  assign \g273434/_0_  = ~n63956 ;
  assign \g273435/_0_  = n63983 ;
  assign \g273436/_0_  = ~n64085 ;
  assign \g273437/_3_  = ~n64117 ;
  assign \g273438/_0_  = ~n64154 ;
  assign \g273439/_0_  = ~n64188 ;
  assign \g273441/_0_  = ~n64223 ;
  assign \g273442/_0_  = ~n64260 ;
  assign \g273443/_0_  = ~n64292 ;
  assign \g273515/_3_  = ~n64325 ;
  assign \g273516/_0_  = ~n64355 ;
  assign \g273517/_0_  = ~n64389 ;
  assign \g273518/_3_  = ~n64424 ;
  assign \g273519/_0_  = ~n64447 ;
  assign \g273520/_0_  = ~n64473 ;
  assign \g273521/_0_  = ~n64496 ;
  assign \g273522/_0_  = ~n64572 ;
  assign \g273557/_0_  = ~n64616 ;
  assign \g273558/_0_  = ~n64648 ;
  assign \g273559/_0_  = ~n64674 ;
  assign \g273560/_0_  = ~n64699 ;
  assign \g273561/_0_  = ~n64724 ;
  assign \g273588/_0_  = ~n64749 ;
  assign \g274960/_3_  = ~n64841 ;
  assign \g275266/_3_  = ~n64940 ;
  assign \g275327/_0_  = ~n65030 ;
  assign \g275396/_0_  = ~n65065 ;
  assign \g275397/_3_  = ~n65155 ;
  assign \g275398/_0_  = ~n65190 ;
  assign \g275455/_0_  = ~n65280 ;
  assign \g275456/_0_  = ~n65313 ;
  assign \g275463/_0_  = ~n65410 ;
  assign \g275510/_3_  = ~n65451 ;
  assign \g275511/_0_  = ~n65484 ;
  assign \g275512/_0_  = n65513 ;
  assign \g275513/_0_  = ~n65544 ;
  assign \g275514/_3_  = ~n65581 ;
  assign \g275515/_0_  = ~n65611 ;
  assign \g275516/_0_  = ~n65699 ;
  assign \g275517/_0_  = ~n65733 ;
  assign \g275518/_0_  = ~n65778 ;
  assign \g275519/_0_  = ~n65801 ;
  assign \g275520/_0_  = ~n65836 ;
  assign \g275521/_0_  = ~n65866 ;
  assign \g275522/_0_  = ~n65902 ;
  assign \g275568/_0_  = ~n65930 ;
  assign \g275569/_0_  = ~n65959 ;
  assign \g275570/_0_  = ~n65984 ;
  assign \g275571/_0_  = ~n66067 ;
  assign \g275572/_3_  = ~n66101 ;
  assign \g275573/_0_  = ~n66123 ;
  assign \g275605/_0_  = ~n66160 ;
  assign \g275606/_0_  = ~n66194 ;
  assign \g275607/_0_  = ~n66219 ;
  assign \g275608/_0_  = ~n66249 ;
  assign \g277189/_0_  = ~n66344 ;
  assign \g277294/_3_  = ~n66441 ;
  assign \g277367/_0_  = ~n66536 ;
  assign \g277456/_0_  = ~n66630 ;
  assign \g277457/_0_  = ~n66723 ;
  assign \g277512/_0_  = ~n66764 ;
  assign \g277513/_0_  = ~n66863 ;
  assign \g277514/_3_  = ~n66953 ;
  assign \g277515/_0_  = ~n66990 ;
  assign \g277516/_0_  = ~n67030 ;
  assign \g277517/_3_  = ~n67059 ;
  assign \g277518/_0_  = ~n67090 ;
  assign \g277519/_0_  = ~n67126 ;
  assign \g277520/_0_  = ~n67155 ;
  assign \g277521/_0_  = ~n67184 ;
  assign \g277594/_0_  = ~n67218 ;
  assign \g277595/_0_  = ~n67248 ;
  assign \g277596/_3_  = ~n67287 ;
  assign \g277597/_0_  = ~n67311 ;
  assign \g277598/_0_  = ~n67339 ;
  assign \g277599/_0_  = ~n67418 ;
  assign \g277600/_0_  = ~n67449 ;
  assign \g277601/_3_  = ~n67483 ;
  assign \g277635/_0_  = ~n67512 ;
  assign \g277636/_0_  = ~n67555 ;
  assign \g277637/_0_  = ~n67586 ;
  assign \g277638/_0_  = ~n67610 ;
  assign \g277639/_0_  = ~n67642 ;
  assign \g277666/_0_  = ~n67667 ;
  assign \g279090/_3_  = ~n67759 ;
  assign \g279330/_0_  = ~n67857 ;
  assign \g279331/_0_  = ~n67947 ;
  assign \g279493/_3_  = ~n68036 ;
  assign \g279494/_0_  = ~n68072 ;
  assign \g279495/_0_  = ~n68108 ;
  assign \g279502/_0_  = ~n68140 ;
  assign \g279503/_0_  = ~n68228 ;
  assign \g279504/_0_  = ~n68321 ;
  assign \g279590/_0_  = ~n68359 ;
  assign \g279591/_0_  = ~n68395 ;
  assign \g279592/_0_  = ~n68426 ;
  assign \g279593/_0_  = ~n68525 ;
  assign \g279594/_3_  = ~n68559 ;
  assign \g279595/_3_  = ~n68596 ;
  assign \g279596/_0_  = ~n68635 ;
  assign \g279597/_0_  = ~n68668 ;
  assign \g279598/_0_  = ~n68694 ;
  assign \g279599/_0_  = ~n68734 ;
  assign \g279600/_0_  = ~n68765 ;
  assign \g279601/_0_  = ~n68791 ;
  assign \g279602/_0_  = n68824 ;
  assign \g279649/_0_  = ~n68910 ;
  assign \g279650/_0_  = ~n68939 ;
  assign \g279651/_0_  = ~n68964 ;
  assign \g279652/_0_  = ~n68987 ;
  assign \g279653/_0_  = ~n69018 ;
  assign \g279654/_3_  = ~n69047 ;
  assign \g279686/_0_  = ~n69084 ;
  assign \g279687/_0_  = ~n69115 ;
  assign \g279688/_0_  = ~n69143 ;
  assign \g279689/_0_  = ~n69168 ;
  assign \g281329/_0_  = ~n69260 ;
  assign \g281394/_0_  = ~n69357 ;
  assign \g281483/_0_  = ~n69446 ;
  assign \g281498/_0_  = ~n69545 ;
  assign \g281532/_0_  = ~n69640 ;
  assign \g281616/_0_  = ~n69741 ;
  assign \g281617/_0_  = ~n69776 ;
  assign \g281618/_0_  = ~n69815 ;
  assign \g281619/_0_  = n69845 ;
  assign \g281620/_0_  = ~n69873 ;
  assign \g281621/_0_  = ~n69903 ;
  assign \g281622/_0_  = ~n69987 ;
  assign \g281623/_3_  = ~n70026 ;
  assign \g281624/_0_  = ~n70061 ;
  assign \g281642/_0_  = ~n70098 ;
  assign \g281643/_0_  = ~n70130 ;
  assign \g281644/_3_  = ~n70171 ;
  assign \g281645/_0_  = ~n70201 ;
  assign \g281696/_0_  = ~n70224 ;
  assign \g281697/_3_  = ~n70258 ;
  assign \g281698/_0_  = ~n70288 ;
  assign \g281699/_0_  = ~n70366 ;
  assign \g281700/_0_  = ~n70395 ;
  assign \g281701/_0_  = ~n70427 ;
  assign \g281702/_3_  = ~n70461 ;
  assign \g281703/_0_  = ~n70486 ;
  assign \g281799/_0_  = ~n70528 ;
  assign \g281800/_0_  = ~n70558 ;
  assign \g281801/_0_  = ~n70587 ;
  assign \g281802/_0_  = ~n70618 ;
  assign \g281803/_0_  = ~n70639 ;
  assign \g281965/_0_  = ~n70664 ;
  assign \g287377/_0_  = ~n70761 ;
  assign \g287867/_0_  = ~n70860 ;
  assign \g287899/_0_  = ~n70956 ;
  assign \g288304/_0_  = ~n70984 ;
  assign \g288334/_0_  = ~n71019 ;
  assign \g288350/_0_  = ~n71116 ;
  assign \g288351/_0_  = ~n71148 ;
  assign \g288352/_3_  = ~n71239 ;
  assign \g288353/_0_  = ~n71329 ;
  assign \g288668/_0_  = ~n71370 ;
  assign \g288669/_0_  = n71398 ;
  assign \g288670/_0_  = ~n71429 ;
  assign \g288671/_0_  = ~n71466 ;
  assign \g288673/_0_  = n71500 ;
  assign \g288674/_3_  = ~n71532 ;
  assign \g288675/_0_  = ~n71621 ;
  assign \g288676/_0_  = ~n71723 ;
  assign \g288677/_0_  = ~n71746 ;
  assign \g288678/_0_  = ~n71784 ;
  assign \g288679/_0_  = ~n71816 ;
  assign \g288680/_3_  = ~n71847 ;
  assign \g288889/_0_  = ~n71874 ;
  assign \g288890/_0_  = ~n71908 ;
  assign \g288891/_0_  = ~n71941 ;
  assign \g288892/_0_  = ~n71964 ;
  assign \g288893/_3_  = ~n71997 ;
  assign \g288894/_0_  = ~n72027 ;
  assign \g288895/_0_  = ~n72059 ;
  assign \g288984/_0_  = ~n72086 ;
  assign \g288985/_0_  = ~n72116 ;
  assign \g288986/_0_  = ~n72143 ;
  assign \g294974/_0_  = ~n72239 ;
  assign \g295054/_0_  = ~n72334 ;
  assign \g295601/_0_  = ~n72428 ;
  assign \g295607/_0_  = ~n72518 ;
  assign \g296036/_0_  = ~n72604 ;
  assign \g296037/_0_  = ~n72696 ;
  assign \g296038/_0_  = ~n72798 ;
  assign \g296039/_0_  = ~n72841 ;
  assign \g296040/_0_  = ~n72873 ;
  assign \g296041/_0_  = ~n72904 ;
  assign \g296042/_0_  = ~n72935 ;
  assign \g296043/_3_  = ~n73027 ;
  assign \g296044/_0_  = ~n73062 ;
  assign \g296045/_0_  = ~n73095 ;
  assign \g296046/_0_  = n73124 ;
  assign \g296047/_0_  = ~n73156 ;
  assign \g296048/_0_  = ~n73187 ;
  assign \g296049/_3_  = ~n73220 ;
  assign \g296522/_3_  = ~n73253 ;
  assign \g296523/_3_  = ~n73276 ;
  assign \g296524/_0_  = ~n73307 ;
  assign \g296525/_0_  = ~n73350 ;
  assign \g296526/_0_  = ~n73386 ;
  assign \g296527/_0_  = ~n73418 ;
  assign \g296528/_3_  = ~n73454 ;
  assign \g296529/_0_  = ~n73484 ;
  assign \g296530/_0_  = ~n73518 ;
  assign \g296531/_0_  = ~n73547 ;
  assign \g297026/_0_  = ~n73571 ;
  assign \g297027/_0_  = ~n73600 ;
  assign \g305620/_3_  = ~n73603 ;
  assign \g305621/_3_  = ~n73606 ;
  assign \g305622/_3_  = ~n73609 ;
  assign \g305623/_3_  = ~n73612 ;
  assign \g305624/_3_  = ~n73615 ;
  assign \g305625/_3_  = ~n73618 ;
  assign \g305626/_3_  = ~n73621 ;
  assign \g305627/_3_  = ~n73624 ;
  assign \g305628/_3_  = ~n73627 ;
  assign \g305629/_3_  = ~n73630 ;
  assign \g305630/_3_  = ~n73633 ;
  assign \g305631/_3_  = ~n73636 ;
  assign \g305632/_3_  = ~n73639 ;
  assign \g305633/_3_  = ~n73642 ;
  assign \g305634/_3_  = ~n73645 ;
  assign \g305635/_3_  = ~n73648 ;
  assign \g305636/_3_  = ~n73651 ;
  assign \g305637/_3_  = ~n73654 ;
  assign \g305638/_3_  = ~n73657 ;
  assign \g305639/_3_  = ~n73660 ;
  assign \g305640/_3_  = ~n73663 ;
  assign \g305641/_3_  = ~n73666 ;
  assign \g305642/_3_  = ~n73669 ;
  assign \g305643/_3_  = ~n73672 ;
  assign \g305644/_3_  = ~n73675 ;
  assign \g305645/_3_  = ~n73678 ;
  assign \g305646/_3_  = ~n73681 ;
  assign \g305647/_3_  = ~n73684 ;
  assign \g305648/_3_  = ~n73687 ;
  assign \g305649/_3_  = ~n73690 ;
  assign \g305650/_3_  = ~n73693 ;
  assign \g305651/_3_  = ~n73696 ;
  assign \g305652/_3_  = ~n73699 ;
  assign \g305653/_3_  = ~n73702 ;
  assign \g305654/_3_  = ~n73705 ;
  assign \g305655/_3_  = ~n73708 ;
  assign \g305656/_3_  = ~n73711 ;
  assign \g305657/_3_  = ~n73714 ;
  assign \g305658/_3_  = ~n73717 ;
  assign \g305659/_3_  = ~n73720 ;
  assign \g305660/_3_  = ~n73723 ;
  assign \g305661/_3_  = ~n73726 ;
  assign \g305662/_3_  = ~n73729 ;
  assign \g305663/_3_  = ~n73732 ;
  assign \g305664/_3_  = ~n73735 ;
  assign \g305665/_3_  = ~n73738 ;
  assign \g305666/_3_  = ~n73741 ;
  assign \g305667/_3_  = ~n73744 ;
  assign \g305668/_3_  = ~n73747 ;
  assign \g305669/_3_  = ~n73750 ;
  assign \g305670/_3_  = ~n73753 ;
  assign \g305671/_3_  = ~n73756 ;
  assign \g305672/_3_  = ~n73759 ;
  assign \g305673/_3_  = ~n73762 ;
  assign \g305674/_3_  = ~n73765 ;
  assign \g305675/_3_  = ~n73768 ;
  assign \g305676/_3_  = ~n73771 ;
  assign \g305677/_3_  = ~n73774 ;
  assign \g305678/_3_  = ~n73777 ;
  assign \g305679/_3_  = ~n73780 ;
  assign \g305680/_3_  = ~n73783 ;
  assign \g305681/_3_  = ~n73786 ;
  assign \g305682/_3_  = ~n73789 ;
  assign \g305683/_3_  = ~n73792 ;
  assign \g305684/_3_  = ~n73795 ;
  assign \g305685/_3_  = ~n73798 ;
  assign \g305686/_3_  = ~n73801 ;
  assign \g305687/_3_  = ~n73804 ;
  assign \g305688/_3_  = ~n73807 ;
  assign \g305689/_3_  = ~n73810 ;
  assign \g305690/_3_  = ~n73813 ;
  assign \g305691/_3_  = ~n73816 ;
  assign \g305692/_3_  = ~n73819 ;
  assign \g305693/_3_  = ~n73822 ;
  assign \g305694/_3_  = ~n73825 ;
  assign \g305695/_3_  = ~n73828 ;
  assign \g305696/_3_  = ~n73831 ;
  assign \g305697/_3_  = ~n73834 ;
  assign \g305698/_3_  = ~n73837 ;
  assign \g305699/_3_  = ~n73840 ;
  assign \g305700/_3_  = ~n73843 ;
  assign \g305701/_3_  = ~n73846 ;
  assign \g305702/_3_  = ~n73849 ;
  assign \g305703/_3_  = ~n73852 ;
  assign \g305704/_3_  = ~n73855 ;
  assign \g305705/_3_  = ~n73858 ;
  assign \g305706/_3_  = ~n73861 ;
  assign \g305707/_3_  = ~n73864 ;
  assign \g305708/_3_  = ~n73867 ;
  assign \g305709/_3_  = ~n73870 ;
  assign \g305710/_3_  = ~n73873 ;
  assign \g305711/_3_  = ~n73876 ;
  assign \g305712/_3_  = ~n73879 ;
  assign \g305713/_3_  = ~n73882 ;
  assign \g305714/_3_  = ~n73885 ;
  assign \g305715/_3_  = ~n73888 ;
  assign \g305716/_3_  = ~n73891 ;
  assign \g305717/_3_  = ~n73894 ;
  assign \g305718/_3_  = ~n73897 ;
  assign \g305719/_3_  = ~n73900 ;
  assign \g305720/_3_  = ~n73903 ;
  assign \g305721/_3_  = ~n73906 ;
  assign \g305722/_3_  = ~n73909 ;
  assign \g305723/_3_  = ~n73912 ;
  assign \g305724/_3_  = ~n73915 ;
  assign \g305725/_3_  = ~n73918 ;
  assign \g305726/_3_  = ~n73921 ;
  assign \g305727/_3_  = ~n73924 ;
  assign \g305728/_3_  = ~n73927 ;
  assign \g305729/_3_  = ~n73930 ;
  assign \g305730/_3_  = ~n73933 ;
  assign \g305731/_3_  = ~n73936 ;
  assign \g321371/_0_  = ~n73962 ;
  assign \g321424/_0_  = ~n73986 ;
  assign \g321474/_3_  = ~n74015 ;
  assign \g321637/_3_  = ~n74040 ;
  assign \g321688/_0_  = ~n74070 ;
  assign \g321712/_0_  = ~n74105 ;
  assign \g321772/_3_  = ~n74134 ;
  assign \g321832/_0_  = ~n74162 ;
  assign \g321999/_0_  = ~n74189 ;
  assign \g322013/_3_  = ~n74215 ;
  assign \g322109/_0_  = ~n74249 ;
  assign \g322184/_0_  = ~n74274 ;
  assign \g322250/_0_  = ~n74307 ;
  assign \g322274/_0_  = n74330 ;
  assign \g322293/_3_  = ~n74355 ;
  assign \g322437/_0_  = ~n74380 ;
  assign \g322537/_3_  = ~n74404 ;
  assign \g322584/_0_  = ~n74436 ;
  assign \g322830/_0_  = ~n74466 ;
  assign \g322871/_0_  = ~n74498 ;
  assign \g322882/_0_  = ~n74530 ;
  assign \g322933/_0_  = ~n74555 ;
  assign \g323004/_0_  = ~n74587 ;
  assign \g323104/_0_  = ~n74609 ;
  assign \g323125/_0_  = ~n74646 ;
  assign \g323138/_3_  = ~n74675 ;
  assign \g323273/_0_  = ~n74706 ;
  assign \u0_desOut_reg[0]/_05_  = ~n74747 ;
  assign \u0_desOut_reg[12]/_05_  = ~n74840 ;
  assign \u0_desOut_reg[14]/_05_  = ~n74879 ;
  assign \u0_desOut_reg[18]/_05_  = ~n74966 ;
  assign \u0_desOut_reg[20]/_05_  = ~n75006 ;
  assign \u0_desOut_reg[24]/_05_  = ~n75039 ;
  assign \u0_desOut_reg[26]/_05_  = ~n75074 ;
  assign \u0_desOut_reg[28]/_05_  = n75151 ;
  assign \u0_desOut_reg[2]/_05_  = ~n75176 ;
  assign \u0_desOut_reg[30]/_05_  = ~n75210 ;
  assign \u0_desOut_reg[32]/_05_  = ~n75239 ;
  assign \u0_desOut_reg[34]/_05_  = ~n75273 ;
  assign \u0_desOut_reg[36]/_05_  = ~n75304 ;
  assign \u0_desOut_reg[42]/_05_  = ~n75346 ;
  assign \u0_desOut_reg[44]/_05_  = ~n75387 ;
  assign \u0_desOut_reg[46]/_05_  = ~n75413 ;
  assign \u0_desOut_reg[48]/_05_  = ~n75446 ;
  assign \u0_desOut_reg[54]/_05_  = ~n75480 ;
  assign \u0_desOut_reg[56]/_05_  = ~n75511 ;
  assign \u0_desOut_reg[62]/_05_  = ~n75535 ;
  assign \u0_desOut_reg[6]/_05_  = ~n75566 ;
  assign \u0_desOut_reg[8]/_05_  = ~n75595 ;
  assign \u1_desOut_reg[0]/_05_  = ~n75686 ;
  assign \u1_desOut_reg[12]/_05_  = ~n75779 ;
  assign \u1_desOut_reg[14]/_05_  = ~n75820 ;
  assign \u1_desOut_reg[16]/_05_  = ~n75861 ;
  assign \u1_desOut_reg[18]/_05_  = ~n75950 ;
  assign \u1_desOut_reg[20]/_05_  = ~n75988 ;
  assign \u1_desOut_reg[22]/_05_  = ~n76024 ;
  assign \u1_desOut_reg[24]/_05_  = ~n76054 ;
  assign \u1_desOut_reg[26]/_05_  = ~n76088 ;
  assign \u1_desOut_reg[28]/_05_  = n76167 ;
  assign \u1_desOut_reg[2]/_05_  = ~n76199 ;
  assign \u1_desOut_reg[30]/_05_  = ~n76231 ;
  assign \u1_desOut_reg[32]/_05_  = ~n76260 ;
  assign \u1_desOut_reg[34]/_05_  = ~n76292 ;
  assign \u1_desOut_reg[36]/_05_  = ~n76321 ;
  assign \u1_desOut_reg[38]/_05_  = ~n76351 ;
  assign \u1_desOut_reg[42]/_05_  = ~n76394 ;
  assign \u1_desOut_reg[44]/_05_  = ~n76432 ;
  assign \u1_desOut_reg[46]/_05_  = ~n76467 ;
  assign \u1_desOut_reg[48]/_05_  = ~n76501 ;
  assign \u1_desOut_reg[4]/_05_  = ~n76525 ;
  assign \u1_desOut_reg[54]/_05_  = ~n76554 ;
  assign \u1_desOut_reg[56]/_05_  = ~n76585 ;
  assign \u1_desOut_reg[58]/_05_  = ~n76618 ;
  assign \u1_desOut_reg[60]/_05_  = ~n76648 ;
  assign \u1_desOut_reg[62]/_05_  = ~n76673 ;
  assign \u1_desOut_reg[6]/_05_  = ~n76705 ;
  assign \u1_desOut_reg[8]/_05_  = ~n76736 ;
  assign \u2_desOut_reg[0]/_05_  = ~n76824 ;
  assign \u2_desOut_reg[10]/_05_  = ~n76906 ;
  assign \u2_desOut_reg[12]/_05_  = ~n76999 ;
  assign \u2_desOut_reg[14]/_05_  = ~n77045 ;
  assign \u2_desOut_reg[16]/_05_  = ~n77142 ;
  assign \u2_desOut_reg[18]/_05_  = ~n77226 ;
  assign \u2_desOut_reg[20]/_05_  = ~n77267 ;
  assign \u2_desOut_reg[22]/_05_  = n77302 ;
  assign \u2_desOut_reg[24]/_05_  = ~n77332 ;
  assign \u2_desOut_reg[26]/_05_  = ~n77368 ;
  assign \u2_desOut_reg[28]/_05_  = n77451 ;
  assign \u2_desOut_reg[2]/_05_  = ~n77537 ;
  assign \u2_desOut_reg[30]/_05_  = ~n77570 ;
  assign \u2_desOut_reg[32]/_05_  = ~n77601 ;
  assign \u2_desOut_reg[34]/_05_  = ~n77639 ;
  assign \u2_desOut_reg[36]/_05_  = ~n77669 ;
  assign \u2_desOut_reg[38]/_05_  = ~n77698 ;
  assign \u2_desOut_reg[40]/_05_  = ~n77784 ;
  assign \u2_desOut_reg[42]/_05_  = ~n77827 ;
  assign \u2_desOut_reg[44]/_05_  = ~n77868 ;
  assign \u2_desOut_reg[46]/_05_  = ~n77903 ;
  assign \u2_desOut_reg[48]/_05_  = ~n77947 ;
  assign \u2_desOut_reg[4]/_05_  = ~n77975 ;
  assign \u2_desOut_reg[50]/_05_  = ~n78007 ;
  assign \u2_desOut_reg[52]/_05_  = ~n78033 ;
  assign \u2_desOut_reg[54]/_05_  = ~n78058 ;
  assign \u2_desOut_reg[56]/_05_  = ~n78090 ;
  assign \u2_desOut_reg[58]/_05_  = ~n78119 ;
  assign \u2_desOut_reg[60]/_05_  = ~n78149 ;
  assign \u2_desOut_reg[62]/_05_  = ~n78174 ;
  assign \u2_desOut_reg[6]/_05_  = ~n78204 ;
  assign \u2_desOut_reg[8]/_05_  = ~n78238 ;
endmodule
