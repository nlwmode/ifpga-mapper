module top( \a[0]  , \a[1]  , \a[2]  , \a[3]  , \a[4]  , \a[5]  , \a[6]  , \a[7]  , \a[8]  , \a[9]  , \a[10]  , \a[11]  , \a[12]  , \a[13]  , \a[14]  , \a[15]  , \a[16]  , \a[17]  , \a[18]  , \a[19]  , \a[20]  , \a[21]  , \a[22]  , \a[23]  , \a[24]  , \a[25]  , \a[26]  , \a[27]  , \a[28]  , \a[29]  , \a[30]  , \a[31]  , \a[32]  , \a[33]  , \a[34]  , \a[35]  , \a[36]  , \a[37]  , \a[38]  , \a[39]  , \a[40]  , \a[41]  , \a[42]  , \a[43]  , \a[44]  , \a[45]  , \a[46]  , \a[47]  , \a[48]  , \a[49]  , \a[50]  , \a[51]  , \a[52]  , \a[53]  , \a[54]  , \a[55]  , \a[56]  , \a[57]  , \a[58]  , \a[59]  , \a[60]  , \a[61]  , \a[62]  , \a[63]  , \a[64]  , \a[65]  , \a[66]  , \a[67]  , \a[68]  , \a[69]  , \a[70]  , \a[71]  , \a[72]  , \a[73]  , \a[74]  , \a[75]  , \a[76]  , \a[77]  , \a[78]  , \a[79]  , \a[80]  , \a[81]  , \a[82]  , \a[83]  , \a[84]  , \a[85]  , \a[86]  , \a[87]  , \a[88]  , \a[89]  , \a[90]  , \a[91]  , \a[92]  , \a[93]  , \a[94]  , \a[95]  , \a[96]  , \a[97]  , \a[98]  , \a[99]  , \a[100]  , \a[101]  , \a[102]  , \a[103]  , \a[104]  , \a[105]  , \a[106]  , \a[107]  , \a[108]  , \a[109]  , \a[110]  , \a[111]  , \a[112]  , \a[113]  , \a[114]  , \a[115]  , \a[116]  , \a[117]  , \a[118]  , \a[119]  , \a[120]  , \a[121]  , \a[122]  , \a[123]  , \a[124]  , \a[125]  , \a[126]  , \a[127]  , \b[0]  , \b[1]  , \b[2]  , \b[3]  , \b[4]  , \b[5]  , \b[6]  , \b[7]  , \b[8]  , \b[9]  , \b[10]  , \b[11]  , \b[12]  , \b[13]  , \b[14]  , \b[15]  , \b[16]  , \b[17]  , \b[18]  , \b[19]  , \b[20]  , \b[21]  , \b[22]  , \b[23]  , \b[24]  , \b[25]  , \b[26]  , \b[27]  , \b[28]  , \b[29]  , \b[30]  , \b[31]  , \b[32]  , \b[33]  , \b[34]  , \b[35]  , \b[36]  , \b[37]  , \b[38]  , \b[39]  , \b[40]  , \b[41]  , \b[42]  , \b[43]  , \b[44]  , \b[45]  , \b[46]  , \b[47]  , \b[48]  , \b[49]  , \b[50]  , \b[51]  , \b[52]  , \b[53]  , \b[54]  , \b[55]  , \b[56]  , \b[57]  , \b[58]  , \b[59]  , \b[60]  , \b[61]  , \b[62]  , \b[63]  , \b[64]  , \b[65]  , \b[66]  , \b[67]  , \b[68]  , \b[69]  , \b[70]  , \b[71]  , \b[72]  , \b[73]  , \b[74]  , \b[75]  , \b[76]  , \b[77]  , \b[78]  , \b[79]  , \b[80]  , \b[81]  , \b[82]  , \b[83]  , \b[84]  , \b[85]  , \b[86]  , \b[87]  , \b[88]  , \b[89]  , \b[90]  , \b[91]  , \b[92]  , \b[93]  , \b[94]  , \b[95]  , \b[96]  , \b[97]  , \b[98]  , \b[99]  , \b[100]  , \b[101]  , \b[102]  , \b[103]  , \b[104]  , \b[105]  , \b[106]  , \b[107]  , \b[108]  , \b[109]  , \b[110]  , \b[111]  , \b[112]  , \b[113]  , \b[114]  , \b[115]  , \b[116]  , \b[117]  , \b[118]  , \b[119]  , \b[120]  , \b[121]  , \b[122]  , \b[123]  , \b[124]  , \b[125]  , \b[126]  , \b[127]  , \f[0]  , \f[1]  , \f[2]  , \f[3]  , \f[4]  , \f[5]  , \f[6]  , \f[7]  , \f[8]  , \f[9]  , \f[10]  , \f[11]  , \f[12]  , \f[13]  , \f[14]  , \f[15]  , \f[16]  , \f[17]  , \f[18]  , \f[19]  , \f[20]  , \f[21]  , \f[22]  , \f[23]  , \f[24]  , \f[25]  , \f[26]  , \f[27]  , \f[28]  , \f[29]  , \f[30]  , \f[31]  , \f[32]  , \f[33]  , \f[34]  , \f[35]  , \f[36]  , \f[37]  , \f[38]  , \f[39]  , \f[40]  , \f[41]  , \f[42]  , \f[43]  , \f[44]  , \f[45]  , \f[46]  , \f[47]  , \f[48]  , \f[49]  , \f[50]  , \f[51]  , \f[52]  , \f[53]  , \f[54]  , \f[55]  , \f[56]  , \f[57]  , \f[58]  , \f[59]  , \f[60]  , \f[61]  , \f[62]  , \f[63]  , \f[64]  , \f[65]  , \f[66]  , \f[67]  , \f[68]  , \f[69]  , \f[70]  , \f[71]  , \f[72]  , \f[73]  , \f[74]  , \f[75]  , \f[76]  , \f[77]  , \f[78]  , \f[79]  , \f[80]  , \f[81]  , \f[82]  , \f[83]  , \f[84]  , \f[85]  , \f[86]  , \f[87]  , \f[88]  , \f[89]  , \f[90]  , \f[91]  , \f[92]  , \f[93]  , \f[94]  , \f[95]  , \f[96]  , \f[97]  , \f[98]  , \f[99]  , \f[100]  , \f[101]  , \f[102]  , \f[103]  , \f[104]  , \f[105]  , \f[106]  , \f[107]  , \f[108]  , \f[109]  , \f[110]  , \f[111]  , \f[112]  , \f[113]  , \f[114]  , \f[115]  , \f[116]  , \f[117]  , \f[118]  , \f[119]  , \f[120]  , \f[121]  , \f[122]  , \f[123]  , \f[124]  , \f[125]  , \f[126]  , \f[127]  , cOut );
  input \a[0]  ;
  input \a[1]  ;
  input \a[2]  ;
  input \a[3]  ;
  input \a[4]  ;
  input \a[5]  ;
  input \a[6]  ;
  input \a[7]  ;
  input \a[8]  ;
  input \a[9]  ;
  input \a[10]  ;
  input \a[11]  ;
  input \a[12]  ;
  input \a[13]  ;
  input \a[14]  ;
  input \a[15]  ;
  input \a[16]  ;
  input \a[17]  ;
  input \a[18]  ;
  input \a[19]  ;
  input \a[20]  ;
  input \a[21]  ;
  input \a[22]  ;
  input \a[23]  ;
  input \a[24]  ;
  input \a[25]  ;
  input \a[26]  ;
  input \a[27]  ;
  input \a[28]  ;
  input \a[29]  ;
  input \a[30]  ;
  input \a[31]  ;
  input \a[32]  ;
  input \a[33]  ;
  input \a[34]  ;
  input \a[35]  ;
  input \a[36]  ;
  input \a[37]  ;
  input \a[38]  ;
  input \a[39]  ;
  input \a[40]  ;
  input \a[41]  ;
  input \a[42]  ;
  input \a[43]  ;
  input \a[44]  ;
  input \a[45]  ;
  input \a[46]  ;
  input \a[47]  ;
  input \a[48]  ;
  input \a[49]  ;
  input \a[50]  ;
  input \a[51]  ;
  input \a[52]  ;
  input \a[53]  ;
  input \a[54]  ;
  input \a[55]  ;
  input \a[56]  ;
  input \a[57]  ;
  input \a[58]  ;
  input \a[59]  ;
  input \a[60]  ;
  input \a[61]  ;
  input \a[62]  ;
  input \a[63]  ;
  input \a[64]  ;
  input \a[65]  ;
  input \a[66]  ;
  input \a[67]  ;
  input \a[68]  ;
  input \a[69]  ;
  input \a[70]  ;
  input \a[71]  ;
  input \a[72]  ;
  input \a[73]  ;
  input \a[74]  ;
  input \a[75]  ;
  input \a[76]  ;
  input \a[77]  ;
  input \a[78]  ;
  input \a[79]  ;
  input \a[80]  ;
  input \a[81]  ;
  input \a[82]  ;
  input \a[83]  ;
  input \a[84]  ;
  input \a[85]  ;
  input \a[86]  ;
  input \a[87]  ;
  input \a[88]  ;
  input \a[89]  ;
  input \a[90]  ;
  input \a[91]  ;
  input \a[92]  ;
  input \a[93]  ;
  input \a[94]  ;
  input \a[95]  ;
  input \a[96]  ;
  input \a[97]  ;
  input \a[98]  ;
  input \a[99]  ;
  input \a[100]  ;
  input \a[101]  ;
  input \a[102]  ;
  input \a[103]  ;
  input \a[104]  ;
  input \a[105]  ;
  input \a[106]  ;
  input \a[107]  ;
  input \a[108]  ;
  input \a[109]  ;
  input \a[110]  ;
  input \a[111]  ;
  input \a[112]  ;
  input \a[113]  ;
  input \a[114]  ;
  input \a[115]  ;
  input \a[116]  ;
  input \a[117]  ;
  input \a[118]  ;
  input \a[119]  ;
  input \a[120]  ;
  input \a[121]  ;
  input \a[122]  ;
  input \a[123]  ;
  input \a[124]  ;
  input \a[125]  ;
  input \a[126]  ;
  input \a[127]  ;
  input \b[0]  ;
  input \b[1]  ;
  input \b[2]  ;
  input \b[3]  ;
  input \b[4]  ;
  input \b[5]  ;
  input \b[6]  ;
  input \b[7]  ;
  input \b[8]  ;
  input \b[9]  ;
  input \b[10]  ;
  input \b[11]  ;
  input \b[12]  ;
  input \b[13]  ;
  input \b[14]  ;
  input \b[15]  ;
  input \b[16]  ;
  input \b[17]  ;
  input \b[18]  ;
  input \b[19]  ;
  input \b[20]  ;
  input \b[21]  ;
  input \b[22]  ;
  input \b[23]  ;
  input \b[24]  ;
  input \b[25]  ;
  input \b[26]  ;
  input \b[27]  ;
  input \b[28]  ;
  input \b[29]  ;
  input \b[30]  ;
  input \b[31]  ;
  input \b[32]  ;
  input \b[33]  ;
  input \b[34]  ;
  input \b[35]  ;
  input \b[36]  ;
  input \b[37]  ;
  input \b[38]  ;
  input \b[39]  ;
  input \b[40]  ;
  input \b[41]  ;
  input \b[42]  ;
  input \b[43]  ;
  input \b[44]  ;
  input \b[45]  ;
  input \b[46]  ;
  input \b[47]  ;
  input \b[48]  ;
  input \b[49]  ;
  input \b[50]  ;
  input \b[51]  ;
  input \b[52]  ;
  input \b[53]  ;
  input \b[54]  ;
  input \b[55]  ;
  input \b[56]  ;
  input \b[57]  ;
  input \b[58]  ;
  input \b[59]  ;
  input \b[60]  ;
  input \b[61]  ;
  input \b[62]  ;
  input \b[63]  ;
  input \b[64]  ;
  input \b[65]  ;
  input \b[66]  ;
  input \b[67]  ;
  input \b[68]  ;
  input \b[69]  ;
  input \b[70]  ;
  input \b[71]  ;
  input \b[72]  ;
  input \b[73]  ;
  input \b[74]  ;
  input \b[75]  ;
  input \b[76]  ;
  input \b[77]  ;
  input \b[78]  ;
  input \b[79]  ;
  input \b[80]  ;
  input \b[81]  ;
  input \b[82]  ;
  input \b[83]  ;
  input \b[84]  ;
  input \b[85]  ;
  input \b[86]  ;
  input \b[87]  ;
  input \b[88]  ;
  input \b[89]  ;
  input \b[90]  ;
  input \b[91]  ;
  input \b[92]  ;
  input \b[93]  ;
  input \b[94]  ;
  input \b[95]  ;
  input \b[96]  ;
  input \b[97]  ;
  input \b[98]  ;
  input \b[99]  ;
  input \b[100]  ;
  input \b[101]  ;
  input \b[102]  ;
  input \b[103]  ;
  input \b[104]  ;
  input \b[105]  ;
  input \b[106]  ;
  input \b[107]  ;
  input \b[108]  ;
  input \b[109]  ;
  input \b[110]  ;
  input \b[111]  ;
  input \b[112]  ;
  input \b[113]  ;
  input \b[114]  ;
  input \b[115]  ;
  input \b[116]  ;
  input \b[117]  ;
  input \b[118]  ;
  input \b[119]  ;
  input \b[120]  ;
  input \b[121]  ;
  input \b[122]  ;
  input \b[123]  ;
  input \b[124]  ;
  input \b[125]  ;
  input \b[126]  ;
  input \b[127]  ;
  output \f[0]  ;
  output \f[1]  ;
  output \f[2]  ;
  output \f[3]  ;
  output \f[4]  ;
  output \f[5]  ;
  output \f[6]  ;
  output \f[7]  ;
  output \f[8]  ;
  output \f[9]  ;
  output \f[10]  ;
  output \f[11]  ;
  output \f[12]  ;
  output \f[13]  ;
  output \f[14]  ;
  output \f[15]  ;
  output \f[16]  ;
  output \f[17]  ;
  output \f[18]  ;
  output \f[19]  ;
  output \f[20]  ;
  output \f[21]  ;
  output \f[22]  ;
  output \f[23]  ;
  output \f[24]  ;
  output \f[25]  ;
  output \f[26]  ;
  output \f[27]  ;
  output \f[28]  ;
  output \f[29]  ;
  output \f[30]  ;
  output \f[31]  ;
  output \f[32]  ;
  output \f[33]  ;
  output \f[34]  ;
  output \f[35]  ;
  output \f[36]  ;
  output \f[37]  ;
  output \f[38]  ;
  output \f[39]  ;
  output \f[40]  ;
  output \f[41]  ;
  output \f[42]  ;
  output \f[43]  ;
  output \f[44]  ;
  output \f[45]  ;
  output \f[46]  ;
  output \f[47]  ;
  output \f[48]  ;
  output \f[49]  ;
  output \f[50]  ;
  output \f[51]  ;
  output \f[52]  ;
  output \f[53]  ;
  output \f[54]  ;
  output \f[55]  ;
  output \f[56]  ;
  output \f[57]  ;
  output \f[58]  ;
  output \f[59]  ;
  output \f[60]  ;
  output \f[61]  ;
  output \f[62]  ;
  output \f[63]  ;
  output \f[64]  ;
  output \f[65]  ;
  output \f[66]  ;
  output \f[67]  ;
  output \f[68]  ;
  output \f[69]  ;
  output \f[70]  ;
  output \f[71]  ;
  output \f[72]  ;
  output \f[73]  ;
  output \f[74]  ;
  output \f[75]  ;
  output \f[76]  ;
  output \f[77]  ;
  output \f[78]  ;
  output \f[79]  ;
  output \f[80]  ;
  output \f[81]  ;
  output \f[82]  ;
  output \f[83]  ;
  output \f[84]  ;
  output \f[85]  ;
  output \f[86]  ;
  output \f[87]  ;
  output \f[88]  ;
  output \f[89]  ;
  output \f[90]  ;
  output \f[91]  ;
  output \f[92]  ;
  output \f[93]  ;
  output \f[94]  ;
  output \f[95]  ;
  output \f[96]  ;
  output \f[97]  ;
  output \f[98]  ;
  output \f[99]  ;
  output \f[100]  ;
  output \f[101]  ;
  output \f[102]  ;
  output \f[103]  ;
  output \f[104]  ;
  output \f[105]  ;
  output \f[106]  ;
  output \f[107]  ;
  output \f[108]  ;
  output \f[109]  ;
  output \f[110]  ;
  output \f[111]  ;
  output \f[112]  ;
  output \f[113]  ;
  output \f[114]  ;
  output \f[115]  ;
  output \f[116]  ;
  output \f[117]  ;
  output \f[118]  ;
  output \f[119]  ;
  output \f[120]  ;
  output \f[121]  ;
  output \f[122]  ;
  output \f[123]  ;
  output \f[124]  ;
  output \f[125]  ;
  output \f[126]  ;
  output \f[127]  ;
  output cOut ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 ;
  assign n257 = \a[0]  & ~\b[0]  ;
  assign n258 = ~\a[0]  & \b[0]  ;
  assign n259 = ~n257 & ~n258 ;
  assign n260 = \a[0]  & \b[0]  ;
  assign n261 = ~\a[1]  & ~\b[1]  ;
  assign n262 = \a[1]  & \b[1]  ;
  assign n263 = ~n261 & ~n262 ;
  assign n264 = n260 & ~n263 ;
  assign n265 = ~n260 & n263 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = n260 & ~n261 ;
  assign n268 = ~n262 & ~n267 ;
  assign n269 = ~\a[2]  & ~\b[2]  ;
  assign n270 = \a[2]  & \b[2]  ;
  assign n271 = ~n269 & ~n270 ;
  assign n272 = n268 & ~n271 ;
  assign n273 = ~n268 & n271 ;
  assign n274 = ~n272 & ~n273 ;
  assign n275 = ~n268 & ~n269 ;
  assign n276 = ~n270 & ~n275 ;
  assign n277 = ~\a[3]  & ~\b[3]  ;
  assign n278 = \a[3]  & \b[3]  ;
  assign n279 = ~n277 & ~n278 ;
  assign n280 = n276 & ~n279 ;
  assign n281 = ~n276 & n279 ;
  assign n282 = ~n280 & ~n281 ;
  assign n283 = ~n276 & ~n277 ;
  assign n284 = ~n278 & ~n283 ;
  assign n285 = ~\a[4]  & ~\b[4]  ;
  assign n286 = \a[4]  & \b[4]  ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = n284 & ~n287 ;
  assign n289 = ~n284 & n287 ;
  assign n290 = ~n288 & ~n289 ;
  assign n291 = ~n284 & ~n285 ;
  assign n292 = ~n286 & ~n291 ;
  assign n293 = ~\a[5]  & ~\b[5]  ;
  assign n294 = \a[5]  & \b[5]  ;
  assign n295 = ~n293 & ~n294 ;
  assign n296 = n292 & ~n295 ;
  assign n297 = ~n292 & n295 ;
  assign n298 = ~n296 & ~n297 ;
  assign n299 = ~n292 & ~n293 ;
  assign n300 = ~n294 & ~n299 ;
  assign n301 = ~\a[6]  & ~\b[6]  ;
  assign n302 = \a[6]  & \b[6]  ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = n300 & ~n303 ;
  assign n305 = ~n300 & n303 ;
  assign n306 = ~n304 & ~n305 ;
  assign n307 = ~n300 & ~n301 ;
  assign n308 = ~n302 & ~n307 ;
  assign n309 = ~\a[7]  & ~\b[7]  ;
  assign n310 = \a[7]  & \b[7]  ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = n308 & ~n311 ;
  assign n313 = ~n308 & n311 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = ~n308 & ~n309 ;
  assign n316 = ~n310 & ~n315 ;
  assign n317 = ~\a[8]  & ~\b[8]  ;
  assign n318 = \a[8]  & \b[8]  ;
  assign n319 = ~n317 & ~n318 ;
  assign n320 = n316 & ~n319 ;
  assign n321 = ~n316 & n319 ;
  assign n322 = ~n320 & ~n321 ;
  assign n323 = ~n316 & ~n317 ;
  assign n324 = ~n318 & ~n323 ;
  assign n325 = ~\a[9]  & ~\b[9]  ;
  assign n326 = \a[9]  & \b[9]  ;
  assign n327 = ~n325 & ~n326 ;
  assign n328 = n324 & ~n327 ;
  assign n329 = ~n324 & n327 ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = ~n324 & ~n325 ;
  assign n332 = ~n326 & ~n331 ;
  assign n333 = ~\a[10]  & ~\b[10]  ;
  assign n334 = \a[10]  & \b[10]  ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = n332 & ~n335 ;
  assign n337 = ~n332 & n335 ;
  assign n338 = ~n336 & ~n337 ;
  assign n339 = ~n332 & ~n333 ;
  assign n340 = ~n334 & ~n339 ;
  assign n341 = ~\a[11]  & ~\b[11]  ;
  assign n342 = \a[11]  & \b[11]  ;
  assign n343 = ~n341 & ~n342 ;
  assign n344 = n340 & ~n343 ;
  assign n345 = ~n340 & n343 ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = ~n340 & ~n341 ;
  assign n348 = ~n342 & ~n347 ;
  assign n349 = ~\a[12]  & ~\b[12]  ;
  assign n350 = \a[12]  & \b[12]  ;
  assign n351 = ~n349 & ~n350 ;
  assign n352 = n348 & ~n351 ;
  assign n353 = ~n348 & n351 ;
  assign n354 = ~n352 & ~n353 ;
  assign n355 = ~n348 & ~n349 ;
  assign n356 = ~n350 & ~n355 ;
  assign n357 = ~\a[13]  & ~\b[13]  ;
  assign n358 = \a[13]  & \b[13]  ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = n356 & ~n359 ;
  assign n361 = ~n356 & n359 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = ~n356 & ~n357 ;
  assign n364 = ~n358 & ~n363 ;
  assign n365 = ~\a[14]  & ~\b[14]  ;
  assign n366 = \a[14]  & \b[14]  ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = n364 & ~n367 ;
  assign n369 = ~n364 & n367 ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = ~n364 & ~n365 ;
  assign n372 = ~n366 & ~n371 ;
  assign n373 = ~\a[15]  & ~\b[15]  ;
  assign n374 = \a[15]  & \b[15]  ;
  assign n375 = ~n373 & ~n374 ;
  assign n376 = n372 & ~n375 ;
  assign n377 = ~n372 & n375 ;
  assign n378 = ~n376 & ~n377 ;
  assign n379 = ~n372 & ~n373 ;
  assign n380 = ~n374 & ~n379 ;
  assign n381 = ~\a[16]  & ~\b[16]  ;
  assign n382 = \a[16]  & \b[16]  ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = n380 & ~n383 ;
  assign n385 = ~n380 & n383 ;
  assign n386 = ~n384 & ~n385 ;
  assign n387 = ~n380 & ~n381 ;
  assign n388 = ~n382 & ~n387 ;
  assign n389 = ~\a[17]  & ~\b[17]  ;
  assign n390 = \a[17]  & \b[17]  ;
  assign n391 = ~n389 & ~n390 ;
  assign n392 = n388 & ~n391 ;
  assign n393 = ~n388 & n391 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = ~n388 & ~n389 ;
  assign n396 = ~n390 & ~n395 ;
  assign n397 = ~\a[18]  & ~\b[18]  ;
  assign n398 = \a[18]  & \b[18]  ;
  assign n399 = ~n397 & ~n398 ;
  assign n400 = n396 & ~n399 ;
  assign n401 = ~n396 & n399 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = ~n396 & ~n397 ;
  assign n404 = ~n398 & ~n403 ;
  assign n405 = ~\a[19]  & ~\b[19]  ;
  assign n406 = \a[19]  & \b[19]  ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = n404 & ~n407 ;
  assign n409 = ~n404 & n407 ;
  assign n410 = ~n408 & ~n409 ;
  assign n411 = ~n404 & ~n405 ;
  assign n412 = ~n406 & ~n411 ;
  assign n413 = ~\a[20]  & ~\b[20]  ;
  assign n414 = \a[20]  & \b[20]  ;
  assign n415 = ~n413 & ~n414 ;
  assign n416 = n412 & ~n415 ;
  assign n417 = ~n412 & n415 ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = ~n412 & ~n413 ;
  assign n420 = ~n414 & ~n419 ;
  assign n421 = ~\a[21]  & ~\b[21]  ;
  assign n422 = \a[21]  & \b[21]  ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = n420 & ~n423 ;
  assign n425 = ~n420 & n423 ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = ~n420 & ~n421 ;
  assign n428 = ~n422 & ~n427 ;
  assign n429 = ~\a[22]  & ~\b[22]  ;
  assign n430 = \a[22]  & \b[22]  ;
  assign n431 = ~n429 & ~n430 ;
  assign n432 = n428 & ~n431 ;
  assign n433 = ~n428 & n431 ;
  assign n434 = ~n432 & ~n433 ;
  assign n435 = ~n428 & ~n429 ;
  assign n436 = ~n430 & ~n435 ;
  assign n437 = ~\a[23]  & ~\b[23]  ;
  assign n438 = \a[23]  & \b[23]  ;
  assign n439 = ~n437 & ~n438 ;
  assign n440 = n436 & ~n439 ;
  assign n441 = ~n436 & n439 ;
  assign n442 = ~n440 & ~n441 ;
  assign n443 = ~n436 & ~n437 ;
  assign n444 = ~n438 & ~n443 ;
  assign n445 = ~\a[24]  & ~\b[24]  ;
  assign n446 = \a[24]  & \b[24]  ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = n444 & ~n447 ;
  assign n449 = ~n444 & n447 ;
  assign n450 = ~n448 & ~n449 ;
  assign n451 = ~n444 & ~n445 ;
  assign n452 = ~n446 & ~n451 ;
  assign n453 = ~\a[25]  & ~\b[25]  ;
  assign n454 = \a[25]  & \b[25]  ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = n452 & ~n455 ;
  assign n457 = ~n452 & n455 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = ~n452 & ~n453 ;
  assign n460 = ~n454 & ~n459 ;
  assign n461 = ~\a[26]  & ~\b[26]  ;
  assign n462 = \a[26]  & \b[26]  ;
  assign n463 = ~n461 & ~n462 ;
  assign n464 = n460 & ~n463 ;
  assign n465 = ~n460 & n463 ;
  assign n466 = ~n464 & ~n465 ;
  assign n467 = ~n460 & ~n461 ;
  assign n468 = ~n462 & ~n467 ;
  assign n469 = ~\a[27]  & ~\b[27]  ;
  assign n470 = \a[27]  & \b[27]  ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = n468 & ~n471 ;
  assign n473 = ~n468 & n471 ;
  assign n474 = ~n472 & ~n473 ;
  assign n475 = ~n468 & ~n469 ;
  assign n476 = ~n470 & ~n475 ;
  assign n477 = ~\a[28]  & ~\b[28]  ;
  assign n478 = \a[28]  & \b[28]  ;
  assign n479 = ~n477 & ~n478 ;
  assign n480 = n476 & ~n479 ;
  assign n481 = ~n476 & n479 ;
  assign n482 = ~n480 & ~n481 ;
  assign n483 = ~n476 & ~n477 ;
  assign n484 = ~n478 & ~n483 ;
  assign n485 = ~\a[29]  & ~\b[29]  ;
  assign n486 = \a[29]  & \b[29]  ;
  assign n487 = ~n485 & ~n486 ;
  assign n488 = n484 & ~n487 ;
  assign n489 = ~n484 & n487 ;
  assign n490 = ~n488 & ~n489 ;
  assign n491 = ~n484 & ~n485 ;
  assign n492 = ~n486 & ~n491 ;
  assign n493 = ~\a[30]  & ~\b[30]  ;
  assign n494 = \a[30]  & \b[30]  ;
  assign n495 = ~n493 & ~n494 ;
  assign n496 = n492 & ~n495 ;
  assign n497 = ~n492 & n495 ;
  assign n498 = ~n496 & ~n497 ;
  assign n499 = ~n492 & ~n493 ;
  assign n500 = ~n494 & ~n499 ;
  assign n501 = ~\a[31]  & ~\b[31]  ;
  assign n502 = \a[31]  & \b[31]  ;
  assign n503 = ~n501 & ~n502 ;
  assign n504 = n500 & ~n503 ;
  assign n505 = ~n500 & n503 ;
  assign n506 = ~n504 & ~n505 ;
  assign n507 = ~n500 & ~n501 ;
  assign n508 = ~n502 & ~n507 ;
  assign n509 = ~\a[32]  & ~\b[32]  ;
  assign n510 = \a[32]  & \b[32]  ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = n508 & ~n511 ;
  assign n513 = ~n508 & n511 ;
  assign n514 = ~n512 & ~n513 ;
  assign n515 = ~n508 & ~n509 ;
  assign n516 = ~n510 & ~n515 ;
  assign n517 = ~\a[33]  & ~\b[33]  ;
  assign n518 = \a[33]  & \b[33]  ;
  assign n519 = ~n517 & ~n518 ;
  assign n520 = n516 & ~n519 ;
  assign n521 = ~n516 & n519 ;
  assign n522 = ~n520 & ~n521 ;
  assign n523 = ~n516 & ~n517 ;
  assign n524 = ~n518 & ~n523 ;
  assign n525 = ~\a[34]  & ~\b[34]  ;
  assign n526 = \a[34]  & \b[34]  ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = n524 & ~n527 ;
  assign n529 = ~n524 & n527 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = ~n524 & ~n525 ;
  assign n532 = ~n526 & ~n531 ;
  assign n533 = ~\a[35]  & ~\b[35]  ;
  assign n534 = \a[35]  & \b[35]  ;
  assign n535 = ~n533 & ~n534 ;
  assign n536 = n532 & ~n535 ;
  assign n537 = ~n532 & n535 ;
  assign n538 = ~n536 & ~n537 ;
  assign n539 = ~n532 & ~n533 ;
  assign n540 = ~n534 & ~n539 ;
  assign n541 = ~\a[36]  & ~\b[36]  ;
  assign n542 = \a[36]  & \b[36]  ;
  assign n543 = ~n541 & ~n542 ;
  assign n544 = n540 & ~n543 ;
  assign n545 = ~n540 & n543 ;
  assign n546 = ~n544 & ~n545 ;
  assign n547 = ~n540 & ~n541 ;
  assign n548 = ~n542 & ~n547 ;
  assign n549 = ~\a[37]  & ~\b[37]  ;
  assign n550 = \a[37]  & \b[37]  ;
  assign n551 = ~n549 & ~n550 ;
  assign n552 = n548 & ~n551 ;
  assign n553 = ~n548 & n551 ;
  assign n554 = ~n552 & ~n553 ;
  assign n555 = ~n548 & ~n549 ;
  assign n556 = ~n550 & ~n555 ;
  assign n557 = ~\a[38]  & ~\b[38]  ;
  assign n558 = \a[38]  & \b[38]  ;
  assign n559 = ~n557 & ~n558 ;
  assign n560 = n556 & ~n559 ;
  assign n561 = ~n556 & n559 ;
  assign n562 = ~n560 & ~n561 ;
  assign n563 = ~n556 & ~n557 ;
  assign n564 = ~n558 & ~n563 ;
  assign n565 = ~\a[39]  & ~\b[39]  ;
  assign n566 = \a[39]  & \b[39]  ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = n564 & ~n567 ;
  assign n569 = ~n564 & n567 ;
  assign n570 = ~n568 & ~n569 ;
  assign n571 = ~n564 & ~n565 ;
  assign n572 = ~n566 & ~n571 ;
  assign n573 = ~\a[40]  & ~\b[40]  ;
  assign n574 = \a[40]  & \b[40]  ;
  assign n575 = ~n573 & ~n574 ;
  assign n576 = n572 & ~n575 ;
  assign n577 = ~n572 & n575 ;
  assign n578 = ~n576 & ~n577 ;
  assign n579 = ~n572 & ~n573 ;
  assign n580 = ~n574 & ~n579 ;
  assign n581 = ~\a[41]  & ~\b[41]  ;
  assign n582 = \a[41]  & \b[41]  ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = n580 & ~n583 ;
  assign n585 = ~n580 & n583 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = ~n580 & ~n581 ;
  assign n588 = ~n582 & ~n587 ;
  assign n589 = ~\a[42]  & ~\b[42]  ;
  assign n590 = \a[42]  & \b[42]  ;
  assign n591 = ~n589 & ~n590 ;
  assign n592 = n588 & ~n591 ;
  assign n593 = ~n588 & n591 ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = ~n588 & ~n589 ;
  assign n596 = ~n590 & ~n595 ;
  assign n597 = ~\a[43]  & ~\b[43]  ;
  assign n598 = \a[43]  & \b[43]  ;
  assign n599 = ~n597 & ~n598 ;
  assign n600 = n596 & ~n599 ;
  assign n601 = ~n596 & n599 ;
  assign n602 = ~n600 & ~n601 ;
  assign n603 = ~n596 & ~n597 ;
  assign n604 = ~n598 & ~n603 ;
  assign n605 = ~\a[44]  & ~\b[44]  ;
  assign n606 = \a[44]  & \b[44]  ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = n604 & ~n607 ;
  assign n609 = ~n604 & n607 ;
  assign n610 = ~n608 & ~n609 ;
  assign n611 = ~n604 & ~n605 ;
  assign n612 = ~n606 & ~n611 ;
  assign n613 = ~\a[45]  & ~\b[45]  ;
  assign n614 = \a[45]  & \b[45]  ;
  assign n615 = ~n613 & ~n614 ;
  assign n616 = n612 & ~n615 ;
  assign n617 = ~n612 & n615 ;
  assign n618 = ~n616 & ~n617 ;
  assign n619 = ~n612 & ~n613 ;
  assign n620 = ~n614 & ~n619 ;
  assign n621 = ~\a[46]  & ~\b[46]  ;
  assign n622 = \a[46]  & \b[46]  ;
  assign n623 = ~n621 & ~n622 ;
  assign n624 = n620 & ~n623 ;
  assign n625 = ~n620 & n623 ;
  assign n626 = ~n624 & ~n625 ;
  assign n627 = ~n620 & ~n621 ;
  assign n628 = ~n622 & ~n627 ;
  assign n629 = ~\a[47]  & ~\b[47]  ;
  assign n630 = \a[47]  & \b[47]  ;
  assign n631 = ~n629 & ~n630 ;
  assign n632 = n628 & ~n631 ;
  assign n633 = ~n628 & n631 ;
  assign n634 = ~n632 & ~n633 ;
  assign n635 = ~n628 & ~n629 ;
  assign n636 = ~n630 & ~n635 ;
  assign n637 = ~\a[48]  & ~\b[48]  ;
  assign n638 = \a[48]  & \b[48]  ;
  assign n639 = ~n637 & ~n638 ;
  assign n640 = n636 & ~n639 ;
  assign n641 = ~n636 & n639 ;
  assign n642 = ~n640 & ~n641 ;
  assign n643 = ~n636 & ~n637 ;
  assign n644 = ~n638 & ~n643 ;
  assign n645 = ~\a[49]  & ~\b[49]  ;
  assign n646 = \a[49]  & \b[49]  ;
  assign n647 = ~n645 & ~n646 ;
  assign n648 = n644 & ~n647 ;
  assign n649 = ~n644 & n647 ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = ~n644 & ~n645 ;
  assign n652 = ~n646 & ~n651 ;
  assign n653 = ~\a[50]  & ~\b[50]  ;
  assign n654 = \a[50]  & \b[50]  ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = n652 & ~n655 ;
  assign n657 = ~n652 & n655 ;
  assign n658 = ~n656 & ~n657 ;
  assign n659 = ~n652 & ~n653 ;
  assign n660 = ~n654 & ~n659 ;
  assign n661 = ~\a[51]  & ~\b[51]  ;
  assign n662 = \a[51]  & \b[51]  ;
  assign n663 = ~n661 & ~n662 ;
  assign n664 = n660 & ~n663 ;
  assign n665 = ~n660 & n663 ;
  assign n666 = ~n664 & ~n665 ;
  assign n667 = ~n660 & ~n661 ;
  assign n668 = ~n662 & ~n667 ;
  assign n669 = ~\a[52]  & ~\b[52]  ;
  assign n670 = \a[52]  & \b[52]  ;
  assign n671 = ~n669 & ~n670 ;
  assign n672 = n668 & ~n671 ;
  assign n673 = ~n668 & n671 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = ~n668 & ~n669 ;
  assign n676 = ~n670 & ~n675 ;
  assign n677 = ~\a[53]  & ~\b[53]  ;
  assign n678 = \a[53]  & \b[53]  ;
  assign n679 = ~n677 & ~n678 ;
  assign n680 = n676 & ~n679 ;
  assign n681 = ~n676 & n679 ;
  assign n682 = ~n680 & ~n681 ;
  assign n683 = ~n676 & ~n677 ;
  assign n684 = ~n678 & ~n683 ;
  assign n685 = ~\a[54]  & ~\b[54]  ;
  assign n686 = \a[54]  & \b[54]  ;
  assign n687 = ~n685 & ~n686 ;
  assign n688 = n684 & ~n687 ;
  assign n689 = ~n684 & n687 ;
  assign n690 = ~n688 & ~n689 ;
  assign n691 = ~n684 & ~n685 ;
  assign n692 = ~n686 & ~n691 ;
  assign n693 = ~\a[55]  & ~\b[55]  ;
  assign n694 = \a[55]  & \b[55]  ;
  assign n695 = ~n693 & ~n694 ;
  assign n696 = n692 & ~n695 ;
  assign n697 = ~n692 & n695 ;
  assign n698 = ~n696 & ~n697 ;
  assign n699 = ~n692 & ~n693 ;
  assign n700 = ~n694 & ~n699 ;
  assign n701 = ~\a[56]  & ~\b[56]  ;
  assign n702 = \a[56]  & \b[56]  ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = n700 & ~n703 ;
  assign n705 = ~n700 & n703 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = ~n700 & ~n701 ;
  assign n708 = ~n702 & ~n707 ;
  assign n709 = ~\a[57]  & ~\b[57]  ;
  assign n710 = \a[57]  & \b[57]  ;
  assign n711 = ~n709 & ~n710 ;
  assign n712 = n708 & ~n711 ;
  assign n713 = ~n708 & n711 ;
  assign n714 = ~n712 & ~n713 ;
  assign n715 = ~n708 & ~n709 ;
  assign n716 = ~n710 & ~n715 ;
  assign n717 = ~\a[58]  & ~\b[58]  ;
  assign n718 = \a[58]  & \b[58]  ;
  assign n719 = ~n717 & ~n718 ;
  assign n720 = n716 & ~n719 ;
  assign n721 = ~n716 & n719 ;
  assign n722 = ~n720 & ~n721 ;
  assign n723 = ~n716 & ~n717 ;
  assign n724 = ~n718 & ~n723 ;
  assign n725 = ~\a[59]  & ~\b[59]  ;
  assign n726 = \a[59]  & \b[59]  ;
  assign n727 = ~n725 & ~n726 ;
  assign n728 = n724 & ~n727 ;
  assign n729 = ~n724 & n727 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = ~n724 & ~n725 ;
  assign n732 = ~n726 & ~n731 ;
  assign n733 = ~\a[60]  & ~\b[60]  ;
  assign n734 = \a[60]  & \b[60]  ;
  assign n735 = ~n733 & ~n734 ;
  assign n736 = n732 & ~n735 ;
  assign n737 = ~n732 & n735 ;
  assign n738 = ~n736 & ~n737 ;
  assign n739 = ~n732 & ~n733 ;
  assign n740 = ~n734 & ~n739 ;
  assign n741 = ~\a[61]  & ~\b[61]  ;
  assign n742 = \a[61]  & \b[61]  ;
  assign n743 = ~n741 & ~n742 ;
  assign n744 = n740 & ~n743 ;
  assign n745 = ~n740 & n743 ;
  assign n746 = ~n744 & ~n745 ;
  assign n747 = ~n740 & ~n741 ;
  assign n748 = ~n742 & ~n747 ;
  assign n749 = ~\a[62]  & ~\b[62]  ;
  assign n750 = \a[62]  & \b[62]  ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = n748 & ~n751 ;
  assign n753 = ~n748 & n751 ;
  assign n754 = ~n752 & ~n753 ;
  assign n755 = ~n748 & ~n749 ;
  assign n756 = ~n750 & ~n755 ;
  assign n757 = ~\a[63]  & ~\b[63]  ;
  assign n758 = \a[63]  & \b[63]  ;
  assign n759 = ~n757 & ~n758 ;
  assign n760 = n756 & ~n759 ;
  assign n761 = ~n756 & n759 ;
  assign n762 = ~n760 & ~n761 ;
  assign n763 = ~n756 & ~n757 ;
  assign n764 = ~n758 & ~n763 ;
  assign n765 = ~\a[64]  & ~\b[64]  ;
  assign n766 = \a[64]  & \b[64]  ;
  assign n767 = ~n765 & ~n766 ;
  assign n768 = n764 & ~n767 ;
  assign n769 = ~n764 & n767 ;
  assign n770 = ~n768 & ~n769 ;
  assign n771 = ~n764 & ~n765 ;
  assign n772 = ~n766 & ~n771 ;
  assign n773 = ~\a[65]  & ~\b[65]  ;
  assign n774 = \a[65]  & \b[65]  ;
  assign n775 = ~n773 & ~n774 ;
  assign n776 = n772 & ~n775 ;
  assign n777 = ~n772 & n775 ;
  assign n778 = ~n776 & ~n777 ;
  assign n779 = ~n772 & ~n773 ;
  assign n780 = ~n774 & ~n779 ;
  assign n781 = ~\a[66]  & ~\b[66]  ;
  assign n782 = \a[66]  & \b[66]  ;
  assign n783 = ~n781 & ~n782 ;
  assign n784 = n780 & ~n783 ;
  assign n785 = ~n780 & n783 ;
  assign n786 = ~n784 & ~n785 ;
  assign n787 = ~n780 & ~n781 ;
  assign n788 = ~n782 & ~n787 ;
  assign n789 = ~\a[67]  & ~\b[67]  ;
  assign n790 = \a[67]  & \b[67]  ;
  assign n791 = ~n789 & ~n790 ;
  assign n792 = n788 & ~n791 ;
  assign n793 = ~n788 & n791 ;
  assign n794 = ~n792 & ~n793 ;
  assign n795 = ~n788 & ~n789 ;
  assign n796 = ~n790 & ~n795 ;
  assign n797 = ~\a[68]  & ~\b[68]  ;
  assign n798 = \a[68]  & \b[68]  ;
  assign n799 = ~n797 & ~n798 ;
  assign n800 = n796 & ~n799 ;
  assign n801 = ~n796 & n799 ;
  assign n802 = ~n800 & ~n801 ;
  assign n803 = ~n796 & ~n797 ;
  assign n804 = ~n798 & ~n803 ;
  assign n805 = ~\a[69]  & ~\b[69]  ;
  assign n806 = \a[69]  & \b[69]  ;
  assign n807 = ~n805 & ~n806 ;
  assign n808 = n804 & ~n807 ;
  assign n809 = ~n804 & n807 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = ~n804 & ~n805 ;
  assign n812 = ~n806 & ~n811 ;
  assign n813 = ~\a[70]  & ~\b[70]  ;
  assign n814 = \a[70]  & \b[70]  ;
  assign n815 = ~n813 & ~n814 ;
  assign n816 = n812 & ~n815 ;
  assign n817 = ~n812 & n815 ;
  assign n818 = ~n816 & ~n817 ;
  assign n819 = ~n812 & ~n813 ;
  assign n820 = ~n814 & ~n819 ;
  assign n821 = ~\a[71]  & ~\b[71]  ;
  assign n822 = \a[71]  & \b[71]  ;
  assign n823 = ~n821 & ~n822 ;
  assign n824 = n820 & ~n823 ;
  assign n825 = ~n820 & n823 ;
  assign n826 = ~n824 & ~n825 ;
  assign n827 = ~n820 & ~n821 ;
  assign n828 = ~n822 & ~n827 ;
  assign n829 = ~\a[72]  & ~\b[72]  ;
  assign n830 = \a[72]  & \b[72]  ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = n828 & ~n831 ;
  assign n833 = ~n828 & n831 ;
  assign n834 = ~n832 & ~n833 ;
  assign n835 = ~n828 & ~n829 ;
  assign n836 = ~n830 & ~n835 ;
  assign n837 = ~\a[73]  & ~\b[73]  ;
  assign n838 = \a[73]  & \b[73]  ;
  assign n839 = ~n837 & ~n838 ;
  assign n840 = n836 & ~n839 ;
  assign n841 = ~n836 & n839 ;
  assign n842 = ~n840 & ~n841 ;
  assign n843 = ~n836 & ~n837 ;
  assign n844 = ~n838 & ~n843 ;
  assign n845 = ~\a[74]  & ~\b[74]  ;
  assign n846 = \a[74]  & \b[74]  ;
  assign n847 = ~n845 & ~n846 ;
  assign n848 = n844 & ~n847 ;
  assign n849 = ~n844 & n847 ;
  assign n850 = ~n848 & ~n849 ;
  assign n851 = ~n844 & ~n845 ;
  assign n852 = ~n846 & ~n851 ;
  assign n853 = ~\a[75]  & ~\b[75]  ;
  assign n854 = \a[75]  & \b[75]  ;
  assign n855 = ~n853 & ~n854 ;
  assign n856 = n852 & ~n855 ;
  assign n857 = ~n852 & n855 ;
  assign n858 = ~n856 & ~n857 ;
  assign n859 = ~n852 & ~n853 ;
  assign n860 = ~n854 & ~n859 ;
  assign n861 = ~\a[76]  & ~\b[76]  ;
  assign n862 = \a[76]  & \b[76]  ;
  assign n863 = ~n861 & ~n862 ;
  assign n864 = n860 & ~n863 ;
  assign n865 = ~n860 & n863 ;
  assign n866 = ~n864 & ~n865 ;
  assign n867 = ~n860 & ~n861 ;
  assign n868 = ~n862 & ~n867 ;
  assign n869 = ~\a[77]  & ~\b[77]  ;
  assign n870 = \a[77]  & \b[77]  ;
  assign n871 = ~n869 & ~n870 ;
  assign n872 = n868 & ~n871 ;
  assign n873 = ~n868 & n871 ;
  assign n874 = ~n872 & ~n873 ;
  assign n875 = ~n868 & ~n869 ;
  assign n876 = ~n870 & ~n875 ;
  assign n877 = ~\a[78]  & ~\b[78]  ;
  assign n878 = \a[78]  & \b[78]  ;
  assign n879 = ~n877 & ~n878 ;
  assign n880 = n876 & ~n879 ;
  assign n881 = ~n876 & n879 ;
  assign n882 = ~n880 & ~n881 ;
  assign n883 = ~n876 & ~n877 ;
  assign n884 = ~n878 & ~n883 ;
  assign n885 = ~\a[79]  & ~\b[79]  ;
  assign n886 = \a[79]  & \b[79]  ;
  assign n887 = ~n885 & ~n886 ;
  assign n888 = n884 & ~n887 ;
  assign n889 = ~n884 & n887 ;
  assign n890 = ~n888 & ~n889 ;
  assign n891 = ~n884 & ~n885 ;
  assign n892 = ~n886 & ~n891 ;
  assign n893 = ~\a[80]  & ~\b[80]  ;
  assign n894 = \a[80]  & \b[80]  ;
  assign n895 = ~n893 & ~n894 ;
  assign n896 = n892 & ~n895 ;
  assign n897 = ~n892 & n895 ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = ~n892 & ~n893 ;
  assign n900 = ~n894 & ~n899 ;
  assign n901 = ~\a[81]  & ~\b[81]  ;
  assign n902 = \a[81]  & \b[81]  ;
  assign n903 = ~n901 & ~n902 ;
  assign n904 = n900 & ~n903 ;
  assign n905 = ~n900 & n903 ;
  assign n906 = ~n904 & ~n905 ;
  assign n907 = ~n900 & ~n901 ;
  assign n908 = ~n902 & ~n907 ;
  assign n909 = ~\a[82]  & ~\b[82]  ;
  assign n910 = \a[82]  & \b[82]  ;
  assign n911 = ~n909 & ~n910 ;
  assign n912 = n908 & ~n911 ;
  assign n913 = ~n908 & n911 ;
  assign n914 = ~n912 & ~n913 ;
  assign n915 = ~n908 & ~n909 ;
  assign n916 = ~n910 & ~n915 ;
  assign n917 = ~\a[83]  & ~\b[83]  ;
  assign n918 = \a[83]  & \b[83]  ;
  assign n919 = ~n917 & ~n918 ;
  assign n920 = n916 & ~n919 ;
  assign n921 = ~n916 & n919 ;
  assign n922 = ~n920 & ~n921 ;
  assign n923 = ~n916 & ~n917 ;
  assign n924 = ~n918 & ~n923 ;
  assign n925 = ~\a[84]  & ~\b[84]  ;
  assign n926 = \a[84]  & \b[84]  ;
  assign n927 = ~n925 & ~n926 ;
  assign n928 = n924 & ~n927 ;
  assign n929 = ~n924 & n927 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = ~n924 & ~n925 ;
  assign n932 = ~n926 & ~n931 ;
  assign n933 = ~\a[85]  & ~\b[85]  ;
  assign n934 = \a[85]  & \b[85]  ;
  assign n935 = ~n933 & ~n934 ;
  assign n936 = n932 & ~n935 ;
  assign n937 = ~n932 & n935 ;
  assign n938 = ~n936 & ~n937 ;
  assign n939 = ~n932 & ~n933 ;
  assign n940 = ~n934 & ~n939 ;
  assign n941 = ~\a[86]  & ~\b[86]  ;
  assign n942 = \a[86]  & \b[86]  ;
  assign n943 = ~n941 & ~n942 ;
  assign n944 = n940 & ~n943 ;
  assign n945 = ~n940 & n943 ;
  assign n946 = ~n944 & ~n945 ;
  assign n947 = ~n940 & ~n941 ;
  assign n948 = ~n942 & ~n947 ;
  assign n949 = ~\a[87]  & ~\b[87]  ;
  assign n950 = \a[87]  & \b[87]  ;
  assign n951 = ~n949 & ~n950 ;
  assign n952 = n948 & ~n951 ;
  assign n953 = ~n948 & n951 ;
  assign n954 = ~n952 & ~n953 ;
  assign n955 = ~n948 & ~n949 ;
  assign n956 = ~n950 & ~n955 ;
  assign n957 = ~\a[88]  & ~\b[88]  ;
  assign n958 = \a[88]  & \b[88]  ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = n956 & ~n959 ;
  assign n961 = ~n956 & n959 ;
  assign n962 = ~n960 & ~n961 ;
  assign n963 = ~n956 & ~n957 ;
  assign n964 = ~n958 & ~n963 ;
  assign n965 = ~\a[89]  & ~\b[89]  ;
  assign n966 = \a[89]  & \b[89]  ;
  assign n967 = ~n965 & ~n966 ;
  assign n968 = n964 & ~n967 ;
  assign n969 = ~n964 & n967 ;
  assign n970 = ~n968 & ~n969 ;
  assign n971 = ~n964 & ~n965 ;
  assign n972 = ~n966 & ~n971 ;
  assign n973 = ~\a[90]  & ~\b[90]  ;
  assign n974 = \a[90]  & \b[90]  ;
  assign n975 = ~n973 & ~n974 ;
  assign n976 = n972 & ~n975 ;
  assign n977 = ~n972 & n975 ;
  assign n978 = ~n976 & ~n977 ;
  assign n979 = ~n972 & ~n973 ;
  assign n980 = ~n974 & ~n979 ;
  assign n981 = ~\a[91]  & ~\b[91]  ;
  assign n982 = \a[91]  & \b[91]  ;
  assign n983 = ~n981 & ~n982 ;
  assign n984 = n980 & ~n983 ;
  assign n985 = ~n980 & n983 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = ~n980 & ~n981 ;
  assign n988 = ~n982 & ~n987 ;
  assign n989 = ~\a[92]  & ~\b[92]  ;
  assign n990 = \a[92]  & \b[92]  ;
  assign n991 = ~n989 & ~n990 ;
  assign n992 = n988 & ~n991 ;
  assign n993 = ~n988 & n991 ;
  assign n994 = ~n992 & ~n993 ;
  assign n995 = ~n988 & ~n989 ;
  assign n996 = ~n990 & ~n995 ;
  assign n997 = ~\a[93]  & ~\b[93]  ;
  assign n998 = \a[93]  & \b[93]  ;
  assign n999 = ~n997 & ~n998 ;
  assign n1000 = n996 & ~n999 ;
  assign n1001 = ~n996 & n999 ;
  assign n1002 = ~n1000 & ~n1001 ;
  assign n1003 = ~n996 & ~n997 ;
  assign n1004 = ~n998 & ~n1003 ;
  assign n1005 = ~\a[94]  & ~\b[94]  ;
  assign n1006 = \a[94]  & \b[94]  ;
  assign n1007 = ~n1005 & ~n1006 ;
  assign n1008 = n1004 & ~n1007 ;
  assign n1009 = ~n1004 & n1007 ;
  assign n1010 = ~n1008 & ~n1009 ;
  assign n1011 = ~n1004 & ~n1005 ;
  assign n1012 = ~n1006 & ~n1011 ;
  assign n1013 = ~\a[95]  & ~\b[95]  ;
  assign n1014 = \a[95]  & \b[95]  ;
  assign n1015 = ~n1013 & ~n1014 ;
  assign n1016 = n1012 & ~n1015 ;
  assign n1017 = ~n1012 & n1015 ;
  assign n1018 = ~n1016 & ~n1017 ;
  assign n1019 = ~n1012 & ~n1013 ;
  assign n1020 = ~n1014 & ~n1019 ;
  assign n1021 = ~\a[96]  & ~\b[96]  ;
  assign n1022 = \a[96]  & \b[96]  ;
  assign n1023 = ~n1021 & ~n1022 ;
  assign n1024 = n1020 & ~n1023 ;
  assign n1025 = ~n1020 & n1023 ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = ~n1020 & ~n1021 ;
  assign n1028 = ~n1022 & ~n1027 ;
  assign n1029 = ~\a[97]  & ~\b[97]  ;
  assign n1030 = \a[97]  & \b[97]  ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = n1028 & ~n1031 ;
  assign n1033 = ~n1028 & n1031 ;
  assign n1034 = ~n1032 & ~n1033 ;
  assign n1035 = ~n1028 & ~n1029 ;
  assign n1036 = ~n1030 & ~n1035 ;
  assign n1037 = ~\a[98]  & ~\b[98]  ;
  assign n1038 = \a[98]  & \b[98]  ;
  assign n1039 = ~n1037 & ~n1038 ;
  assign n1040 = n1036 & ~n1039 ;
  assign n1041 = ~n1036 & n1039 ;
  assign n1042 = ~n1040 & ~n1041 ;
  assign n1043 = ~n1036 & ~n1037 ;
  assign n1044 = ~n1038 & ~n1043 ;
  assign n1045 = ~\a[99]  & ~\b[99]  ;
  assign n1046 = \a[99]  & \b[99]  ;
  assign n1047 = ~n1045 & ~n1046 ;
  assign n1048 = n1044 & ~n1047 ;
  assign n1049 = ~n1044 & n1047 ;
  assign n1050 = ~n1048 & ~n1049 ;
  assign n1051 = ~n1044 & ~n1045 ;
  assign n1052 = ~n1046 & ~n1051 ;
  assign n1053 = ~\a[100]  & ~\b[100]  ;
  assign n1054 = \a[100]  & \b[100]  ;
  assign n1055 = ~n1053 & ~n1054 ;
  assign n1056 = n1052 & ~n1055 ;
  assign n1057 = ~n1052 & n1055 ;
  assign n1058 = ~n1056 & ~n1057 ;
  assign n1059 = ~n1052 & ~n1053 ;
  assign n1060 = ~n1054 & ~n1059 ;
  assign n1061 = ~\a[101]  & ~\b[101]  ;
  assign n1062 = \a[101]  & \b[101]  ;
  assign n1063 = ~n1061 & ~n1062 ;
  assign n1064 = n1060 & ~n1063 ;
  assign n1065 = ~n1060 & n1063 ;
  assign n1066 = ~n1064 & ~n1065 ;
  assign n1067 = ~n1060 & ~n1061 ;
  assign n1068 = ~n1062 & ~n1067 ;
  assign n1069 = ~\a[102]  & ~\b[102]  ;
  assign n1070 = \a[102]  & \b[102]  ;
  assign n1071 = ~n1069 & ~n1070 ;
  assign n1072 = n1068 & ~n1071 ;
  assign n1073 = ~n1068 & n1071 ;
  assign n1074 = ~n1072 & ~n1073 ;
  assign n1075 = ~n1068 & ~n1069 ;
  assign n1076 = ~n1070 & ~n1075 ;
  assign n1077 = ~\a[103]  & ~\b[103]  ;
  assign n1078 = \a[103]  & \b[103]  ;
  assign n1079 = ~n1077 & ~n1078 ;
  assign n1080 = n1076 & ~n1079 ;
  assign n1081 = ~n1076 & n1079 ;
  assign n1082 = ~n1080 & ~n1081 ;
  assign n1083 = ~n1076 & ~n1077 ;
  assign n1084 = ~n1078 & ~n1083 ;
  assign n1085 = ~\a[104]  & ~\b[104]  ;
  assign n1086 = \a[104]  & \b[104]  ;
  assign n1087 = ~n1085 & ~n1086 ;
  assign n1088 = n1084 & ~n1087 ;
  assign n1089 = ~n1084 & n1087 ;
  assign n1090 = ~n1088 & ~n1089 ;
  assign n1091 = ~n1084 & ~n1085 ;
  assign n1092 = ~n1086 & ~n1091 ;
  assign n1093 = ~\a[105]  & ~\b[105]  ;
  assign n1094 = \a[105]  & \b[105]  ;
  assign n1095 = ~n1093 & ~n1094 ;
  assign n1096 = n1092 & ~n1095 ;
  assign n1097 = ~n1092 & n1095 ;
  assign n1098 = ~n1096 & ~n1097 ;
  assign n1099 = ~n1092 & ~n1093 ;
  assign n1100 = ~n1094 & ~n1099 ;
  assign n1101 = ~\a[106]  & ~\b[106]  ;
  assign n1102 = \a[106]  & \b[106]  ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = n1100 & ~n1103 ;
  assign n1105 = ~n1100 & n1103 ;
  assign n1106 = ~n1104 & ~n1105 ;
  assign n1107 = ~n1100 & ~n1101 ;
  assign n1108 = ~n1102 & ~n1107 ;
  assign n1109 = ~\a[107]  & ~\b[107]  ;
  assign n1110 = \a[107]  & \b[107]  ;
  assign n1111 = ~n1109 & ~n1110 ;
  assign n1112 = n1108 & ~n1111 ;
  assign n1113 = ~n1108 & n1111 ;
  assign n1114 = ~n1112 & ~n1113 ;
  assign n1115 = ~n1108 & ~n1109 ;
  assign n1116 = ~n1110 & ~n1115 ;
  assign n1117 = ~\a[108]  & ~\b[108]  ;
  assign n1118 = \a[108]  & \b[108]  ;
  assign n1119 = ~n1117 & ~n1118 ;
  assign n1120 = n1116 & ~n1119 ;
  assign n1121 = ~n1116 & n1119 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = ~n1116 & ~n1117 ;
  assign n1124 = ~n1118 & ~n1123 ;
  assign n1125 = ~\a[109]  & ~\b[109]  ;
  assign n1126 = \a[109]  & \b[109]  ;
  assign n1127 = ~n1125 & ~n1126 ;
  assign n1128 = n1124 & ~n1127 ;
  assign n1129 = ~n1124 & n1127 ;
  assign n1130 = ~n1128 & ~n1129 ;
  assign n1131 = ~n1124 & ~n1125 ;
  assign n1132 = ~n1126 & ~n1131 ;
  assign n1133 = ~\a[110]  & ~\b[110]  ;
  assign n1134 = \a[110]  & \b[110]  ;
  assign n1135 = ~n1133 & ~n1134 ;
  assign n1136 = n1132 & ~n1135 ;
  assign n1137 = ~n1132 & n1135 ;
  assign n1138 = ~n1136 & ~n1137 ;
  assign n1139 = ~n1132 & ~n1133 ;
  assign n1140 = ~n1134 & ~n1139 ;
  assign n1141 = ~\a[111]  & ~\b[111]  ;
  assign n1142 = \a[111]  & \b[111]  ;
  assign n1143 = ~n1141 & ~n1142 ;
  assign n1144 = n1140 & ~n1143 ;
  assign n1145 = ~n1140 & n1143 ;
  assign n1146 = ~n1144 & ~n1145 ;
  assign n1147 = ~n1140 & ~n1141 ;
  assign n1148 = ~n1142 & ~n1147 ;
  assign n1149 = ~\a[112]  & ~\b[112]  ;
  assign n1150 = \a[112]  & \b[112]  ;
  assign n1151 = ~n1149 & ~n1150 ;
  assign n1152 = n1148 & ~n1151 ;
  assign n1153 = ~n1148 & n1151 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = ~n1148 & ~n1149 ;
  assign n1156 = ~n1150 & ~n1155 ;
  assign n1157 = ~\a[113]  & ~\b[113]  ;
  assign n1158 = \a[113]  & \b[113]  ;
  assign n1159 = ~n1157 & ~n1158 ;
  assign n1160 = n1156 & ~n1159 ;
  assign n1161 = ~n1156 & n1159 ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1163 = ~n1156 & ~n1157 ;
  assign n1164 = ~n1158 & ~n1163 ;
  assign n1165 = ~\a[114]  & ~\b[114]  ;
  assign n1166 = \a[114]  & \b[114]  ;
  assign n1167 = ~n1165 & ~n1166 ;
  assign n1168 = n1164 & ~n1167 ;
  assign n1169 = ~n1164 & n1167 ;
  assign n1170 = ~n1168 & ~n1169 ;
  assign n1171 = ~n1164 & ~n1165 ;
  assign n1172 = ~n1166 & ~n1171 ;
  assign n1173 = ~\a[115]  & ~\b[115]  ;
  assign n1174 = \a[115]  & \b[115]  ;
  assign n1175 = ~n1173 & ~n1174 ;
  assign n1176 = n1172 & ~n1175 ;
  assign n1177 = ~n1172 & n1175 ;
  assign n1178 = ~n1176 & ~n1177 ;
  assign n1179 = ~n1172 & ~n1173 ;
  assign n1180 = ~n1174 & ~n1179 ;
  assign n1181 = ~\a[116]  & ~\b[116]  ;
  assign n1182 = \a[116]  & \b[116]  ;
  assign n1183 = ~n1181 & ~n1182 ;
  assign n1184 = n1180 & ~n1183 ;
  assign n1185 = ~n1180 & n1183 ;
  assign n1186 = ~n1184 & ~n1185 ;
  assign n1187 = ~n1180 & ~n1181 ;
  assign n1188 = ~n1182 & ~n1187 ;
  assign n1189 = ~\a[117]  & ~\b[117]  ;
  assign n1190 = \a[117]  & \b[117]  ;
  assign n1191 = ~n1189 & ~n1190 ;
  assign n1192 = n1188 & ~n1191 ;
  assign n1193 = ~n1188 & n1191 ;
  assign n1194 = ~n1192 & ~n1193 ;
  assign n1195 = ~n1188 & ~n1189 ;
  assign n1196 = ~n1190 & ~n1195 ;
  assign n1197 = ~\a[118]  & ~\b[118]  ;
  assign n1198 = \a[118]  & \b[118]  ;
  assign n1199 = ~n1197 & ~n1198 ;
  assign n1200 = n1196 & ~n1199 ;
  assign n1201 = ~n1196 & n1199 ;
  assign n1202 = ~n1200 & ~n1201 ;
  assign n1203 = ~n1196 & ~n1197 ;
  assign n1204 = ~n1198 & ~n1203 ;
  assign n1205 = ~\a[119]  & ~\b[119]  ;
  assign n1206 = \a[119]  & \b[119]  ;
  assign n1207 = ~n1205 & ~n1206 ;
  assign n1208 = n1204 & ~n1207 ;
  assign n1209 = ~n1204 & n1207 ;
  assign n1210 = ~n1208 & ~n1209 ;
  assign n1211 = ~n1204 & ~n1205 ;
  assign n1212 = ~n1206 & ~n1211 ;
  assign n1213 = ~\a[120]  & ~\b[120]  ;
  assign n1214 = \a[120]  & \b[120]  ;
  assign n1215 = ~n1213 & ~n1214 ;
  assign n1216 = n1212 & ~n1215 ;
  assign n1217 = ~n1212 & n1215 ;
  assign n1218 = ~n1216 & ~n1217 ;
  assign n1219 = ~n1212 & ~n1213 ;
  assign n1220 = ~n1214 & ~n1219 ;
  assign n1221 = ~\a[121]  & ~\b[121]  ;
  assign n1222 = \a[121]  & \b[121]  ;
  assign n1223 = ~n1221 & ~n1222 ;
  assign n1224 = n1220 & ~n1223 ;
  assign n1225 = ~n1220 & n1223 ;
  assign n1226 = ~n1224 & ~n1225 ;
  assign n1227 = ~n1220 & ~n1221 ;
  assign n1228 = ~n1222 & ~n1227 ;
  assign n1229 = ~\a[122]  & ~\b[122]  ;
  assign n1230 = \a[122]  & \b[122]  ;
  assign n1231 = ~n1229 & ~n1230 ;
  assign n1232 = n1228 & ~n1231 ;
  assign n1233 = ~n1228 & n1231 ;
  assign n1234 = ~n1232 & ~n1233 ;
  assign n1235 = ~n1228 & ~n1229 ;
  assign n1236 = ~n1230 & ~n1235 ;
  assign n1237 = ~\a[123]  & ~\b[123]  ;
  assign n1238 = \a[123]  & \b[123]  ;
  assign n1239 = ~n1237 & ~n1238 ;
  assign n1240 = n1236 & ~n1239 ;
  assign n1241 = ~n1236 & n1239 ;
  assign n1242 = ~n1240 & ~n1241 ;
  assign n1243 = ~n1236 & ~n1237 ;
  assign n1244 = ~n1238 & ~n1243 ;
  assign n1245 = ~\a[124]  & ~\b[124]  ;
  assign n1246 = \a[124]  & \b[124]  ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = n1244 & ~n1247 ;
  assign n1249 = ~n1244 & n1247 ;
  assign n1250 = ~n1248 & ~n1249 ;
  assign n1251 = ~n1244 & ~n1245 ;
  assign n1252 = ~n1246 & ~n1251 ;
  assign n1253 = ~\a[125]  & ~\b[125]  ;
  assign n1254 = \a[125]  & \b[125]  ;
  assign n1255 = ~n1253 & ~n1254 ;
  assign n1256 = n1252 & ~n1255 ;
  assign n1257 = ~n1252 & n1255 ;
  assign n1258 = ~n1256 & ~n1257 ;
  assign n1259 = ~n1252 & ~n1253 ;
  assign n1260 = ~n1254 & ~n1259 ;
  assign n1261 = ~\a[126]  & ~\b[126]  ;
  assign n1262 = \a[126]  & \b[126]  ;
  assign n1263 = ~n1261 & ~n1262 ;
  assign n1264 = n1260 & ~n1263 ;
  assign n1265 = ~n1260 & n1263 ;
  assign n1266 = ~n1264 & ~n1265 ;
  assign n1267 = ~n1260 & ~n1261 ;
  assign n1268 = ~n1262 & ~n1267 ;
  assign n1269 = ~\a[127]  & ~\b[127]  ;
  assign n1270 = \a[127]  & \b[127]  ;
  assign n1271 = ~n1269 & ~n1270 ;
  assign n1272 = n1268 & ~n1271 ;
  assign n1273 = ~n1268 & n1271 ;
  assign n1274 = ~n1272 & ~n1273 ;
  assign n1275 = ~n1268 & ~n1269 ;
  assign n1276 = ~n1270 & ~n1275 ;
  assign \f[0]  = ~n259 ;
  assign \f[1]  = ~n266 ;
  assign \f[2]  = n274 ;
  assign \f[3]  = n282 ;
  assign \f[4]  = n290 ;
  assign \f[5]  = n298 ;
  assign \f[6]  = n306 ;
  assign \f[7]  = n314 ;
  assign \f[8]  = n322 ;
  assign \f[9]  = n330 ;
  assign \f[10]  = n338 ;
  assign \f[11]  = n346 ;
  assign \f[12]  = n354 ;
  assign \f[13]  = n362 ;
  assign \f[14]  = n370 ;
  assign \f[15]  = n378 ;
  assign \f[16]  = n386 ;
  assign \f[17]  = n394 ;
  assign \f[18]  = n402 ;
  assign \f[19]  = n410 ;
  assign \f[20]  = n418 ;
  assign \f[21]  = n426 ;
  assign \f[22]  = n434 ;
  assign \f[23]  = n442 ;
  assign \f[24]  = n450 ;
  assign \f[25]  = n458 ;
  assign \f[26]  = n466 ;
  assign \f[27]  = n474 ;
  assign \f[28]  = n482 ;
  assign \f[29]  = n490 ;
  assign \f[30]  = n498 ;
  assign \f[31]  = n506 ;
  assign \f[32]  = n514 ;
  assign \f[33]  = n522 ;
  assign \f[34]  = n530 ;
  assign \f[35]  = n538 ;
  assign \f[36]  = n546 ;
  assign \f[37]  = n554 ;
  assign \f[38]  = n562 ;
  assign \f[39]  = n570 ;
  assign \f[40]  = n578 ;
  assign \f[41]  = n586 ;
  assign \f[42]  = n594 ;
  assign \f[43]  = n602 ;
  assign \f[44]  = n610 ;
  assign \f[45]  = n618 ;
  assign \f[46]  = n626 ;
  assign \f[47]  = n634 ;
  assign \f[48]  = n642 ;
  assign \f[49]  = n650 ;
  assign \f[50]  = n658 ;
  assign \f[51]  = n666 ;
  assign \f[52]  = n674 ;
  assign \f[53]  = n682 ;
  assign \f[54]  = n690 ;
  assign \f[55]  = n698 ;
  assign \f[56]  = n706 ;
  assign \f[57]  = n714 ;
  assign \f[58]  = n722 ;
  assign \f[59]  = n730 ;
  assign \f[60]  = n738 ;
  assign \f[61]  = n746 ;
  assign \f[62]  = n754 ;
  assign \f[63]  = n762 ;
  assign \f[64]  = n770 ;
  assign \f[65]  = n778 ;
  assign \f[66]  = n786 ;
  assign \f[67]  = n794 ;
  assign \f[68]  = n802 ;
  assign \f[69]  = n810 ;
  assign \f[70]  = n818 ;
  assign \f[71]  = n826 ;
  assign \f[72]  = n834 ;
  assign \f[73]  = n842 ;
  assign \f[74]  = n850 ;
  assign \f[75]  = n858 ;
  assign \f[76]  = n866 ;
  assign \f[77]  = n874 ;
  assign \f[78]  = n882 ;
  assign \f[79]  = n890 ;
  assign \f[80]  = n898 ;
  assign \f[81]  = n906 ;
  assign \f[82]  = n914 ;
  assign \f[83]  = n922 ;
  assign \f[84]  = n930 ;
  assign \f[85]  = n938 ;
  assign \f[86]  = n946 ;
  assign \f[87]  = n954 ;
  assign \f[88]  = n962 ;
  assign \f[89]  = n970 ;
  assign \f[90]  = n978 ;
  assign \f[91]  = n986 ;
  assign \f[92]  = n994 ;
  assign \f[93]  = n1002 ;
  assign \f[94]  = n1010 ;
  assign \f[95]  = n1018 ;
  assign \f[96]  = n1026 ;
  assign \f[97]  = n1034 ;
  assign \f[98]  = n1042 ;
  assign \f[99]  = n1050 ;
  assign \f[100]  = n1058 ;
  assign \f[101]  = n1066 ;
  assign \f[102]  = n1074 ;
  assign \f[103]  = n1082 ;
  assign \f[104]  = n1090 ;
  assign \f[105]  = n1098 ;
  assign \f[106]  = n1106 ;
  assign \f[107]  = n1114 ;
  assign \f[108]  = n1122 ;
  assign \f[109]  = n1130 ;
  assign \f[110]  = n1138 ;
  assign \f[111]  = n1146 ;
  assign \f[112]  = n1154 ;
  assign \f[113]  = n1162 ;
  assign \f[114]  = n1170 ;
  assign \f[115]  = n1178 ;
  assign \f[116]  = n1186 ;
  assign \f[117]  = n1194 ;
  assign \f[118]  = n1202 ;
  assign \f[119]  = n1210 ;
  assign \f[120]  = n1218 ;
  assign \f[121]  = n1226 ;
  assign \f[122]  = n1234 ;
  assign \f[123]  = n1242 ;
  assign \f[124]  = n1250 ;
  assign \f[125]  = n1258 ;
  assign \f[126]  = n1266 ;
  assign \f[127]  = n1274 ;
  assign cOut = ~n1276 ;
endmodule
