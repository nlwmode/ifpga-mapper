module top( \g108_reg/NET0131  , \g109_pad  , \g1212_reg/NET0131  , \g1218_reg/NET0131  , \g1223_reg/NET0131  , \g1227_reg/NET0131  , \g1231_reg/NET0131  , \g1235_reg/NET0131  , \g1240_reg/NET0131  , \g1245_reg/NET0131  , \g1250_reg/NET0131  , \g1255_reg/NET0131  , \g1260_reg/NET0131  , \g1265_reg/NET0131  , \g1270_reg/NET0131  , \g1275_reg/NET0131  , \g1280_reg/NET0131  , \g1284_reg/NET0131  , \g1289_reg/NET0131  , \g1292_reg/NET0131  , \g1296_reg/NET0131  , \g1300_reg/NET0131  , \g1304_reg/NET0131  , \g1336_reg/NET0131  , \g1341_reg/NET0131  , \g1346_reg/NET0131  , \g1351_reg/NET0131  , \g1361_reg/NET0131  , \g1362_reg/NET0131  , \g1365_reg/NET0131  , \g1368_reg/NET0131  , \g1371_reg/NET0131  , \g1374_reg/NET0131  , \g1377_reg/NET0131  , \g1380_reg/NET0131  , \g1383_reg/NET0131  , \g1386_reg/NET0131  , \g1389_reg/NET0131  , \g1397_reg/NET0131  , \g1400_reg/NET0131  , \g1615_reg/NET0131  , \g1618_reg/NET0131  , \g1621_reg/NET0131  , \g1624_reg/NET0131  , \g1627_reg/NET0131  , \g1630_reg/NET0131  , \g1633_reg/NET0131  , \g1636_reg/NET0131  , \g1718_reg/NET0131  , \g186_reg/NET0131  , \g192_reg/NET0131  , \g197_reg/NET0131  , \g201_reg/NET0131  , \g207_reg/NET0131  , \g213_reg/NET0131  , \g219_reg/NET0131  , \g225_reg/NET0131  , \g231_reg/NET0131  , \g2355_pad  , \g237_reg/NET0131  , \g243_reg/NET0131  , \g248_reg/NET0131  , \g3007_pad  , \g305_reg/NET0131  , \g3069_pad  , \g309_reg/NET0131  , \g312_reg/NET0131  , \g315_reg/NET0131  , \g318_reg/NET0131  , \g321_reg/NET0131  , \g324_reg/NET0131  , \g327_reg/NET0131  , \g330_reg/NET0131  , \g333_reg/NET0131  , \g369_reg/NET0131  , \g374_reg/NET0131  , \g378_reg/NET0131  , \g382_reg/NET0131  , \g386_reg/NET0131  , \g391_reg/NET0131  , \g396_reg/NET0131  , \g401_reg/NET0131  , \g406_reg/NET0131  , \g411_reg/NET0131  , \g416_reg/NET0131  , \g4173_pad  , \g4174_pad  , \g4175_pad  , \g4176_pad  , \g4177_pad  , \g4178_pad  , \g4179_pad  , \g4180_pad  , \g4181_pad  , \g421_reg/NET0131  , \g426_reg/NET0131  , \g431_reg/NET0131  , \g435_reg/NET0131  , \g440_reg/NET0131  , \g444_reg/NET0131  , \g448_reg/NET0131  , \g452_reg/NET0131  , \g546_reg/NET0131  , \g549_reg/NET0131  , \g554_reg/NET0131  , \g557_reg/NET0131  , \g560_reg/NET0131  , \g563_reg/NET0131  , \g566_reg/NET0131  , \g569_reg/NET0131  , \g572_reg/NET0131  , \g575_reg/NET0131  , \g741_pad  , \g742_pad  , \g743_pad  , \g744_pad  , \g757_reg/NET0131  , \g876_reg/NET0131  , \g971_reg/NET0131  , \g976_reg/NET0131  , \g981_reg/NET0131  , \g986_reg/NET0131  , \g21280/_0_  , \g21281/_0_  , \g21282/_0_  , \g21307/_0_  , \g21322/_0_  , \g21333/_0_  , \g21334/_0_  , \g21338/_0_  , \g21350/_0_  , \g21355/_0_  , \g21356/_0_  , \g21357/_0_  , \g21358/_1_  , \g21359/_0_  , \g21370/_0_  , \g21371/_0_  , \g21378/_0_  , \g21379/_0_  , \g21380/_1_  , \g21381/_0_  , \g21390/_0_  , \g21394/_0_  , \g21396/_0_  , \g21397/_0_  , \g21398/_1_  , \g21412/_0_  , \g21413/_0_  , \g21419/_0_  , \g21420/_00_  , \g21421/_00_  , \g21424/_0_  , \g21425/_0_  , \g21426/_1_  , \g21437/_0_  , \g21444/_0_  , \g21450/_0_  , \g21455/_0_  , \g21457/_0_  , \g21458/_1_  , \g21459/_0_  , \g21470/_0_  , \g21486/_0_  , \g21487/_0_  , \g21495/_0_  , \g21498/_1_  , \g21499/_0_  , \g21500/_0_  , \g21502/_0_  , \g21503/_0_  , \g21508/_0_  , \g21509/_0_  , \g21510/_0_  , \g21511/_0_  , \g21515/_0_  , \g21520/_0_  , \g21523/_0_  , \g21524/_0_  , \g21525/_0_  , \g21538/_0_  , \g21544/_0_  , \g21550/_1_  , \g21562/_0_  , \g21563/_0_  , \g21584/_0_  , \g21591/_0_  , \g21593/_0_  , \g21601/_3_  , \g21603/_3_  , \g21605/_3_  , \g21607/_3_  , \g21609/_3_  , \g21611/_3_  , \g21613/_3_  , \g21615/_3_  , \g21617/_3_  , \g21619/_3_  , \g21621/_3_  , \g21623/_3_  , \g21625/_3_  , \g21627/_3_  , \g21640/_0_  , \g21641/_0_  , \g21642/_0_  , \g21693/_0_  , \g21694/_0_  , \g21735/_2_  , \g21745/_2_  , \g21796/_0_  , \g21799/_0_  , \g21803/_0_  , \g21812/_0_  , \g21814/_0_  , \g21816/_0_  , \g21828/_0_  , \g22203/_0_  , \g22260/_1_  , \g22317/_0_  , \g22339/_0_  , \g22392/_0_  , \g22395/_1_  , \g2601_pad  , \g27_dup/_0_  , \g5816_pad  );
  input \g108_reg/NET0131  ;
  input \g109_pad  ;
  input \g1212_reg/NET0131  ;
  input \g1218_reg/NET0131  ;
  input \g1223_reg/NET0131  ;
  input \g1227_reg/NET0131  ;
  input \g1231_reg/NET0131  ;
  input \g1235_reg/NET0131  ;
  input \g1240_reg/NET0131  ;
  input \g1245_reg/NET0131  ;
  input \g1250_reg/NET0131  ;
  input \g1255_reg/NET0131  ;
  input \g1260_reg/NET0131  ;
  input \g1265_reg/NET0131  ;
  input \g1270_reg/NET0131  ;
  input \g1275_reg/NET0131  ;
  input \g1280_reg/NET0131  ;
  input \g1284_reg/NET0131  ;
  input \g1289_reg/NET0131  ;
  input \g1292_reg/NET0131  ;
  input \g1296_reg/NET0131  ;
  input \g1300_reg/NET0131  ;
  input \g1304_reg/NET0131  ;
  input \g1336_reg/NET0131  ;
  input \g1341_reg/NET0131  ;
  input \g1346_reg/NET0131  ;
  input \g1351_reg/NET0131  ;
  input \g1361_reg/NET0131  ;
  input \g1362_reg/NET0131  ;
  input \g1365_reg/NET0131  ;
  input \g1368_reg/NET0131  ;
  input \g1371_reg/NET0131  ;
  input \g1374_reg/NET0131  ;
  input \g1377_reg/NET0131  ;
  input \g1380_reg/NET0131  ;
  input \g1383_reg/NET0131  ;
  input \g1386_reg/NET0131  ;
  input \g1389_reg/NET0131  ;
  input \g1397_reg/NET0131  ;
  input \g1400_reg/NET0131  ;
  input \g1615_reg/NET0131  ;
  input \g1618_reg/NET0131  ;
  input \g1621_reg/NET0131  ;
  input \g1624_reg/NET0131  ;
  input \g1627_reg/NET0131  ;
  input \g1630_reg/NET0131  ;
  input \g1633_reg/NET0131  ;
  input \g1636_reg/NET0131  ;
  input \g1718_reg/NET0131  ;
  input \g186_reg/NET0131  ;
  input \g192_reg/NET0131  ;
  input \g197_reg/NET0131  ;
  input \g201_reg/NET0131  ;
  input \g207_reg/NET0131  ;
  input \g213_reg/NET0131  ;
  input \g219_reg/NET0131  ;
  input \g225_reg/NET0131  ;
  input \g231_reg/NET0131  ;
  input \g2355_pad  ;
  input \g237_reg/NET0131  ;
  input \g243_reg/NET0131  ;
  input \g248_reg/NET0131  ;
  input \g3007_pad  ;
  input \g305_reg/NET0131  ;
  input \g3069_pad  ;
  input \g309_reg/NET0131  ;
  input \g312_reg/NET0131  ;
  input \g315_reg/NET0131  ;
  input \g318_reg/NET0131  ;
  input \g321_reg/NET0131  ;
  input \g324_reg/NET0131  ;
  input \g327_reg/NET0131  ;
  input \g330_reg/NET0131  ;
  input \g333_reg/NET0131  ;
  input \g369_reg/NET0131  ;
  input \g374_reg/NET0131  ;
  input \g378_reg/NET0131  ;
  input \g382_reg/NET0131  ;
  input \g386_reg/NET0131  ;
  input \g391_reg/NET0131  ;
  input \g396_reg/NET0131  ;
  input \g401_reg/NET0131  ;
  input \g406_reg/NET0131  ;
  input \g411_reg/NET0131  ;
  input \g416_reg/NET0131  ;
  input \g4173_pad  ;
  input \g4174_pad  ;
  input \g4175_pad  ;
  input \g4176_pad  ;
  input \g4177_pad  ;
  input \g4178_pad  ;
  input \g4179_pad  ;
  input \g4180_pad  ;
  input \g4181_pad  ;
  input \g421_reg/NET0131  ;
  input \g426_reg/NET0131  ;
  input \g431_reg/NET0131  ;
  input \g435_reg/NET0131  ;
  input \g440_reg/NET0131  ;
  input \g444_reg/NET0131  ;
  input \g448_reg/NET0131  ;
  input \g452_reg/NET0131  ;
  input \g546_reg/NET0131  ;
  input \g549_reg/NET0131  ;
  input \g554_reg/NET0131  ;
  input \g557_reg/NET0131  ;
  input \g560_reg/NET0131  ;
  input \g563_reg/NET0131  ;
  input \g566_reg/NET0131  ;
  input \g569_reg/NET0131  ;
  input \g572_reg/NET0131  ;
  input \g575_reg/NET0131  ;
  input \g741_pad  ;
  input \g742_pad  ;
  input \g743_pad  ;
  input \g744_pad  ;
  input \g757_reg/NET0131  ;
  input \g876_reg/NET0131  ;
  input \g971_reg/NET0131  ;
  input \g976_reg/NET0131  ;
  input \g981_reg/NET0131  ;
  input \g986_reg/NET0131  ;
  output \g21280/_0_  ;
  output \g21281/_0_  ;
  output \g21282/_0_  ;
  output \g21307/_0_  ;
  output \g21322/_0_  ;
  output \g21333/_0_  ;
  output \g21334/_0_  ;
  output \g21338/_0_  ;
  output \g21350/_0_  ;
  output \g21355/_0_  ;
  output \g21356/_0_  ;
  output \g21357/_0_  ;
  output \g21358/_1_  ;
  output \g21359/_0_  ;
  output \g21370/_0_  ;
  output \g21371/_0_  ;
  output \g21378/_0_  ;
  output \g21379/_0_  ;
  output \g21380/_1_  ;
  output \g21381/_0_  ;
  output \g21390/_0_  ;
  output \g21394/_0_  ;
  output \g21396/_0_  ;
  output \g21397/_0_  ;
  output \g21398/_1_  ;
  output \g21412/_0_  ;
  output \g21413/_0_  ;
  output \g21419/_0_  ;
  output \g21420/_00_  ;
  output \g21421/_00_  ;
  output \g21424/_0_  ;
  output \g21425/_0_  ;
  output \g21426/_1_  ;
  output \g21437/_0_  ;
  output \g21444/_0_  ;
  output \g21450/_0_  ;
  output \g21455/_0_  ;
  output \g21457/_0_  ;
  output \g21458/_1_  ;
  output \g21459/_0_  ;
  output \g21470/_0_  ;
  output \g21486/_0_  ;
  output \g21487/_0_  ;
  output \g21495/_0_  ;
  output \g21498/_1_  ;
  output \g21499/_0_  ;
  output \g21500/_0_  ;
  output \g21502/_0_  ;
  output \g21503/_0_  ;
  output \g21508/_0_  ;
  output \g21509/_0_  ;
  output \g21510/_0_  ;
  output \g21511/_0_  ;
  output \g21515/_0_  ;
  output \g21520/_0_  ;
  output \g21523/_0_  ;
  output \g21524/_0_  ;
  output \g21525/_0_  ;
  output \g21538/_0_  ;
  output \g21544/_0_  ;
  output \g21550/_1_  ;
  output \g21562/_0_  ;
  output \g21563/_0_  ;
  output \g21584/_0_  ;
  output \g21591/_0_  ;
  output \g21593/_0_  ;
  output \g21601/_3_  ;
  output \g21603/_3_  ;
  output \g21605/_3_  ;
  output \g21607/_3_  ;
  output \g21609/_3_  ;
  output \g21611/_3_  ;
  output \g21613/_3_  ;
  output \g21615/_3_  ;
  output \g21617/_3_  ;
  output \g21619/_3_  ;
  output \g21621/_3_  ;
  output \g21623/_3_  ;
  output \g21625/_3_  ;
  output \g21627/_3_  ;
  output \g21640/_0_  ;
  output \g21641/_0_  ;
  output \g21642/_0_  ;
  output \g21693/_0_  ;
  output \g21694/_0_  ;
  output \g21735/_2_  ;
  output \g21745/_2_  ;
  output \g21796/_0_  ;
  output \g21799/_0_  ;
  output \g21803/_0_  ;
  output \g21812/_0_  ;
  output \g21814/_0_  ;
  output \g21816/_0_  ;
  output \g21828/_0_  ;
  output \g22203/_0_  ;
  output \g22260/_1_  ;
  output \g22317/_0_  ;
  output \g22339/_0_  ;
  output \g22392/_0_  ;
  output \g22395/_1_  ;
  output \g2601_pad  ;
  output \g27_dup/_0_  ;
  output \g5816_pad  ;
  wire n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 ;
  assign n123 = \g369_reg/NET0131  & \g374_reg/NET0131  ;
  assign n124 = \g378_reg/NET0131  & n123 ;
  assign n125 = \g382_reg/NET0131  & n124 ;
  assign n150 = ~\g396_reg/NET0131  & ~\g401_reg/NET0131  ;
  assign n151 = ~\g406_reg/NET0131  & ~\g411_reg/NET0131  ;
  assign n157 = n150 & n151 ;
  assign n148 = ~\g431_reg/NET0131  & ~\g435_reg/NET0131  ;
  assign n149 = ~\g386_reg/NET0131  & ~\g391_reg/NET0131  ;
  assign n158 = n148 & n149 ;
  assign n159 = n157 & n158 ;
  assign n154 = ~\g444_reg/NET0131  & ~\g448_reg/NET0131  ;
  assign n155 = ~\g452_reg/NET0131  & n154 ;
  assign n152 = ~\g416_reg/NET0131  & ~\g421_reg/NET0131  ;
  assign n153 = ~\g426_reg/NET0131  & ~\g440_reg/NET0131  ;
  assign n156 = n152 & n153 ;
  assign n160 = n155 & n156 ;
  assign n161 = n159 & n160 ;
  assign n162 = \g431_reg/NET0131  & \g435_reg/NET0131  ;
  assign n163 = ~n148 & ~n162 ;
  assign n164 = ~n161 & ~n163 ;
  assign n166 = \g305_reg/NET0131  & n164 ;
  assign n165 = ~\g305_reg/NET0131  & ~n164 ;
  assign n142 = ~\g315_reg/NET0131  & ~\g426_reg/NET0131  ;
  assign n143 = \g315_reg/NET0131  & \g426_reg/NET0131  ;
  assign n144 = ~n142 & ~n143 ;
  assign n134 = ~\g324_reg/NET0131  & ~\g396_reg/NET0131  ;
  assign n135 = \g324_reg/NET0131  & \g396_reg/NET0131  ;
  assign n136 = ~n134 & ~n135 ;
  assign n137 = ~\g312_reg/NET0131  & ~\g421_reg/NET0131  ;
  assign n138 = \g312_reg/NET0131  & \g421_reg/NET0131  ;
  assign n139 = ~n137 & ~n138 ;
  assign n175 = ~n136 & ~n139 ;
  assign n176 = ~n144 & n175 ;
  assign n141 = ~\g330_reg/NET0131  & \g406_reg/NET0131  ;
  assign n145 = \g318_reg/NET0131  & ~\g386_reg/NET0131  ;
  assign n170 = ~n141 & ~n145 ;
  assign n146 = ~\g318_reg/NET0131  & \g386_reg/NET0131  ;
  assign n147 = \g321_reg/NET0131  & ~\g391_reg/NET0131  ;
  assign n171 = ~n146 & ~n147 ;
  assign n172 = n170 & n171 ;
  assign n128 = ~\g321_reg/NET0131  & \g391_reg/NET0131  ;
  assign n129 = ~\g333_reg/NET0131  & \g411_reg/NET0131  ;
  assign n168 = ~n128 & ~n129 ;
  assign n130 = \g309_reg/NET0131  & ~\g416_reg/NET0131  ;
  assign n140 = \g330_reg/NET0131  & ~\g406_reg/NET0131  ;
  assign n169 = ~n130 & ~n140 ;
  assign n173 = n168 & n169 ;
  assign n131 = ~\g327_reg/NET0131  & ~\g401_reg/NET0131  ;
  assign n132 = \g327_reg/NET0131  & \g401_reg/NET0131  ;
  assign n133 = ~n131 & ~n132 ;
  assign n126 = ~\g309_reg/NET0131  & \g416_reg/NET0131  ;
  assign n127 = \g333_reg/NET0131  & ~\g411_reg/NET0131  ;
  assign n167 = ~n126 & ~n127 ;
  assign n174 = ~n133 & n167 ;
  assign n177 = n173 & n174 ;
  assign n178 = n172 & n177 ;
  assign n179 = n176 & n178 ;
  assign n180 = ~n165 & n179 ;
  assign n181 = ~n166 & n180 ;
  assign n182 = n125 & ~n181 ;
  assign n183 = \g3007_pad  & ~\g876_reg/NET0131  ;
  assign n184 = \g1212_reg/NET0131  & ~\g757_reg/NET0131  ;
  assign n185 = ~n183 & n184 ;
  assign n186 = \g109_pad  & ~n185 ;
  assign n187 = ~n182 & n186 ;
  assign n188 = \g976_reg/NET0131  & n187 ;
  assign n189 = \g971_reg/NET0131  & \g976_reg/NET0131  ;
  assign n190 = ~\g971_reg/NET0131  & ~\g976_reg/NET0131  ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = n186 & n191 ;
  assign n193 = n182 & n192 ;
  assign n194 = ~n188 & ~n193 ;
  assign n195 = \g981_reg/NET0131  & n187 ;
  assign n196 = \g981_reg/NET0131  & n189 ;
  assign n197 = ~\g981_reg/NET0131  & ~n189 ;
  assign n198 = ~n196 & ~n197 ;
  assign n199 = n186 & n198 ;
  assign n200 = n182 & n199 ;
  assign n201 = ~n195 & ~n200 ;
  assign n202 = \g986_reg/NET0131  & n187 ;
  assign n204 = \g986_reg/NET0131  & n196 ;
  assign n203 = ~\g986_reg/NET0131  & ~n196 ;
  assign n205 = n186 & ~n203 ;
  assign n206 = ~n204 & n205 ;
  assign n207 = n182 & n206 ;
  assign n208 = ~n202 & ~n207 ;
  assign n215 = ~\g1362_reg/NET0131  & ~\g1365_reg/NET0131  ;
  assign n216 = ~\g1368_reg/NET0131  & ~\g1371_reg/NET0131  ;
  assign n229 = n215 & n216 ;
  assign n209 = ~\g1386_reg/NET0131  & ~\g1389_reg/NET0131  ;
  assign n212 = ~\g197_reg/NET0131  & ~\g201_reg/NET0131  ;
  assign n230 = n209 & n212 ;
  assign n231 = n229 & n230 ;
  assign n219 = ~\g1397_reg/NET0131  & ~\g1400_reg/NET0131  ;
  assign n220 = ~\g186_reg/NET0131  & ~\g192_reg/NET0131  ;
  assign n227 = n219 & n220 ;
  assign n217 = ~\g1374_reg/NET0131  & ~\g1377_reg/NET0131  ;
  assign n218 = ~\g1380_reg/NET0131  & ~\g1383_reg/NET0131  ;
  assign n228 = n217 & n218 ;
  assign n232 = n227 & n228 ;
  assign n223 = ~\g231_reg/NET0131  & ~\g237_reg/NET0131  ;
  assign n224 = ~\g243_reg/NET0131  & ~\g248_reg/NET0131  ;
  assign n225 = n223 & n224 ;
  assign n221 = ~\g207_reg/NET0131  & ~\g213_reg/NET0131  ;
  assign n222 = ~\g219_reg/NET0131  & ~\g225_reg/NET0131  ;
  assign n226 = n221 & n222 ;
  assign n233 = n225 & n226 ;
  assign n234 = n232 & n233 ;
  assign n235 = n231 & n234 ;
  assign n210 = \g1386_reg/NET0131  & \g1389_reg/NET0131  ;
  assign n211 = ~n209 & ~n210 ;
  assign n213 = \g197_reg/NET0131  & \g201_reg/NET0131  ;
  assign n214 = ~n212 & ~n213 ;
  assign n236 = ~n211 & ~n214 ;
  assign n237 = ~n235 & n236 ;
  assign n238 = n211 & n214 ;
  assign n239 = \g109_pad  & ~n238 ;
  assign n240 = ~n237 & n239 ;
  assign n241 = ~\g2355_pad  & \g557_reg/NET0131  ;
  assign n242 = \g213_reg/NET0131  & \g2355_pad  ;
  assign n243 = ~n241 & ~n242 ;
  assign n244 = ~\g2355_pad  & \g546_reg/NET0131  ;
  assign n245 = \g186_reg/NET0131  & \g2355_pad  ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = \g1615_reg/NET0131  & ~\g2355_pad  ;
  assign n248 = ~n242 & ~n247 ;
  assign n249 = ~\g1718_reg/NET0131  & ~n248 ;
  assign n250 = ~\g2355_pad  & \g560_reg/NET0131  ;
  assign n251 = \g219_reg/NET0131  & \g2355_pad  ;
  assign n252 = ~n250 & ~n251 ;
  assign n253 = \g1618_reg/NET0131  & ~\g2355_pad  ;
  assign n254 = ~n245 & ~n253 ;
  assign n255 = ~\g1718_reg/NET0131  & ~n254 ;
  assign n256 = ~\g2355_pad  & \g554_reg/NET0131  ;
  assign n257 = \g207_reg/NET0131  & \g2355_pad  ;
  assign n258 = ~n256 & ~n257 ;
  assign n259 = \g1621_reg/NET0131  & ~\g2355_pad  ;
  assign n260 = ~n251 & ~n259 ;
  assign n261 = ~\g1718_reg/NET0131  & ~n260 ;
  assign n262 = \g109_pad  & \g186_reg/NET0131  ;
  assign n263 = ~\g2355_pad  & \g563_reg/NET0131  ;
  assign n264 = \g225_reg/NET0131  & \g2355_pad  ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = \g109_pad  & \g1383_reg/NET0131  ;
  assign n267 = ~\g1718_reg/NET0131  & ~n257 ;
  assign n268 = \g1624_reg/NET0131  & ~\g2355_pad  ;
  assign n269 = ~n264 & ~n268 ;
  assign n270 = ~\g1718_reg/NET0131  & ~n269 ;
  assign n271 = \g109_pad  & \g207_reg/NET0131  ;
  assign n272 = ~\g2355_pad  & \g566_reg/NET0131  ;
  assign n273 = \g231_reg/NET0131  & \g2355_pad  ;
  assign n274 = ~n272 & ~n273 ;
  assign n275 = \g109_pad  & \g1380_reg/NET0131  ;
  assign n276 = \g1627_reg/NET0131  & ~\g2355_pad  ;
  assign n277 = ~n273 & ~n276 ;
  assign n278 = ~\g1718_reg/NET0131  & ~n277 ;
  assign n279 = ~\g2355_pad  & \g569_reg/NET0131  ;
  assign n280 = \g2355_pad  & \g237_reg/NET0131  ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = \g109_pad  & \g213_reg/NET0131  ;
  assign n283 = \g4173_pad  & \g4174_pad  ;
  assign n284 = \g4175_pad  & n283 ;
  assign n285 = \g4176_pad  & n284 ;
  assign n286 = \g4177_pad  & n285 ;
  assign n287 = \g4178_pad  & n286 ;
  assign n288 = \g4179_pad  & n287 ;
  assign n289 = \g4180_pad  & n288 ;
  assign n291 = \g4181_pad  & n289 ;
  assign n292 = ~\g1718_reg/NET0131  & ~n291 ;
  assign n290 = ~\g4181_pad  & ~n289 ;
  assign n293 = \g109_pad  & ~n290 ;
  assign n294 = n292 & n293 ;
  assign n295 = \g109_pad  & \g1377_reg/NET0131  ;
  assign n296 = \g1630_reg/NET0131  & ~\g2355_pad  ;
  assign n297 = ~n280 & ~n296 ;
  assign n298 = ~\g1718_reg/NET0131  & ~n297 ;
  assign n302 = ~\g1240_reg/NET0131  & ~\g1245_reg/NET0131  ;
  assign n303 = ~\g1255_reg/NET0131  & ~\g1260_reg/NET0131  ;
  assign n304 = ~\g1270_reg/NET0131  & n303 ;
  assign n305 = n302 & n304 ;
  assign n299 = ~\g1235_reg/NET0131  & ~\g1250_reg/NET0131  ;
  assign n300 = ~\g1265_reg/NET0131  & ~\g1275_reg/NET0131  ;
  assign n301 = n299 & n300 ;
  assign n306 = ~\g1292_reg/NET0131  & ~\g1296_reg/NET0131  ;
  assign n307 = ~\g1300_reg/NET0131  & ~\g1304_reg/NET0131  ;
  assign n308 = n306 & n307 ;
  assign n309 = n301 & n308 ;
  assign n310 = n305 & n309 ;
  assign n311 = ~\g1280_reg/NET0131  & ~n310 ;
  assign n312 = ~\g1284_reg/NET0131  & ~n311 ;
  assign n313 = ~\g1280_reg/NET0131  & \g1284_reg/NET0131  ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = n301 & n305 ;
  assign n316 = n314 & n315 ;
  assign n317 = ~\g1212_reg/NET0131  & \g1289_reg/NET0131  ;
  assign n318 = \g1218_reg/NET0131  & \g1223_reg/NET0131  ;
  assign n319 = \g1227_reg/NET0131  & n318 ;
  assign n320 = n317 & n319 ;
  assign n321 = \g1231_reg/NET0131  & n320 ;
  assign n322 = ~n316 & n321 ;
  assign n323 = ~\g1361_reg/NET0131  & \g3069_pad  ;
  assign n324 = ~\g108_reg/NET0131  & \g1212_reg/NET0131  ;
  assign n325 = ~n323 & n324 ;
  assign n326 = \g109_pad  & ~n325 ;
  assign n327 = ~n322 & n326 ;
  assign n328 = \g1346_reg/NET0131  & n327 ;
  assign n329 = n322 & n326 ;
  assign n330 = \g1336_reg/NET0131  & \g1341_reg/NET0131  ;
  assign n331 = ~\g1346_reg/NET0131  & ~n330 ;
  assign n332 = \g1346_reg/NET0131  & n330 ;
  assign n333 = ~n331 & ~n332 ;
  assign n334 = n329 & n333 ;
  assign n335 = ~n328 & ~n334 ;
  assign n336 = \g1351_reg/NET0131  & n327 ;
  assign n337 = ~\g1351_reg/NET0131  & ~n332 ;
  assign n338 = \g1351_reg/NET0131  & n332 ;
  assign n339 = ~n337 & ~n338 ;
  assign n340 = n329 & n339 ;
  assign n341 = ~n336 & ~n340 ;
  assign n342 = ~\g2355_pad  & \g572_reg/NET0131  ;
  assign n343 = \g2355_pad  & \g243_reg/NET0131  ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = \g109_pad  & \g219_reg/NET0131  ;
  assign n347 = ~\g4180_pad  & ~n288 ;
  assign n346 = \g109_pad  & ~\g1718_reg/NET0131  ;
  assign n348 = ~n289 & n346 ;
  assign n349 = ~n347 & n348 ;
  assign n350 = \g109_pad  & \g1371_reg/NET0131  ;
  assign n351 = \g1633_reg/NET0131  & ~\g2355_pad  ;
  assign n352 = ~\g1718_reg/NET0131  & ~n343 ;
  assign n353 = ~n351 & n352 ;
  assign n354 = \g109_pad  & \g225_reg/NET0131  ;
  assign n355 = ~\g4179_pad  & ~n287 ;
  assign n356 = ~n288 & n346 ;
  assign n357 = ~n355 & n356 ;
  assign n358 = ~\g2355_pad  & \g575_reg/NET0131  ;
  assign n359 = \g2355_pad  & \g248_reg/NET0131  ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = \g109_pad  & \g1368_reg/NET0131  ;
  assign n362 = \g1636_reg/NET0131  & ~\g2355_pad  ;
  assign n363 = ~\g1718_reg/NET0131  & ~n359 ;
  assign n364 = ~n362 & n363 ;
  assign n365 = ~\g4178_pad  & ~n286 ;
  assign n366 = ~n287 & n346 ;
  assign n367 = ~n365 & n366 ;
  assign n368 = \g109_pad  & \g231_reg/NET0131  ;
  assign n370 = \g1231_reg/NET0131  & n319 ;
  assign n371 = n317 & ~n370 ;
  assign n373 = ~\g1218_reg/NET0131  & ~n371 ;
  assign n369 = \g109_pad  & ~\g1212_reg/NET0131  ;
  assign n372 = \g1218_reg/NET0131  & n371 ;
  assign n374 = n369 & ~n372 ;
  assign n375 = ~n373 & n374 ;
  assign n377 = \g1223_reg/NET0131  & n372 ;
  assign n376 = ~\g1223_reg/NET0131  & ~n372 ;
  assign n378 = n369 & ~n376 ;
  assign n379 = ~n377 & n378 ;
  assign n380 = ~\g1227_reg/NET0131  & ~n318 ;
  assign n381 = \g109_pad  & ~n319 ;
  assign n382 = ~n380 & n381 ;
  assign n383 = n371 & n382 ;
  assign n384 = \g1227_reg/NET0131  & n369 ;
  assign n385 = ~n371 & n384 ;
  assign n386 = ~n383 & ~n385 ;
  assign n387 = ~\g1231_reg/NET0131  & ~n320 ;
  assign n388 = n369 & ~n387 ;
  assign n389 = \g369_reg/NET0131  & ~n125 ;
  assign n390 = n369 & ~n389 ;
  assign n391 = ~\g369_reg/NET0131  & ~\g374_reg/NET0131  ;
  assign n392 = ~n123 & ~n391 ;
  assign n393 = ~n125 & ~n392 ;
  assign n394 = n369 & ~n393 ;
  assign n395 = ~\g382_reg/NET0131  & n124 ;
  assign n396 = ~\g378_reg/NET0131  & ~n123 ;
  assign n397 = n369 & ~n396 ;
  assign n398 = ~n395 & n397 ;
  assign n399 = ~\g382_reg/NET0131  & ~n124 ;
  assign n400 = n369 & ~n399 ;
  assign n401 = \g109_pad  & ~n317 ;
  assign n402 = \g1275_reg/NET0131  & n401 ;
  assign n403 = ~n314 & n321 ;
  assign n404 = ~n402 & ~n403 ;
  assign n405 = ~\g4177_pad  & ~n285 ;
  assign n406 = ~n286 & n346 ;
  assign n407 = ~n405 & n406 ;
  assign n408 = \g109_pad  & \g1365_reg/NET0131  ;
  assign n409 = ~\g2355_pad  & \g549_reg/NET0131  ;
  assign n410 = \g192_reg/NET0131  & \g2355_pad  ;
  assign n411 = ~n409 & ~n410 ;
  assign n412 = ~\g201_reg/NET0131  & \g2355_pad  ;
  assign n413 = \g109_pad  & \g237_reg/NET0131  ;
  assign n414 = ~\g4176_pad  & ~n284 ;
  assign n415 = ~n285 & n346 ;
  assign n416 = ~n414 & n415 ;
  assign n417 = ~\g1718_reg/NET0131  & ~n410 ;
  assign n418 = \g109_pad  & \g1362_reg/NET0131  ;
  assign n419 = ~\g4173_pad  & ~\g4174_pad  ;
  assign n420 = ~n283 & n346 ;
  assign n421 = ~n419 & n420 ;
  assign n422 = \g1275_reg/NET0131  & n317 ;
  assign n423 = \g1235_reg/NET0131  & n401 ;
  assign n424 = ~n422 & ~n423 ;
  assign n425 = \g1235_reg/NET0131  & n317 ;
  assign n426 = \g1240_reg/NET0131  & n401 ;
  assign n427 = ~n425 & ~n426 ;
  assign n428 = \g1240_reg/NET0131  & n317 ;
  assign n429 = \g1245_reg/NET0131  & n401 ;
  assign n430 = ~n428 & ~n429 ;
  assign n431 = \g1245_reg/NET0131  & n317 ;
  assign n432 = \g1250_reg/NET0131  & n401 ;
  assign n433 = ~n431 & ~n432 ;
  assign n434 = \g1250_reg/NET0131  & n317 ;
  assign n435 = \g1255_reg/NET0131  & n401 ;
  assign n436 = ~n434 & ~n435 ;
  assign n437 = \g1255_reg/NET0131  & n317 ;
  assign n438 = \g1260_reg/NET0131  & n401 ;
  assign n439 = ~n437 & ~n438 ;
  assign n440 = \g1260_reg/NET0131  & n317 ;
  assign n441 = \g1265_reg/NET0131  & n401 ;
  assign n442 = ~n440 & ~n441 ;
  assign n443 = \g1265_reg/NET0131  & n317 ;
  assign n444 = \g1270_reg/NET0131  & n401 ;
  assign n445 = ~n443 & ~n444 ;
  assign n446 = \g1284_reg/NET0131  & n317 ;
  assign n447 = \g1280_reg/NET0131  & n401 ;
  assign n448 = ~n446 & ~n447 ;
  assign n449 = \g1292_reg/NET0131  & n317 ;
  assign n450 = \g1284_reg/NET0131  & n401 ;
  assign n451 = ~n449 & ~n450 ;
  assign n452 = \g1296_reg/NET0131  & n317 ;
  assign n453 = \g1292_reg/NET0131  & n401 ;
  assign n454 = ~n452 & ~n453 ;
  assign n455 = \g1300_reg/NET0131  & n317 ;
  assign n456 = \g1296_reg/NET0131  & n401 ;
  assign n457 = ~n455 & ~n456 ;
  assign n458 = \g1304_reg/NET0131  & n317 ;
  assign n459 = \g1300_reg/NET0131  & n401 ;
  assign n460 = ~n458 & ~n459 ;
  assign n461 = \g1270_reg/NET0131  & n317 ;
  assign n462 = \g1304_reg/NET0131  & n401 ;
  assign n463 = ~n461 & ~n462 ;
  assign n464 = \g109_pad  & \g243_reg/NET0131  ;
  assign n465 = ~\g4173_pad  & n346 ;
  assign n466 = ~\g4175_pad  & ~n283 ;
  assign n467 = ~n284 & n346 ;
  assign n468 = ~n466 & n467 ;
  assign n469 = \g109_pad  & \g1400_reg/NET0131  ;
  assign n470 = ~\g1212_reg/NET0131  & ~\g1289_reg/NET0131  ;
  assign n471 = \g109_pad  & \g741_pad  ;
  assign n472 = \g742_pad  & n471 ;
  assign n473 = \g109_pad  & \g743_pad  ;
  assign n474 = \g744_pad  & n473 ;
  assign n475 = \g109_pad  & \g1374_reg/NET0131  ;
  assign n476 = \g109_pad  & \g197_reg/NET0131  ;
  assign n477 = \g109_pad  & \g201_reg/NET0131  ;
  assign n478 = \g109_pad  & \g1389_reg/NET0131  ;
  assign n479 = \g109_pad  & \g1397_reg/NET0131  ;
  assign n480 = \g109_pad  & \g192_reg/NET0131  ;
  assign n481 = \g109_pad  & \g248_reg/NET0131  ;
  assign n482 = \g1718_reg/NET0131  & n291 ;
  assign n483 = ~n292 & ~n482 ;
  assign n485 = \g971_reg/NET0131  & n182 ;
  assign n484 = ~\g971_reg/NET0131  & ~n182 ;
  assign n486 = n186 & ~n484 ;
  assign n487 = ~n485 & n486 ;
  assign n488 = ~\g1336_reg/NET0131  & n329 ;
  assign n489 = \g1336_reg/NET0131  & n327 ;
  assign n490 = ~n488 & ~n489 ;
  assign n491 = \g1341_reg/NET0131  & n327 ;
  assign n492 = ~\g1336_reg/NET0131  & ~\g1341_reg/NET0131  ;
  assign n493 = ~n330 & ~n492 ;
  assign n494 = n329 & n493 ;
  assign n495 = ~n491 & ~n494 ;
  assign n496 = n125 & ~n164 ;
  assign n497 = \g305_reg/NET0131  & ~n125 ;
  assign n498 = ~n496 & ~n497 ;
  assign \g21280/_0_  = ~n194 ;
  assign \g21281/_0_  = ~n201 ;
  assign \g21282/_0_  = ~n208 ;
  assign \g21307/_0_  = n240 ;
  assign \g21322/_0_  = ~n243 ;
  assign \g21333/_0_  = ~n246 ;
  assign \g21334/_0_  = n249 ;
  assign \g21338/_0_  = ~n252 ;
  assign \g21350/_0_  = n255 ;
  assign \g21355/_0_  = ~n258 ;
  assign \g21356/_0_  = n261 ;
  assign \g21357/_0_  = n262 ;
  assign \g21358/_1_  = n245 ;
  assign \g21359/_0_  = ~n265 ;
  assign \g21370/_0_  = n266 ;
  assign \g21371/_0_  = ~n267 ;
  assign \g21378/_0_  = n270 ;
  assign \g21379/_0_  = n271 ;
  assign \g21380/_1_  = n257 ;
  assign \g21381/_0_  = ~n274 ;
  assign \g21390/_0_  = n275 ;
  assign \g21394/_0_  = n278 ;
  assign \g21396/_0_  = ~n281 ;
  assign \g21397/_0_  = n282 ;
  assign \g21398/_1_  = n242 ;
  assign \g21412/_0_  = n294 ;
  assign \g21413/_0_  = n295 ;
  assign \g21419/_0_  = n298 ;
  assign \g21420/_00_  = ~n335 ;
  assign \g21421/_00_  = ~n341 ;
  assign \g21424/_0_  = ~n344 ;
  assign \g21425/_0_  = n345 ;
  assign \g21426/_1_  = n251 ;
  assign \g21437/_0_  = n349 ;
  assign \g21444/_0_  = n350 ;
  assign \g21450/_0_  = ~n353 ;
  assign \g21455/_0_  = n354 ;
  assign \g21457/_0_  = n357 ;
  assign \g21458/_1_  = n264 ;
  assign \g21459/_0_  = ~n360 ;
  assign \g21470/_0_  = n361 ;
  assign \g21486/_0_  = ~n364 ;
  assign \g21487/_0_  = n367 ;
  assign \g21495/_0_  = n368 ;
  assign \g21498/_1_  = n273 ;
  assign \g21499/_0_  = n375 ;
  assign \g21500/_0_  = n379 ;
  assign \g21502/_0_  = ~n386 ;
  assign \g21503/_0_  = n388 ;
  assign \g21508/_0_  = n390 ;
  assign \g21509/_0_  = n394 ;
  assign \g21510/_0_  = n398 ;
  assign \g21511/_0_  = n400 ;
  assign \g21515/_0_  = ~n404 ;
  assign \g21520/_0_  = n407 ;
  assign \g21523/_0_  = n408 ;
  assign \g21524/_0_  = ~n411 ;
  assign \g21525/_0_  = n412 ;
  assign \g21538/_0_  = n280 ;
  assign \g21544/_0_  = n413 ;
  assign \g21550/_1_  = n204 ;
  assign \g21562/_0_  = n416 ;
  assign \g21563/_0_  = ~n417 ;
  assign \g21584/_0_  = n338 ;
  assign \g21591/_0_  = n418 ;
  assign \g21593/_0_  = n421 ;
  assign \g21601/_3_  = ~n424 ;
  assign \g21603/_3_  = ~n427 ;
  assign \g21605/_3_  = ~n430 ;
  assign \g21607/_3_  = ~n433 ;
  assign \g21609/_3_  = ~n436 ;
  assign \g21611/_3_  = ~n439 ;
  assign \g21613/_3_  = ~n442 ;
  assign \g21615/_3_  = ~n445 ;
  assign \g21617/_3_  = ~n448 ;
  assign \g21619/_3_  = ~n451 ;
  assign \g21621/_3_  = ~n454 ;
  assign \g21623/_3_  = ~n457 ;
  assign \g21625/_3_  = ~n460 ;
  assign \g21627/_3_  = ~n463 ;
  assign \g21640/_0_  = n464 ;
  assign \g21641/_0_  = n465 ;
  assign \g21642/_0_  = n468 ;
  assign \g21693/_0_  = n469 ;
  assign \g21694/_0_  = ~n470 ;
  assign \g21735/_2_  = n472 ;
  assign \g21745/_2_  = n474 ;
  assign \g21796/_0_  = n475 ;
  assign \g21799/_0_  = n476 ;
  assign \g21803/_0_  = n477 ;
  assign \g21812/_0_  = n478 ;
  assign \g21814/_0_  = n479 ;
  assign \g21816/_0_  = n480 ;
  assign \g21828/_0_  = n481 ;
  assign \g22203/_0_  = n483 ;
  assign \g22260/_1_  = n182 ;
  assign \g22317/_0_  = n487 ;
  assign \g22339/_0_  = ~n490 ;
  assign \g22392/_0_  = ~n495 ;
  assign \g22395/_1_  = n322 ;
  assign \g2601_pad  = 1'b0 ;
  assign \g27_dup/_0_  = ~n498 ;
  assign \g5816_pad  = ~1'b0 ;
endmodule
