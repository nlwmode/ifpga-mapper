module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G1_pad , \G22_reg/NET0131 , \G23_reg/NET0131 , \G24_reg/NET0131 , \G25_reg/NET0131 , \G26_reg/NET0131 , \G27_reg/NET0131 , \G28_reg/NET0131 , \G29_reg/NET0131 , \G2_pad , \G30_reg/NET0131 , \G31_reg/NET0131 , \G32_reg/NET0131 , \G33_reg/NET0131 , \G34_reg/NET0131 , \G35_reg/NET0131 , \G36_reg/NET0131 , \G37_reg/NET0131 , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G43_reg/NET0131 , \G44_reg/NET0131 , \G45_reg/NET0131 , \G46_reg/NET0131 , \G47_reg/NET0131 , \G48_reg/NET0131 , \G49_reg/NET0131 , \G4_pad , \G50_reg/NET0131 , \G51_reg/NET0131 , \G52_reg/NET0131 , \G53_reg/NET0131 , \G55_reg/NET0131 , \G56_reg/NET0131 , \G57_reg/NET0131 , \G58_reg/NET0131 , \G59_reg/NET0131 , \G5_pad , \G60_reg/NET0131 , \G61_reg/NET0131 , \G62_reg/NET0131 , \G63_reg/NET0131 , \G64_reg/NET0131 , \G65_reg/NET0131 , \G66_reg/NET0131 , \G67_reg/NET0131 , \G68_reg/NET0131 , \G69_reg/NET0131 , \G6_pad , \G70_reg/NET0131 , \G71_reg/NET0131 , \G72_reg/NET0131 , \G73_reg/NET0131 , \G74_reg/NET0131 , \G75_reg/NET0131 , \G76_reg/NET0131 , \G77_reg/NET0131 , \G78_reg/NET0131 , \G79_reg/NET0131 , \G7_pad , \G80_reg/NET0131 , \G81_reg/NET0131 , \G82_reg/NET0131 , \G83_reg/NET0131 , \G84_reg/NET0131 , \G85_reg/NET0131 , \G86_reg/NET0131 , \G87_reg/NET0131 , \G88_reg/NET0131 , \G89_reg/NET0131 , \G8_pad , \G90_reg/NET0131 , \G91_reg/NET0131 , \G92_reg/NET0131 , \G94_reg/NET0131 , \G9_pad , \G701BF_pad , \G702_pad , \G727_pad , \_al_n0 , \_al_n1 , \g2503/_0_ , \g2514/_0_ , \g2516/_0_ , \g2542/_0_ , \g2549/_0_ , \g2553/_0_ , \g2554/_0_ , \g2570/_0_ , \g2574/_0_ , \g2576/_0_ , \g2583/_0_ , \g2588/_0_ , \g2602/_0_ , \g2603/_0_ , \g2604/_0_ , \g2605/_0_ , \g2611/_0_ , \g2614/_0_ , \g2615/_0_ , \g2644/_0_ , \g2657/_0_ , \g2663/_0_ , \g2664/_0_ , \g2666/_0_ , \g2672/_0_ , \g2678/_0_ , \g2681/_0_ , \g2696/_00_ , \g2698/_0_ , \g2699/_0_ , \g2700/_00_ , \g2717/_0_ , \g2719/_0_ , \g2723/_0_ , \g2726/_3_ , \g2735/_0_ , \g2737/_0_ , \g2740/_0_ , \g2785/_0_ , \g2786/_0_ , \g2787/_1__syn_2 , \g2790/_1__syn_2 , \g2798/_2_ , \g2801/_0_ , \g2841/_0_ , \g2844/_0_ , \g2845/_0_ , \g2846/_0_ , \g2860/_0_ , \g2861/_0_ , \g2862/_0_ , \g2864/_0_ , \g2882/_3_ , \g2883/_3_ , \g2887/_3_ , \g2906/_0_ , \g2911/_0_ , \g3282/_0_ , \g3406/_0_ , \g3409/_0_ , \g3506/_0_ , \g3685/_3_ , \g3694/_0_ , \g3743/_0_ , \g3753/_0_ , \g3785/_0_ , \g3835/_0_ , \g3946/_2_ , \g3976/_0_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G1_pad  ;
	input \G22_reg/NET0131  ;
	input \G23_reg/NET0131  ;
	input \G24_reg/NET0131  ;
	input \G25_reg/NET0131  ;
	input \G26_reg/NET0131  ;
	input \G27_reg/NET0131  ;
	input \G28_reg/NET0131  ;
	input \G29_reg/NET0131  ;
	input \G2_pad  ;
	input \G30_reg/NET0131  ;
	input \G31_reg/NET0131  ;
	input \G32_reg/NET0131  ;
	input \G33_reg/NET0131  ;
	input \G34_reg/NET0131  ;
	input \G35_reg/NET0131  ;
	input \G36_reg/NET0131  ;
	input \G37_reg/NET0131  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G43_reg/NET0131  ;
	input \G44_reg/NET0131  ;
	input \G45_reg/NET0131  ;
	input \G46_reg/NET0131  ;
	input \G47_reg/NET0131  ;
	input \G48_reg/NET0131  ;
	input \G49_reg/NET0131  ;
	input \G4_pad  ;
	input \G50_reg/NET0131  ;
	input \G51_reg/NET0131  ;
	input \G52_reg/NET0131  ;
	input \G53_reg/NET0131  ;
	input \G55_reg/NET0131  ;
	input \G56_reg/NET0131  ;
	input \G57_reg/NET0131  ;
	input \G58_reg/NET0131  ;
	input \G59_reg/NET0131  ;
	input \G5_pad  ;
	input \G60_reg/NET0131  ;
	input \G61_reg/NET0131  ;
	input \G62_reg/NET0131  ;
	input \G63_reg/NET0131  ;
	input \G64_reg/NET0131  ;
	input \G65_reg/NET0131  ;
	input \G66_reg/NET0131  ;
	input \G67_reg/NET0131  ;
	input \G68_reg/NET0131  ;
	input \G69_reg/NET0131  ;
	input \G6_pad  ;
	input \G70_reg/NET0131  ;
	input \G71_reg/NET0131  ;
	input \G72_reg/NET0131  ;
	input \G73_reg/NET0131  ;
	input \G74_reg/NET0131  ;
	input \G75_reg/NET0131  ;
	input \G76_reg/NET0131  ;
	input \G77_reg/NET0131  ;
	input \G78_reg/NET0131  ;
	input \G79_reg/NET0131  ;
	input \G7_pad  ;
	input \G80_reg/NET0131  ;
	input \G81_reg/NET0131  ;
	input \G82_reg/NET0131  ;
	input \G83_reg/NET0131  ;
	input \G84_reg/NET0131  ;
	input \G85_reg/NET0131  ;
	input \G86_reg/NET0131  ;
	input \G87_reg/NET0131  ;
	input \G88_reg/NET0131  ;
	input \G89_reg/NET0131  ;
	input \G8_pad  ;
	input \G90_reg/NET0131  ;
	input \G91_reg/NET0131  ;
	input \G92_reg/NET0131  ;
	input \G94_reg/NET0131  ;
	input \G9_pad  ;
	output \G701BF_pad  ;
	output \G702_pad  ;
	output \G727_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g2503/_0_  ;
	output \g2514/_0_  ;
	output \g2516/_0_  ;
	output \g2542/_0_  ;
	output \g2549/_0_  ;
	output \g2553/_0_  ;
	output \g2554/_0_  ;
	output \g2570/_0_  ;
	output \g2574/_0_  ;
	output \g2576/_0_  ;
	output \g2583/_0_  ;
	output \g2588/_0_  ;
	output \g2602/_0_  ;
	output \g2603/_0_  ;
	output \g2604/_0_  ;
	output \g2605/_0_  ;
	output \g2611/_0_  ;
	output \g2614/_0_  ;
	output \g2615/_0_  ;
	output \g2644/_0_  ;
	output \g2657/_0_  ;
	output \g2663/_0_  ;
	output \g2664/_0_  ;
	output \g2666/_0_  ;
	output \g2672/_0_  ;
	output \g2678/_0_  ;
	output \g2681/_0_  ;
	output \g2696/_00_  ;
	output \g2698/_0_  ;
	output \g2699/_0_  ;
	output \g2700/_00_  ;
	output \g2717/_0_  ;
	output \g2719/_0_  ;
	output \g2723/_0_  ;
	output \g2726/_3_  ;
	output \g2735/_0_  ;
	output \g2737/_0_  ;
	output \g2740/_0_  ;
	output \g2785/_0_  ;
	output \g2786/_0_  ;
	output \g2787/_1__syn_2  ;
	output \g2790/_1__syn_2  ;
	output \g2798/_2_  ;
	output \g2801/_0_  ;
	output \g2841/_0_  ;
	output \g2844/_0_  ;
	output \g2845/_0_  ;
	output \g2846/_0_  ;
	output \g2860/_0_  ;
	output \g2861/_0_  ;
	output \g2862/_0_  ;
	output \g2864/_0_  ;
	output \g2882/_3_  ;
	output \g2883/_3_  ;
	output \g2887/_3_  ;
	output \g2906/_0_  ;
	output \g2911/_0_  ;
	output \g3282/_0_  ;
	output \g3406/_0_  ;
	output \g3409/_0_  ;
	output \g3506/_0_  ;
	output \g3685/_3_  ;
	output \g3694/_0_  ;
	output \g3743/_0_  ;
	output \g3753/_0_  ;
	output \g3785/_0_  ;
	output \g3835/_0_  ;
	output \g3946/_2_  ;
	output \g3976/_0_  ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w266_ ;
	wire _w9_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w127_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w100_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\G15_pad ,
		_w9_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\G4_pad ,
		\G90_reg/NET0131 ,
		_w91_
	);
	LUT4 #(
		.INIT('h1130)
	) name2 (
		\G64_reg/NET0131 ,
		\G84_reg/NET0131 ,
		\G8_pad ,
		\G90_reg/NET0131 ,
		_w92_
	);
	LUT4 #(
		.INIT('h2203)
	) name3 (
		\G64_reg/NET0131 ,
		\G85_reg/NET0131 ,
		\G8_pad ,
		\G90_reg/NET0131 ,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\G78_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w94_
	);
	LUT4 #(
		.INIT('h5455)
	) name5 (
		_w91_,
		_w92_,
		_w93_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\G3_pad ,
		\G90_reg/NET0131 ,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\G77_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w97_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name8 (
		_w92_,
		_w93_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\G45_reg/NET0131 ,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\G2_pad ,
		\G90_reg/NET0131 ,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\G76_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w101_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name12 (
		_w92_,
		_w93_,
		_w100_,
		_w101_,
		_w102_
	);
	LUT4 #(
		.INIT('h153f)
	) name13 (
		\G44_reg/NET0131 ,
		\G45_reg/NET0131 ,
		_w98_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\G0_pad ,
		\G90_reg/NET0131 ,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\G74_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w105_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name16 (
		_w92_,
		_w93_,
		_w104_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\G1_pad ,
		\G90_reg/NET0131 ,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\G75_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w108_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name19 (
		_w92_,
		_w93_,
		_w107_,
		_w108_,
		_w109_
	);
	LUT4 #(
		.INIT('h135f)
	) name20 (
		\G42_reg/NET0131 ,
		\G43_reg/NET0131 ,
		_w106_,
		_w109_,
		_w110_
	);
	LUT4 #(
		.INIT('hfca8)
	) name21 (
		\G43_reg/NET0131 ,
		\G44_reg/NET0131 ,
		_w102_,
		_w109_,
		_w111_
	);
	LUT4 #(
		.INIT('h1511)
	) name22 (
		_w99_,
		_w103_,
		_w110_,
		_w111_,
		_w112_
	);
	LUT3 #(
		.INIT('he8)
	) name23 (
		\G46_reg/NET0131 ,
		_w95_,
		_w112_,
		_w113_
	);
	LUT4 #(
		.INIT('h0040)
	) name24 (
		\G24_reg/NET0131 ,
		\G25_reg/NET0131 ,
		\G26_reg/NET0131 ,
		\G27_reg/NET0131 ,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\G28_reg/NET0131 ,
		_w114_,
		_w115_
	);
	LUT4 #(
		.INIT('h1700)
	) name26 (
		\G46_reg/NET0131 ,
		_w95_,
		_w112_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		\G29_reg/NET0131 ,
		\G30_reg/NET0131 ,
		_w117_
	);
	LUT4 #(
		.INIT('h0080)
	) name28 (
		\G31_reg/NET0131 ,
		\G32_reg/NET0131 ,
		\G33_reg/NET0131 ,
		\G34_reg/NET0131 ,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w117_,
		_w118_,
		_w119_
	);
	LUT3 #(
		.INIT('h2a)
	) name30 (
		\G92_reg/NET0131 ,
		_w116_,
		_w119_,
		_w120_
	);
	LUT4 #(
		.INIT('h0001)
	) name31 (
		\G79_reg/NET0131 ,
		\G80_reg/NET0131 ,
		\G81_reg/NET0131 ,
		\G82_reg/NET0131 ,
		_w121_
	);
	LUT4 #(
		.INIT('h8421)
	) name32 (
		\G74_reg/NET0131 ,
		\G77_reg/NET0131 ,
		\G79_reg/NET0131 ,
		\G82_reg/NET0131 ,
		_w122_
	);
	LUT4 #(
		.INIT('h8421)
	) name33 (
		\G75_reg/NET0131 ,
		\G76_reg/NET0131 ,
		\G80_reg/NET0131 ,
		\G81_reg/NET0131 ,
		_w123_
	);
	LUT4 #(
		.INIT('h9000)
	) name34 (
		\G78_reg/NET0131 ,
		_w121_,
		_w122_,
		_w123_,
		_w124_
	);
	LUT3 #(
		.INIT('h02)
	) name35 (
		\G16_pad ,
		\G66_reg/NET0131 ,
		\G83_reg/NET0131 ,
		_w125_
	);
	LUT3 #(
		.INIT('h2a)
	) name36 (
		\G90_reg/NET0131 ,
		_w124_,
		_w125_,
		_w126_
	);
	LUT4 #(
		.INIT('h00d5)
	) name37 (
		\G92_reg/NET0131 ,
		_w116_,
		_w119_,
		_w126_,
		_w127_
	);
	LUT4 #(
		.INIT('h0888)
	) name38 (
		\G91_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w116_,
		_w119_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		\G36_reg/NET0131 ,
		\G37_reg/NET0131 ,
		_w129_
	);
	LUT4 #(
		.INIT('h0888)
	) name40 (
		\G38_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w124_,
		_w125_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT3 #(
		.INIT('h10)
	) name42 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w132_
	);
	LUT4 #(
		.INIT('hef00)
	) name43 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w133_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\G58_reg/NET0131 ,
		_w133_,
		_w134_
	);
	LUT3 #(
		.INIT('h80)
	) name45 (
		_w129_,
		_w130_,
		_w134_,
		_w135_
	);
	LUT4 #(
		.INIT('h7077)
	) name46 (
		\G58_reg/NET0131 ,
		_w127_,
		_w128_,
		_w135_,
		_w136_
	);
	LUT3 #(
		.INIT('hc4)
	) name47 (
		\G59_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\G53_reg/NET0131 ,
		\G61_reg/NET0131 ,
		_w138_
	);
	LUT3 #(
		.INIT('h80)
	) name49 (
		\G53_reg/NET0131 ,
		\G61_reg/NET0131 ,
		\G62_reg/NET0131 ,
		_w139_
	);
	LUT4 #(
		.INIT('h3b00)
	) name50 (
		\G59_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w136_,
		_w139_,
		_w140_
	);
	LUT4 #(
		.INIT('hd500)
	) name51 (
		\G92_reg/NET0131 ,
		_w116_,
		_w119_,
		_w132_,
		_w141_
	);
	LUT3 #(
		.INIT('hd0)
	) name52 (
		\G92_reg/NET0131 ,
		_w116_,
		_w119_,
		_w142_
	);
	LUT4 #(
		.INIT('ha200)
	) name53 (
		\G87_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w116_,
		_w119_,
		_w143_
	);
	LUT3 #(
		.INIT('h45)
	) name54 (
		\G90_reg/NET0131 ,
		\G94_reg/NET0131 ,
		_w116_,
		_w144_
	);
	LUT4 #(
		.INIT('h0700)
	) name55 (
		\G88_reg/NET0131 ,
		_w141_,
		_w143_,
		_w144_,
		_w145_
	);
	LUT3 #(
		.INIT('h70)
	) name56 (
		\G89_reg/NET0131 ,
		_w140_,
		_w145_,
		_w146_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name57 (
		\G67_reg/NET0131 ,
		\G68_reg/NET0131 ,
		\G71_reg/NET0131 ,
		\G72_reg/NET0131 ,
		_w147_
	);
	LUT2 #(
		.INIT('h9)
	) name58 (
		\G69_reg/NET0131 ,
		\G73_reg/NET0131 ,
		_w148_
	);
	LUT4 #(
		.INIT('haf23)
	) name59 (
		\G67_reg/NET0131 ,
		\G68_reg/NET0131 ,
		\G71_reg/NET0131 ,
		\G72_reg/NET0131 ,
		_w149_
	);
	LUT4 #(
		.INIT('h5556)
	) name60 (
		\G70_reg/NET0131 ,
		\G71_reg/NET0131 ,
		\G72_reg/NET0131 ,
		\G73_reg/NET0131 ,
		_w150_
	);
	LUT4 #(
		.INIT('h8000)
	) name61 (
		_w147_,
		_w148_,
		_w149_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\G14_pad ,
		_w151_,
		_w152_
	);
	LUT3 #(
		.INIT('h31)
	) name63 (
		\G14_pad ,
		\G90_reg/NET0131 ,
		_w151_,
		_w153_
	);
	LUT4 #(
		.INIT('h3b00)
	) name64 (
		\G59_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w136_,
		_w138_,
		_w154_
	);
	LUT4 #(
		.INIT('h8288)
	) name65 (
		\G14_pad ,
		\G62_reg/NET0131 ,
		_w137_,
		_w138_,
		_w155_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name66 (
		\G53_reg/NET0131 ,
		\G59_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w136_,
		_w156_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name67 (
		\G51_reg/NET0131 ,
		\G59_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w136_,
		_w157_
	);
	LUT4 #(
		.INIT('ha565)
	) name68 (
		\G51_reg/NET0131 ,
		\G59_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w136_,
		_w158_
	);
	LUT3 #(
		.INIT('h20)
	) name69 (
		\G14_pad ,
		_w156_,
		_w158_,
		_w159_
	);
	LUT4 #(
		.INIT('h002a)
	) name70 (
		\G14_pad ,
		\G52_reg/NET0131 ,
		_w157_,
		_w156_,
		_w160_
	);
	LUT4 #(
		.INIT('h0028)
	) name71 (
		\G14_pad ,
		\G52_reg/NET0131 ,
		_w157_,
		_w156_,
		_w161_
	);
	LUT4 #(
		.INIT('h5010)
	) name72 (
		\G38_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w129_,
		_w141_,
		_w162_
	);
	LUT3 #(
		.INIT('hd0)
	) name73 (
		\G92_reg/NET0131 ,
		_w116_,
		_w117_,
		_w163_
	);
	LUT4 #(
		.INIT('ha200)
	) name74 (
		\G31_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w116_,
		_w117_,
		_w164_
	);
	LUT3 #(
		.INIT('h80)
	) name75 (
		\G32_reg/NET0131 ,
		\G33_reg/NET0131 ,
		\G34_reg/NET0131 ,
		_w165_
	);
	LUT4 #(
		.INIT('hc444)
	) name76 (
		\G90_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w124_,
		_w125_,
		_w166_
	);
	LUT4 #(
		.INIT('h4055)
	) name77 (
		_w124_,
		_w164_,
		_w165_,
		_w166_,
		_w167_
	);
	LUT3 #(
		.INIT('hd0)
	) name78 (
		_w126_,
		_w162_,
		_w167_,
		_w168_
	);
	LUT4 #(
		.INIT('h038b)
	) name79 (
		\G14_pad ,
		\G90_reg/NET0131 ,
		\G9_pad ,
		_w151_,
		_w169_
	);
	LUT4 #(
		.INIT('ha200)
	) name80 (
		\G74_reg/NET0131 ,
		_w126_,
		_w162_,
		_w167_,
		_w170_
	);
	LUT3 #(
		.INIT('h48)
	) name81 (
		\G74_reg/NET0131 ,
		_w169_,
		_w168_,
		_w171_
	);
	LUT4 #(
		.INIT('h0323)
	) name82 (
		\G91_reg/NET0131 ,
		_w127_,
		_w131_,
		_w141_,
		_w172_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\G57_reg/NET0131 ,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\G14_pad ,
		_w136_,
		_w174_
	);
	LUT3 #(
		.INIT('h48)
	) name85 (
		\G58_reg/NET0131 ,
		_w174_,
		_w173_,
		_w175_
	);
	LUT4 #(
		.INIT('h8020)
	) name86 (
		\G14_pad ,
		\G57_reg/NET0131 ,
		_w136_,
		_w172_,
		_w176_
	);
	LUT3 #(
		.INIT('h82)
	) name87 (
		\G14_pad ,
		\G59_reg/NET0131 ,
		_w136_,
		_w177_
	);
	LUT4 #(
		.INIT('ha565)
	) name88 (
		\G38_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w129_,
		_w141_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\G14_pad ,
		_w178_,
		_w179_
	);
	LUT4 #(
		.INIT('h2232)
	) name90 (
		\G36_reg/NET0131 ,
		\G37_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w141_,
		_w180_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name91 (
		\G14_pad ,
		\G91_reg/NET0131 ,
		_w129_,
		_w141_,
		_w181_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w180_,
		_w181_,
		_w182_
	);
	LUT4 #(
		.INIT('h2282)
	) name93 (
		\G14_pad ,
		\G36_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w141_,
		_w183_
	);
	LUT4 #(
		.INIT('h5111)
	) name94 (
		\G39_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w116_,
		_w119_,
		_w184_
	);
	LUT3 #(
		.INIT('h23)
	) name95 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		\G14_pad ,
		_w141_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT3 #(
		.INIT('h28)
	) name98 (
		\G14_pad ,
		\G40_reg/NET0131 ,
		_w184_,
		_w188_
	);
	LUT4 #(
		.INIT('ha222)
	) name99 (
		\G39_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w116_,
		_w119_,
		_w189_
	);
	LUT4 #(
		.INIT('h1050)
	) name100 (
		\G47_reg/NET0131 ,
		\G56_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w189_,
		_w190_
	);
	LUT4 #(
		.INIT('h4505)
	) name101 (
		\G12_pad ,
		\G56_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w189_,
		_w191_
	);
	LUT3 #(
		.INIT('h02)
	) name102 (
		\G14_pad ,
		_w191_,
		_w190_,
		_w192_
	);
	LUT4 #(
		.INIT('h1050)
	) name103 (
		\G49_reg/NET0131 ,
		\G56_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w189_,
		_w193_
	);
	LUT4 #(
		.INIT('h4505)
	) name104 (
		\G48_reg/NET0131 ,
		\G56_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w189_,
		_w194_
	);
	LUT3 #(
		.INIT('h02)
	) name105 (
		\G14_pad ,
		_w194_,
		_w193_,
		_w195_
	);
	LUT4 #(
		.INIT('h1050)
	) name106 (
		\G48_reg/NET0131 ,
		\G56_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w189_,
		_w196_
	);
	LUT4 #(
		.INIT('h4505)
	) name107 (
		\G47_reg/NET0131 ,
		\G56_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w189_,
		_w197_
	);
	LUT3 #(
		.INIT('h02)
	) name108 (
		\G14_pad ,
		_w197_,
		_w196_,
		_w198_
	);
	LUT4 #(
		.INIT('h1050)
	) name109 (
		\G50_reg/NET0131 ,
		\G56_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w189_,
		_w199_
	);
	LUT4 #(
		.INIT('h4505)
	) name110 (
		\G49_reg/NET0131 ,
		\G56_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w189_,
		_w200_
	);
	LUT3 #(
		.INIT('h02)
	) name111 (
		\G14_pad ,
		_w200_,
		_w199_,
		_w201_
	);
	LUT4 #(
		.INIT('h08a0)
	) name112 (
		\G14_pad ,
		\G55_reg/NET0131 ,
		\G56_reg/NET0131 ,
		_w189_,
		_w202_
	);
	LUT4 #(
		.INIT('h0288)
	) name113 (
		\G14_pad ,
		\G55_reg/NET0131 ,
		\G56_reg/NET0131 ,
		_w189_,
		_w203_
	);
	LUT3 #(
		.INIT('h82)
	) name114 (
		\G14_pad ,
		\G39_reg/NET0131 ,
		_w120_,
		_w204_
	);
	LUT4 #(
		.INIT('h70f0)
	) name115 (
		\G32_reg/NET0131 ,
		\G33_reg/NET0131 ,
		\G34_reg/NET0131 ,
		_w164_,
		_w205_
	);
	LUT3 #(
		.INIT('ha8)
	) name116 (
		\G14_pad ,
		_w142_,
		_w205_,
		_w206_
	);
	LUT4 #(
		.INIT('h28a0)
	) name117 (
		\G14_pad ,
		\G32_reg/NET0131 ,
		\G33_reg/NET0131 ,
		_w164_,
		_w207_
	);
	LUT4 #(
		.INIT('h2232)
	) name118 (
		\G29_reg/NET0131 ,
		\G30_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w116_,
		_w208_
	);
	LUT4 #(
		.INIT('h08aa)
	) name119 (
		\G14_pad ,
		\G92_reg/NET0131 ,
		_w116_,
		_w117_,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w208_,
		_w209_,
		_w210_
	);
	LUT3 #(
		.INIT('h28)
	) name121 (
		\G14_pad ,
		\G32_reg/NET0131 ,
		_w164_,
		_w211_
	);
	LUT4 #(
		.INIT('h2282)
	) name122 (
		\G14_pad ,
		\G29_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w116_,
		_w212_
	);
	LUT3 #(
		.INIT('h28)
	) name123 (
		\G14_pad ,
		\G31_reg/NET0131 ,
		_w163_,
		_w213_
	);
	LUT4 #(
		.INIT('h1700)
	) name124 (
		\G46_reg/NET0131 ,
		_w95_,
		_w112_,
		_w114_,
		_w214_
	);
	LUT4 #(
		.INIT('h8288)
	) name125 (
		\G14_pad ,
		\G28_reg/NET0131 ,
		_w113_,
		_w114_,
		_w215_
	);
	LUT4 #(
		.INIT('h0115)
	) name126 (
		\G24_reg/NET0131 ,
		\G46_reg/NET0131 ,
		_w95_,
		_w112_,
		_w216_
	);
	LUT4 #(
		.INIT('h70f0)
	) name127 (
		\G25_reg/NET0131 ,
		\G26_reg/NET0131 ,
		\G27_reg/NET0131 ,
		_w216_,
		_w217_
	);
	LUT3 #(
		.INIT('ha8)
	) name128 (
		\G14_pad ,
		_w214_,
		_w217_,
		_w218_
	);
	LUT3 #(
		.INIT('h28)
	) name129 (
		\G14_pad ,
		\G25_reg/NET0131 ,
		_w216_,
		_w219_
	);
	LUT4 #(
		.INIT('h28a0)
	) name130 (
		\G14_pad ,
		\G25_reg/NET0131 ,
		\G26_reg/NET0131 ,
		_w216_,
		_w220_
	);
	LUT4 #(
		.INIT('h566a)
	) name131 (
		\G24_reg/NET0131 ,
		\G46_reg/NET0131 ,
		_w95_,
		_w112_,
		_w221_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		\G14_pad ,
		_w221_,
		_w222_
	);
	LUT4 #(
		.INIT('he222)
	) name133 (
		\G6_pad ,
		\G90_reg/NET0131 ,
		_w124_,
		_w125_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		\G5_pad ,
		\G90_reg/NET0131 ,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		\G83_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w225_
	);
	LUT3 #(
		.INIT('h13)
	) name136 (
		_w124_,
		_w224_,
		_w225_,
		_w226_
	);
	LUT4 #(
		.INIT('hfca8)
	) name137 (
		\G45_reg/NET0131 ,
		\G46_reg/NET0131 ,
		_w95_,
		_w98_,
		_w227_
	);
	LUT4 #(
		.INIT('h3f2a)
	) name138 (
		\G42_reg/NET0131 ,
		\G46_reg/NET0131 ,
		_w95_,
		_w106_,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w227_,
		_w228_,
		_w229_
	);
	LUT3 #(
		.INIT('h80)
	) name140 (
		_w103_,
		_w110_,
		_w111_,
		_w230_
	);
	LUT3 #(
		.INIT('h5c)
	) name141 (
		\G34_reg/NET0131 ,
		\G35_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w231_
	);
	LUT4 #(
		.INIT('hd500)
	) name142 (
		\G90_reg/NET0131 ,
		_w124_,
		_w125_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w130_,
		_w232_,
		_w233_
	);
	LUT4 #(
		.INIT('h00ea)
	) name144 (
		_w226_,
		_w229_,
		_w230_,
		_w233_,
		_w234_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name145 (
		\G59_reg/NET0131 ,
		\G62_reg/NET0131 ,
		\G90_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		\G35_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		_w235_,
		_w236_,
		_w237_
	);
	LUT3 #(
		.INIT('h2a)
	) name148 (
		\G14_pad ,
		_w223_,
		_w237_,
		_w238_
	);
	LUT4 #(
		.INIT('hcd00)
	) name149 (
		_w113_,
		_w223_,
		_w234_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\G15_pad ,
		\G22_reg/NET0131 ,
		_w240_
	);
	LUT3 #(
		.INIT('hd8)
	) name151 (
		\G15_pad ,
		\G22_reg/NET0131 ,
		\G23_reg/NET0131 ,
		_w241_
	);
	LUT4 #(
		.INIT('h8000)
	) name152 (
		\G47_reg/NET0131 ,
		\G48_reg/NET0131 ,
		\G49_reg/NET0131 ,
		\G50_reg/NET0131 ,
		_w242_
	);
	LUT4 #(
		.INIT('h0800)
	) name153 (
		\G42_reg/NET0131 ,
		\G43_reg/NET0131 ,
		_w241_,
		_w242_,
		_w243_
	);
	LUT3 #(
		.INIT('h80)
	) name154 (
		\G44_reg/NET0131 ,
		\G45_reg/NET0131 ,
		_w243_,
		_w244_
	);
	LUT4 #(
		.INIT('h03a3)
	) name155 (
		\G14_pad ,
		\G7_pad ,
		\G90_reg/NET0131 ,
		_w151_,
		_w245_
	);
	LUT3 #(
		.INIT('h48)
	) name156 (
		\G46_reg/NET0131 ,
		_w245_,
		_w244_,
		_w246_
	);
	LUT4 #(
		.INIT('haaa8)
	) name157 (
		\G14_pad ,
		\G63_reg/NET0131 ,
		_w130_,
		_w232_,
		_w247_
	);
	LUT3 #(
		.INIT('h6c)
	) name158 (
		\G44_reg/NET0131 ,
		\G45_reg/NET0131 ,
		_w243_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w245_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\G14_pad ,
		\G83_reg/NET0131 ,
		_w250_
	);
	LUT3 #(
		.INIT('h10)
	) name161 (
		_w92_,
		_w93_,
		_w250_,
		_w251_
	);
	LUT3 #(
		.INIT('he0)
	) name162 (
		_w130_,
		_w232_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h6)
	) name163 (
		\G44_reg/NET0131 ,
		_w243_,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w245_,
		_w253_,
		_w254_
	);
	LUT3 #(
		.INIT('h9a)
	) name165 (
		\G42_reg/NET0131 ,
		_w241_,
		_w242_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		_w245_,
		_w255_,
		_w256_
	);
	LUT4 #(
		.INIT('hc6cc)
	) name167 (
		\G42_reg/NET0131 ,
		\G43_reg/NET0131 ,
		_w241_,
		_w242_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w245_,
		_w257_,
		_w258_
	);
	LUT4 #(
		.INIT('h88a0)
	) name169 (
		\G14_pad ,
		\G63_reg/NET0131 ,
		\G64_reg/NET0131 ,
		_w151_,
		_w259_
	);
	LUT4 #(
		.INIT('h88a0)
	) name170 (
		\G14_pad ,
		\G65_reg/NET0131 ,
		\G66_reg/NET0131 ,
		_w151_,
		_w260_
	);
	LUT3 #(
		.INIT('hd5)
	) name171 (
		\G14_pad ,
		\G90_reg/NET0131 ,
		_w151_,
		_w261_
	);
	LUT3 #(
		.INIT('hd5)
	) name172 (
		\G14_pad ,
		\G91_reg/NET0131 ,
		_w151_,
		_w262_
	);
	LUT3 #(
		.INIT('ha8)
	) name173 (
		\G14_pad ,
		\G65_reg/NET0131 ,
		_w151_,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\G13_pad ,
		\G14_pad ,
		_w264_
	);
	LUT3 #(
		.INIT('hc8)
	) name175 (
		\G10_pad ,
		\G86_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w265_
	);
	LUT2 #(
		.INIT('hd)
	) name176 (
		_w264_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		_w240_,
		_w242_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\G15_pad ,
		\G47_reg/NET0131 ,
		_w268_
	);
	LUT3 #(
		.INIT('h01)
	) name179 (
		\G48_reg/NET0131 ,
		\G49_reg/NET0131 ,
		\G50_reg/NET0131 ,
		_w269_
	);
	LUT3 #(
		.INIT('h2a)
	) name180 (
		\G22_reg/NET0131 ,
		_w268_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('he)
	) name181 (
		_w267_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		\G10_pad ,
		\G92_reg/NET0131 ,
		_w272_
	);
	LUT4 #(
		.INIT('hf351)
	) name183 (
		\G10_pad ,
		\G13_pad ,
		\G86_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w273_
	);
	LUT3 #(
		.INIT('h75)
	) name184 (
		_w264_,
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\G10_pad ,
		\G90_reg/NET0131 ,
		_w275_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name186 (
		\G10_pad ,
		\G13_pad ,
		\G86_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w276_
	);
	LUT3 #(
		.INIT('h75)
	) name187 (
		_w264_,
		_w275_,
		_w276_,
		_w277_
	);
	LUT4 #(
		.INIT('h40c8)
	) name188 (
		\G11_pad ,
		\G14_pad ,
		\G87_reg/NET0131 ,
		\G94_reg/NET0131 ,
		_w278_
	);
	LUT4 #(
		.INIT('hc480)
	) name189 (
		\G11_pad ,
		\G14_pad ,
		\G87_reg/NET0131 ,
		\G88_reg/NET0131 ,
		_w279_
	);
	LUT4 #(
		.INIT('hc480)
	) name190 (
		\G11_pad ,
		\G14_pad ,
		\G88_reg/NET0131 ,
		\G89_reg/NET0131 ,
		_w280_
	);
	LUT4 #(
		.INIT('h4c08)
	) name191 (
		\G11_pad ,
		\G14_pad ,
		\G89_reg/NET0131 ,
		\G94_reg/NET0131 ,
		_w281_
	);
	LUT3 #(
		.INIT('hca)
	) name192 (
		\G1_pad ,
		\G4_pad ,
		\G63_reg/NET0131 ,
		_w282_
	);
	LUT3 #(
		.INIT('hca)
	) name193 (
		\G0_pad ,
		\G3_pad ,
		\G63_reg/NET0131 ,
		_w283_
	);
	LUT3 #(
		.INIT('hca)
	) name194 (
		\G2_pad ,
		\G5_pad ,
		\G63_reg/NET0131 ,
		_w284_
	);
	LUT2 #(
		.INIT('h2)
	) name195 (
		\G14_pad ,
		\G35_reg/NET0131 ,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\G74_reg/NET0131 ,
		\G75_reg/NET0131 ,
		_w286_
	);
	LUT4 #(
		.INIT('hd000)
	) name197 (
		_w126_,
		_w162_,
		_w167_,
		_w286_,
		_w287_
	);
	LUT3 #(
		.INIT('h80)
	) name198 (
		\G76_reg/NET0131 ,
		\G77_reg/NET0131 ,
		_w287_,
		_w288_
	);
	LUT3 #(
		.INIT('h48)
	) name199 (
		\G78_reg/NET0131 ,
		_w169_,
		_w288_,
		_w289_
	);
	LUT4 #(
		.INIT('h00c8)
	) name200 (
		\G75_reg/NET0131 ,
		_w169_,
		_w170_,
		_w287_,
		_w290_
	);
	LUT4 #(
		.INIT('haaa2)
	) name201 (
		\G83_reg/NET0131 ,
		_w124_,
		_w130_,
		_w232_,
		_w291_
	);
	LUT4 #(
		.INIT('h002f)
	) name202 (
		_w126_,
		_w162_,
		_w167_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		_w169_,
		_w292_,
		_w293_
	);
	LUT4 #(
		.INIT('h60c0)
	) name204 (
		\G76_reg/NET0131 ,
		\G77_reg/NET0131 ,
		_w169_,
		_w287_,
		_w294_
	);
	LUT4 #(
		.INIT('h7f00)
	) name205 (
		\G53_reg/NET0131 ,
		\G61_reg/NET0131 ,
		\G62_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w295_
	);
	LUT4 #(
		.INIT('hccc4)
	) name206 (
		\G59_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w136_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\G67_reg/NET0131 ,
		\G68_reg/NET0131 ,
		_w297_
	);
	LUT4 #(
		.INIT('hc060)
	) name208 (
		\G67_reg/NET0131 ,
		\G68_reg/NET0131 ,
		_w152_,
		_w296_,
		_w298_
	);
	LUT2 #(
		.INIT('h2)
	) name209 (
		\G14_pad ,
		_w154_,
		_w299_
	);
	LUT4 #(
		.INIT('h0208)
	) name210 (
		\G14_pad ,
		\G60_reg/NET0131 ,
		_w154_,
		_w156_,
		_w300_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\G14_pad ,
		\G53_reg/NET0131 ,
		_w301_
	);
	LUT3 #(
		.INIT('h80)
	) name212 (
		\G52_reg/NET0131 ,
		_w157_,
		_w301_,
		_w302_
	);
	LUT3 #(
		.INIT('hf8)
	) name213 (
		\G53_reg/NET0131 ,
		_w160_,
		_w302_,
		_w303_
	);
	LUT3 #(
		.INIT('h13)
	) name214 (
		\G60_reg/NET0131 ,
		\G61_reg/NET0131 ,
		_w156_,
		_w304_
	);
	LUT2 #(
		.INIT('h2)
	) name215 (
		_w299_,
		_w304_,
		_w305_
	);
	LUT3 #(
		.INIT('h48)
	) name216 (
		\G76_reg/NET0131 ,
		_w169_,
		_w287_,
		_w306_
	);
	LUT3 #(
		.INIT('h84)
	) name217 (
		\G67_reg/NET0131 ,
		_w152_,
		_w296_,
		_w307_
	);
	LUT3 #(
		.INIT('h20)
	) name218 (
		\G69_reg/NET0131 ,
		_w296_,
		_w297_,
		_w308_
	);
	LUT4 #(
		.INIT('h8488)
	) name219 (
		\G69_reg/NET0131 ,
		_w152_,
		_w296_,
		_w297_,
		_w309_
	);
	LUT3 #(
		.INIT('h48)
	) name220 (
		\G70_reg/NET0131 ,
		_w152_,
		_w308_,
		_w310_
	);
	assign \G701BF_pad  = _w9_ ;
	assign \G702_pad  = _w146_ ;
	assign \G727_pad  = _w153_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g2503/_0_  = _w155_ ;
	assign \g2514/_0_  = _w159_ ;
	assign \g2516/_0_  = _w161_ ;
	assign \g2542/_0_  = _w171_ ;
	assign \g2549/_0_  = _w175_ ;
	assign \g2553/_0_  = _w176_ ;
	assign \g2554/_0_  = _w177_ ;
	assign \g2570/_0_  = _w179_ ;
	assign \g2574/_0_  = _w182_ ;
	assign \g2576/_0_  = _w183_ ;
	assign \g2583/_0_  = _w187_ ;
	assign \g2588/_0_  = _w188_ ;
	assign \g2602/_0_  = _w192_ ;
	assign \g2603/_0_  = _w195_ ;
	assign \g2604/_0_  = _w198_ ;
	assign \g2605/_0_  = _w201_ ;
	assign \g2611/_0_  = _w202_ ;
	assign \g2614/_0_  = _w203_ ;
	assign \g2615/_0_  = _w204_ ;
	assign \g2644/_0_  = _w206_ ;
	assign \g2657/_0_  = _w207_ ;
	assign \g2663/_0_  = _w210_ ;
	assign \g2664/_0_  = _w211_ ;
	assign \g2666/_0_  = _w212_ ;
	assign \g2672/_0_  = _w213_ ;
	assign \g2678/_0_  = _w215_ ;
	assign \g2681/_0_  = _w218_ ;
	assign \g2696/_00_  = _w219_ ;
	assign \g2698/_0_  = _w220_ ;
	assign \g2699/_0_  = _w222_ ;
	assign \g2700/_00_  = _w239_ ;
	assign \g2717/_0_  = _w246_ ;
	assign \g2719/_0_  = _w247_ ;
	assign \g2723/_0_  = _w249_ ;
	assign \g2726/_3_  = _w252_ ;
	assign \g2735/_0_  = _w254_ ;
	assign \g2737/_0_  = _w256_ ;
	assign \g2740/_0_  = _w258_ ;
	assign \g2785/_0_  = _w259_ ;
	assign \g2786/_0_  = _w260_ ;
	assign \g2787/_1__syn_2  = _w261_ ;
	assign \g2790/_1__syn_2  = _w262_ ;
	assign \g2798/_2_  = _w241_ ;
	assign \g2801/_0_  = _w263_ ;
	assign \g2841/_0_  = _w266_ ;
	assign \g2844/_0_  = _w271_ ;
	assign \g2845/_0_  = _w274_ ;
	assign \g2846/_0_  = _w277_ ;
	assign \g2860/_0_  = _w278_ ;
	assign \g2861/_0_  = _w279_ ;
	assign \g2862/_0_  = _w280_ ;
	assign \g2864/_0_  = _w281_ ;
	assign \g2882/_3_  = _w282_ ;
	assign \g2883/_3_  = _w283_ ;
	assign \g2887/_3_  = _w284_ ;
	assign \g2906/_0_  = _w285_ ;
	assign \g2911/_0_  = _w264_ ;
	assign \g3282/_0_  = _w289_ ;
	assign \g3406/_0_  = _w290_ ;
	assign \g3409/_0_  = _w293_ ;
	assign \g3506/_0_  = _w294_ ;
	assign \g3685/_3_  = _w298_ ;
	assign \g3694/_0_  = _w300_ ;
	assign \g3743/_0_  = _w303_ ;
	assign \g3753/_0_  = _w305_ ;
	assign \g3785/_0_  = _w306_ ;
	assign \g3835/_0_  = _w307_ ;
	assign \g3946/_2_  = _w309_ ;
	assign \g3976/_0_  = _w310_ ;
endmodule;