module top (\B_reg/NET0131 , \IR_reg[0]/NET0131 , \IR_reg[10]/NET0131 , \IR_reg[11]/NET0131 , \IR_reg[12]/NET0131 , \IR_reg[13]/NET0131 , \IR_reg[14]/NET0131 , \IR_reg[15]/NET0131 , \IR_reg[16]/NET0131 , \IR_reg[17]/NET0131 , \IR_reg[18]/NET0131 , \IR_reg[19]/NET0131 , \IR_reg[1]/NET0131 , \IR_reg[20]/NET0131 , \IR_reg[21]/NET0131 , \IR_reg[22]/NET0131 , \IR_reg[23]/NET0131 , \IR_reg[24]/NET0131 , \IR_reg[25]/NET0131 , \IR_reg[26]/NET0131 , \IR_reg[27]/NET0131 , \IR_reg[28]/NET0131 , \IR_reg[29]/NET0131 , \IR_reg[2]/NET0131 , \IR_reg[30]/NET0131 , \IR_reg[31]/NET0131 , \IR_reg[3]/NET0131 , \IR_reg[4]/NET0131 , \IR_reg[5]/NET0131 , \IR_reg[6]/NET0131 , \IR_reg[7]/NET0131 , \IR_reg[8]/NET0131 , \IR_reg[9]/NET0131 , \addr[0]_pad , \addr[10]_pad , \addr[11]_pad , \addr[12]_pad , \addr[13]_pad , \addr[14]_pad , \addr[15]_pad , \addr[16]_pad , \addr[17]_pad , \addr[18]_pad , \addr[19]_pad , \addr[1]_pad , \addr[2]_pad , \addr[3]_pad , \addr[4]_pad , \addr[5]_pad , \addr[6]_pad , \addr[7]_pad , \addr[8]_pad , \addr[9]_pad , \d_reg[0]/NET0131 , \d_reg[1]/NET0131 , \datai[0]_pad , \datai[10]_pad , \datai[11]_pad , \datai[12]_pad , \datai[13]_pad , \datai[14]_pad , \datai[15]_pad , \datai[16]_pad , \datai[17]_pad , \datai[18]_pad , \datai[19]_pad , \datai[1]_pad , \datai[20]_pad , \datai[21]_pad , \datai[22]_pad , \datai[23]_pad , \datai[24]_pad , \datai[25]_pad , \datai[26]_pad , \datai[27]_pad , \datai[28]_pad , \datai[29]_pad , \datai[2]_pad , \datai[30]_pad , \datai[31]_pad , \datai[3]_pad , \datai[4]_pad , \datai[5]_pad , \datai[6]_pad , \datai[7]_pad , \datai[8]_pad , \datai[9]_pad , \datao[15]_pad , \datao[28]_pad , \datao[8]_pad , \reg0_reg[0]/NET0131 , \reg0_reg[10]/NET0131 , \reg0_reg[11]/NET0131 , \reg0_reg[12]/NET0131 , \reg0_reg[13]/NET0131 , \reg0_reg[14]/NET0131 , \reg0_reg[15]/NET0131 , \reg0_reg[16]/NET0131 , \reg0_reg[17]/NET0131 , \reg0_reg[18]/NET0131 , \reg0_reg[19]/NET0131 , \reg0_reg[1]/NET0131 , \reg0_reg[20]/NET0131 , \reg0_reg[21]/NET0131 , \reg0_reg[22]/NET0131 , \reg0_reg[23]/NET0131 , \reg0_reg[24]/NET0131 , \reg0_reg[25]/NET0131 , \reg0_reg[26]/NET0131 , \reg0_reg[27]/NET0131 , \reg0_reg[28]/NET0131 , \reg0_reg[29]/NET0131 , \reg0_reg[2]/NET0131 , \reg0_reg[30]/NET0131 , \reg0_reg[31]/NET0131 , \reg0_reg[3]/NET0131 , \reg0_reg[4]/NET0131 , \reg0_reg[5]/NET0131 , \reg0_reg[6]/NET0131 , \reg0_reg[7]/NET0131 , \reg0_reg[8]/NET0131 , \reg0_reg[9]/NET0131 , \reg1_reg[0]/NET0131 , \reg1_reg[10]/NET0131 , \reg1_reg[11]/NET0131 , \reg1_reg[12]/NET0131 , \reg1_reg[13]/NET0131 , \reg1_reg[14]/NET0131 , \reg1_reg[15]/NET0131 , \reg1_reg[16]/NET0131 , \reg1_reg[17]/NET0131 , \reg1_reg[18]/NET0131 , \reg1_reg[19]/NET0131 , \reg1_reg[1]/NET0131 , \reg1_reg[20]/NET0131 , \reg1_reg[21]/NET0131 , \reg1_reg[22]/NET0131 , \reg1_reg[23]/NET0131 , \reg1_reg[24]/NET0131 , \reg1_reg[25]/NET0131 , \reg1_reg[26]/NET0131 , \reg1_reg[27]/NET0131 , \reg1_reg[28]/NET0131 , \reg1_reg[29]/NET0131 , \reg1_reg[2]/NET0131 , \reg1_reg[30]/NET0131 , \reg1_reg[31]/NET0131 , \reg1_reg[3]/NET0131 , \reg1_reg[4]/NET0131 , \reg1_reg[5]/NET0131 , \reg1_reg[6]/NET0131 , \reg1_reg[7]/NET0131 , \reg1_reg[8]/NET0131 , \reg1_reg[9]/NET0131 , \reg2_reg[0]/NET0131 , \reg2_reg[10]/NET0131 , \reg2_reg[11]/NET0131 , \reg2_reg[12]/NET0131 , \reg2_reg[13]/NET0131 , \reg2_reg[14]/NET0131 , \reg2_reg[15]/NET0131 , \reg2_reg[16]/NET0131 , \reg2_reg[17]/NET0131 , \reg2_reg[18]/NET0131 , \reg2_reg[19]/NET0131 , \reg2_reg[1]/NET0131 , \reg2_reg[20]/NET0131 , \reg2_reg[21]/NET0131 , \reg2_reg[22]/NET0131 , \reg2_reg[23]/NET0131 , \reg2_reg[24]/NET0131 , \reg2_reg[25]/NET0131 , \reg2_reg[26]/NET0131 , \reg2_reg[27]/NET0131 , \reg2_reg[28]/NET0131 , \reg2_reg[29]/NET0131 , \reg2_reg[2]/NET0131 , \reg2_reg[30]/NET0131 , \reg2_reg[31]/NET0131 , \reg2_reg[3]/NET0131 , \reg2_reg[4]/NET0131 , \reg2_reg[5]/NET0131 , \reg2_reg[6]/NET0131 , \reg2_reg[7]/NET0131 , \reg2_reg[8]/NET0131 , \reg2_reg[9]/NET0131 , \reg3_reg[0]/NET0131 , \reg3_reg[10]/NET0131 , \reg3_reg[11]/NET0131 , \reg3_reg[12]/NET0131 , \reg3_reg[13]/NET0131 , \reg3_reg[14]/NET0131 , \reg3_reg[15]/NET0131 , \reg3_reg[16]/NET0131 , \reg3_reg[17]/NET0131 , \reg3_reg[18]/NET0131 , \reg3_reg[19]/NET0131 , \reg3_reg[1]/NET0131 , \reg3_reg[20]/NET0131 , \reg3_reg[21]/NET0131 , \reg3_reg[22]/NET0131 , \reg3_reg[23]/NET0131 , \reg3_reg[24]/NET0131 , \reg3_reg[25]/NET0131 , \reg3_reg[26]/NET0131 , \reg3_reg[27]/NET0131 , \reg3_reg[28]/NET0131 , \reg3_reg[2]/NET0131 , \reg3_reg[3]/NET0131 , \reg3_reg[4]/NET0131 , \reg3_reg[5]/NET0131 , \reg3_reg[6]/NET0131 , \reg3_reg[7]/NET0131 , \reg3_reg[8]/NET0131 , \reg3_reg[9]/NET0131 , \state_reg[0]/NET0131 , \_al_n0 , \_al_n1 , \g22/_0_ , \g32_dup/_0_ , \g35904/_0_ , \g35905/_0_ , \g35906/_0_ , \g35907/_0_ , \g35908/_0_ , \g35909/_0_ , \g35910/_0_ , \g35911/_0_ , \g35932/_0_ , \g35955/_0_ , \g35956/_0_ , \g35957/_0_ , \g35962/_0_ , \g35967/_0_ , \g35968/_0_ , \g35971/_0_ , \g35972/_0_ , \g35973/_0_ , \g35974/_0_ , \g35975/_0_ , \g35976/_0_ , \g35977/_0_ , \g35978/_0_ , \g36015/_0_ , \g36016/_0_ , \g36018/_0_ , \g36022/_0_ , \g36023/_0_ , \g36025/_0_ , \g36029/_0_ , \g36030/_0_ , \g36031/_0_ , \g36032/_0_ , \g36033/_0_ , \g36034/_0_ , \g36035/_0_ , \g36036/_0_ , \g36038/_0_ , \g36039/_0_ , \g36040/_0_ , \g36041/_0_ , \g36073/_0_ , \g36087/_0_ , \g36091/_0_ , \g36092/_0_ , \g36093/_0_ , \g36094/_0_ , \g36096/_0_ , \g36097/_0_ , \g36098/_0_ , \g36099/_0_ , \g36100/_0_ , \g36101/_0_ , \g36102/_0_ , \g36103/_0_ , \g36104/_0_ , \g36105/_0_ , \g36106/_0_ , \g36107/_0_ , \g36108/_0_ , \g36109/_0_ , \g36110/_0_ , \g36111/_0_ , \g36112/_0_ , \g36113/_0_ , \g36165/_0_ , \g36169/_0_ , \g36170/_0_ , \g36171/_0_ , \g36172/_0_ , \g36198/_0_ , \g36199/_0_ , \g36200/_0_ , \g36201/_0_ , \g36202/_0_ , \g36203/_0_ , \g36205/_0_ , \g36206/_0_ , \g36207/_0_ , \g36208/_0_ , \g36209/_0_ , \g36240/_0_ , \g36281/_0_ , \g36282/_0_ , \g36283/_0_ , \g36284/_0_ , \g36285/_0_ , \g36286/_0_ , \g36287/_0_ , \g36288/_0_ , \g36289/_0_ , \g36290/_0_ , \g36291/_0_ , \g36292/_0_ , \g36293/_0_ , \g36294/_0_ , \g36295/_0_ , \g36296/_0_ , \g36297/_0_ , \g36298/_0_ , \g36330/_0_ , \g36385/_0_ , \g36390/_0_ , \g36391/_0_ , \g36392/_0_ , \g36393/_0_ , \g36394/_0_ , \g36470/_0_ , \g36471/_0_ , \g36472/_0_ , \g36473/_0_ , \g36474/_0_ , \g36475/_0_ , \g38/_0_ , \g38399/_0_ , \g38400/_0_ , \g39639/_0_ , \g39641/_0_ , \g39644/_0_ , \g39647/_0_ , \g39648/_0_ , \g39650/_0_ , \g39654/_0_ , \g39658/_0_ , \g39660/_0_ , \g39662/_0_ , \g39663/_0_ , \g39665/_0_ , \g39666/_0_ , \g39667/_0_ , \g39730/_0_ , \g39796/_0_ , \g39930/_0_ , \g39931/_0_ , \g39932/_0_ , \g40045/_0_ , \g40150/u3_syn_4 , \g40608/_0_ , \g41017/u3_syn_4 , \g42159/_0_ , \g42169/_0_ , \g42174/_0_ , \g42483/_0_ , \g42736/_0_ , \g42746/_0_ , \g42755/_0_ , \g42767/_0_ , \g42776/_0_ , \g42871_dup/_1_ , \g42908/_0_ , \g42938/_0_ , \g42969/_0_ , \g43022/_0_ , \g44035/_1__syn_2 , \g44227/_3_ , \g44260/_3_ , \g44261/_3_ , \g44262/_3_ , \g44311/_3_ , \g44378/_3_ , \g44379/_3_ , \g44383/_3_ , \g44384/_3_ , \g44385/_3_ , \g44386/_3_ , \g44390/_3_ , \g44391/_3_ , \g44492/_3_ , \g44493/_3_ , \g44494/_3_ , \g44495/_3_ , \g44496/_3_ , \g44497/_3_ , \g44498/_3_ , \g44499/_3_ , \g44575/_3_ , \g44589/_3_ , \g44596/_3_ , \g44615/_3_ , \g44795/_3_ , \g44803/_3_ , \g44804/_3_ , \g44888/_3_ , \g44889/_3_ , \g45004/_3_ , \g46129/_0_ , \g46133/_0_ , \g46265/_2_ , \g46313/_0_ , \g46372/_0_ , \g46377/_0_ , \g46399/_0_ , \g46405/_0_ , \g46427/_0_ , \g46461/_0_ , \g46526/_0_ , \g46576/_0_ , \g46608/_0_ , \g46697/_0_ , \g46778/_0_ , \g47007/_0_ , \g47023/_0_ , \g47077/_1_ , \g47097/_0_ , \g47109/_1_ , \g47142_dup/_1_ , \g47256/_0_ , \g47328/_0_ , \g47373/_0_ , \g47465/_0_ , \g47518/_0_ , \g47556/_1_ , \g56/_0_ , \state_reg[0]/NET0131_syn_2 );
	input \B_reg/NET0131  ;
	input \IR_reg[0]/NET0131  ;
	input \IR_reg[10]/NET0131  ;
	input \IR_reg[11]/NET0131  ;
	input \IR_reg[12]/NET0131  ;
	input \IR_reg[13]/NET0131  ;
	input \IR_reg[14]/NET0131  ;
	input \IR_reg[15]/NET0131  ;
	input \IR_reg[16]/NET0131  ;
	input \IR_reg[17]/NET0131  ;
	input \IR_reg[18]/NET0131  ;
	input \IR_reg[19]/NET0131  ;
	input \IR_reg[1]/NET0131  ;
	input \IR_reg[20]/NET0131  ;
	input \IR_reg[21]/NET0131  ;
	input \IR_reg[22]/NET0131  ;
	input \IR_reg[23]/NET0131  ;
	input \IR_reg[24]/NET0131  ;
	input \IR_reg[25]/NET0131  ;
	input \IR_reg[26]/NET0131  ;
	input \IR_reg[27]/NET0131  ;
	input \IR_reg[28]/NET0131  ;
	input \IR_reg[29]/NET0131  ;
	input \IR_reg[2]/NET0131  ;
	input \IR_reg[30]/NET0131  ;
	input \IR_reg[31]/NET0131  ;
	input \IR_reg[3]/NET0131  ;
	input \IR_reg[4]/NET0131  ;
	input \IR_reg[5]/NET0131  ;
	input \IR_reg[6]/NET0131  ;
	input \IR_reg[7]/NET0131  ;
	input \IR_reg[8]/NET0131  ;
	input \IR_reg[9]/NET0131  ;
	input \addr[0]_pad  ;
	input \addr[10]_pad  ;
	input \addr[11]_pad  ;
	input \addr[12]_pad  ;
	input \addr[13]_pad  ;
	input \addr[14]_pad  ;
	input \addr[15]_pad  ;
	input \addr[16]_pad  ;
	input \addr[17]_pad  ;
	input \addr[18]_pad  ;
	input \addr[19]_pad  ;
	input \addr[1]_pad  ;
	input \addr[2]_pad  ;
	input \addr[3]_pad  ;
	input \addr[4]_pad  ;
	input \addr[5]_pad  ;
	input \addr[6]_pad  ;
	input \addr[7]_pad  ;
	input \addr[8]_pad  ;
	input \addr[9]_pad  ;
	input \d_reg[0]/NET0131  ;
	input \d_reg[1]/NET0131  ;
	input \datai[0]_pad  ;
	input \datai[10]_pad  ;
	input \datai[11]_pad  ;
	input \datai[12]_pad  ;
	input \datai[13]_pad  ;
	input \datai[14]_pad  ;
	input \datai[15]_pad  ;
	input \datai[16]_pad  ;
	input \datai[17]_pad  ;
	input \datai[18]_pad  ;
	input \datai[19]_pad  ;
	input \datai[1]_pad  ;
	input \datai[20]_pad  ;
	input \datai[21]_pad  ;
	input \datai[22]_pad  ;
	input \datai[23]_pad  ;
	input \datai[24]_pad  ;
	input \datai[25]_pad  ;
	input \datai[26]_pad  ;
	input \datai[27]_pad  ;
	input \datai[28]_pad  ;
	input \datai[29]_pad  ;
	input \datai[2]_pad  ;
	input \datai[30]_pad  ;
	input \datai[31]_pad  ;
	input \datai[3]_pad  ;
	input \datai[4]_pad  ;
	input \datai[5]_pad  ;
	input \datai[6]_pad  ;
	input \datai[7]_pad  ;
	input \datai[8]_pad  ;
	input \datai[9]_pad  ;
	input \datao[15]_pad  ;
	input \datao[28]_pad  ;
	input \datao[8]_pad  ;
	input \reg0_reg[0]/NET0131  ;
	input \reg0_reg[10]/NET0131  ;
	input \reg0_reg[11]/NET0131  ;
	input \reg0_reg[12]/NET0131  ;
	input \reg0_reg[13]/NET0131  ;
	input \reg0_reg[14]/NET0131  ;
	input \reg0_reg[15]/NET0131  ;
	input \reg0_reg[16]/NET0131  ;
	input \reg0_reg[17]/NET0131  ;
	input \reg0_reg[18]/NET0131  ;
	input \reg0_reg[19]/NET0131  ;
	input \reg0_reg[1]/NET0131  ;
	input \reg0_reg[20]/NET0131  ;
	input \reg0_reg[21]/NET0131  ;
	input \reg0_reg[22]/NET0131  ;
	input \reg0_reg[23]/NET0131  ;
	input \reg0_reg[24]/NET0131  ;
	input \reg0_reg[25]/NET0131  ;
	input \reg0_reg[26]/NET0131  ;
	input \reg0_reg[27]/NET0131  ;
	input \reg0_reg[28]/NET0131  ;
	input \reg0_reg[29]/NET0131  ;
	input \reg0_reg[2]/NET0131  ;
	input \reg0_reg[30]/NET0131  ;
	input \reg0_reg[31]/NET0131  ;
	input \reg0_reg[3]/NET0131  ;
	input \reg0_reg[4]/NET0131  ;
	input \reg0_reg[5]/NET0131  ;
	input \reg0_reg[6]/NET0131  ;
	input \reg0_reg[7]/NET0131  ;
	input \reg0_reg[8]/NET0131  ;
	input \reg0_reg[9]/NET0131  ;
	input \reg1_reg[0]/NET0131  ;
	input \reg1_reg[10]/NET0131  ;
	input \reg1_reg[11]/NET0131  ;
	input \reg1_reg[12]/NET0131  ;
	input \reg1_reg[13]/NET0131  ;
	input \reg1_reg[14]/NET0131  ;
	input \reg1_reg[15]/NET0131  ;
	input \reg1_reg[16]/NET0131  ;
	input \reg1_reg[17]/NET0131  ;
	input \reg1_reg[18]/NET0131  ;
	input \reg1_reg[19]/NET0131  ;
	input \reg1_reg[1]/NET0131  ;
	input \reg1_reg[20]/NET0131  ;
	input \reg1_reg[21]/NET0131  ;
	input \reg1_reg[22]/NET0131  ;
	input \reg1_reg[23]/NET0131  ;
	input \reg1_reg[24]/NET0131  ;
	input \reg1_reg[25]/NET0131  ;
	input \reg1_reg[26]/NET0131  ;
	input \reg1_reg[27]/NET0131  ;
	input \reg1_reg[28]/NET0131  ;
	input \reg1_reg[29]/NET0131  ;
	input \reg1_reg[2]/NET0131  ;
	input \reg1_reg[30]/NET0131  ;
	input \reg1_reg[31]/NET0131  ;
	input \reg1_reg[3]/NET0131  ;
	input \reg1_reg[4]/NET0131  ;
	input \reg1_reg[5]/NET0131  ;
	input \reg1_reg[6]/NET0131  ;
	input \reg1_reg[7]/NET0131  ;
	input \reg1_reg[8]/NET0131  ;
	input \reg1_reg[9]/NET0131  ;
	input \reg2_reg[0]/NET0131  ;
	input \reg2_reg[10]/NET0131  ;
	input \reg2_reg[11]/NET0131  ;
	input \reg2_reg[12]/NET0131  ;
	input \reg2_reg[13]/NET0131  ;
	input \reg2_reg[14]/NET0131  ;
	input \reg2_reg[15]/NET0131  ;
	input \reg2_reg[16]/NET0131  ;
	input \reg2_reg[17]/NET0131  ;
	input \reg2_reg[18]/NET0131  ;
	input \reg2_reg[19]/NET0131  ;
	input \reg2_reg[1]/NET0131  ;
	input \reg2_reg[20]/NET0131  ;
	input \reg2_reg[21]/NET0131  ;
	input \reg2_reg[22]/NET0131  ;
	input \reg2_reg[23]/NET0131  ;
	input \reg2_reg[24]/NET0131  ;
	input \reg2_reg[25]/NET0131  ;
	input \reg2_reg[26]/NET0131  ;
	input \reg2_reg[27]/NET0131  ;
	input \reg2_reg[28]/NET0131  ;
	input \reg2_reg[29]/NET0131  ;
	input \reg2_reg[2]/NET0131  ;
	input \reg2_reg[30]/NET0131  ;
	input \reg2_reg[31]/NET0131  ;
	input \reg2_reg[3]/NET0131  ;
	input \reg2_reg[4]/NET0131  ;
	input \reg2_reg[5]/NET0131  ;
	input \reg2_reg[6]/NET0131  ;
	input \reg2_reg[7]/NET0131  ;
	input \reg2_reg[8]/NET0131  ;
	input \reg2_reg[9]/NET0131  ;
	input \reg3_reg[0]/NET0131  ;
	input \reg3_reg[10]/NET0131  ;
	input \reg3_reg[11]/NET0131  ;
	input \reg3_reg[12]/NET0131  ;
	input \reg3_reg[13]/NET0131  ;
	input \reg3_reg[14]/NET0131  ;
	input \reg3_reg[15]/NET0131  ;
	input \reg3_reg[16]/NET0131  ;
	input \reg3_reg[17]/NET0131  ;
	input \reg3_reg[18]/NET0131  ;
	input \reg3_reg[19]/NET0131  ;
	input \reg3_reg[1]/NET0131  ;
	input \reg3_reg[20]/NET0131  ;
	input \reg3_reg[21]/NET0131  ;
	input \reg3_reg[22]/NET0131  ;
	input \reg3_reg[23]/NET0131  ;
	input \reg3_reg[24]/NET0131  ;
	input \reg3_reg[25]/NET0131  ;
	input \reg3_reg[26]/NET0131  ;
	input \reg3_reg[27]/NET0131  ;
	input \reg3_reg[28]/NET0131  ;
	input \reg3_reg[2]/NET0131  ;
	input \reg3_reg[3]/NET0131  ;
	input \reg3_reg[4]/NET0131  ;
	input \reg3_reg[5]/NET0131  ;
	input \reg3_reg[6]/NET0131  ;
	input \reg3_reg[7]/NET0131  ;
	input \reg3_reg[8]/NET0131  ;
	input \reg3_reg[9]/NET0131  ;
	input \state_reg[0]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g22/_0_  ;
	output \g32_dup/_0_  ;
	output \g35904/_0_  ;
	output \g35905/_0_  ;
	output \g35906/_0_  ;
	output \g35907/_0_  ;
	output \g35908/_0_  ;
	output \g35909/_0_  ;
	output \g35910/_0_  ;
	output \g35911/_0_  ;
	output \g35932/_0_  ;
	output \g35955/_0_  ;
	output \g35956/_0_  ;
	output \g35957/_0_  ;
	output \g35962/_0_  ;
	output \g35967/_0_  ;
	output \g35968/_0_  ;
	output \g35971/_0_  ;
	output \g35972/_0_  ;
	output \g35973/_0_  ;
	output \g35974/_0_  ;
	output \g35975/_0_  ;
	output \g35976/_0_  ;
	output \g35977/_0_  ;
	output \g35978/_0_  ;
	output \g36015/_0_  ;
	output \g36016/_0_  ;
	output \g36018/_0_  ;
	output \g36022/_0_  ;
	output \g36023/_0_  ;
	output \g36025/_0_  ;
	output \g36029/_0_  ;
	output \g36030/_0_  ;
	output \g36031/_0_  ;
	output \g36032/_0_  ;
	output \g36033/_0_  ;
	output \g36034/_0_  ;
	output \g36035/_0_  ;
	output \g36036/_0_  ;
	output \g36038/_0_  ;
	output \g36039/_0_  ;
	output \g36040/_0_  ;
	output \g36041/_0_  ;
	output \g36073/_0_  ;
	output \g36087/_0_  ;
	output \g36091/_0_  ;
	output \g36092/_0_  ;
	output \g36093/_0_  ;
	output \g36094/_0_  ;
	output \g36096/_0_  ;
	output \g36097/_0_  ;
	output \g36098/_0_  ;
	output \g36099/_0_  ;
	output \g36100/_0_  ;
	output \g36101/_0_  ;
	output \g36102/_0_  ;
	output \g36103/_0_  ;
	output \g36104/_0_  ;
	output \g36105/_0_  ;
	output \g36106/_0_  ;
	output \g36107/_0_  ;
	output \g36108/_0_  ;
	output \g36109/_0_  ;
	output \g36110/_0_  ;
	output \g36111/_0_  ;
	output \g36112/_0_  ;
	output \g36113/_0_  ;
	output \g36165/_0_  ;
	output \g36169/_0_  ;
	output \g36170/_0_  ;
	output \g36171/_0_  ;
	output \g36172/_0_  ;
	output \g36198/_0_  ;
	output \g36199/_0_  ;
	output \g36200/_0_  ;
	output \g36201/_0_  ;
	output \g36202/_0_  ;
	output \g36203/_0_  ;
	output \g36205/_0_  ;
	output \g36206/_0_  ;
	output \g36207/_0_  ;
	output \g36208/_0_  ;
	output \g36209/_0_  ;
	output \g36240/_0_  ;
	output \g36281/_0_  ;
	output \g36282/_0_  ;
	output \g36283/_0_  ;
	output \g36284/_0_  ;
	output \g36285/_0_  ;
	output \g36286/_0_  ;
	output \g36287/_0_  ;
	output \g36288/_0_  ;
	output \g36289/_0_  ;
	output \g36290/_0_  ;
	output \g36291/_0_  ;
	output \g36292/_0_  ;
	output \g36293/_0_  ;
	output \g36294/_0_  ;
	output \g36295/_0_  ;
	output \g36296/_0_  ;
	output \g36297/_0_  ;
	output \g36298/_0_  ;
	output \g36330/_0_  ;
	output \g36385/_0_  ;
	output \g36390/_0_  ;
	output \g36391/_0_  ;
	output \g36392/_0_  ;
	output \g36393/_0_  ;
	output \g36394/_0_  ;
	output \g36470/_0_  ;
	output \g36471/_0_  ;
	output \g36472/_0_  ;
	output \g36473/_0_  ;
	output \g36474/_0_  ;
	output \g36475/_0_  ;
	output \g38/_0_  ;
	output \g38399/_0_  ;
	output \g38400/_0_  ;
	output \g39639/_0_  ;
	output \g39641/_0_  ;
	output \g39644/_0_  ;
	output \g39647/_0_  ;
	output \g39648/_0_  ;
	output \g39650/_0_  ;
	output \g39654/_0_  ;
	output \g39658/_0_  ;
	output \g39660/_0_  ;
	output \g39662/_0_  ;
	output \g39663/_0_  ;
	output \g39665/_0_  ;
	output \g39666/_0_  ;
	output \g39667/_0_  ;
	output \g39730/_0_  ;
	output \g39796/_0_  ;
	output \g39930/_0_  ;
	output \g39931/_0_  ;
	output \g39932/_0_  ;
	output \g40045/_0_  ;
	output \g40150/u3_syn_4  ;
	output \g40608/_0_  ;
	output \g41017/u3_syn_4  ;
	output \g42159/_0_  ;
	output \g42169/_0_  ;
	output \g42174/_0_  ;
	output \g42483/_0_  ;
	output \g42736/_0_  ;
	output \g42746/_0_  ;
	output \g42755/_0_  ;
	output \g42767/_0_  ;
	output \g42776/_0_  ;
	output \g42871_dup/_1_  ;
	output \g42908/_0_  ;
	output \g42938/_0_  ;
	output \g42969/_0_  ;
	output \g43022/_0_  ;
	output \g44035/_1__syn_2  ;
	output \g44227/_3_  ;
	output \g44260/_3_  ;
	output \g44261/_3_  ;
	output \g44262/_3_  ;
	output \g44311/_3_  ;
	output \g44378/_3_  ;
	output \g44379/_3_  ;
	output \g44383/_3_  ;
	output \g44384/_3_  ;
	output \g44385/_3_  ;
	output \g44386/_3_  ;
	output \g44390/_3_  ;
	output \g44391/_3_  ;
	output \g44492/_3_  ;
	output \g44493/_3_  ;
	output \g44494/_3_  ;
	output \g44495/_3_  ;
	output \g44496/_3_  ;
	output \g44497/_3_  ;
	output \g44498/_3_  ;
	output \g44499/_3_  ;
	output \g44575/_3_  ;
	output \g44589/_3_  ;
	output \g44596/_3_  ;
	output \g44615/_3_  ;
	output \g44795/_3_  ;
	output \g44803/_3_  ;
	output \g44804/_3_  ;
	output \g44888/_3_  ;
	output \g44889/_3_  ;
	output \g45004/_3_  ;
	output \g46129/_0_  ;
	output \g46133/_0_  ;
	output \g46265/_2_  ;
	output \g46313/_0_  ;
	output \g46372/_0_  ;
	output \g46377/_0_  ;
	output \g46399/_0_  ;
	output \g46405/_0_  ;
	output \g46427/_0_  ;
	output \g46461/_0_  ;
	output \g46526/_0_  ;
	output \g46576/_0_  ;
	output \g46608/_0_  ;
	output \g46697/_0_  ;
	output \g46778/_0_  ;
	output \g47007/_0_  ;
	output \g47023/_0_  ;
	output \g47077/_1_  ;
	output \g47097/_0_  ;
	output \g47109/_1_  ;
	output \g47142_dup/_1_  ;
	output \g47256/_0_  ;
	output \g47328/_0_  ;
	output \g47373/_0_  ;
	output \g47465/_0_  ;
	output \g47518/_0_  ;
	output \g47556/_1_  ;
	output \g56/_0_  ;
	output \state_reg[0]/NET0131_syn_2  ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\state_reg[0]/NET0131 ,
		_w218_
	);
	LUT4 #(
		.INIT('h8000)
	) name1 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		\reg3_reg[5]/NET0131 ,
		\reg3_reg[6]/NET0131 ,
		_w219_
	);
	LUT4 #(
		.INIT('h8000)
	) name2 (
		\reg3_reg[7]/NET0131 ,
		\reg3_reg[8]/NET0131 ,
		\reg3_reg[9]/NET0131 ,
		_w219_,
		_w220_
	);
	LUT4 #(
		.INIT('h8000)
	) name3 (
		\reg3_reg[10]/NET0131 ,
		\reg3_reg[11]/NET0131 ,
		\reg3_reg[12]/NET0131 ,
		_w220_,
		_w221_
	);
	LUT4 #(
		.INIT('h8000)
	) name4 (
		\reg3_reg[13]/NET0131 ,
		\reg3_reg[14]/NET0131 ,
		\reg3_reg[15]/NET0131 ,
		\reg3_reg[16]/NET0131 ,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w221_,
		_w222_,
		_w223_
	);
	LUT3 #(
		.INIT('h6a)
	) name6 (
		\reg3_reg[17]/NET0131 ,
		_w221_,
		_w222_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\IR_reg[14]/NET0131 ,
		\IR_reg[15]/NET0131 ,
		_w226_
	);
	LUT4 #(
		.INIT('h0001)
	) name9 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[2]/NET0131 ,
		\IR_reg[3]/NET0131 ,
		_w227_
	);
	LUT3 #(
		.INIT('h01)
	) name10 (
		\IR_reg[5]/NET0131 ,
		\IR_reg[6]/NET0131 ,
		\IR_reg[7]/NET0131 ,
		_w228_
	);
	LUT3 #(
		.INIT('h40)
	) name11 (
		\IR_reg[4]/NET0131 ,
		_w227_,
		_w228_,
		_w229_
	);
	LUT4 #(
		.INIT('h0001)
	) name12 (
		\IR_reg[10]/NET0131 ,
		\IR_reg[11]/NET0131 ,
		\IR_reg[8]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\IR_reg[12]/NET0131 ,
		_w230_,
		_w231_
	);
	LUT3 #(
		.INIT('h10)
	) name14 (
		\IR_reg[12]/NET0131 ,
		\IR_reg[13]/NET0131 ,
		_w230_,
		_w232_
	);
	LUT3 #(
		.INIT('h80)
	) name15 (
		_w226_,
		_w229_,
		_w232_,
		_w233_
	);
	LUT4 #(
		.INIT('h0001)
	) name16 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[17]/NET0131 ,
		\IR_reg[18]/NET0131 ,
		\IR_reg[19]/NET0131 ,
		_w234_
	);
	LUT4 #(
		.INIT('h8000)
	) name17 (
		_w226_,
		_w229_,
		_w232_,
		_w234_,
		_w235_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name18 (
		\IR_reg[22]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w225_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h6)
	) name19 (
		\IR_reg[23]/NET0131 ,
		_w236_,
		_w237_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name20 (
		\IR_reg[31]/NET0131 ,
		_w226_,
		_w229_,
		_w232_,
		_w238_
	);
	LUT4 #(
		.INIT('h0001)
	) name21 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		\IR_reg[22]/NET0131 ,
		\IR_reg[23]/NET0131 ,
		_w239_
	);
	LUT3 #(
		.INIT('h2a)
	) name22 (
		\IR_reg[31]/NET0131 ,
		_w234_,
		_w239_,
		_w240_
	);
	LUT3 #(
		.INIT('h56)
	) name23 (
		\IR_reg[24]/NET0131 ,
		_w238_,
		_w240_,
		_w241_
	);
	LUT4 #(
		.INIT('h0001)
	) name24 (
		\IR_reg[14]/NET0131 ,
		\IR_reg[15]/NET0131 ,
		\IR_reg[24]/NET0131 ,
		\IR_reg[25]/NET0131 ,
		_w242_
	);
	LUT3 #(
		.INIT('h80)
	) name25 (
		_w234_,
		_w239_,
		_w242_,
		_w243_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name26 (
		\IR_reg[31]/NET0131 ,
		_w229_,
		_w232_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h9)
	) name27 (
		\IR_reg[26]/NET0131 ,
		_w244_,
		_w245_
	);
	LUT4 #(
		.INIT('h0001)
	) name28 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[14]/NET0131 ,
		\IR_reg[15]/NET0131 ,
		\IR_reg[24]/NET0131 ,
		_w246_
	);
	LUT3 #(
		.INIT('h80)
	) name29 (
		_w234_,
		_w239_,
		_w246_,
		_w247_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name30 (
		\IR_reg[31]/NET0131 ,
		_w229_,
		_w231_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h9)
	) name31 (
		\IR_reg[25]/NET0131 ,
		_w248_,
		_w249_
	);
	LUT4 #(
		.INIT('h1428)
	) name32 (
		\IR_reg[25]/NET0131 ,
		\IR_reg[26]/NET0131 ,
		_w244_,
		_w248_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w241_,
		_w250_,
		_w251_
	);
	LUT4 #(
		.INIT('h9000)
	) name34 (
		\IR_reg[23]/NET0131 ,
		_w236_,
		_w241_,
		_w250_,
		_w252_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w224_,
		_w252_,
		_w253_
	);
	LUT4 #(
		.INIT('h0999)
	) name36 (
		\IR_reg[23]/NET0131 ,
		_w236_,
		_w241_,
		_w250_,
		_w254_
	);
	LUT4 #(
		.INIT('h8882)
	) name37 (
		\B_reg/NET0131 ,
		\IR_reg[24]/NET0131 ,
		_w238_,
		_w240_,
		_w255_
	);
	LUT4 #(
		.INIT('h3222)
	) name38 (
		\d_reg[0]/NET0131 ,
		_w245_,
		_w249_,
		_w255_,
		_w256_
	);
	LUT3 #(
		.INIT('h41)
	) name39 (
		\B_reg/NET0131 ,
		\IR_reg[25]/NET0131 ,
		_w248_,
		_w257_
	);
	LUT3 #(
		.INIT('hc8)
	) name40 (
		_w245_,
		_w241_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('he)
	) name41 (
		_w256_,
		_w258_,
		_w259_
	);
	LUT4 #(
		.INIT('h6669)
	) name42 (
		\B_reg/NET0131 ,
		\IR_reg[24]/NET0131 ,
		_w238_,
		_w240_,
		_w260_
	);
	LUT4 #(
		.INIT('h2e3e)
	) name43 (
		\d_reg[1]/NET0131 ,
		_w245_,
		_w249_,
		_w260_,
		_w261_
	);
	LUT3 #(
		.INIT('he0)
	) name44 (
		_w256_,
		_w258_,
		_w261_,
		_w262_
	);
	LUT4 #(
		.INIT('h02aa)
	) name45 (
		_w224_,
		_w256_,
		_w258_,
		_w261_,
		_w263_
	);
	LUT4 #(
		.INIT('h0001)
	) name46 (
		\IR_reg[24]/NET0131 ,
		\IR_reg[25]/NET0131 ,
		\IR_reg[26]/NET0131 ,
		\IR_reg[27]/NET0131 ,
		_w264_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name47 (
		\IR_reg[31]/NET0131 ,
		_w234_,
		_w239_,
		_w264_,
		_w265_
	);
	LUT3 #(
		.INIT('h56)
	) name48 (
		\IR_reg[28]/NET0131 ,
		_w238_,
		_w265_,
		_w266_
	);
	LUT4 #(
		.INIT('h0001)
	) name49 (
		\IR_reg[25]/NET0131 ,
		\IR_reg[26]/NET0131 ,
		\IR_reg[27]/NET0131 ,
		\IR_reg[28]/NET0131 ,
		_w267_
	);
	LUT4 #(
		.INIT('h8000)
	) name50 (
		_w229_,
		_w231_,
		_w247_,
		_w267_,
		_w268_
	);
	LUT3 #(
		.INIT('ha6)
	) name51 (
		\IR_reg[29]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w268_,
		_w269_
	);
	LUT4 #(
		.INIT('h0001)
	) name52 (
		\IR_reg[26]/NET0131 ,
		\IR_reg[27]/NET0131 ,
		\IR_reg[28]/NET0131 ,
		\IR_reg[29]/NET0131 ,
		_w270_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\IR_reg[31]/NET0131 ,
		_w270_,
		_w271_
	);
	LUT3 #(
		.INIT('h56)
	) name54 (
		\IR_reg[30]/NET0131 ,
		_w244_,
		_w271_,
		_w272_
	);
	LUT4 #(
		.INIT('hf35f)
	) name55 (
		\reg1_reg[2]/NET0131 ,
		\reg2_reg[2]/NET0131 ,
		_w269_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w269_,
		_w272_,
		_w274_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name57 (
		\reg0_reg[2]/NET0131 ,
		\reg3_reg[2]/NET0131 ,
		_w269_,
		_w272_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w273_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h7)
	) name59 (
		_w273_,
		_w275_,
		_w277_
	);
	LUT4 #(
		.INIT('hff35)
	) name60 (
		\reg0_reg[1]/NET0131 ,
		\reg1_reg[1]/NET0131 ,
		_w269_,
		_w272_,
		_w278_
	);
	LUT4 #(
		.INIT('h35ff)
	) name61 (
		\reg2_reg[1]/NET0131 ,
		\reg3_reg[1]/NET0131 ,
		_w269_,
		_w272_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w278_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h7)
	) name63 (
		_w278_,
		_w279_,
		_w281_
	);
	LUT4 #(
		.INIT('hff35)
	) name64 (
		\reg0_reg[0]/NET0131 ,
		\reg1_reg[0]/NET0131 ,
		_w269_,
		_w272_,
		_w282_
	);
	LUT4 #(
		.INIT('h35ff)
	) name65 (
		\reg2_reg[0]/NET0131 ,
		\reg3_reg[0]/NET0131 ,
		_w269_,
		_w272_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w282_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h7)
	) name67 (
		_w282_,
		_w283_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\reg3_reg[17]/NET0131 ,
		\reg3_reg[18]/NET0131 ,
		_w286_
	);
	LUT3 #(
		.INIT('h80)
	) name69 (
		_w221_,
		_w222_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\reg3_reg[19]/NET0131 ,
		\reg3_reg[20]/NET0131 ,
		_w288_
	);
	LUT3 #(
		.INIT('h80)
	) name71 (
		\reg3_reg[19]/NET0131 ,
		\reg3_reg[20]/NET0131 ,
		\reg3_reg[21]/NET0131 ,
		_w289_
	);
	LUT4 #(
		.INIT('h8000)
	) name72 (
		\reg3_reg[19]/NET0131 ,
		\reg3_reg[20]/NET0131 ,
		\reg3_reg[21]/NET0131 ,
		\reg3_reg[22]/NET0131 ,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\reg3_reg[23]/NET0131 ,
		_w290_,
		_w291_
	);
	LUT3 #(
		.INIT('h80)
	) name74 (
		\reg3_reg[23]/NET0131 ,
		\reg3_reg[24]/NET0131 ,
		_w290_,
		_w292_
	);
	LUT4 #(
		.INIT('h8000)
	) name75 (
		_w221_,
		_w222_,
		_w286_,
		_w292_,
		_w293_
	);
	LUT4 #(
		.INIT('h8000)
	) name76 (
		\reg3_reg[25]/NET0131 ,
		\reg3_reg[26]/NET0131 ,
		\reg3_reg[27]/NET0131 ,
		\reg3_reg[28]/NET0131 ,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w293_,
		_w294_,
		_w295_
	);
	LUT4 #(
		.INIT('h8000)
	) name78 (
		_w269_,
		_w272_,
		_w293_,
		_w294_,
		_w296_
	);
	LUT3 #(
		.INIT('h02)
	) name79 (
		\reg0_reg[31]/NET0131 ,
		_w269_,
		_w272_,
		_w297_
	);
	LUT4 #(
		.INIT('hf35f)
	) name80 (
		\reg1_reg[31]/NET0131 ,
		\reg2_reg[31]/NET0131 ,
		_w269_,
		_w272_,
		_w298_
	);
	LUT3 #(
		.INIT('h10)
	) name81 (
		_w296_,
		_w297_,
		_w298_,
		_w299_
	);
	LUT3 #(
		.INIT('hef)
	) name82 (
		_w296_,
		_w297_,
		_w298_,
		_w300_
	);
	LUT4 #(
		.INIT('h0001)
	) name83 (
		_w276_,
		_w280_,
		_w284_,
		_w299_,
		_w301_
	);
	LUT4 #(
		.INIT('hc5ff)
	) name84 (
		\reg2_reg[3]/NET0131 ,
		\reg3_reg[3]/NET0131 ,
		_w269_,
		_w272_,
		_w302_
	);
	LUT4 #(
		.INIT('hff35)
	) name85 (
		\reg0_reg[3]/NET0131 ,
		\reg1_reg[3]/NET0131 ,
		_w269_,
		_w272_,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		_w302_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h7)
	) name87 (
		_w302_,
		_w303_,
		_w305_
	);
	LUT2 #(
		.INIT('h6)
	) name88 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		_w306_
	);
	LUT4 #(
		.INIT('h37f7)
	) name89 (
		\reg1_reg[4]/NET0131 ,
		_w269_,
		_w272_,
		_w306_,
		_w307_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name90 (
		\reg0_reg[4]/NET0131 ,
		\reg2_reg[4]/NET0131 ,
		_w269_,
		_w272_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w307_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h7)
	) name92 (
		_w307_,
		_w308_,
		_w310_
	);
	LUT4 #(
		.INIT('h0777)
	) name93 (
		_w302_,
		_w303_,
		_w307_,
		_w308_,
		_w311_
	);
	LUT4 #(
		.INIT('hff35)
	) name94 (
		\reg0_reg[6]/NET0131 ,
		\reg1_reg[6]/NET0131 ,
		_w269_,
		_w272_,
		_w312_
	);
	LUT4 #(
		.INIT('h7f80)
	) name95 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		\reg3_reg[5]/NET0131 ,
		\reg3_reg[6]/NET0131 ,
		_w313_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name96 (
		\reg2_reg[6]/NET0131 ,
		_w269_,
		_w272_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w312_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h7)
	) name98 (
		_w312_,
		_w314_,
		_w316_
	);
	LUT3 #(
		.INIT('h78)
	) name99 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		\reg3_reg[5]/NET0131 ,
		_w317_
	);
	LUT4 #(
		.INIT('h37f7)
	) name100 (
		\reg1_reg[5]/NET0131 ,
		_w269_,
		_w272_,
		_w317_,
		_w318_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name101 (
		\reg0_reg[5]/NET0131 ,
		\reg2_reg[5]/NET0131 ,
		_w269_,
		_w272_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w318_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h7)
	) name103 (
		_w318_,
		_w319_,
		_w321_
	);
	LUT4 #(
		.INIT('h0777)
	) name104 (
		_w312_,
		_w314_,
		_w318_,
		_w319_,
		_w322_
	);
	LUT4 #(
		.INIT('hff35)
	) name105 (
		\reg0_reg[7]/NET0131 ,
		\reg1_reg[7]/NET0131 ,
		_w269_,
		_w272_,
		_w323_
	);
	LUT2 #(
		.INIT('h6)
	) name106 (
		\reg3_reg[7]/NET0131 ,
		_w219_,
		_w324_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name107 (
		\reg2_reg[7]/NET0131 ,
		_w269_,
		_w272_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w323_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h7)
	) name109 (
		_w323_,
		_w325_,
		_w327_
	);
	LUT4 #(
		.INIT('hff35)
	) name110 (
		\reg0_reg[8]/NET0131 ,
		\reg1_reg[8]/NET0131 ,
		_w269_,
		_w272_,
		_w328_
	);
	LUT3 #(
		.INIT('h6c)
	) name111 (
		\reg3_reg[7]/NET0131 ,
		\reg3_reg[8]/NET0131 ,
		_w219_,
		_w329_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name112 (
		\reg2_reg[8]/NET0131 ,
		_w269_,
		_w272_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w328_,
		_w330_,
		_w331_
	);
	LUT4 #(
		.INIT('hff35)
	) name114 (
		\reg0_reg[9]/NET0131 ,
		\reg1_reg[9]/NET0131 ,
		_w269_,
		_w272_,
		_w332_
	);
	LUT4 #(
		.INIT('h78f0)
	) name115 (
		\reg3_reg[7]/NET0131 ,
		\reg3_reg[8]/NET0131 ,
		\reg3_reg[9]/NET0131 ,
		_w219_,
		_w333_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name116 (
		\reg2_reg[9]/NET0131 ,
		_w269_,
		_w272_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		_w332_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h7)
	) name118 (
		_w332_,
		_w334_,
		_w336_
	);
	LUT4 #(
		.INIT('h0777)
	) name119 (
		_w328_,
		_w330_,
		_w332_,
		_w334_,
		_w337_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w326_,
		_w337_,
		_w338_
	);
	LUT4 #(
		.INIT('h8000)
	) name121 (
		_w301_,
		_w311_,
		_w322_,
		_w338_,
		_w339_
	);
	LUT4 #(
		.INIT('h78f0)
	) name122 (
		\reg3_reg[10]/NET0131 ,
		\reg3_reg[11]/NET0131 ,
		\reg3_reg[12]/NET0131 ,
		_w220_,
		_w340_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name123 (
		\reg2_reg[12]/NET0131 ,
		_w269_,
		_w272_,
		_w340_,
		_w341_
	);
	LUT4 #(
		.INIT('hff35)
	) name124 (
		\reg0_reg[12]/NET0131 ,
		\reg1_reg[12]/NET0131 ,
		_w269_,
		_w272_,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w341_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h7)
	) name126 (
		_w341_,
		_w342_,
		_w344_
	);
	LUT4 #(
		.INIT('hff35)
	) name127 (
		\reg0_reg[11]/NET0131 ,
		\reg1_reg[11]/NET0131 ,
		_w269_,
		_w272_,
		_w345_
	);
	LUT3 #(
		.INIT('h6c)
	) name128 (
		\reg3_reg[10]/NET0131 ,
		\reg3_reg[11]/NET0131 ,
		_w220_,
		_w346_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name129 (
		\reg2_reg[11]/NET0131 ,
		_w269_,
		_w272_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w345_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h7)
	) name131 (
		_w345_,
		_w347_,
		_w349_
	);
	LUT4 #(
		.INIT('hf35f)
	) name132 (
		\reg1_reg[10]/NET0131 ,
		\reg2_reg[10]/NET0131 ,
		_w269_,
		_w272_,
		_w350_
	);
	LUT2 #(
		.INIT('h6)
	) name133 (
		\reg3_reg[10]/NET0131 ,
		_w220_,
		_w351_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name134 (
		\reg0_reg[10]/NET0131 ,
		_w269_,
		_w272_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w350_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h7)
	) name136 (
		_w350_,
		_w352_,
		_w354_
	);
	LUT4 #(
		.INIT('h0777)
	) name137 (
		_w345_,
		_w347_,
		_w350_,
		_w352_,
		_w355_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		_w343_,
		_w355_,
		_w356_
	);
	LUT4 #(
		.INIT('h8000)
	) name139 (
		\reg3_reg[13]/NET0131 ,
		\reg3_reg[14]/NET0131 ,
		\reg3_reg[15]/NET0131 ,
		_w221_,
		_w357_
	);
	LUT3 #(
		.INIT('h32)
	) name140 (
		\reg3_reg[16]/NET0131 ,
		_w223_,
		_w357_,
		_w358_
	);
	LUT3 #(
		.INIT('h02)
	) name141 (
		\reg0_reg[16]/NET0131 ,
		_w269_,
		_w272_,
		_w359_
	);
	LUT4 #(
		.INIT('hf35f)
	) name142 (
		\reg1_reg[16]/NET0131 ,
		\reg2_reg[16]/NET0131 ,
		_w269_,
		_w272_,
		_w360_
	);
	LUT4 #(
		.INIT('h1300)
	) name143 (
		_w274_,
		_w359_,
		_w358_,
		_w360_,
		_w361_
	);
	LUT4 #(
		.INIT('hecff)
	) name144 (
		_w274_,
		_w359_,
		_w358_,
		_w360_,
		_w362_
	);
	LUT3 #(
		.INIT('h6c)
	) name145 (
		\reg3_reg[13]/NET0131 ,
		\reg3_reg[14]/NET0131 ,
		_w221_,
		_w363_
	);
	LUT3 #(
		.INIT('h80)
	) name146 (
		_w269_,
		_w272_,
		_w363_,
		_w364_
	);
	LUT3 #(
		.INIT('h20)
	) name147 (
		\reg2_reg[14]/NET0131 ,
		_w269_,
		_w272_,
		_w365_
	);
	LUT4 #(
		.INIT('hff35)
	) name148 (
		\reg0_reg[14]/NET0131 ,
		\reg1_reg[14]/NET0131 ,
		_w269_,
		_w272_,
		_w366_
	);
	LUT3 #(
		.INIT('h10)
	) name149 (
		_w365_,
		_w364_,
		_w366_,
		_w367_
	);
	LUT3 #(
		.INIT('hef)
	) name150 (
		_w365_,
		_w364_,
		_w366_,
		_w368_
	);
	LUT2 #(
		.INIT('h6)
	) name151 (
		\reg3_reg[13]/NET0131 ,
		_w221_,
		_w369_
	);
	LUT4 #(
		.INIT('h37f7)
	) name152 (
		\reg1_reg[13]/NET0131 ,
		_w269_,
		_w272_,
		_w369_,
		_w370_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name153 (
		\reg0_reg[13]/NET0131 ,
		\reg2_reg[13]/NET0131 ,
		_w269_,
		_w272_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		_w370_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h7)
	) name155 (
		_w370_,
		_w371_,
		_w373_
	);
	LUT4 #(
		.INIT('h78f0)
	) name156 (
		\reg3_reg[13]/NET0131 ,
		\reg3_reg[14]/NET0131 ,
		\reg3_reg[15]/NET0131 ,
		_w221_,
		_w374_
	);
	LUT3 #(
		.INIT('h80)
	) name157 (
		_w269_,
		_w272_,
		_w374_,
		_w375_
	);
	LUT3 #(
		.INIT('h20)
	) name158 (
		\reg2_reg[15]/NET0131 ,
		_w269_,
		_w272_,
		_w376_
	);
	LUT4 #(
		.INIT('hff35)
	) name159 (
		\reg0_reg[15]/NET0131 ,
		\reg1_reg[15]/NET0131 ,
		_w269_,
		_w272_,
		_w377_
	);
	LUT3 #(
		.INIT('h10)
	) name160 (
		_w376_,
		_w375_,
		_w377_,
		_w378_
	);
	LUT4 #(
		.INIT('h0001)
	) name161 (
		_w372_,
		_w378_,
		_w367_,
		_w361_,
		_w379_
	);
	LUT3 #(
		.INIT('h80)
	) name162 (
		_w339_,
		_w356_,
		_w379_,
		_w380_
	);
	LUT3 #(
		.INIT('h80)
	) name163 (
		_w224_,
		_w269_,
		_w272_,
		_w381_
	);
	LUT3 #(
		.INIT('h02)
	) name164 (
		\reg0_reg[17]/NET0131 ,
		_w269_,
		_w272_,
		_w382_
	);
	LUT4 #(
		.INIT('hf35f)
	) name165 (
		\reg1_reg[17]/NET0131 ,
		\reg2_reg[17]/NET0131 ,
		_w269_,
		_w272_,
		_w383_
	);
	LUT3 #(
		.INIT('h10)
	) name166 (
		_w382_,
		_w381_,
		_w383_,
		_w384_
	);
	LUT3 #(
		.INIT('hef)
	) name167 (
		_w382_,
		_w381_,
		_w383_,
		_w385_
	);
	LUT4 #(
		.INIT('h0080)
	) name168 (
		_w339_,
		_w356_,
		_w379_,
		_w384_,
		_w386_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name169 (
		\reg3_reg[17]/NET0131 ,
		\reg3_reg[18]/NET0131 ,
		_w221_,
		_w222_,
		_w387_
	);
	LUT3 #(
		.INIT('h80)
	) name170 (
		_w269_,
		_w272_,
		_w387_,
		_w388_
	);
	LUT3 #(
		.INIT('h20)
	) name171 (
		\reg2_reg[18]/NET0131 ,
		_w269_,
		_w272_,
		_w389_
	);
	LUT4 #(
		.INIT('hff35)
	) name172 (
		\reg0_reg[18]/NET0131 ,
		\reg1_reg[18]/NET0131 ,
		_w269_,
		_w272_,
		_w390_
	);
	LUT3 #(
		.INIT('h10)
	) name173 (
		_w389_,
		_w388_,
		_w390_,
		_w391_
	);
	LUT3 #(
		.INIT('hef)
	) name174 (
		_w389_,
		_w388_,
		_w390_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w384_,
		_w391_,
		_w393_
	);
	LUT4 #(
		.INIT('h8000)
	) name176 (
		_w339_,
		_w356_,
		_w379_,
		_w393_,
		_w394_
	);
	LUT4 #(
		.INIT('h5510)
	) name177 (
		_w266_,
		_w386_,
		_w391_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w266_,
		_w361_,
		_w396_
	);
	LUT4 #(
		.INIT('h3331)
	) name179 (
		_w262_,
		_w263_,
		_w395_,
		_w396_,
		_w397_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name180 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w235_,
		_w398_
	);
	LUT3 #(
		.INIT('ha6)
	) name181 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w235_,
		_w399_
	);
	LUT4 #(
		.INIT('h4424)
	) name182 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w235_,
		_w400_
	);
	LUT4 #(
		.INIT('h5999)
	) name183 (
		\IR_reg[22]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w225_,
		_w235_,
		_w401_
	);
	LUT4 #(
		.INIT('hfe00)
	) name184 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[17]/NET0131 ,
		\IR_reg[18]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w402_
	);
	LUT3 #(
		.INIT('h56)
	) name185 (
		\IR_reg[19]/NET0131 ,
		_w238_,
		_w402_,
		_w403_
	);
	LUT3 #(
		.INIT('h10)
	) name186 (
		_w401_,
		_w403_,
		_w400_,
		_w404_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		_w397_,
		_w404_,
		_w405_
	);
	LUT3 #(
		.INIT('he0)
	) name188 (
		\IR_reg[25]/NET0131 ,
		\IR_reg[26]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w406_
	);
	LUT3 #(
		.INIT('h56)
	) name189 (
		\IR_reg[27]/NET0131 ,
		_w248_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w266_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w409_
	);
	LUT3 #(
		.INIT('h56)
	) name192 (
		\IR_reg[17]/NET0131 ,
		_w238_,
		_w409_,
		_w410_
	);
	LUT4 #(
		.INIT('haba8)
	) name193 (
		\datai[17]_pad ,
		_w266_,
		_w407_,
		_w410_,
		_w411_
	);
	LUT4 #(
		.INIT('h0100)
	) name194 (
		_w411_,
		_w382_,
		_w381_,
		_w383_,
		_w412_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name195 (
		_w411_,
		_w382_,
		_w381_,
		_w383_,
		_w413_
	);
	LUT4 #(
		.INIT('h5655)
	) name196 (
		_w411_,
		_w382_,
		_w381_,
		_w383_,
		_w414_
	);
	LUT4 #(
		.INIT('h1000)
	) name197 (
		\IR_reg[4]/NET0131 ,
		\IR_reg[8]/NET0131 ,
		_w227_,
		_w228_,
		_w415_
	);
	LUT3 #(
		.INIT('hc8)
	) name198 (
		\IR_reg[10]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		_w416_
	);
	LUT4 #(
		.INIT('h55a6)
	) name199 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w415_,
		_w416_,
		_w417_
	);
	LUT4 #(
		.INIT('h5457)
	) name200 (
		\datai[11]_pad ,
		_w266_,
		_w407_,
		_w417_,
		_w418_
	);
	LUT3 #(
		.INIT('h08)
	) name201 (
		_w345_,
		_w347_,
		_w418_,
		_w419_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name202 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		_w227_,
		_w228_,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\IR_reg[31]/NET0131 ,
		_w230_,
		_w421_
	);
	LUT3 #(
		.INIT('h56)
	) name204 (
		\IR_reg[12]/NET0131 ,
		_w420_,
		_w421_,
		_w422_
	);
	LUT4 #(
		.INIT('h5457)
	) name205 (
		\datai[12]_pad ,
		_w266_,
		_w407_,
		_w422_,
		_w423_
	);
	LUT3 #(
		.INIT('h08)
	) name206 (
		_w341_,
		_w342_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w419_,
		_w424_,
		_w425_
	);
	LUT4 #(
		.INIT('h6a66)
	) name208 (
		\IR_reg[10]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		_w415_,
		_w426_
	);
	LUT4 #(
		.INIT('h5457)
	) name209 (
		\datai[10]_pad ,
		_w266_,
		_w407_,
		_w426_,
		_w427_
	);
	LUT3 #(
		.INIT('h08)
	) name210 (
		_w350_,
		_w352_,
		_w427_,
		_w428_
	);
	LUT3 #(
		.INIT('h70)
	) name211 (
		_w350_,
		_w352_,
		_w427_,
		_w429_
	);
	LUT3 #(
		.INIT('h39)
	) name212 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		_w415_,
		_w430_
	);
	LUT4 #(
		.INIT('h5754)
	) name213 (
		\datai[9]_pad ,
		_w266_,
		_w407_,
		_w430_,
		_w431_
	);
	LUT3 #(
		.INIT('h70)
	) name214 (
		_w332_,
		_w334_,
		_w431_,
		_w432_
	);
	LUT3 #(
		.INIT('h54)
	) name215 (
		_w428_,
		_w429_,
		_w432_,
		_w433_
	);
	LUT3 #(
		.INIT('h70)
	) name216 (
		_w341_,
		_w342_,
		_w423_,
		_w434_
	);
	LUT3 #(
		.INIT('h70)
	) name217 (
		_w345_,
		_w347_,
		_w418_,
		_w435_
	);
	LUT3 #(
		.INIT('h54)
	) name218 (
		_w424_,
		_w434_,
		_w435_,
		_w436_
	);
	LUT3 #(
		.INIT('h07)
	) name219 (
		_w425_,
		_w433_,
		_w436_,
		_w437_
	);
	LUT4 #(
		.INIT('h5999)
	) name220 (
		\IR_reg[14]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w229_,
		_w232_,
		_w438_
	);
	LUT4 #(
		.INIT('h5754)
	) name221 (
		\datai[14]_pad ,
		_w266_,
		_w407_,
		_w438_,
		_w439_
	);
	LUT4 #(
		.INIT('h0010)
	) name222 (
		_w365_,
		_w364_,
		_w366_,
		_w439_,
		_w440_
	);
	LUT4 #(
		.INIT('ha666)
	) name223 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w229_,
		_w231_,
		_w441_
	);
	LUT4 #(
		.INIT('h5457)
	) name224 (
		\datai[13]_pad ,
		_w266_,
		_w407_,
		_w441_,
		_w442_
	);
	LUT3 #(
		.INIT('h08)
	) name225 (
		_w370_,
		_w371_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		_w440_,
		_w443_,
		_w444_
	);
	LUT3 #(
		.INIT('ha6)
	) name227 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w233_,
		_w445_
	);
	LUT4 #(
		.INIT('h5457)
	) name228 (
		\datai[16]_pad ,
		_w266_,
		_w407_,
		_w445_,
		_w446_
	);
	LUT4 #(
		.INIT('h7333)
	) name229 (
		\IR_reg[14]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w229_,
		_w232_,
		_w447_
	);
	LUT2 #(
		.INIT('h9)
	) name230 (
		\IR_reg[15]/NET0131 ,
		_w447_,
		_w448_
	);
	LUT4 #(
		.INIT('haba8)
	) name231 (
		\datai[15]_pad ,
		_w266_,
		_w407_,
		_w448_,
		_w449_
	);
	LUT4 #(
		.INIT('h1000)
	) name232 (
		_w376_,
		_w375_,
		_w377_,
		_w449_,
		_w450_
	);
	LUT3 #(
		.INIT('h0d)
	) name233 (
		_w361_,
		_w446_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w444_,
		_w451_,
		_w452_
	);
	LUT4 #(
		.INIT('hef00)
	) name235 (
		_w365_,
		_w364_,
		_w366_,
		_w439_,
		_w453_
	);
	LUT3 #(
		.INIT('h70)
	) name236 (
		_w370_,
		_w371_,
		_w442_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w453_,
		_w454_,
		_w455_
	);
	LUT3 #(
		.INIT('h54)
	) name238 (
		_w440_,
		_w453_,
		_w454_,
		_w456_
	);
	LUT4 #(
		.INIT('h00ef)
	) name239 (
		_w376_,
		_w375_,
		_w377_,
		_w449_,
		_w457_
	);
	LUT3 #(
		.INIT('hd4)
	) name240 (
		_w361_,
		_w446_,
		_w457_,
		_w458_
	);
	LUT3 #(
		.INIT('h07)
	) name241 (
		_w451_,
		_w456_,
		_w458_,
		_w459_
	);
	LUT3 #(
		.INIT('hb0)
	) name242 (
		_w437_,
		_w452_,
		_w459_,
		_w460_
	);
	LUT3 #(
		.INIT('h08)
	) name243 (
		_w332_,
		_w334_,
		_w431_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w428_,
		_w461_,
		_w462_
	);
	LUT4 #(
		.INIT('h0001)
	) name245 (
		_w419_,
		_w424_,
		_w428_,
		_w461_,
		_w463_
	);
	LUT3 #(
		.INIT('ha8)
	) name246 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[5]/NET0131 ,
		\IR_reg[6]/NET0131 ,
		_w464_
	);
	LUT4 #(
		.INIT('h0075)
	) name247 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		_w227_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h9)
	) name248 (
		\IR_reg[7]/NET0131 ,
		_w465_,
		_w466_
	);
	LUT4 #(
		.INIT('h5457)
	) name249 (
		\datai[7]_pad ,
		_w266_,
		_w407_,
		_w466_,
		_w467_
	);
	LUT3 #(
		.INIT('h08)
	) name250 (
		_w323_,
		_w325_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h6)
	) name251 (
		\IR_reg[8]/NET0131 ,
		_w420_,
		_w469_
	);
	LUT4 #(
		.INIT('h5457)
	) name252 (
		\datai[8]_pad ,
		_w266_,
		_w407_,
		_w469_,
		_w470_
	);
	LUT3 #(
		.INIT('h08)
	) name253 (
		_w328_,
		_w330_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		_w468_,
		_w471_,
		_w472_
	);
	LUT4 #(
		.INIT('h5755)
	) name255 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		\IR_reg[5]/NET0131 ,
		_w227_,
		_w473_
	);
	LUT2 #(
		.INIT('h9)
	) name256 (
		\IR_reg[6]/NET0131 ,
		_w473_,
		_w474_
	);
	LUT4 #(
		.INIT('h5457)
	) name257 (
		\datai[6]_pad ,
		_w266_,
		_w407_,
		_w474_,
		_w475_
	);
	LUT3 #(
		.INIT('h08)
	) name258 (
		_w312_,
		_w314_,
		_w475_,
		_w476_
	);
	LUT3 #(
		.INIT('h70)
	) name259 (
		_w312_,
		_w314_,
		_w475_,
		_w477_
	);
	LUT4 #(
		.INIT('h785a)
	) name260 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		\IR_reg[5]/NET0131 ,
		_w227_,
		_w478_
	);
	LUT4 #(
		.INIT('h5457)
	) name261 (
		\datai[5]_pad ,
		_w266_,
		_w407_,
		_w478_,
		_w479_
	);
	LUT3 #(
		.INIT('h70)
	) name262 (
		_w318_,
		_w319_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w477_,
		_w480_,
		_w481_
	);
	LUT3 #(
		.INIT('h54)
	) name264 (
		_w476_,
		_w477_,
		_w480_,
		_w482_
	);
	LUT3 #(
		.INIT('h70)
	) name265 (
		_w328_,
		_w330_,
		_w470_,
		_w483_
	);
	LUT3 #(
		.INIT('h70)
	) name266 (
		_w323_,
		_w325_,
		_w467_,
		_w484_
	);
	LUT3 #(
		.INIT('h54)
	) name267 (
		_w471_,
		_w483_,
		_w484_,
		_w485_
	);
	LUT3 #(
		.INIT('h07)
	) name268 (
		_w472_,
		_w482_,
		_w485_,
		_w486_
	);
	LUT3 #(
		.INIT('h39)
	) name269 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		_w227_,
		_w487_
	);
	LUT4 #(
		.INIT('h5754)
	) name270 (
		\datai[4]_pad ,
		_w266_,
		_w407_,
		_w487_,
		_w488_
	);
	LUT3 #(
		.INIT('h08)
	) name271 (
		_w307_,
		_w308_,
		_w488_,
		_w489_
	);
	LUT3 #(
		.INIT('h6c)
	) name272 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w490_
	);
	LUT4 #(
		.INIT('h5457)
	) name273 (
		\datai[1]_pad ,
		_w266_,
		_w407_,
		_w490_,
		_w491_
	);
	LUT3 #(
		.INIT('h08)
	) name274 (
		_w278_,
		_w279_,
		_w491_,
		_w492_
	);
	LUT4 #(
		.INIT('h3335)
	) name275 (
		\IR_reg[0]/NET0131 ,
		\datai[0]_pad ,
		_w266_,
		_w407_,
		_w493_
	);
	LUT3 #(
		.INIT('h08)
	) name276 (
		_w282_,
		_w283_,
		_w493_,
		_w494_
	);
	LUT3 #(
		.INIT('h70)
	) name277 (
		_w278_,
		_w279_,
		_w491_,
		_w495_
	);
	LUT4 #(
		.INIT('he10f)
	) name278 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[2]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w496_
	);
	LUT4 #(
		.INIT('h5754)
	) name279 (
		\datai[2]_pad ,
		_w266_,
		_w407_,
		_w496_,
		_w497_
	);
	LUT3 #(
		.INIT('h70)
	) name280 (
		_w273_,
		_w275_,
		_w497_,
		_w498_
	);
	LUT4 #(
		.INIT('h00b2)
	) name281 (
		_w280_,
		_w491_,
		_w494_,
		_w498_,
		_w499_
	);
	LUT4 #(
		.INIT('h01ff)
	) name282 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[2]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w500_
	);
	LUT2 #(
		.INIT('h9)
	) name283 (
		\IR_reg[3]/NET0131 ,
		_w500_,
		_w501_
	);
	LUT4 #(
		.INIT('h5457)
	) name284 (
		\datai[3]_pad ,
		_w266_,
		_w407_,
		_w501_,
		_w502_
	);
	LUT3 #(
		.INIT('h08)
	) name285 (
		_w302_,
		_w303_,
		_w502_,
		_w503_
	);
	LUT3 #(
		.INIT('h08)
	) name286 (
		_w273_,
		_w275_,
		_w497_,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w503_,
		_w504_,
		_w505_
	);
	LUT3 #(
		.INIT('h70)
	) name288 (
		_w302_,
		_w303_,
		_w502_,
		_w506_
	);
	LUT3 #(
		.INIT('h70)
	) name289 (
		_w307_,
		_w308_,
		_w488_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w506_,
		_w507_,
		_w508_
	);
	LUT4 #(
		.INIT('h1055)
	) name291 (
		_w489_,
		_w499_,
		_w505_,
		_w508_,
		_w509_
	);
	LUT3 #(
		.INIT('h08)
	) name292 (
		_w318_,
		_w319_,
		_w479_,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w476_,
		_w510_,
		_w511_
	);
	LUT4 #(
		.INIT('h0001)
	) name294 (
		_w468_,
		_w471_,
		_w476_,
		_w510_,
		_w512_
	);
	LUT4 #(
		.INIT('ha222)
	) name295 (
		_w463_,
		_w486_,
		_w509_,
		_w512_,
		_w513_
	);
	LUT4 #(
		.INIT('h65a5)
	) name296 (
		_w414_,
		_w452_,
		_w460_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		_w401_,
		_w398_,
		_w515_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w401_,
		_w398_,
		_w516_
	);
	LUT2 #(
		.INIT('h9)
	) name299 (
		_w401_,
		_w398_,
		_w517_
	);
	LUT4 #(
		.INIT('h9180)
	) name300 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w518_
	);
	LUT4 #(
		.INIT('h2e00)
	) name301 (
		_w224_,
		_w262_,
		_w514_,
		_w518_,
		_w519_
	);
	LUT4 #(
		.INIT('h0200)
	) name302 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w520_
	);
	LUT4 #(
		.INIT('h001f)
	) name303 (
		_w256_,
		_w258_,
		_w261_,
		_w520_,
		_w521_
	);
	LUT4 #(
		.INIT('h2220)
	) name304 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w522_
	);
	LUT3 #(
		.INIT('h40)
	) name305 (
		_w521_,
		_w522_,
		_w411_,
		_w523_
	);
	LUT4 #(
		.INIT('h4440)
	) name306 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w524_
	);
	LUT3 #(
		.INIT('h20)
	) name307 (
		_w401_,
		_w398_,
		_w399_,
		_w525_
	);
	LUT4 #(
		.INIT('h1f00)
	) name308 (
		_w256_,
		_w258_,
		_w261_,
		_w525_,
		_w526_
	);
	LUT3 #(
		.INIT('ha8)
	) name309 (
		_w224_,
		_w524_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w523_,
		_w527_,
		_w528_
	);
	LUT4 #(
		.INIT('h0010)
	) name311 (
		_w376_,
		_w375_,
		_w377_,
		_w449_,
		_w529_
	);
	LUT3 #(
		.INIT('h07)
	) name312 (
		_w361_,
		_w446_,
		_w529_,
		_w530_
	);
	LUT4 #(
		.INIT('h00ef)
	) name313 (
		_w365_,
		_w364_,
		_w366_,
		_w439_,
		_w531_
	);
	LUT4 #(
		.INIT('h1000)
	) name314 (
		_w365_,
		_w364_,
		_w366_,
		_w439_,
		_w532_
	);
	LUT3 #(
		.INIT('h07)
	) name315 (
		_w370_,
		_w371_,
		_w442_,
		_w533_
	);
	LUT3 #(
		.INIT('h45)
	) name316 (
		_w531_,
		_w532_,
		_w533_,
		_w534_
	);
	LUT4 #(
		.INIT('hef00)
	) name317 (
		_w376_,
		_w375_,
		_w377_,
		_w449_,
		_w535_
	);
	LUT3 #(
		.INIT('h71)
	) name318 (
		_w361_,
		_w446_,
		_w535_,
		_w536_
	);
	LUT3 #(
		.INIT('h0d)
	) name319 (
		_w530_,
		_w534_,
		_w536_,
		_w537_
	);
	LUT3 #(
		.INIT('h80)
	) name320 (
		_w370_,
		_w371_,
		_w442_,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w532_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w530_,
		_w539_,
		_w540_
	);
	LUT3 #(
		.INIT('h80)
	) name323 (
		_w345_,
		_w347_,
		_w418_,
		_w541_
	);
	LUT3 #(
		.INIT('h80)
	) name324 (
		_w341_,
		_w342_,
		_w423_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w541_,
		_w542_,
		_w543_
	);
	LUT3 #(
		.INIT('h80)
	) name326 (
		_w350_,
		_w352_,
		_w427_,
		_w544_
	);
	LUT3 #(
		.INIT('h07)
	) name327 (
		_w350_,
		_w352_,
		_w427_,
		_w545_
	);
	LUT3 #(
		.INIT('h07)
	) name328 (
		_w332_,
		_w334_,
		_w431_,
		_w546_
	);
	LUT3 #(
		.INIT('h54)
	) name329 (
		_w544_,
		_w545_,
		_w546_,
		_w547_
	);
	LUT3 #(
		.INIT('h07)
	) name330 (
		_w341_,
		_w342_,
		_w423_,
		_w548_
	);
	LUT3 #(
		.INIT('h07)
	) name331 (
		_w345_,
		_w347_,
		_w418_,
		_w549_
	);
	LUT3 #(
		.INIT('h23)
	) name332 (
		_w542_,
		_w548_,
		_w549_,
		_w550_
	);
	LUT3 #(
		.INIT('h70)
	) name333 (
		_w543_,
		_w547_,
		_w550_,
		_w551_
	);
	LUT3 #(
		.INIT('ha2)
	) name334 (
		_w537_,
		_w540_,
		_w551_,
		_w552_
	);
	LUT3 #(
		.INIT('h80)
	) name335 (
		_w332_,
		_w334_,
		_w431_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w544_,
		_w553_,
		_w554_
	);
	LUT4 #(
		.INIT('h0001)
	) name337 (
		_w541_,
		_w542_,
		_w544_,
		_w553_,
		_w555_
	);
	LUT3 #(
		.INIT('h80)
	) name338 (
		_w328_,
		_w330_,
		_w470_,
		_w556_
	);
	LUT3 #(
		.INIT('h80)
	) name339 (
		_w323_,
		_w325_,
		_w467_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w556_,
		_w557_,
		_w558_
	);
	LUT3 #(
		.INIT('h07)
	) name341 (
		_w312_,
		_w314_,
		_w475_,
		_w559_
	);
	LUT3 #(
		.INIT('h80)
	) name342 (
		_w312_,
		_w314_,
		_w475_,
		_w560_
	);
	LUT3 #(
		.INIT('h07)
	) name343 (
		_w318_,
		_w319_,
		_w479_,
		_w561_
	);
	LUT3 #(
		.INIT('h45)
	) name344 (
		_w559_,
		_w560_,
		_w561_,
		_w562_
	);
	LUT3 #(
		.INIT('h07)
	) name345 (
		_w328_,
		_w330_,
		_w470_,
		_w563_
	);
	LUT3 #(
		.INIT('h07)
	) name346 (
		_w323_,
		_w325_,
		_w467_,
		_w564_
	);
	LUT3 #(
		.INIT('h54)
	) name347 (
		_w556_,
		_w563_,
		_w564_,
		_w565_
	);
	LUT3 #(
		.INIT('h0d)
	) name348 (
		_w558_,
		_w562_,
		_w565_,
		_w566_
	);
	LUT3 #(
		.INIT('h07)
	) name349 (
		_w273_,
		_w275_,
		_w497_,
		_w567_
	);
	LUT3 #(
		.INIT('h07)
	) name350 (
		_w278_,
		_w279_,
		_w491_,
		_w568_
	);
	LUT3 #(
		.INIT('h80)
	) name351 (
		_w278_,
		_w279_,
		_w491_,
		_w569_
	);
	LUT3 #(
		.INIT('h07)
	) name352 (
		_w282_,
		_w283_,
		_w493_,
		_w570_
	);
	LUT3 #(
		.INIT('h45)
	) name353 (
		_w568_,
		_w569_,
		_w570_,
		_w571_
	);
	LUT4 #(
		.INIT('h080e)
	) name354 (
		_w280_,
		_w491_,
		_w567_,
		_w570_,
		_w572_
	);
	LUT3 #(
		.INIT('h80)
	) name355 (
		_w302_,
		_w303_,
		_w502_,
		_w573_
	);
	LUT3 #(
		.INIT('h80)
	) name356 (
		_w273_,
		_w275_,
		_w497_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w573_,
		_w574_,
		_w575_
	);
	LUT3 #(
		.INIT('h80)
	) name358 (
		_w307_,
		_w308_,
		_w488_,
		_w576_
	);
	LUT3 #(
		.INIT('h01)
	) name359 (
		_w573_,
		_w574_,
		_w576_,
		_w577_
	);
	LUT3 #(
		.INIT('h07)
	) name360 (
		_w307_,
		_w308_,
		_w488_,
		_w578_
	);
	LUT3 #(
		.INIT('h07)
	) name361 (
		_w302_,
		_w303_,
		_w502_,
		_w579_
	);
	LUT3 #(
		.INIT('h54)
	) name362 (
		_w576_,
		_w578_,
		_w579_,
		_w580_
	);
	LUT3 #(
		.INIT('h80)
	) name363 (
		_w318_,
		_w319_,
		_w479_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w560_,
		_w581_,
		_w582_
	);
	LUT4 #(
		.INIT('h0001)
	) name365 (
		_w556_,
		_w557_,
		_w560_,
		_w581_,
		_w583_
	);
	LUT4 #(
		.INIT('hf400)
	) name366 (
		_w572_,
		_w577_,
		_w580_,
		_w583_,
		_w584_
	);
	LUT4 #(
		.INIT('h8808)
	) name367 (
		_w540_,
		_w555_,
		_w566_,
		_w584_,
		_w585_
	);
	LUT4 #(
		.INIT('h2282)
	) name368 (
		_w262_,
		_w414_,
		_w552_,
		_w585_,
		_w586_
	);
	LUT4 #(
		.INIT('h0819)
	) name369 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w587_
	);
	LUT3 #(
		.INIT('he0)
	) name370 (
		_w263_,
		_w586_,
		_w587_,
		_w588_
	);
	LUT3 #(
		.INIT('h80)
	) name371 (
		_w491_,
		_w493_,
		_w497_,
		_w589_
	);
	LUT4 #(
		.INIT('h8000)
	) name372 (
		_w491_,
		_w493_,
		_w497_,
		_w502_,
		_w590_
	);
	LUT3 #(
		.INIT('h80)
	) name373 (
		_w479_,
		_w488_,
		_w590_,
		_w591_
	);
	LUT4 #(
		.INIT('h8000)
	) name374 (
		_w475_,
		_w479_,
		_w488_,
		_w590_,
		_w592_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w431_,
		_w470_,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		_w418_,
		_w427_,
		_w594_
	);
	LUT4 #(
		.INIT('h8000)
	) name377 (
		_w418_,
		_w423_,
		_w427_,
		_w442_,
		_w595_
	);
	LUT4 #(
		.INIT('h8000)
	) name378 (
		_w467_,
		_w592_,
		_w593_,
		_w595_,
		_w596_
	);
	LUT4 #(
		.INIT('h0800)
	) name379 (
		_w439_,
		_w446_,
		_w449_,
		_w596_,
		_w597_
	);
	LUT4 #(
		.INIT('h0040)
	) name380 (
		_w411_,
		_w439_,
		_w446_,
		_w449_,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		_w596_,
		_w598_,
		_w599_
	);
	LUT4 #(
		.INIT('h00a2)
	) name382 (
		_w262_,
		_w411_,
		_w597_,
		_w599_,
		_w600_
	);
	LUT4 #(
		.INIT('h0002)
	) name383 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w601_
	);
	LUT3 #(
		.INIT('he0)
	) name384 (
		_w263_,
		_w600_,
		_w601_,
		_w602_
	);
	LUT4 #(
		.INIT('h0100)
	) name385 (
		_w519_,
		_w588_,
		_w602_,
		_w528_,
		_w603_
	);
	LUT4 #(
		.INIT('h1511)
	) name386 (
		_w253_,
		_w254_,
		_w405_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		\reg3_reg[17]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w605_
	);
	LUT3 #(
		.INIT('h48)
	) name388 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w606_
	);
	LUT4 #(
		.INIT('h4080)
	) name389 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w224_,
		_w236_,
		_w607_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		_w605_,
		_w607_,
		_w608_
	);
	LUT3 #(
		.INIT('h2f)
	) name391 (
		\state_reg[0]/NET0131 ,
		_w604_,
		_w608_,
		_w609_
	);
	LUT4 #(
		.INIT('h8000)
	) name392 (
		_w221_,
		_w222_,
		_w286_,
		_w290_,
		_w610_
	);
	LUT4 #(
		.INIT('h8000)
	) name393 (
		_w221_,
		_w222_,
		_w286_,
		_w291_,
		_w611_
	);
	LUT3 #(
		.INIT('h6a)
	) name394 (
		\reg3_reg[23]/NET0131 ,
		_w287_,
		_w290_,
		_w612_
	);
	LUT3 #(
		.INIT('h20)
	) name395 (
		\reg2_reg[23]/NET0131 ,
		_w269_,
		_w272_,
		_w613_
	);
	LUT4 #(
		.INIT('hff35)
	) name396 (
		\reg0_reg[23]/NET0131 ,
		\reg1_reg[23]/NET0131 ,
		_w269_,
		_w272_,
		_w614_
	);
	LUT4 #(
		.INIT('h1300)
	) name397 (
		_w274_,
		_w613_,
		_w612_,
		_w614_,
		_w615_
	);
	LUT4 #(
		.INIT('hecff)
	) name398 (
		_w274_,
		_w613_,
		_w612_,
		_w614_,
		_w616_
	);
	LUT4 #(
		.INIT('h8000)
	) name399 (
		\reg3_reg[25]/NET0131 ,
		\reg3_reg[26]/NET0131 ,
		\reg3_reg[27]/NET0131 ,
		_w293_,
		_w617_
	);
	LUT2 #(
		.INIT('h6)
	) name400 (
		\reg3_reg[28]/NET0131 ,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		_w262_,
		_w618_,
		_w619_
	);
	LUT3 #(
		.INIT('ha8)
	) name402 (
		\datai[27]_pad ,
		_w266_,
		_w407_,
		_w620_
	);
	LUT4 #(
		.INIT('h78f0)
	) name403 (
		\reg3_reg[25]/NET0131 ,
		\reg3_reg[26]/NET0131 ,
		\reg3_reg[27]/NET0131 ,
		_w293_,
		_w621_
	);
	LUT3 #(
		.INIT('h20)
	) name404 (
		\reg2_reg[27]/NET0131 ,
		_w269_,
		_w272_,
		_w622_
	);
	LUT4 #(
		.INIT('hff35)
	) name405 (
		\reg0_reg[27]/NET0131 ,
		\reg1_reg[27]/NET0131 ,
		_w269_,
		_w272_,
		_w623_
	);
	LUT4 #(
		.INIT('h1300)
	) name406 (
		_w274_,
		_w622_,
		_w621_,
		_w623_,
		_w624_
	);
	LUT4 #(
		.INIT('hecff)
	) name407 (
		_w274_,
		_w622_,
		_w621_,
		_w623_,
		_w625_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		_w620_,
		_w624_,
		_w626_
	);
	LUT3 #(
		.INIT('ha8)
	) name409 (
		\datai[26]_pad ,
		_w266_,
		_w407_,
		_w627_
	);
	LUT3 #(
		.INIT('h6c)
	) name410 (
		\reg3_reg[25]/NET0131 ,
		\reg3_reg[26]/NET0131 ,
		_w293_,
		_w628_
	);
	LUT3 #(
		.INIT('h02)
	) name411 (
		\reg0_reg[26]/NET0131 ,
		_w269_,
		_w272_,
		_w629_
	);
	LUT4 #(
		.INIT('hf35f)
	) name412 (
		\reg1_reg[26]/NET0131 ,
		\reg2_reg[26]/NET0131 ,
		_w269_,
		_w272_,
		_w630_
	);
	LUT4 #(
		.INIT('h1300)
	) name413 (
		_w274_,
		_w629_,
		_w628_,
		_w630_,
		_w631_
	);
	LUT4 #(
		.INIT('hecff)
	) name414 (
		_w274_,
		_w629_,
		_w628_,
		_w630_,
		_w632_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		_w627_,
		_w631_,
		_w633_
	);
	LUT4 #(
		.INIT('h0777)
	) name416 (
		_w620_,
		_w624_,
		_w627_,
		_w631_,
		_w634_
	);
	LUT3 #(
		.INIT('ha8)
	) name417 (
		\datai[25]_pad ,
		_w266_,
		_w407_,
		_w635_
	);
	LUT2 #(
		.INIT('h6)
	) name418 (
		\reg3_reg[25]/NET0131 ,
		_w293_,
		_w636_
	);
	LUT4 #(
		.INIT('h4080)
	) name419 (
		\reg3_reg[25]/NET0131 ,
		_w269_,
		_w272_,
		_w293_,
		_w637_
	);
	LUT3 #(
		.INIT('h20)
	) name420 (
		\reg2_reg[25]/NET0131 ,
		_w269_,
		_w272_,
		_w638_
	);
	LUT4 #(
		.INIT('hff35)
	) name421 (
		\reg0_reg[25]/NET0131 ,
		\reg1_reg[25]/NET0131 ,
		_w269_,
		_w272_,
		_w639_
	);
	LUT3 #(
		.INIT('h10)
	) name422 (
		_w638_,
		_w637_,
		_w639_,
		_w640_
	);
	LUT3 #(
		.INIT('hef)
	) name423 (
		_w638_,
		_w637_,
		_w639_,
		_w641_
	);
	LUT4 #(
		.INIT('h0200)
	) name424 (
		_w635_,
		_w638_,
		_w637_,
		_w639_,
		_w642_
	);
	LUT3 #(
		.INIT('ha8)
	) name425 (
		\datai[24]_pad ,
		_w266_,
		_w407_,
		_w643_
	);
	LUT3 #(
		.INIT('h32)
	) name426 (
		\reg3_reg[24]/NET0131 ,
		_w293_,
		_w611_,
		_w644_
	);
	LUT3 #(
		.INIT('h20)
	) name427 (
		\reg2_reg[24]/NET0131 ,
		_w269_,
		_w272_,
		_w645_
	);
	LUT4 #(
		.INIT('hff35)
	) name428 (
		\reg0_reg[24]/NET0131 ,
		\reg1_reg[24]/NET0131 ,
		_w269_,
		_w272_,
		_w646_
	);
	LUT4 #(
		.INIT('h1300)
	) name429 (
		_w274_,
		_w645_,
		_w644_,
		_w646_,
		_w647_
	);
	LUT4 #(
		.INIT('hecff)
	) name430 (
		_w274_,
		_w645_,
		_w644_,
		_w646_,
		_w648_
	);
	LUT3 #(
		.INIT('h15)
	) name431 (
		_w642_,
		_w643_,
		_w647_,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		_w634_,
		_w649_,
		_w650_
	);
	LUT3 #(
		.INIT('ha8)
	) name433 (
		\datai[23]_pad ,
		_w266_,
		_w407_,
		_w651_
	);
	LUT3 #(
		.INIT('ha8)
	) name434 (
		\datai[22]_pad ,
		_w266_,
		_w407_,
		_w652_
	);
	LUT4 #(
		.INIT('h8000)
	) name435 (
		_w221_,
		_w222_,
		_w286_,
		_w289_,
		_w653_
	);
	LUT3 #(
		.INIT('h32)
	) name436 (
		\reg3_reg[22]/NET0131 ,
		_w610_,
		_w653_,
		_w654_
	);
	LUT3 #(
		.INIT('h08)
	) name437 (
		\reg1_reg[22]/NET0131 ,
		_w269_,
		_w272_,
		_w655_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name438 (
		\reg0_reg[22]/NET0131 ,
		\reg2_reg[22]/NET0131 ,
		_w269_,
		_w272_,
		_w656_
	);
	LUT4 #(
		.INIT('h1300)
	) name439 (
		_w274_,
		_w655_,
		_w654_,
		_w656_,
		_w657_
	);
	LUT4 #(
		.INIT('hecff)
	) name440 (
		_w274_,
		_w655_,
		_w654_,
		_w656_,
		_w658_
	);
	LUT4 #(
		.INIT('h0777)
	) name441 (
		_w615_,
		_w651_,
		_w652_,
		_w657_,
		_w659_
	);
	LUT3 #(
		.INIT('ha8)
	) name442 (
		\datai[21]_pad ,
		_w266_,
		_w407_,
		_w660_
	);
	LUT4 #(
		.INIT('h8000)
	) name443 (
		_w221_,
		_w222_,
		_w286_,
		_w288_,
		_w661_
	);
	LUT3 #(
		.INIT('h32)
	) name444 (
		\reg3_reg[21]/NET0131 ,
		_w653_,
		_w661_,
		_w662_
	);
	LUT3 #(
		.INIT('h20)
	) name445 (
		\reg2_reg[21]/NET0131 ,
		_w269_,
		_w272_,
		_w663_
	);
	LUT4 #(
		.INIT('hff35)
	) name446 (
		\reg0_reg[21]/NET0131 ,
		\reg1_reg[21]/NET0131 ,
		_w269_,
		_w272_,
		_w664_
	);
	LUT4 #(
		.INIT('h1300)
	) name447 (
		_w274_,
		_w663_,
		_w662_,
		_w664_,
		_w665_
	);
	LUT4 #(
		.INIT('hecff)
	) name448 (
		_w274_,
		_w663_,
		_w662_,
		_w664_,
		_w666_
	);
	LUT3 #(
		.INIT('ha8)
	) name449 (
		\datai[20]_pad ,
		_w266_,
		_w407_,
		_w667_
	);
	LUT3 #(
		.INIT('h6c)
	) name450 (
		\reg3_reg[19]/NET0131 ,
		\reg3_reg[20]/NET0131 ,
		_w287_,
		_w668_
	);
	LUT3 #(
		.INIT('h08)
	) name451 (
		\reg1_reg[20]/NET0131 ,
		_w269_,
		_w272_,
		_w669_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name452 (
		\reg0_reg[20]/NET0131 ,
		\reg2_reg[20]/NET0131 ,
		_w269_,
		_w272_,
		_w670_
	);
	LUT4 #(
		.INIT('h1300)
	) name453 (
		_w274_,
		_w669_,
		_w668_,
		_w670_,
		_w671_
	);
	LUT4 #(
		.INIT('hecff)
	) name454 (
		_w274_,
		_w669_,
		_w668_,
		_w670_,
		_w672_
	);
	LUT4 #(
		.INIT('h0777)
	) name455 (
		_w660_,
		_w665_,
		_w667_,
		_w671_,
		_w673_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		_w659_,
		_w673_,
		_w674_
	);
	LUT4 #(
		.INIT('h8000)
	) name457 (
		_w634_,
		_w649_,
		_w659_,
		_w673_,
		_w675_
	);
	LUT3 #(
		.INIT('he0)
	) name458 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[17]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w676_
	);
	LUT3 #(
		.INIT('h56)
	) name459 (
		\IR_reg[18]/NET0131 ,
		_w238_,
		_w676_,
		_w677_
	);
	LUT4 #(
		.INIT('haba8)
	) name460 (
		\datai[18]_pad ,
		_w266_,
		_w407_,
		_w677_,
		_w678_
	);
	LUT4 #(
		.INIT('h1000)
	) name461 (
		_w389_,
		_w388_,
		_w390_,
		_w678_,
		_w679_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name462 (
		\reg3_reg[19]/NET0131 ,
		_w221_,
		_w222_,
		_w286_,
		_w680_
	);
	LUT3 #(
		.INIT('h80)
	) name463 (
		_w269_,
		_w272_,
		_w680_,
		_w681_
	);
	LUT3 #(
		.INIT('h02)
	) name464 (
		\reg0_reg[19]/NET0131 ,
		_w269_,
		_w272_,
		_w682_
	);
	LUT4 #(
		.INIT('hf35f)
	) name465 (
		\reg1_reg[19]/NET0131 ,
		\reg2_reg[19]/NET0131 ,
		_w269_,
		_w272_,
		_w683_
	);
	LUT3 #(
		.INIT('h10)
	) name466 (
		_w682_,
		_w681_,
		_w683_,
		_w684_
	);
	LUT3 #(
		.INIT('hef)
	) name467 (
		_w682_,
		_w681_,
		_w683_,
		_w685_
	);
	LUT4 #(
		.INIT('h5553)
	) name468 (
		\datai[19]_pad ,
		_w403_,
		_w266_,
		_w407_,
		_w686_
	);
	LUT4 #(
		.INIT('h0010)
	) name469 (
		_w682_,
		_w681_,
		_w683_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w679_,
		_w687_,
		_w688_
	);
	LUT4 #(
		.INIT('h0200)
	) name471 (
		_w411_,
		_w382_,
		_w381_,
		_w383_,
		_w689_
	);
	LUT3 #(
		.INIT('h0d)
	) name472 (
		_w361_,
		_w446_,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w688_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w419_,
		_w428_,
		_w692_
	);
	LUT3 #(
		.INIT('h32)
	) name475 (
		_w432_,
		_w461_,
		_w483_,
		_w693_
	);
	LUT3 #(
		.INIT('h0b)
	) name476 (
		_w419_,
		_w429_,
		_w435_,
		_w694_
	);
	LUT3 #(
		.INIT('h70)
	) name477 (
		_w692_,
		_w693_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w468_,
		_w476_,
		_w696_
	);
	LUT3 #(
		.INIT('hb2)
	) name479 (
		_w280_,
		_w491_,
		_w494_,
		_w697_
	);
	LUT3 #(
		.INIT('h32)
	) name480 (
		_w498_,
		_w503_,
		_w506_,
		_w698_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w489_,
		_w510_,
		_w699_
	);
	LUT4 #(
		.INIT('hf200)
	) name482 (
		_w505_,
		_w697_,
		_w698_,
		_w699_,
		_w700_
	);
	LUT3 #(
		.INIT('h0e)
	) name483 (
		_w480_,
		_w507_,
		_w510_,
		_w701_
	);
	LUT3 #(
		.INIT('h0b)
	) name484 (
		_w468_,
		_w477_,
		_w484_,
		_w702_
	);
	LUT3 #(
		.INIT('h70)
	) name485 (
		_w696_,
		_w701_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w461_,
		_w471_,
		_w704_
	);
	LUT4 #(
		.INIT('h0001)
	) name487 (
		_w419_,
		_w428_,
		_w461_,
		_w471_,
		_w705_
	);
	LUT4 #(
		.INIT('h8f00)
	) name488 (
		_w696_,
		_w700_,
		_w703_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		_w440_,
		_w450_,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w424_,
		_w443_,
		_w708_
	);
	LUT4 #(
		.INIT('h0001)
	) name491 (
		_w424_,
		_w440_,
		_w443_,
		_w450_,
		_w709_
	);
	LUT4 #(
		.INIT('ha200)
	) name492 (
		_w691_,
		_w695_,
		_w706_,
		_w709_,
		_w710_
	);
	LUT3 #(
		.INIT('h0d)
	) name493 (
		_w434_,
		_w443_,
		_w454_,
		_w711_
	);
	LUT3 #(
		.INIT('h54)
	) name494 (
		_w450_,
		_w453_,
		_w457_,
		_w712_
	);
	LUT3 #(
		.INIT('h0d)
	) name495 (
		_w707_,
		_w711_,
		_w712_,
		_w713_
	);
	LUT4 #(
		.INIT('h5455)
	) name496 (
		_w411_,
		_w382_,
		_w381_,
		_w383_,
		_w714_
	);
	LUT4 #(
		.INIT('h0f04)
	) name497 (
		_w361_,
		_w446_,
		_w689_,
		_w714_,
		_w715_
	);
	LUT4 #(
		.INIT('hef00)
	) name498 (
		_w682_,
		_w681_,
		_w683_,
		_w686_,
		_w716_
	);
	LUT4 #(
		.INIT('h00ef)
	) name499 (
		_w389_,
		_w388_,
		_w390_,
		_w678_,
		_w717_
	);
	LUT3 #(
		.INIT('h54)
	) name500 (
		_w687_,
		_w716_,
		_w717_,
		_w718_
	);
	LUT3 #(
		.INIT('h07)
	) name501 (
		_w688_,
		_w715_,
		_w718_,
		_w719_
	);
	LUT3 #(
		.INIT('hd0)
	) name502 (
		_w691_,
		_w713_,
		_w719_,
		_w720_
	);
	LUT4 #(
		.INIT('h1117)
	) name503 (
		_w660_,
		_w665_,
		_w667_,
		_w671_,
		_w721_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w615_,
		_w651_,
		_w722_
	);
	LUT4 #(
		.INIT('heee8)
	) name505 (
		_w615_,
		_w651_,
		_w652_,
		_w657_,
		_w723_
	);
	LUT3 #(
		.INIT('h70)
	) name506 (
		_w659_,
		_w721_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w620_,
		_w624_,
		_w725_
	);
	LUT4 #(
		.INIT('heee0)
	) name508 (
		_w620_,
		_w624_,
		_w627_,
		_w631_,
		_w726_
	);
	LUT4 #(
		.INIT('h5455)
	) name509 (
		_w635_,
		_w638_,
		_w637_,
		_w639_,
		_w727_
	);
	LUT3 #(
		.INIT('h0e)
	) name510 (
		_w643_,
		_w647_,
		_w727_,
		_w728_
	);
	LUT4 #(
		.INIT('h5501)
	) name511 (
		_w642_,
		_w643_,
		_w647_,
		_w727_,
		_w729_
	);
	LUT4 #(
		.INIT('h1505)
	) name512 (
		_w626_,
		_w633_,
		_w726_,
		_w729_,
		_w730_
	);
	LUT3 #(
		.INIT('h0d)
	) name513 (
		_w650_,
		_w724_,
		_w730_,
		_w731_
	);
	LUT4 #(
		.INIT('h7500)
	) name514 (
		_w675_,
		_w710_,
		_w720_,
		_w731_,
		_w732_
	);
	LUT3 #(
		.INIT('ha8)
	) name515 (
		\datai[28]_pad ,
		_w266_,
		_w407_,
		_w733_
	);
	LUT3 #(
		.INIT('h48)
	) name516 (
		\reg3_reg[28]/NET0131 ,
		_w274_,
		_w617_,
		_w734_
	);
	LUT3 #(
		.INIT('h20)
	) name517 (
		\reg2_reg[28]/NET0131 ,
		_w269_,
		_w272_,
		_w735_
	);
	LUT4 #(
		.INIT('hff35)
	) name518 (
		\reg0_reg[28]/NET0131 ,
		\reg1_reg[28]/NET0131 ,
		_w269_,
		_w272_,
		_w736_
	);
	LUT2 #(
		.INIT('h4)
	) name519 (
		_w735_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name520 (
		_w734_,
		_w737_,
		_w738_
	);
	LUT3 #(
		.INIT('h10)
	) name521 (
		_w733_,
		_w734_,
		_w737_,
		_w739_
	);
	LUT3 #(
		.INIT('h8a)
	) name522 (
		_w733_,
		_w734_,
		_w737_,
		_w740_
	);
	LUT3 #(
		.INIT('h65)
	) name523 (
		_w733_,
		_w734_,
		_w737_,
		_w741_
	);
	LUT4 #(
		.INIT('h3113)
	) name524 (
		_w262_,
		_w619_,
		_w732_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w538_,
		_w542_,
		_w743_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		_w529_,
		_w532_,
		_w744_
	);
	LUT4 #(
		.INIT('h0001)
	) name527 (
		_w529_,
		_w532_,
		_w538_,
		_w542_,
		_w745_
	);
	LUT3 #(
		.INIT('h13)
	) name528 (
		_w361_,
		_w412_,
		_w446_,
		_w746_
	);
	LUT4 #(
		.INIT('h1000)
	) name529 (
		_w682_,
		_w681_,
		_w683_,
		_w686_,
		_w747_
	);
	LUT4 #(
		.INIT('h0010)
	) name530 (
		_w389_,
		_w388_,
		_w390_,
		_w678_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w747_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h8)
	) name532 (
		_w746_,
		_w749_,
		_w750_
	);
	LUT3 #(
		.INIT('h80)
	) name533 (
		_w745_,
		_w746_,
		_w749_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		_w541_,
		_w544_,
		_w752_
	);
	LUT3 #(
		.INIT('h32)
	) name535 (
		_w546_,
		_w553_,
		_w563_,
		_w753_
	);
	LUT3 #(
		.INIT('h0b)
	) name536 (
		_w541_,
		_w545_,
		_w549_,
		_w754_
	);
	LUT3 #(
		.INIT('h70)
	) name537 (
		_w752_,
		_w753_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w557_,
		_w560_,
		_w756_
	);
	LUT3 #(
		.INIT('h32)
	) name539 (
		_w567_,
		_w573_,
		_w579_,
		_w757_
	);
	LUT3 #(
		.INIT('h0b)
	) name540 (
		_w571_,
		_w575_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w581_,
		_w576_,
		_w759_
	);
	LUT4 #(
		.INIT('hf400)
	) name542 (
		_w571_,
		_w575_,
		_w757_,
		_w759_,
		_w760_
	);
	LUT3 #(
		.INIT('h45)
	) name543 (
		_w561_,
		_w581_,
		_w578_,
		_w761_
	);
	LUT3 #(
		.INIT('h0b)
	) name544 (
		_w557_,
		_w559_,
		_w564_,
		_w762_
	);
	LUT3 #(
		.INIT('hd0)
	) name545 (
		_w756_,
		_w761_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		_w553_,
		_w556_,
		_w764_
	);
	LUT4 #(
		.INIT('h0001)
	) name547 (
		_w541_,
		_w544_,
		_w553_,
		_w556_,
		_w765_
	);
	LUT4 #(
		.INIT('h8f00)
	) name548 (
		_w756_,
		_w760_,
		_w763_,
		_w765_,
		_w766_
	);
	LUT3 #(
		.INIT('h45)
	) name549 (
		_w533_,
		_w538_,
		_w548_,
		_w767_
	);
	LUT3 #(
		.INIT('h0b)
	) name550 (
		_w529_,
		_w531_,
		_w535_,
		_w768_
	);
	LUT3 #(
		.INIT('hd0)
	) name551 (
		_w744_,
		_w767_,
		_w768_,
		_w769_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name552 (
		_w361_,
		_w412_,
		_w413_,
		_w446_,
		_w770_
	);
	LUT4 #(
		.INIT('h00ef)
	) name553 (
		_w682_,
		_w681_,
		_w683_,
		_w686_,
		_w771_
	);
	LUT4 #(
		.INIT('hef00)
	) name554 (
		_w389_,
		_w388_,
		_w390_,
		_w678_,
		_w772_
	);
	LUT3 #(
		.INIT('h23)
	) name555 (
		_w747_,
		_w771_,
		_w772_,
		_w773_
	);
	LUT3 #(
		.INIT('hd0)
	) name556 (
		_w749_,
		_w770_,
		_w773_,
		_w774_
	);
	LUT3 #(
		.INIT('hd0)
	) name557 (
		_w750_,
		_w769_,
		_w774_,
		_w775_
	);
	LUT4 #(
		.INIT('h5d00)
	) name558 (
		_w751_,
		_w755_,
		_w766_,
		_w775_,
		_w776_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name559 (
		_w660_,
		_w665_,
		_w667_,
		_w671_,
		_w777_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name560 (
		_w615_,
		_w651_,
		_w652_,
		_w657_,
		_w778_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		_w777_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		_w627_,
		_w631_,
		_w780_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name563 (
		_w620_,
		_w624_,
		_w627_,
		_w631_,
		_w781_
	);
	LUT4 #(
		.INIT('h0100)
	) name564 (
		_w635_,
		_w638_,
		_w637_,
		_w639_,
		_w782_
	);
	LUT3 #(
		.INIT('h0b)
	) name565 (
		_w643_,
		_w647_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h8)
	) name566 (
		_w781_,
		_w783_,
		_w784_
	);
	LUT4 #(
		.INIT('h8000)
	) name567 (
		_w777_,
		_w778_,
		_w781_,
		_w783_,
		_w785_
	);
	LUT4 #(
		.INIT('hdd4d)
	) name568 (
		_w660_,
		_w665_,
		_w667_,
		_w671_,
		_w786_
	);
	LUT4 #(
		.INIT('hbb2b)
	) name569 (
		_w615_,
		_w651_,
		_w652_,
		_w657_,
		_w787_
	);
	LUT3 #(
		.INIT('hd0)
	) name570 (
		_w778_,
		_w786_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h2)
	) name571 (
		_w620_,
		_w624_,
		_w789_
	);
	LUT2 #(
		.INIT('h2)
	) name572 (
		_w627_,
		_w631_,
		_w790_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name573 (
		_w635_,
		_w638_,
		_w637_,
		_w639_,
		_w791_
	);
	LUT4 #(
		.INIT('h00fd)
	) name574 (
		_w643_,
		_w647_,
		_w782_,
		_w791_,
		_w792_
	);
	LUT4 #(
		.INIT('h1311)
	) name575 (
		_w781_,
		_w789_,
		_w790_,
		_w792_,
		_w793_
	);
	LUT3 #(
		.INIT('hd0)
	) name576 (
		_w784_,
		_w788_,
		_w793_,
		_w794_
	);
	LUT4 #(
		.INIT('h65aa)
	) name577 (
		_w741_,
		_w776_,
		_w785_,
		_w794_,
		_w795_
	);
	LUT4 #(
		.INIT('h40c8)
	) name578 (
		_w262_,
		_w587_,
		_w618_,
		_w795_,
		_w796_
	);
	LUT4 #(
		.INIT('h111f)
	) name579 (
		\datai[25]_pad ,
		\datai[26]_pad ,
		_w266_,
		_w407_,
		_w797_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		_w678_,
		_w686_,
		_w798_
	);
	LUT3 #(
		.INIT('h80)
	) name581 (
		_w596_,
		_w598_,
		_w798_,
		_w799_
	);
	LUT4 #(
		.INIT('h111f)
	) name582 (
		\datai[21]_pad ,
		\datai[22]_pad ,
		_w266_,
		_w407_,
		_w800_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		_w667_,
		_w800_,
		_w801_
	);
	LUT3 #(
		.INIT('h10)
	) name584 (
		_w651_,
		_w667_,
		_w800_,
		_w802_
	);
	LUT4 #(
		.INIT('h0100)
	) name585 (
		_w643_,
		_w651_,
		_w667_,
		_w800_,
		_w803_
	);
	LUT4 #(
		.INIT('h8000)
	) name586 (
		_w596_,
		_w598_,
		_w798_,
		_w803_,
		_w804_
	);
	LUT4 #(
		.INIT('h111f)
	) name587 (
		\datai[27]_pad ,
		\datai[28]_pad ,
		_w266_,
		_w407_,
		_w805_
	);
	LUT2 #(
		.INIT('h8)
	) name588 (
		_w797_,
		_w805_,
		_w806_
	);
	LUT4 #(
		.INIT('h6333)
	) name589 (
		_w620_,
		_w733_,
		_w797_,
		_w804_,
		_w807_
	);
	LUT4 #(
		.INIT('hc840)
	) name590 (
		_w262_,
		_w601_,
		_w618_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name591 (
		_w657_,
		_w665_,
		_w809_
	);
	LUT4 #(
		.INIT('h0001)
	) name592 (
		_w615_,
		_w657_,
		_w665_,
		_w671_,
		_w810_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		_w647_,
		_w684_,
		_w811_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		_w810_,
		_w811_,
		_w812_
	);
	LUT3 #(
		.INIT('h40)
	) name595 (
		_w640_,
		_w810_,
		_w811_,
		_w813_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w624_,
		_w631_,
		_w814_
	);
	LUT4 #(
		.INIT('h1011)
	) name597 (
		_w384_,
		_w391_,
		_w734_,
		_w737_,
		_w815_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		_w814_,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		_w813_,
		_w816_,
		_w817_
	);
	LUT3 #(
		.INIT('h08)
	) name600 (
		\reg1_reg[29]/NET0131 ,
		_w269_,
		_w272_,
		_w818_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name601 (
		\reg0_reg[29]/NET0131 ,
		\reg2_reg[29]/NET0131 ,
		_w269_,
		_w272_,
		_w819_
	);
	LUT3 #(
		.INIT('h10)
	) name602 (
		_w296_,
		_w818_,
		_w819_,
		_w820_
	);
	LUT3 #(
		.INIT('hef)
	) name603 (
		_w296_,
		_w818_,
		_w819_,
		_w821_
	);
	LUT4 #(
		.INIT('h4015)
	) name604 (
		_w266_,
		_w380_,
		_w817_,
		_w820_,
		_w822_
	);
	LUT2 #(
		.INIT('h2)
	) name605 (
		_w266_,
		_w624_,
		_w823_
	);
	LUT4 #(
		.INIT('h1113)
	) name606 (
		_w262_,
		_w619_,
		_w822_,
		_w823_,
		_w824_
	);
	LUT3 #(
		.INIT('he0)
	) name607 (
		_w524_,
		_w526_,
		_w618_,
		_w825_
	);
	LUT3 #(
		.INIT('h40)
	) name608 (
		_w521_,
		_w522_,
		_w733_,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		_w825_,
		_w826_,
		_w827_
	);
	LUT4 #(
		.INIT('h3100)
	) name610 (
		_w404_,
		_w808_,
		_w824_,
		_w827_,
		_w828_
	);
	LUT4 #(
		.INIT('h0d00)
	) name611 (
		_w518_,
		_w742_,
		_w796_,
		_w828_,
		_w829_
	);
	LUT3 #(
		.INIT('h48)
	) name612 (
		\reg3_reg[28]/NET0131 ,
		_w252_,
		_w617_,
		_w830_
	);
	LUT4 #(
		.INIT('haa08)
	) name613 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w829_,
		_w830_,
		_w831_
	);
	LUT4 #(
		.INIT('h9d5d)
	) name614 (
		\reg3_reg[28]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w237_,
		_w617_,
		_w832_
	);
	LUT2 #(
		.INIT('hb)
	) name615 (
		_w831_,
		_w832_,
		_w833_
	);
	LUT4 #(
		.INIT('h1f00)
	) name616 (
		_w256_,
		_w258_,
		_w261_,
		_w621_,
		_w834_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		_w412_,
		_w748_,
		_w835_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		_w530_,
		_w835_,
		_w836_
	);
	LUT4 #(
		.INIT('haa20)
	) name619 (
		_w582_,
		_w572_,
		_w577_,
		_w580_,
		_w837_
	);
	LUT4 #(
		.INIT('h0001)
	) name620 (
		_w544_,
		_w553_,
		_w556_,
		_w557_,
		_w838_
	);
	LUT3 #(
		.INIT('h15)
	) name621 (
		_w547_,
		_w554_,
		_w565_,
		_w839_
	);
	LUT4 #(
		.INIT('h2f00)
	) name622 (
		_w562_,
		_w837_,
		_w838_,
		_w839_,
		_w840_
	);
	LUT4 #(
		.INIT('h0001)
	) name623 (
		_w532_,
		_w538_,
		_w541_,
		_w542_,
		_w841_
	);
	LUT3 #(
		.INIT('ha2)
	) name624 (
		_w534_,
		_w539_,
		_w550_,
		_w842_
	);
	LUT3 #(
		.INIT('h0d)
	) name625 (
		_w413_,
		_w748_,
		_w772_,
		_w843_
	);
	LUT3 #(
		.INIT('h70)
	) name626 (
		_w536_,
		_w835_,
		_w843_,
		_w844_
	);
	LUT3 #(
		.INIT('hd0)
	) name627 (
		_w836_,
		_w842_,
		_w844_,
		_w845_
	);
	LUT4 #(
		.INIT('hdf00)
	) name628 (
		_w836_,
		_w840_,
		_w841_,
		_w845_,
		_w846_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name629 (
		_w652_,
		_w657_,
		_w660_,
		_w665_,
		_w847_
	);
	LUT3 #(
		.INIT('h0b)
	) name630 (
		_w667_,
		_w671_,
		_w747_,
		_w848_
	);
	LUT2 #(
		.INIT('h8)
	) name631 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT4 #(
		.INIT('hcf45)
	) name632 (
		_w615_,
		_w643_,
		_w647_,
		_w651_,
		_w850_
	);
	LUT3 #(
		.INIT('h0b)
	) name633 (
		_w627_,
		_w631_,
		_w782_,
		_w851_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		_w850_,
		_w851_,
		_w852_
	);
	LUT4 #(
		.INIT('h8000)
	) name635 (
		_w847_,
		_w848_,
		_w850_,
		_w851_,
		_w853_
	);
	LUT3 #(
		.INIT('h4d)
	) name636 (
		_w667_,
		_w671_,
		_w771_,
		_w854_
	);
	LUT4 #(
		.INIT('hdd4d)
	) name637 (
		_w652_,
		_w657_,
		_w660_,
		_w665_,
		_w855_
	);
	LUT3 #(
		.INIT('hd0)
	) name638 (
		_w847_,
		_w854_,
		_w855_,
		_w856_
	);
	LUT3 #(
		.INIT('h0d)
	) name639 (
		_w627_,
		_w631_,
		_w791_,
		_w857_
	);
	LUT4 #(
		.INIT('hb2f3)
	) name640 (
		_w615_,
		_w643_,
		_w647_,
		_w651_,
		_w858_
	);
	LUT4 #(
		.INIT('h0515)
	) name641 (
		_w780_,
		_w782_,
		_w857_,
		_w858_,
		_w859_
	);
	LUT3 #(
		.INIT('h0d)
	) name642 (
		_w852_,
		_w856_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h9)
	) name643 (
		_w620_,
		_w624_,
		_w861_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name644 (
		_w846_,
		_w853_,
		_w860_,
		_w861_,
		_w862_
	);
	LUT4 #(
		.INIT('h40c8)
	) name645 (
		_w262_,
		_w587_,
		_w621_,
		_w862_,
		_w863_
	);
	LUT4 #(
		.INIT('h0001)
	) name646 (
		_w428_,
		_w461_,
		_w468_,
		_w471_,
		_w864_
	);
	LUT4 #(
		.INIT('hea00)
	) name647 (
		_w482_,
		_w509_,
		_w511_,
		_w864_,
		_w865_
	);
	LUT3 #(
		.INIT('h15)
	) name648 (
		_w433_,
		_w462_,
		_w485_,
		_w866_
	);
	LUT2 #(
		.INIT('h1)
	) name649 (
		_w679_,
		_w689_,
		_w867_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		_w451_,
		_w867_,
		_w868_
	);
	LUT4 #(
		.INIT('h0001)
	) name651 (
		_w419_,
		_w424_,
		_w440_,
		_w443_,
		_w869_
	);
	LUT3 #(
		.INIT('h80)
	) name652 (
		_w451_,
		_w867_,
		_w869_,
		_w870_
	);
	LUT3 #(
		.INIT('h07)
	) name653 (
		_w436_,
		_w444_,
		_w456_,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w714_,
		_w717_,
		_w872_
	);
	LUT3 #(
		.INIT('h54)
	) name655 (
		_w679_,
		_w714_,
		_w717_,
		_w873_
	);
	LUT3 #(
		.INIT('h07)
	) name656 (
		_w458_,
		_w867_,
		_w873_,
		_w874_
	);
	LUT3 #(
		.INIT('hd0)
	) name657 (
		_w868_,
		_w871_,
		_w874_,
		_w875_
	);
	LUT4 #(
		.INIT('h4f00)
	) name658 (
		_w865_,
		_w866_,
		_w870_,
		_w875_,
		_w876_
	);
	LUT3 #(
		.INIT('h07)
	) name659 (
		_w667_,
		_w671_,
		_w687_,
		_w877_
	);
	LUT4 #(
		.INIT('h0777)
	) name660 (
		_w652_,
		_w657_,
		_w660_,
		_w665_,
		_w878_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		_w877_,
		_w878_,
		_w879_
	);
	LUT4 #(
		.INIT('h153f)
	) name662 (
		_w615_,
		_w643_,
		_w647_,
		_w651_,
		_w880_
	);
	LUT3 #(
		.INIT('h07)
	) name663 (
		_w627_,
		_w631_,
		_w642_,
		_w881_
	);
	LUT2 #(
		.INIT('h8)
	) name664 (
		_w880_,
		_w881_,
		_w882_
	);
	LUT4 #(
		.INIT('h8000)
	) name665 (
		_w877_,
		_w878_,
		_w880_,
		_w881_,
		_w883_
	);
	LUT3 #(
		.INIT('h0e)
	) name666 (
		_w667_,
		_w671_,
		_w716_,
		_w884_
	);
	LUT3 #(
		.INIT('h71)
	) name667 (
		_w667_,
		_w671_,
		_w716_,
		_w885_
	);
	LUT4 #(
		.INIT('heee0)
	) name668 (
		_w652_,
		_w657_,
		_w660_,
		_w665_,
		_w886_
	);
	LUT4 #(
		.INIT('h1117)
	) name669 (
		_w652_,
		_w657_,
		_w660_,
		_w665_,
		_w887_
	);
	LUT3 #(
		.INIT('h07)
	) name670 (
		_w878_,
		_w885_,
		_w887_,
		_w888_
	);
	LUT3 #(
		.INIT('h0e)
	) name671 (
		_w627_,
		_w631_,
		_w727_,
		_w889_
	);
	LUT3 #(
		.INIT('h71)
	) name672 (
		_w627_,
		_w631_,
		_w727_,
		_w890_
	);
	LUT4 #(
		.INIT('hfce8)
	) name673 (
		_w615_,
		_w643_,
		_w647_,
		_w651_,
		_w891_
	);
	LUT3 #(
		.INIT('h31)
	) name674 (
		_w881_,
		_w890_,
		_w891_,
		_w892_
	);
	LUT3 #(
		.INIT('hd0)
	) name675 (
		_w882_,
		_w888_,
		_w892_,
		_w893_
	);
	LUT4 #(
		.INIT('h9a55)
	) name676 (
		_w861_,
		_w876_,
		_w883_,
		_w893_,
		_w894_
	);
	LUT4 #(
		.INIT('h40c8)
	) name677 (
		_w262_,
		_w518_,
		_w621_,
		_w894_,
		_w895_
	);
	LUT3 #(
		.INIT('h01)
	) name678 (
		_w384_,
		_w391_,
		_w684_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name679 (
		_w379_,
		_w896_,
		_w897_
	);
	LUT3 #(
		.INIT('h80)
	) name680 (
		_w339_,
		_w356_,
		_w897_,
		_w898_
	);
	LUT4 #(
		.INIT('h8000)
	) name681 (
		_w339_,
		_w356_,
		_w810_,
		_w897_,
		_w899_
	);
	LUT4 #(
		.INIT('h0001)
	) name682 (
		_w624_,
		_w631_,
		_w640_,
		_w647_,
		_w900_
	);
	LUT4 #(
		.INIT('h1444)
	) name683 (
		_w266_,
		_w738_,
		_w899_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		_w266_,
		_w631_,
		_w902_
	);
	LUT4 #(
		.INIT('h3331)
	) name685 (
		_w262_,
		_w834_,
		_w901_,
		_w902_,
		_w903_
	);
	LUT4 #(
		.INIT('h8222)
	) name686 (
		_w601_,
		_w620_,
		_w797_,
		_w804_,
		_w904_
	);
	LUT4 #(
		.INIT('h2022)
	) name687 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w905_
	);
	LUT4 #(
		.INIT('h1f00)
	) name688 (
		_w256_,
		_w258_,
		_w261_,
		_w905_,
		_w906_
	);
	LUT3 #(
		.INIT('hc8)
	) name689 (
		_w524_,
		_w621_,
		_w906_,
		_w907_
	);
	LUT3 #(
		.INIT('h40)
	) name690 (
		_w521_,
		_w522_,
		_w620_,
		_w908_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		_w907_,
		_w908_,
		_w909_
	);
	LUT3 #(
		.INIT('h70)
	) name692 (
		_w262_,
		_w904_,
		_w909_,
		_w910_
	);
	LUT3 #(
		.INIT('hd0)
	) name693 (
		_w404_,
		_w903_,
		_w910_,
		_w911_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name694 (
		_w254_,
		_w863_,
		_w895_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h8)
	) name695 (
		_w252_,
		_w621_,
		_w913_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		\reg3_reg[27]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w914_
	);
	LUT3 #(
		.INIT('h07)
	) name697 (
		_w606_,
		_w621_,
		_w914_,
		_w915_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name698 (
		\state_reg[0]/NET0131 ,
		_w912_,
		_w913_,
		_w915_,
		_w916_
	);
	LUT3 #(
		.INIT('h01)
	) name699 (
		_w256_,
		_w258_,
		_w261_,
		_w917_
	);
	LUT4 #(
		.INIT('h0c88)
	) name700 (
		\reg0_reg[27]/NET0131 ,
		_w587_,
		_w862_,
		_w917_,
		_w918_
	);
	LUT4 #(
		.INIT('h0c88)
	) name701 (
		\reg0_reg[27]/NET0131 ,
		_w518_,
		_w894_,
		_w917_,
		_w919_
	);
	LUT3 #(
		.INIT('h02)
	) name702 (
		_w404_,
		_w901_,
		_w902_,
		_w920_
	);
	LUT2 #(
		.INIT('h8)
	) name703 (
		_w525_,
		_w620_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w904_,
		_w921_,
		_w922_
	);
	LUT4 #(
		.INIT('hfe00)
	) name705 (
		_w256_,
		_w258_,
		_w261_,
		_w525_,
		_w923_
	);
	LUT4 #(
		.INIT('hb9bf)
	) name706 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w924_
	);
	LUT4 #(
		.INIT('h0006)
	) name707 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w925_
	);
	LUT4 #(
		.INIT('hfe00)
	) name708 (
		_w256_,
		_w258_,
		_w261_,
		_w925_,
		_w926_
	);
	LUT4 #(
		.INIT('haa8a)
	) name709 (
		\reg0_reg[27]/NET0131 ,
		_w923_,
		_w924_,
		_w926_,
		_w927_
	);
	LUT4 #(
		.INIT('h0075)
	) name710 (
		_w917_,
		_w920_,
		_w922_,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name711 (
		_w254_,
		_w918_,
		_w919_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		\reg0_reg[27]/NET0131 ,
		_w252_,
		_w930_
	);
	LUT3 #(
		.INIT('h84)
	) name713 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w931_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name714 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[27]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w932_
	);
	LUT4 #(
		.INIT('hffa8)
	) name715 (
		\state_reg[0]/NET0131 ,
		_w929_,
		_w930_,
		_w932_,
		_w933_
	);
	LUT4 #(
		.INIT('hc355)
	) name716 (
		\reg0_reg[28]/NET0131 ,
		_w732_,
		_w741_,
		_w917_,
		_w934_
	);
	LUT4 #(
		.INIT('h0c88)
	) name717 (
		\reg0_reg[28]/NET0131 ,
		_w587_,
		_w795_,
		_w917_,
		_w935_
	);
	LUT2 #(
		.INIT('h8)
	) name718 (
		_w601_,
		_w807_,
		_w936_
	);
	LUT2 #(
		.INIT('h8)
	) name719 (
		_w525_,
		_w733_,
		_w937_
	);
	LUT4 #(
		.INIT('h0057)
	) name720 (
		_w404_,
		_w822_,
		_w823_,
		_w937_,
		_w938_
	);
	LUT4 #(
		.INIT('haa8a)
	) name721 (
		\reg0_reg[28]/NET0131 ,
		_w923_,
		_w924_,
		_w926_,
		_w939_
	);
	LUT4 #(
		.INIT('h0075)
	) name722 (
		_w917_,
		_w936_,
		_w938_,
		_w939_,
		_w940_
	);
	LUT4 #(
		.INIT('h0d00)
	) name723 (
		_w518_,
		_w934_,
		_w935_,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h8)
	) name724 (
		\reg0_reg[28]/NET0131 ,
		_w252_,
		_w942_
	);
	LUT4 #(
		.INIT('haa08)
	) name725 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w941_,
		_w942_,
		_w943_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name726 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[28]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w944_
	);
	LUT2 #(
		.INIT('he)
	) name727 (
		_w943_,
		_w944_,
		_w945_
	);
	LUT3 #(
		.INIT('h0e)
	) name728 (
		_w256_,
		_w258_,
		_w261_,
		_w946_
	);
	LUT4 #(
		.INIT('h0c88)
	) name729 (
		\reg1_reg[27]/NET0131 ,
		_w587_,
		_w862_,
		_w946_,
		_w947_
	);
	LUT4 #(
		.INIT('h0c88)
	) name730 (
		\reg1_reg[27]/NET0131 ,
		_w518_,
		_w894_,
		_w946_,
		_w948_
	);
	LUT4 #(
		.INIT('hf100)
	) name731 (
		_w256_,
		_w258_,
		_w261_,
		_w905_,
		_w949_
	);
	LUT4 #(
		.INIT('hf100)
	) name732 (
		_w256_,
		_w258_,
		_w261_,
		_w404_,
		_w950_
	);
	LUT4 #(
		.INIT('haaa2)
	) name733 (
		\reg1_reg[27]/NET0131 ,
		_w924_,
		_w949_,
		_w950_,
		_w951_
	);
	LUT4 #(
		.INIT('h004f)
	) name734 (
		_w920_,
		_w922_,
		_w946_,
		_w951_,
		_w952_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name735 (
		_w254_,
		_w947_,
		_w948_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h8)
	) name736 (
		\reg1_reg[27]/NET0131 ,
		_w252_,
		_w954_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name737 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[27]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w955_
	);
	LUT4 #(
		.INIT('hffa8)
	) name738 (
		\state_reg[0]/NET0131 ,
		_w953_,
		_w954_,
		_w955_,
		_w956_
	);
	LUT4 #(
		.INIT('hc355)
	) name739 (
		\reg1_reg[28]/NET0131 ,
		_w732_,
		_w741_,
		_w946_,
		_w957_
	);
	LUT4 #(
		.INIT('h0c88)
	) name740 (
		\reg1_reg[28]/NET0131 ,
		_w587_,
		_w795_,
		_w946_,
		_w958_
	);
	LUT4 #(
		.INIT('hf100)
	) name741 (
		_w256_,
		_w258_,
		_w261_,
		_w525_,
		_w959_
	);
	LUT4 #(
		.INIT('hf100)
	) name742 (
		_w256_,
		_w258_,
		_w261_,
		_w601_,
		_w960_
	);
	LUT3 #(
		.INIT('h02)
	) name743 (
		_w924_,
		_w959_,
		_w960_,
		_w961_
	);
	LUT4 #(
		.INIT('h0002)
	) name744 (
		_w924_,
		_w950_,
		_w959_,
		_w960_,
		_w962_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		\reg1_reg[28]/NET0131 ,
		_w962_,
		_w963_
	);
	LUT4 #(
		.INIT('h004f)
	) name746 (
		_w936_,
		_w938_,
		_w946_,
		_w963_,
		_w964_
	);
	LUT4 #(
		.INIT('h0d00)
	) name747 (
		_w518_,
		_w957_,
		_w958_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h8)
	) name748 (
		\reg1_reg[28]/NET0131 ,
		_w252_,
		_w966_
	);
	LUT4 #(
		.INIT('haa08)
	) name749 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w965_,
		_w966_,
		_w967_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name750 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[28]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w968_
	);
	LUT2 #(
		.INIT('he)
	) name751 (
		_w967_,
		_w968_,
		_w969_
	);
	LUT3 #(
		.INIT('h10)
	) name752 (
		_w256_,
		_w258_,
		_w261_,
		_w970_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name753 (
		\reg2_reg[27]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w971_
	);
	LUT4 #(
		.INIT('h0c88)
	) name754 (
		\reg2_reg[27]/NET0131 ,
		_w587_,
		_w862_,
		_w970_,
		_w972_
	);
	LUT4 #(
		.INIT('h0c88)
	) name755 (
		\reg2_reg[27]/NET0131 ,
		_w518_,
		_w894_,
		_w970_,
		_w973_
	);
	LUT4 #(
		.INIT('hfc55)
	) name756 (
		\reg2_reg[27]/NET0131 ,
		_w901_,
		_w902_,
		_w970_,
		_w974_
	);
	LUT4 #(
		.INIT('h9500)
	) name757 (
		_w620_,
		_w797_,
		_w804_,
		_w970_,
		_w975_
	);
	LUT4 #(
		.INIT('hef00)
	) name758 (
		_w256_,
		_w258_,
		_w261_,
		_w525_,
		_w976_
	);
	LUT3 #(
		.INIT('ha8)
	) name759 (
		\reg2_reg[27]/NET0131 ,
		_w524_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		_w520_,
		_w621_,
		_w978_
	);
	LUT3 #(
		.INIT('h07)
	) name761 (
		_w921_,
		_w970_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h4)
	) name762 (
		_w977_,
		_w979_,
		_w980_
	);
	LUT4 #(
		.INIT('h5700)
	) name763 (
		_w601_,
		_w971_,
		_w975_,
		_w980_,
		_w981_
	);
	LUT3 #(
		.INIT('hd0)
	) name764 (
		_w404_,
		_w974_,
		_w981_,
		_w982_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name765 (
		_w254_,
		_w972_,
		_w973_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		\reg2_reg[27]/NET0131 ,
		_w252_,
		_w984_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name767 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[27]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w985_
	);
	LUT4 #(
		.INIT('hffa8)
	) name768 (
		\state_reg[0]/NET0131 ,
		_w983_,
		_w984_,
		_w985_,
		_w986_
	);
	LUT4 #(
		.INIT('hc355)
	) name769 (
		\reg2_reg[28]/NET0131 ,
		_w732_,
		_w741_,
		_w970_,
		_w987_
	);
	LUT4 #(
		.INIT('h0c88)
	) name770 (
		\reg2_reg[28]/NET0131 ,
		_w587_,
		_w795_,
		_w970_,
		_w988_
	);
	LUT3 #(
		.INIT('h48)
	) name771 (
		\reg3_reg[28]/NET0131 ,
		_w520_,
		_w617_,
		_w989_
	);
	LUT4 #(
		.INIT('hef00)
	) name772 (
		_w256_,
		_w258_,
		_w261_,
		_w404_,
		_w990_
	);
	LUT4 #(
		.INIT('hef00)
	) name773 (
		_w256_,
		_w258_,
		_w261_,
		_w601_,
		_w991_
	);
	LUT4 #(
		.INIT('h0001)
	) name774 (
		_w524_,
		_w976_,
		_w990_,
		_w991_,
		_w992_
	);
	LUT3 #(
		.INIT('h31)
	) name775 (
		\reg2_reg[28]/NET0131 ,
		_w989_,
		_w992_,
		_w993_
	);
	LUT4 #(
		.INIT('h4f00)
	) name776 (
		_w936_,
		_w938_,
		_w970_,
		_w993_,
		_w994_
	);
	LUT4 #(
		.INIT('h0d00)
	) name777 (
		_w518_,
		_w987_,
		_w988_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h8)
	) name778 (
		\reg2_reg[28]/NET0131 ,
		_w252_,
		_w996_
	);
	LUT4 #(
		.INIT('haa08)
	) name779 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w995_,
		_w996_,
		_w997_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name780 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[28]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w998_
	);
	LUT2 #(
		.INIT('he)
	) name781 (
		_w997_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h8)
	) name782 (
		_w252_,
		_w374_,
		_w1000_
	);
	LUT4 #(
		.INIT('h1f00)
	) name783 (
		_w256_,
		_w258_,
		_w261_,
		_w374_,
		_w1001_
	);
	LUT4 #(
		.INIT('h0008)
	) name784 (
		_w339_,
		_w356_,
		_w372_,
		_w367_,
		_w1002_
	);
	LUT4 #(
		.INIT('h0703)
	) name785 (
		_w378_,
		_w361_,
		_w380_,
		_w1002_,
		_w1003_
	);
	LUT4 #(
		.INIT('h2a08)
	) name786 (
		_w262_,
		_w266_,
		_w367_,
		_w1003_,
		_w1004_
	);
	LUT3 #(
		.INIT('ha8)
	) name787 (
		_w404_,
		_w1001_,
		_w1004_,
		_w1005_
	);
	LUT4 #(
		.INIT('h10ef)
	) name788 (
		_w376_,
		_w375_,
		_w377_,
		_w449_,
		_w1006_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name789 (
		_w840_,
		_w841_,
		_w842_,
		_w1006_,
		_w1007_
	);
	LUT4 #(
		.INIT('h40e0)
	) name790 (
		_w262_,
		_w374_,
		_w587_,
		_w1007_,
		_w1008_
	);
	LUT4 #(
		.INIT('h4f00)
	) name791 (
		_w865_,
		_w866_,
		_w869_,
		_w871_,
		_w1009_
	);
	LUT4 #(
		.INIT('h3113)
	) name792 (
		_w262_,
		_w1001_,
		_w1006_,
		_w1009_,
		_w1010_
	);
	LUT4 #(
		.INIT('h820a)
	) name793 (
		_w262_,
		_w439_,
		_w449_,
		_w596_,
		_w1011_
	);
	LUT3 #(
		.INIT('h40)
	) name794 (
		_w521_,
		_w522_,
		_w449_,
		_w1012_
	);
	LUT3 #(
		.INIT('ha8)
	) name795 (
		_w374_,
		_w524_,
		_w526_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name796 (
		_w1012_,
		_w1013_,
		_w1014_
	);
	LUT4 #(
		.INIT('h5700)
	) name797 (
		_w601_,
		_w1001_,
		_w1011_,
		_w1014_,
		_w1015_
	);
	LUT4 #(
		.INIT('h0d00)
	) name798 (
		_w518_,
		_w1010_,
		_w1008_,
		_w1015_,
		_w1016_
	);
	LUT4 #(
		.INIT('h1311)
	) name799 (
		_w254_,
		_w1000_,
		_w1005_,
		_w1016_,
		_w1017_
	);
	LUT4 #(
		.INIT('h4800)
	) name800 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w374_,
		_w1018_
	);
	LUT2 #(
		.INIT('h2)
	) name801 (
		\reg3_reg[15]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1019_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		_w1018_,
		_w1019_,
		_w1020_
	);
	LUT3 #(
		.INIT('h2f)
	) name803 (
		\state_reg[0]/NET0131 ,
		_w1017_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h8)
	) name804 (
		_w252_,
		_w346_,
		_w1022_
	);
	LUT4 #(
		.INIT('h1f00)
	) name805 (
		_w256_,
		_w258_,
		_w261_,
		_w346_,
		_w1023_
	);
	LUT3 #(
		.INIT('h78)
	) name806 (
		_w345_,
		_w347_,
		_w418_,
		_w1024_
	);
	LUT4 #(
		.INIT('h8a20)
	) name807 (
		_w262_,
		_w865_,
		_w866_,
		_w1024_,
		_w1025_
	);
	LUT4 #(
		.INIT('h8000)
	) name808 (
		_w427_,
		_w467_,
		_w592_,
		_w593_,
		_w1026_
	);
	LUT4 #(
		.INIT('h8000)
	) name809 (
		_w467_,
		_w592_,
		_w593_,
		_w594_,
		_w1027_
	);
	LUT4 #(
		.INIT('h00a8)
	) name810 (
		_w262_,
		_w418_,
		_w1026_,
		_w1027_,
		_w1028_
	);
	LUT3 #(
		.INIT('h04)
	) name811 (
		_w521_,
		_w522_,
		_w418_,
		_w1029_
	);
	LUT3 #(
		.INIT('ha8)
	) name812 (
		_w346_,
		_w524_,
		_w526_,
		_w1030_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		_w1029_,
		_w1030_,
		_w1031_
	);
	LUT4 #(
		.INIT('h5700)
	) name814 (
		_w601_,
		_w1023_,
		_w1028_,
		_w1031_,
		_w1032_
	);
	LUT4 #(
		.INIT('h5700)
	) name815 (
		_w518_,
		_w1023_,
		_w1025_,
		_w1032_,
		_w1033_
	);
	LUT4 #(
		.INIT('h1450)
	) name816 (
		_w266_,
		_w339_,
		_w343_,
		_w355_,
		_w1034_
	);
	LUT3 #(
		.INIT('h80)
	) name817 (
		_w266_,
		_w350_,
		_w352_,
		_w1035_
	);
	LUT4 #(
		.INIT('h3331)
	) name818 (
		_w262_,
		_w1023_,
		_w1034_,
		_w1035_,
		_w1036_
	);
	LUT4 #(
		.INIT('h070d)
	) name819 (
		_w262_,
		_w840_,
		_w1023_,
		_w1024_,
		_w1037_
	);
	LUT4 #(
		.INIT('hf531)
	) name820 (
		_w404_,
		_w587_,
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT4 #(
		.INIT('h3111)
	) name821 (
		_w254_,
		_w1022_,
		_w1033_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h2)
	) name822 (
		\reg3_reg[11]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1040_
	);
	LUT4 #(
		.INIT('h4800)
	) name823 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w346_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w1040_,
		_w1041_,
		_w1042_
	);
	LUT3 #(
		.INIT('h2f)
	) name825 (
		\state_reg[0]/NET0131 ,
		_w1039_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h8)
	) name826 (
		_w252_,
		_w340_,
		_w1044_
	);
	LUT4 #(
		.INIT('h1f00)
	) name827 (
		_w256_,
		_w258_,
		_w261_,
		_w340_,
		_w1045_
	);
	LUT3 #(
		.INIT('h78)
	) name828 (
		_w341_,
		_w342_,
		_w423_,
		_w1046_
	);
	LUT4 #(
		.INIT('ha208)
	) name829 (
		_w262_,
		_w695_,
		_w706_,
		_w1046_,
		_w1047_
	);
	LUT4 #(
		.INIT('h00d7)
	) name830 (
		_w262_,
		_w423_,
		_w1027_,
		_w1045_,
		_w1048_
	);
	LUT3 #(
		.INIT('h04)
	) name831 (
		_w521_,
		_w522_,
		_w423_,
		_w1049_
	);
	LUT3 #(
		.INIT('ha8)
	) name832 (
		_w340_,
		_w524_,
		_w526_,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		_w1049_,
		_w1050_,
		_w1051_
	);
	LUT3 #(
		.INIT('hd0)
	) name834 (
		_w601_,
		_w1048_,
		_w1051_,
		_w1052_
	);
	LUT4 #(
		.INIT('h5700)
	) name835 (
		_w518_,
		_w1045_,
		_w1047_,
		_w1052_,
		_w1053_
	);
	LUT4 #(
		.INIT('h08a2)
	) name836 (
		_w262_,
		_w755_,
		_w766_,
		_w1046_,
		_w1054_
	);
	LUT3 #(
		.INIT('ha8)
	) name837 (
		_w587_,
		_w1045_,
		_w1054_,
		_w1055_
	);
	LUT4 #(
		.INIT('h1540)
	) name838 (
		_w266_,
		_w339_,
		_w356_,
		_w372_,
		_w1056_
	);
	LUT3 #(
		.INIT('h80)
	) name839 (
		_w266_,
		_w345_,
		_w347_,
		_w1057_
	);
	LUT4 #(
		.INIT('h3331)
	) name840 (
		_w262_,
		_w1045_,
		_w1056_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h2)
	) name841 (
		_w404_,
		_w1058_,
		_w1059_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name842 (
		_w254_,
		_w1055_,
		_w1059_,
		_w1053_,
		_w1060_
	);
	LUT4 #(
		.INIT('h4800)
	) name843 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w340_,
		_w1061_
	);
	LUT2 #(
		.INIT('h2)
	) name844 (
		\reg3_reg[12]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w1061_,
		_w1062_,
		_w1063_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name846 (
		\state_reg[0]/NET0131 ,
		_w1044_,
		_w1060_,
		_w1063_,
		_w1064_
	);
	LUT4 #(
		.INIT('h1f00)
	) name847 (
		_w256_,
		_w258_,
		_w261_,
		_w680_,
		_w1065_
	);
	LUT4 #(
		.INIT('hef10)
	) name848 (
		_w682_,
		_w681_,
		_w683_,
		_w686_,
		_w1066_
	);
	LUT4 #(
		.INIT('h070d)
	) name849 (
		_w262_,
		_w846_,
		_w1065_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		_w587_,
		_w1067_,
		_w1068_
	);
	LUT4 #(
		.INIT('h0d07)
	) name851 (
		_w262_,
		_w876_,
		_w1065_,
		_w1066_,
		_w1069_
	);
	LUT4 #(
		.INIT('h0800)
	) name852 (
		_w339_,
		_w356_,
		_w671_,
		_w897_,
		_w1070_
	);
	LUT4 #(
		.INIT('h870f)
	) name853 (
		_w339_,
		_w356_,
		_w671_,
		_w897_,
		_w1071_
	);
	LUT4 #(
		.INIT('h0200)
	) name854 (
		_w266_,
		_w389_,
		_w388_,
		_w390_,
		_w1072_
	);
	LUT2 #(
		.INIT('h2)
	) name855 (
		_w404_,
		_w1072_,
		_w1073_
	);
	LUT3 #(
		.INIT('he0)
	) name856 (
		_w266_,
		_w1071_,
		_w1073_,
		_w1074_
	);
	LUT4 #(
		.INIT('h00f7)
	) name857 (
		_w596_,
		_w598_,
		_w678_,
		_w686_,
		_w1075_
	);
	LUT4 #(
		.INIT('h70f0)
	) name858 (
		_w596_,
		_w598_,
		_w601_,
		_w798_,
		_w1076_
	);
	LUT2 #(
		.INIT('h4)
	) name859 (
		_w1075_,
		_w1076_,
		_w1077_
	);
	LUT4 #(
		.INIT('h1f00)
	) name860 (
		_w256_,
		_w258_,
		_w261_,
		_w925_,
		_w1078_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name861 (
		_w524_,
		_w526_,
		_w680_,
		_w1078_,
		_w1079_
	);
	LUT3 #(
		.INIT('h04)
	) name862 (
		_w521_,
		_w522_,
		_w686_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name863 (
		_w1079_,
		_w1080_,
		_w1081_
	);
	LUT4 #(
		.INIT('h5700)
	) name864 (
		_w262_,
		_w1074_,
		_w1077_,
		_w1081_,
		_w1082_
	);
	LUT3 #(
		.INIT('hd0)
	) name865 (
		_w518_,
		_w1069_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		_w252_,
		_w680_,
		_w1084_
	);
	LUT4 #(
		.INIT('h0075)
	) name867 (
		_w254_,
		_w1068_,
		_w1083_,
		_w1084_,
		_w1085_
	);
	LUT4 #(
		.INIT('h4800)
	) name868 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w680_,
		_w1086_
	);
	LUT2 #(
		.INIT('h2)
	) name869 (
		\reg3_reg[19]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		_w1086_,
		_w1087_,
		_w1088_
	);
	LUT3 #(
		.INIT('h2f)
	) name871 (
		\state_reg[0]/NET0131 ,
		_w1085_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h8)
	) name872 (
		_w252_,
		_w644_,
		_w1090_
	);
	LUT4 #(
		.INIT('h1f00)
	) name873 (
		_w256_,
		_w258_,
		_w261_,
		_w644_,
		_w1091_
	);
	LUT2 #(
		.INIT('h9)
	) name874 (
		_w643_,
		_w647_,
		_w1092_
	);
	LUT4 #(
		.INIT('h80aa)
	) name875 (
		_w745_,
		_w752_,
		_w753_,
		_w754_,
		_w1093_
	);
	LUT4 #(
		.INIT('h50d0)
	) name876 (
		_w750_,
		_w769_,
		_w774_,
		_w1093_,
		_w1094_
	);
	LUT4 #(
		.INIT('h80f0)
	) name877 (
		_w751_,
		_w766_,
		_w779_,
		_w1094_,
		_w1095_
	);
	LUT4 #(
		.INIT('h0a82)
	) name878 (
		_w262_,
		_w788_,
		_w1092_,
		_w1095_,
		_w1096_
	);
	LUT3 #(
		.INIT('ha8)
	) name879 (
		_w587_,
		_w1091_,
		_w1096_,
		_w1097_
	);
	LUT3 #(
		.INIT('h80)
	) name880 (
		_w659_,
		_w673_,
		_w709_,
		_w1098_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		_w691_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		_w706_,
		_w1099_,
		_w1100_
	);
	LUT4 #(
		.INIT('h8f00)
	) name883 (
		_w692_,
		_w693_,
		_w694_,
		_w709_,
		_w1101_
	);
	LUT4 #(
		.INIT('h50d0)
	) name884 (
		_w691_,
		_w713_,
		_w719_,
		_w1101_,
		_w1102_
	);
	LUT3 #(
		.INIT('hc4)
	) name885 (
		_w674_,
		_w724_,
		_w1102_,
		_w1103_
	);
	LUT4 #(
		.INIT('h8288)
	) name886 (
		_w262_,
		_w1092_,
		_w1100_,
		_w1103_,
		_w1104_
	);
	LUT3 #(
		.INIT('ha8)
	) name887 (
		_w518_,
		_w1091_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h2)
	) name888 (
		_w266_,
		_w615_,
		_w1106_
	);
	LUT4 #(
		.INIT('h4105)
	) name889 (
		_w266_,
		_w394_,
		_w640_,
		_w812_,
		_w1107_
	);
	LUT4 #(
		.INIT('h1113)
	) name890 (
		_w262_,
		_w1091_,
		_w1106_,
		_w1107_,
		_w1108_
	);
	LUT4 #(
		.INIT('h8222)
	) name891 (
		_w262_,
		_w643_,
		_w799_,
		_w802_,
		_w1109_
	);
	LUT3 #(
		.INIT('h40)
	) name892 (
		_w521_,
		_w522_,
		_w643_,
		_w1110_
	);
	LUT3 #(
		.INIT('he0)
	) name893 (
		_w524_,
		_w526_,
		_w644_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name894 (
		_w1110_,
		_w1111_,
		_w1112_
	);
	LUT4 #(
		.INIT('h5700)
	) name895 (
		_w601_,
		_w1091_,
		_w1109_,
		_w1112_,
		_w1113_
	);
	LUT3 #(
		.INIT('hd0)
	) name896 (
		_w404_,
		_w1108_,
		_w1113_,
		_w1114_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name897 (
		_w254_,
		_w1097_,
		_w1105_,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h2)
	) name898 (
		\reg3_reg[24]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1116_
	);
	LUT3 #(
		.INIT('h07)
	) name899 (
		_w606_,
		_w644_,
		_w1116_,
		_w1117_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name900 (
		\state_reg[0]/NET0131 ,
		_w1090_,
		_w1115_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h8)
	) name901 (
		_w252_,
		_w612_,
		_w1119_
	);
	LUT4 #(
		.INIT('h1f00)
	) name902 (
		_w256_,
		_w258_,
		_w261_,
		_w612_,
		_w1120_
	);
	LUT2 #(
		.INIT('h9)
	) name903 (
		_w615_,
		_w651_,
		_w1121_
	);
	LUT4 #(
		.INIT('h8000)
	) name904 (
		_w530_,
		_w835_,
		_w847_,
		_w848_,
		_w1122_
	);
	LUT4 #(
		.INIT('h4f00)
	) name905 (
		_w840_,
		_w841_,
		_w842_,
		_w1122_,
		_w1123_
	);
	LUT3 #(
		.INIT('hb0)
	) name906 (
		_w844_,
		_w849_,
		_w856_,
		_w1124_
	);
	LUT4 #(
		.INIT('h2822)
	) name907 (
		_w262_,
		_w1121_,
		_w1123_,
		_w1124_,
		_w1125_
	);
	LUT3 #(
		.INIT('ha8)
	) name908 (
		_w587_,
		_w1120_,
		_w1125_,
		_w1126_
	);
	LUT4 #(
		.INIT('h8000)
	) name909 (
		_w451_,
		_w867_,
		_w877_,
		_w878_,
		_w1127_
	);
	LUT3 #(
		.INIT('hb0)
	) name910 (
		_w874_,
		_w879_,
		_w888_,
		_w1128_
	);
	LUT4 #(
		.INIT('h9c33)
	) name911 (
		_w1009_,
		_w1121_,
		_w1127_,
		_w1128_,
		_w1129_
	);
	LUT4 #(
		.INIT('h40c8)
	) name912 (
		_w262_,
		_w518_,
		_w612_,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name913 (
		_w266_,
		_w657_,
		_w1131_
	);
	LUT4 #(
		.INIT('h00eb)
	) name914 (
		_w266_,
		_w647_,
		_w899_,
		_w1131_,
		_w1132_
	);
	LUT4 #(
		.INIT('hc840)
	) name915 (
		_w262_,
		_w404_,
		_w612_,
		_w1132_,
		_w1133_
	);
	LUT4 #(
		.INIT('h8000)
	) name916 (
		_w596_,
		_w598_,
		_w798_,
		_w801_,
		_w1134_
	);
	LUT4 #(
		.INIT('h8222)
	) name917 (
		_w262_,
		_w651_,
		_w799_,
		_w801_,
		_w1135_
	);
	LUT3 #(
		.INIT('h40)
	) name918 (
		_w521_,
		_w522_,
		_w651_,
		_w1136_
	);
	LUT3 #(
		.INIT('he0)
	) name919 (
		_w524_,
		_w526_,
		_w612_,
		_w1137_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w1136_,
		_w1137_,
		_w1138_
	);
	LUT4 #(
		.INIT('h5700)
	) name921 (
		_w601_,
		_w1120_,
		_w1135_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h4)
	) name922 (
		_w1133_,
		_w1139_,
		_w1140_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name923 (
		_w254_,
		_w1130_,
		_w1126_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h2)
	) name924 (
		\reg3_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1142_
	);
	LUT3 #(
		.INIT('h07)
	) name925 (
		_w606_,
		_w612_,
		_w1142_,
		_w1143_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name926 (
		\state_reg[0]/NET0131 ,
		_w1119_,
		_w1141_,
		_w1143_,
		_w1144_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name927 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[15]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1145_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		\reg0_reg[15]/NET0131 ,
		_w252_,
		_w1146_
	);
	LUT4 #(
		.INIT('haaa8)
	) name929 (
		\reg0_reg[15]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1147_
	);
	LUT4 #(
		.INIT('h7020)
	) name930 (
		_w266_,
		_w367_,
		_w917_,
		_w1003_,
		_w1148_
	);
	LUT3 #(
		.INIT('ha8)
	) name931 (
		_w404_,
		_w1147_,
		_w1148_,
		_w1149_
	);
	LUT4 #(
		.INIT('h08c8)
	) name932 (
		\reg0_reg[15]/NET0131 ,
		_w587_,
		_w917_,
		_w1007_,
		_w1150_
	);
	LUT4 #(
		.INIT('hd11d)
	) name933 (
		\reg0_reg[15]/NET0131 ,
		_w917_,
		_w1006_,
		_w1009_,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name934 (
		_w449_,
		_w525_,
		_w1152_
	);
	LUT4 #(
		.INIT('h9300)
	) name935 (
		_w439_,
		_w449_,
		_w596_,
		_w601_,
		_w1153_
	);
	LUT4 #(
		.INIT('hfe00)
	) name936 (
		_w256_,
		_w258_,
		_w261_,
		_w601_,
		_w1154_
	);
	LUT3 #(
		.INIT('h04)
	) name937 (
		_w923_,
		_w924_,
		_w1154_,
		_w1155_
	);
	LUT4 #(
		.INIT('haa8a)
	) name938 (
		\reg0_reg[15]/NET0131 ,
		_w923_,
		_w924_,
		_w1154_,
		_w1156_
	);
	LUT4 #(
		.INIT('h0057)
	) name939 (
		_w917_,
		_w1152_,
		_w1153_,
		_w1156_,
		_w1157_
	);
	LUT4 #(
		.INIT('h0d00)
	) name940 (
		_w518_,
		_w1151_,
		_w1150_,
		_w1157_,
		_w1158_
	);
	LUT4 #(
		.INIT('h1311)
	) name941 (
		_w254_,
		_w1146_,
		_w1149_,
		_w1158_,
		_w1159_
	);
	LUT3 #(
		.INIT('hce)
	) name942 (
		\state_reg[0]/NET0131 ,
		_w1145_,
		_w1159_,
		_w1160_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name943 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1161_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		\reg0_reg[23]/NET0131 ,
		_w252_,
		_w1162_
	);
	LUT4 #(
		.INIT('haaa8)
	) name945 (
		\reg0_reg[23]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1163_
	);
	LUT4 #(
		.INIT('h2822)
	) name946 (
		_w917_,
		_w1121_,
		_w1123_,
		_w1124_,
		_w1164_
	);
	LUT3 #(
		.INIT('ha8)
	) name947 (
		_w587_,
		_w1163_,
		_w1164_,
		_w1165_
	);
	LUT4 #(
		.INIT('h08c8)
	) name948 (
		\reg0_reg[23]/NET0131 ,
		_w518_,
		_w917_,
		_w1129_,
		_w1166_
	);
	LUT4 #(
		.INIT('hc808)
	) name949 (
		\reg0_reg[23]/NET0131 ,
		_w404_,
		_w917_,
		_w1132_,
		_w1167_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		_w525_,
		_w651_,
		_w1168_
	);
	LUT4 #(
		.INIT('h8222)
	) name951 (
		_w601_,
		_w651_,
		_w799_,
		_w801_,
		_w1169_
	);
	LUT4 #(
		.INIT('haa8a)
	) name952 (
		\reg0_reg[23]/NET0131 ,
		_w923_,
		_w924_,
		_w1154_,
		_w1170_
	);
	LUT4 #(
		.INIT('h0057)
	) name953 (
		_w917_,
		_w1168_,
		_w1169_,
		_w1170_,
		_w1171_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w1167_,
		_w1171_,
		_w1172_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name955 (
		_w254_,
		_w1166_,
		_w1165_,
		_w1172_,
		_w1173_
	);
	LUT4 #(
		.INIT('heeec)
	) name956 (
		\state_reg[0]/NET0131 ,
		_w1161_,
		_w1162_,
		_w1173_,
		_w1174_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name957 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[24]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1175_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		\reg0_reg[24]/NET0131 ,
		_w252_,
		_w1176_
	);
	LUT4 #(
		.INIT('h8288)
	) name959 (
		_w518_,
		_w1092_,
		_w1100_,
		_w1103_,
		_w1177_
	);
	LUT3 #(
		.INIT('ha8)
	) name960 (
		_w404_,
		_w1106_,
		_w1107_,
		_w1178_
	);
	LUT4 #(
		.INIT('h8222)
	) name961 (
		_w601_,
		_w643_,
		_w799_,
		_w802_,
		_w1179_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		_w525_,
		_w643_,
		_w1180_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w1179_,
		_w1180_,
		_w1181_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name964 (
		_w917_,
		_w1178_,
		_w1177_,
		_w1181_,
		_w1182_
	);
	LUT4 #(
		.INIT('h6e7b)
	) name965 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w1183_
	);
	LUT4 #(
		.INIT('h00fe)
	) name966 (
		_w256_,
		_w258_,
		_w261_,
		_w1183_,
		_w1184_
	);
	LUT4 #(
		.INIT('h0004)
	) name967 (
		_w923_,
		_w924_,
		_w1154_,
		_w1184_,
		_w1185_
	);
	LUT2 #(
		.INIT('h2)
	) name968 (
		\reg0_reg[24]/NET0131 ,
		_w1185_,
		_w1186_
	);
	LUT4 #(
		.INIT('hc048)
	) name969 (
		_w788_,
		_w917_,
		_w1092_,
		_w1095_,
		_w1187_
	);
	LUT4 #(
		.INIT('h5554)
	) name970 (
		\reg0_reg[24]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1188_
	);
	LUT2 #(
		.INIT('h2)
	) name971 (
		_w587_,
		_w1188_,
		_w1189_
	);
	LUT3 #(
		.INIT('h45)
	) name972 (
		_w1186_,
		_w1187_,
		_w1189_,
		_w1190_
	);
	LUT4 #(
		.INIT('h1311)
	) name973 (
		_w254_,
		_w1176_,
		_w1182_,
		_w1190_,
		_w1191_
	);
	LUT3 #(
		.INIT('hce)
	) name974 (
		\state_reg[0]/NET0131 ,
		_w1175_,
		_w1191_,
		_w1192_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name975 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[15]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name976 (
		\reg1_reg[15]/NET0131 ,
		_w252_,
		_w1194_
	);
	LUT4 #(
		.INIT('haa02)
	) name977 (
		\reg1_reg[15]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1195_
	);
	LUT4 #(
		.INIT('h7020)
	) name978 (
		_w266_,
		_w367_,
		_w946_,
		_w1003_,
		_w1196_
	);
	LUT3 #(
		.INIT('ha8)
	) name979 (
		_w404_,
		_w1195_,
		_w1196_,
		_w1197_
	);
	LUT4 #(
		.INIT('h08c8)
	) name980 (
		\reg1_reg[15]/NET0131 ,
		_w587_,
		_w946_,
		_w1007_,
		_w1198_
	);
	LUT4 #(
		.INIT('hd11d)
	) name981 (
		\reg1_reg[15]/NET0131 ,
		_w946_,
		_w1006_,
		_w1009_,
		_w1199_
	);
	LUT3 #(
		.INIT('ha2)
	) name982 (
		\reg1_reg[15]/NET0131 ,
		_w924_,
		_w949_,
		_w1200_
	);
	LUT4 #(
		.INIT('h0057)
	) name983 (
		_w946_,
		_w1152_,
		_w1153_,
		_w1200_,
		_w1201_
	);
	LUT4 #(
		.INIT('h0d00)
	) name984 (
		_w518_,
		_w1199_,
		_w1198_,
		_w1201_,
		_w1202_
	);
	LUT4 #(
		.INIT('h1311)
	) name985 (
		_w254_,
		_w1194_,
		_w1197_,
		_w1202_,
		_w1203_
	);
	LUT3 #(
		.INIT('hce)
	) name986 (
		\state_reg[0]/NET0131 ,
		_w1193_,
		_w1203_,
		_w1204_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name987 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1205_
	);
	LUT2 #(
		.INIT('h8)
	) name988 (
		\reg1_reg[23]/NET0131 ,
		_w252_,
		_w1206_
	);
	LUT4 #(
		.INIT('haa02)
	) name989 (
		\reg1_reg[23]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1207_
	);
	LUT4 #(
		.INIT('h2822)
	) name990 (
		_w946_,
		_w1121_,
		_w1123_,
		_w1124_,
		_w1208_
	);
	LUT3 #(
		.INIT('ha8)
	) name991 (
		_w587_,
		_w1207_,
		_w1208_,
		_w1209_
	);
	LUT4 #(
		.INIT('h08c8)
	) name992 (
		\reg1_reg[23]/NET0131 ,
		_w518_,
		_w946_,
		_w1129_,
		_w1210_
	);
	LUT4 #(
		.INIT('hc808)
	) name993 (
		\reg1_reg[23]/NET0131 ,
		_w404_,
		_w946_,
		_w1132_,
		_w1211_
	);
	LUT3 #(
		.INIT('ha2)
	) name994 (
		\reg1_reg[23]/NET0131 ,
		_w924_,
		_w949_,
		_w1212_
	);
	LUT4 #(
		.INIT('h0057)
	) name995 (
		_w946_,
		_w1168_,
		_w1169_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		_w1211_,
		_w1213_,
		_w1214_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name997 (
		_w254_,
		_w1210_,
		_w1209_,
		_w1214_,
		_w1215_
	);
	LUT4 #(
		.INIT('heeec)
	) name998 (
		\state_reg[0]/NET0131 ,
		_w1205_,
		_w1206_,
		_w1215_,
		_w1216_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name999 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[24]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1217_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		\reg1_reg[24]/NET0131 ,
		_w252_,
		_w1218_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1001 (
		_w946_,
		_w1178_,
		_w1177_,
		_w1181_,
		_w1219_
	);
	LUT4 #(
		.INIT('hf100)
	) name1002 (
		_w256_,
		_w258_,
		_w261_,
		_w518_,
		_w1220_
	);
	LUT4 #(
		.INIT('h0002)
	) name1003 (
		_w924_,
		_w949_,
		_w950_,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h2)
	) name1004 (
		\reg1_reg[24]/NET0131 ,
		_w1221_,
		_w1222_
	);
	LUT4 #(
		.INIT('hc048)
	) name1005 (
		_w788_,
		_w946_,
		_w1092_,
		_w1095_,
		_w1223_
	);
	LUT4 #(
		.INIT('h5501)
	) name1006 (
		\reg1_reg[24]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1224_
	);
	LUT2 #(
		.INIT('h2)
	) name1007 (
		_w587_,
		_w1224_,
		_w1225_
	);
	LUT3 #(
		.INIT('h45)
	) name1008 (
		_w1222_,
		_w1223_,
		_w1225_,
		_w1226_
	);
	LUT4 #(
		.INIT('h1311)
	) name1009 (
		_w254_,
		_w1218_,
		_w1219_,
		_w1226_,
		_w1227_
	);
	LUT3 #(
		.INIT('hce)
	) name1010 (
		\state_reg[0]/NET0131 ,
		_w1217_,
		_w1227_,
		_w1228_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1011 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[15]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name1012 (
		\reg2_reg[15]/NET0131 ,
		_w252_,
		_w1230_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1013 (
		\reg2_reg[15]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1231_
	);
	LUT4 #(
		.INIT('h7020)
	) name1014 (
		_w266_,
		_w367_,
		_w970_,
		_w1003_,
		_w1232_
	);
	LUT3 #(
		.INIT('ha8)
	) name1015 (
		_w404_,
		_w1231_,
		_w1232_,
		_w1233_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1016 (
		\reg2_reg[15]/NET0131 ,
		_w587_,
		_w970_,
		_w1007_,
		_w1234_
	);
	LUT4 #(
		.INIT('hd11d)
	) name1017 (
		\reg2_reg[15]/NET0131 ,
		_w970_,
		_w1006_,
		_w1009_,
		_w1235_
	);
	LUT2 #(
		.INIT('h8)
	) name1018 (
		_w520_,
		_w374_,
		_w1236_
	);
	LUT4 #(
		.INIT('hef00)
	) name1019 (
		_w256_,
		_w258_,
		_w261_,
		_w905_,
		_w1237_
	);
	LUT4 #(
		.INIT('h0507)
	) name1020 (
		\reg2_reg[15]/NET0131 ,
		_w524_,
		_w1236_,
		_w1237_,
		_w1238_
	);
	LUT4 #(
		.INIT('h5700)
	) name1021 (
		_w970_,
		_w1152_,
		_w1153_,
		_w1238_,
		_w1239_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1022 (
		_w518_,
		_w1235_,
		_w1234_,
		_w1239_,
		_w1240_
	);
	LUT4 #(
		.INIT('h1311)
	) name1023 (
		_w254_,
		_w1230_,
		_w1233_,
		_w1240_,
		_w1241_
	);
	LUT3 #(
		.INIT('hce)
	) name1024 (
		\state_reg[0]/NET0131 ,
		_w1229_,
		_w1241_,
		_w1242_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1025 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1243_
	);
	LUT2 #(
		.INIT('h8)
	) name1026 (
		\reg2_reg[23]/NET0131 ,
		_w252_,
		_w1244_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1027 (
		\reg2_reg[23]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1245_
	);
	LUT4 #(
		.INIT('h2822)
	) name1028 (
		_w970_,
		_w1121_,
		_w1123_,
		_w1124_,
		_w1246_
	);
	LUT3 #(
		.INIT('ha8)
	) name1029 (
		_w587_,
		_w1245_,
		_w1246_,
		_w1247_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1030 (
		\reg2_reg[23]/NET0131 ,
		_w518_,
		_w970_,
		_w1129_,
		_w1248_
	);
	LUT4 #(
		.INIT('hc808)
	) name1031 (
		\reg2_reg[23]/NET0131 ,
		_w404_,
		_w970_,
		_w1132_,
		_w1249_
	);
	LUT2 #(
		.INIT('h8)
	) name1032 (
		_w520_,
		_w612_,
		_w1250_
	);
	LUT4 #(
		.INIT('h0057)
	) name1033 (
		\reg2_reg[23]/NET0131 ,
		_w524_,
		_w1237_,
		_w1250_,
		_w1251_
	);
	LUT4 #(
		.INIT('h5700)
	) name1034 (
		_w970_,
		_w1168_,
		_w1169_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h4)
	) name1035 (
		_w1249_,
		_w1252_,
		_w1253_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1036 (
		_w254_,
		_w1248_,
		_w1247_,
		_w1253_,
		_w1254_
	);
	LUT4 #(
		.INIT('heeec)
	) name1037 (
		\state_reg[0]/NET0131 ,
		_w1243_,
		_w1244_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name1038 (
		\reg2_reg[29]/NET0131 ,
		_w252_,
		_w1256_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1039 (
		\reg2_reg[29]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1257_
	);
	LUT3 #(
		.INIT('h8a)
	) name1040 (
		_w266_,
		_w734_,
		_w737_,
		_w1258_
	);
	LUT4 #(
		.INIT('h1000)
	) name1041 (
		_w738_,
		_w820_,
		_w899_,
		_w900_,
		_w1259_
	);
	LUT3 #(
		.INIT('h02)
	) name1042 (
		\reg0_reg[30]/NET0131 ,
		_w269_,
		_w272_,
		_w1260_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1043 (
		\reg1_reg[30]/NET0131 ,
		\reg2_reg[30]/NET0131 ,
		_w269_,
		_w272_,
		_w1261_
	);
	LUT3 #(
		.INIT('h10)
	) name1044 (
		_w296_,
		_w1260_,
		_w1261_,
		_w1262_
	);
	LUT3 #(
		.INIT('hef)
	) name1045 (
		_w296_,
		_w1260_,
		_w1261_,
		_w1263_
	);
	LUT3 #(
		.INIT('hec)
	) name1046 (
		\B_reg/NET0131 ,
		_w266_,
		_w407_,
		_w1264_
	);
	LUT4 #(
		.INIT('h4554)
	) name1047 (
		_w1258_,
		_w1264_,
		_w1259_,
		_w1262_,
		_w1265_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1048 (
		\reg2_reg[29]/NET0131 ,
		_w404_,
		_w970_,
		_w1265_,
		_w1266_
	);
	LUT3 #(
		.INIT('ha8)
	) name1049 (
		\datai[29]_pad ,
		_w266_,
		_w407_,
		_w1267_
	);
	LUT4 #(
		.INIT('h1000)
	) name1050 (
		_w296_,
		_w818_,
		_w819_,
		_w1267_,
		_w1268_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1051 (
		_w296_,
		_w818_,
		_w819_,
		_w1267_,
		_w1269_
	);
	LUT4 #(
		.INIT('hef10)
	) name1052 (
		_w296_,
		_w818_,
		_w819_,
		_w1267_,
		_w1270_
	);
	LUT3 #(
		.INIT('h80)
	) name1053 (
		_w463_,
		_w509_,
		_w512_,
		_w1271_
	);
	LUT4 #(
		.INIT('haa80)
	) name1054 (
		_w463_,
		_w472_,
		_w482_,
		_w485_,
		_w1272_
	);
	LUT2 #(
		.INIT('h2)
	) name1055 (
		_w437_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h8)
	) name1056 (
		_w867_,
		_w877_,
		_w1274_
	);
	LUT4 #(
		.INIT('h8000)
	) name1057 (
		_w444_,
		_w451_,
		_w867_,
		_w877_,
		_w1275_
	);
	LUT3 #(
		.INIT('h07)
	) name1058 (
		_w873_,
		_w877_,
		_w885_,
		_w1276_
	);
	LUT3 #(
		.INIT('hb0)
	) name1059 (
		_w459_,
		_w1274_,
		_w1276_,
		_w1277_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1060 (
		_w1271_,
		_w1273_,
		_w1275_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		_w878_,
		_w880_,
		_w1279_
	);
	LUT3 #(
		.INIT('h20)
	) name1062 (
		_w733_,
		_w734_,
		_w737_,
		_w1280_
	);
	LUT3 #(
		.INIT('h04)
	) name1063 (
		_w626_,
		_w881_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		_w1279_,
		_w1281_,
		_w1282_
	);
	LUT3 #(
		.INIT('h70)
	) name1065 (
		_w880_,
		_w887_,
		_w891_,
		_w1283_
	);
	LUT3 #(
		.INIT('h04)
	) name1066 (
		_w626_,
		_w890_,
		_w1280_,
		_w1284_
	);
	LUT3 #(
		.INIT('hd4)
	) name1067 (
		_w725_,
		_w733_,
		_w738_,
		_w1285_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1068 (
		_w1281_,
		_w1283_,
		_w1284_,
		_w1285_,
		_w1286_
	);
	LUT4 #(
		.INIT('h9a55)
	) name1069 (
		_w1270_,
		_w1278_,
		_w1282_,
		_w1286_,
		_w1287_
	);
	LUT4 #(
		.INIT('hc808)
	) name1070 (
		\reg2_reg[29]/NET0131 ,
		_w518_,
		_w970_,
		_w1287_,
		_w1288_
	);
	LUT4 #(
		.INIT('h22a2)
	) name1071 (
		_w551_,
		_w555_,
		_w566_,
		_w584_,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name1072 (
		_w835_,
		_w848_,
		_w1290_
	);
	LUT4 #(
		.INIT('h8000)
	) name1073 (
		_w530_,
		_w539_,
		_w835_,
		_w848_,
		_w1291_
	);
	LUT3 #(
		.INIT('hb0)
	) name1074 (
		_w843_,
		_w848_,
		_w854_,
		_w1292_
	);
	LUT3 #(
		.INIT('hb0)
	) name1075 (
		_w537_,
		_w1290_,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h8)
	) name1076 (
		_w847_,
		_w850_,
		_w1294_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1077 (
		_w733_,
		_w734_,
		_w737_,
		_w782_,
		_w1295_
	);
	LUT2 #(
		.INIT('h8)
	) name1078 (
		_w781_,
		_w1295_,
		_w1296_
	);
	LUT4 #(
		.INIT('h8000)
	) name1079 (
		_w781_,
		_w847_,
		_w850_,
		_w1295_,
		_w1297_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1080 (
		_w1289_,
		_w1291_,
		_w1293_,
		_w1297_,
		_w1298_
	);
	LUT4 #(
		.INIT('h5054)
	) name1081 (
		_w739_,
		_w781_,
		_w789_,
		_w857_,
		_w1299_
	);
	LUT3 #(
		.INIT('hd0)
	) name1082 (
		_w850_,
		_w855_,
		_w858_,
		_w1300_
	);
	LUT4 #(
		.INIT('h0051)
	) name1083 (
		_w740_,
		_w1296_,
		_w1300_,
		_w1299_,
		_w1301_
	);
	LUT4 #(
		.INIT('h8288)
	) name1084 (
		_w970_,
		_w1270_,
		_w1298_,
		_w1301_,
		_w1302_
	);
	LUT4 #(
		.INIT('h8070)
	) name1085 (
		_w804_,
		_w806_,
		_w970_,
		_w1267_,
		_w1303_
	);
	LUT3 #(
		.INIT('ha8)
	) name1086 (
		\reg2_reg[29]/NET0131 ,
		_w524_,
		_w976_,
		_w1304_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		_w520_,
		_w295_,
		_w1305_
	);
	LUT2 #(
		.INIT('h8)
	) name1088 (
		_w525_,
		_w1267_,
		_w1306_
	);
	LUT3 #(
		.INIT('h13)
	) name1089 (
		_w970_,
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT2 #(
		.INIT('h4)
	) name1090 (
		_w1304_,
		_w1307_,
		_w1308_
	);
	LUT4 #(
		.INIT('h5700)
	) name1091 (
		_w601_,
		_w1257_,
		_w1303_,
		_w1308_,
		_w1309_
	);
	LUT4 #(
		.INIT('h5700)
	) name1092 (
		_w587_,
		_w1257_,
		_w1302_,
		_w1309_,
		_w1310_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1093 (
		_w254_,
		_w1266_,
		_w1288_,
		_w1310_,
		_w1311_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1094 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[29]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1312_
	);
	LUT4 #(
		.INIT('hffa8)
	) name1095 (
		\state_reg[0]/NET0131 ,
		_w1256_,
		_w1311_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h8)
	) name1096 (
		_w252_,
		_w363_,
		_w1314_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1097 (
		_w256_,
		_w258_,
		_w261_,
		_w363_,
		_w1315_
	);
	LUT3 #(
		.INIT('h80)
	) name1098 (
		_w266_,
		_w370_,
		_w371_,
		_w1316_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1099 (
		_w266_,
		_w378_,
		_w1002_,
		_w1316_,
		_w1317_
	);
	LUT4 #(
		.INIT('he040)
	) name1100 (
		_w262_,
		_w363_,
		_w404_,
		_w1317_,
		_w1318_
	);
	LUT4 #(
		.INIT('h10ef)
	) name1101 (
		_w365_,
		_w364_,
		_w366_,
		_w439_,
		_w1319_
	);
	LUT4 #(
		.INIT('h0001)
	) name1102 (
		_w553_,
		_w556_,
		_w557_,
		_w560_,
		_w1320_
	);
	LUT3 #(
		.INIT('h45)
	) name1103 (
		_w753_,
		_w762_,
		_w764_,
		_w1321_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1104 (
		_w760_,
		_w761_,
		_w1320_,
		_w1321_,
		_w1322_
	);
	LUT4 #(
		.INIT('h0001)
	) name1105 (
		_w538_,
		_w541_,
		_w542_,
		_w544_,
		_w1323_
	);
	LUT3 #(
		.INIT('hd0)
	) name1106 (
		_w743_,
		_w754_,
		_w767_,
		_w1324_
	);
	LUT4 #(
		.INIT('h65aa)
	) name1107 (
		_w1319_,
		_w1322_,
		_w1323_,
		_w1324_,
		_w1325_
	);
	LUT4 #(
		.INIT('he040)
	) name1108 (
		_w262_,
		_w363_,
		_w587_,
		_w1325_,
		_w1326_
	);
	LUT3 #(
		.INIT('h8a)
	) name1109 (
		_w711_,
		_w694_,
		_w708_,
		_w1327_
	);
	LUT4 #(
		.INIT('h0001)
	) name1110 (
		_w419_,
		_w424_,
		_w428_,
		_w443_,
		_w1328_
	);
	LUT3 #(
		.INIT('h45)
	) name1111 (
		_w693_,
		_w702_,
		_w704_,
		_w1329_
	);
	LUT4 #(
		.INIT('h0001)
	) name1112 (
		_w461_,
		_w468_,
		_w471_,
		_w476_,
		_w1330_
	);
	LUT4 #(
		.INIT('h10f0)
	) name1113 (
		_w700_,
		_w701_,
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT4 #(
		.INIT('h5da2)
	) name1114 (
		_w1327_,
		_w1328_,
		_w1331_,
		_w1319_,
		_w1332_
	);
	LUT4 #(
		.INIT('h40e0)
	) name1115 (
		_w262_,
		_w363_,
		_w518_,
		_w1332_,
		_w1333_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1116 (
		_w262_,
		_w439_,
		_w596_,
		_w1315_,
		_w1334_
	);
	LUT3 #(
		.INIT('h04)
	) name1117 (
		_w521_,
		_w522_,
		_w439_,
		_w1335_
	);
	LUT3 #(
		.INIT('ha8)
	) name1118 (
		_w363_,
		_w524_,
		_w526_,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name1119 (
		_w1335_,
		_w1336_,
		_w1337_
	);
	LUT3 #(
		.INIT('hd0)
	) name1120 (
		_w601_,
		_w1334_,
		_w1337_,
		_w1338_
	);
	LUT4 #(
		.INIT('h0100)
	) name1121 (
		_w1318_,
		_w1333_,
		_w1326_,
		_w1338_,
		_w1339_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1122 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1314_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h2)
	) name1123 (
		\reg3_reg[14]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1341_
	);
	LUT4 #(
		.INIT('h4800)
	) name1124 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w363_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name1125 (
		_w1341_,
		_w1342_,
		_w1343_
	);
	LUT2 #(
		.INIT('hb)
	) name1126 (
		_w1340_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h8)
	) name1127 (
		_w252_,
		_w358_,
		_w1345_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1128 (
		_w256_,
		_w258_,
		_w261_,
		_w358_,
		_w1346_
	);
	LUT2 #(
		.INIT('h9)
	) name1129 (
		_w361_,
		_w446_,
		_w1347_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1130 (
		_w745_,
		_w755_,
		_w766_,
		_w769_,
		_w1348_
	);
	LUT4 #(
		.INIT('h3113)
	) name1131 (
		_w262_,
		_w1346_,
		_w1347_,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h2)
	) name1132 (
		_w587_,
		_w1349_,
		_w1350_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1133 (
		_w713_,
		_w695_,
		_w706_,
		_w709_,
		_w1351_
	);
	LUT4 #(
		.INIT('h1331)
	) name1134 (
		_w262_,
		_w1346_,
		_w1347_,
		_w1351_,
		_w1352_
	);
	LUT4 #(
		.INIT('h807f)
	) name1135 (
		_w339_,
		_w356_,
		_w379_,
		_w384_,
		_w1353_
	);
	LUT4 #(
		.INIT('h2a08)
	) name1136 (
		_w262_,
		_w266_,
		_w378_,
		_w1353_,
		_w1354_
	);
	LUT3 #(
		.INIT('ha8)
	) name1137 (
		_w404_,
		_w1346_,
		_w1354_,
		_w1355_
	);
	LUT4 #(
		.INIT('hc6cc)
	) name1138 (
		_w439_,
		_w446_,
		_w449_,
		_w596_,
		_w1356_
	);
	LUT4 #(
		.INIT('he040)
	) name1139 (
		_w262_,
		_w358_,
		_w601_,
		_w1356_,
		_w1357_
	);
	LUT3 #(
		.INIT('h04)
	) name1140 (
		_w521_,
		_w522_,
		_w446_,
		_w1358_
	);
	LUT3 #(
		.INIT('ha8)
	) name1141 (
		_w358_,
		_w524_,
		_w526_,
		_w1359_
	);
	LUT2 #(
		.INIT('h1)
	) name1142 (
		_w1358_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h4)
	) name1143 (
		_w1357_,
		_w1360_,
		_w1361_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1144 (
		_w518_,
		_w1352_,
		_w1355_,
		_w1361_,
		_w1362_
	);
	LUT4 #(
		.INIT('h1311)
	) name1145 (
		_w254_,
		_w1345_,
		_w1350_,
		_w1362_,
		_w1363_
	);
	LUT2 #(
		.INIT('h2)
	) name1146 (
		\reg3_reg[16]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1364_
	);
	LUT3 #(
		.INIT('h07)
	) name1147 (
		_w606_,
		_w358_,
		_w1364_,
		_w1365_
	);
	LUT3 #(
		.INIT('h2f)
	) name1148 (
		\state_reg[0]/NET0131 ,
		_w1363_,
		_w1365_,
		_w1366_
	);
	LUT2 #(
		.INIT('h8)
	) name1149 (
		_w252_,
		_w324_,
		_w1367_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1150 (
		_w256_,
		_w258_,
		_w261_,
		_w324_,
		_w1368_
	);
	LUT4 #(
		.INIT('h0080)
	) name1151 (
		_w301_,
		_w311_,
		_w322_,
		_w326_,
		_w1369_
	);
	LUT3 #(
		.INIT('h80)
	) name1152 (
		_w266_,
		_w312_,
		_w314_,
		_w1370_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1153 (
		_w266_,
		_w331_,
		_w1369_,
		_w1370_,
		_w1371_
	);
	LUT4 #(
		.INIT('he040)
	) name1154 (
		_w262_,
		_w324_,
		_w404_,
		_w1371_,
		_w1372_
	);
	LUT3 #(
		.INIT('h78)
	) name1155 (
		_w323_,
		_w325_,
		_w467_,
		_w1373_
	);
	LUT4 #(
		.INIT('h15ea)
	) name1156 (
		_w482_,
		_w509_,
		_w511_,
		_w1373_,
		_w1374_
	);
	LUT4 #(
		.INIT('h40e0)
	) name1157 (
		_w262_,
		_w324_,
		_w518_,
		_w1374_,
		_w1375_
	);
	LUT4 #(
		.INIT('h08a2)
	) name1158 (
		_w262_,
		_w562_,
		_w837_,
		_w1373_,
		_w1376_
	);
	LUT4 #(
		.INIT('h2800)
	) name1159 (
		_w262_,
		_w467_,
		_w592_,
		_w601_,
		_w1377_
	);
	LUT3 #(
		.INIT('ha8)
	) name1160 (
		_w324_,
		_w524_,
		_w906_,
		_w1378_
	);
	LUT3 #(
		.INIT('h04)
	) name1161 (
		_w521_,
		_w522_,
		_w467_,
		_w1379_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		_w1378_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h4)
	) name1163 (
		_w1377_,
		_w1380_,
		_w1381_
	);
	LUT4 #(
		.INIT('h5700)
	) name1164 (
		_w587_,
		_w1368_,
		_w1376_,
		_w1381_,
		_w1382_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1165 (
		_w254_,
		_w1372_,
		_w1375_,
		_w1382_,
		_w1383_
	);
	LUT2 #(
		.INIT('h2)
	) name1166 (
		\reg3_reg[7]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1384_
	);
	LUT4 #(
		.INIT('h4800)
	) name1167 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w324_,
		_w1385_
	);
	LUT2 #(
		.INIT('h1)
	) name1168 (
		_w1384_,
		_w1385_,
		_w1386_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1169 (
		\state_reg[0]/NET0131 ,
		_w1367_,
		_w1383_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h8)
	) name1170 (
		_w252_,
		_w668_,
		_w1388_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1171 (
		_w256_,
		_w258_,
		_w261_,
		_w668_,
		_w1389_
	);
	LUT2 #(
		.INIT('h9)
	) name1172 (
		_w667_,
		_w671_,
		_w1390_
	);
	LUT4 #(
		.INIT('h8a20)
	) name1173 (
		_w262_,
		_w710_,
		_w720_,
		_w1390_,
		_w1391_
	);
	LUT3 #(
		.INIT('ha8)
	) name1174 (
		_w518_,
		_w1389_,
		_w1391_,
		_w1392_
	);
	LUT4 #(
		.INIT('h0200)
	) name1175 (
		_w266_,
		_w682_,
		_w681_,
		_w683_,
		_w1393_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1176 (
		_w266_,
		_w665_,
		_w1070_,
		_w1393_,
		_w1394_
	);
	LUT4 #(
		.INIT('hc840)
	) name1177 (
		_w262_,
		_w404_,
		_w668_,
		_w1394_,
		_w1395_
	);
	LUT4 #(
		.INIT('h070d)
	) name1178 (
		_w262_,
		_w776_,
		_w1389_,
		_w1390_,
		_w1396_
	);
	LUT4 #(
		.INIT('h0800)
	) name1179 (
		_w596_,
		_w598_,
		_w667_,
		_w798_,
		_w1397_
	);
	LUT4 #(
		.INIT('h870f)
	) name1180 (
		_w596_,
		_w598_,
		_w667_,
		_w798_,
		_w1398_
	);
	LUT4 #(
		.INIT('hc840)
	) name1181 (
		_w262_,
		_w601_,
		_w668_,
		_w1398_,
		_w1399_
	);
	LUT3 #(
		.INIT('h40)
	) name1182 (
		_w521_,
		_w522_,
		_w667_,
		_w1400_
	);
	LUT3 #(
		.INIT('he0)
	) name1183 (
		_w524_,
		_w526_,
		_w668_,
		_w1401_
	);
	LUT2 #(
		.INIT('h1)
	) name1184 (
		_w1400_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h4)
	) name1185 (
		_w1399_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1186 (
		_w587_,
		_w1396_,
		_w1395_,
		_w1403_,
		_w1404_
	);
	LUT4 #(
		.INIT('h1311)
	) name1187 (
		_w254_,
		_w1388_,
		_w1392_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h2)
	) name1188 (
		\reg3_reg[20]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1406_
	);
	LUT3 #(
		.INIT('h07)
	) name1189 (
		_w606_,
		_w668_,
		_w1406_,
		_w1407_
	);
	LUT3 #(
		.INIT('h2f)
	) name1190 (
		\state_reg[0]/NET0131 ,
		_w1405_,
		_w1407_,
		_w1408_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1191 (
		_w256_,
		_w258_,
		_w261_,
		_w520_,
		_w1409_
	);
	LUT2 #(
		.INIT('h8)
	) name1192 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1410_
	);
	LUT3 #(
		.INIT('h08)
	) name1193 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w524_,
		_w1411_
	);
	LUT3 #(
		.INIT('h8a)
	) name1194 (
		\reg2_reg[31]/NET0131 ,
		_w1409_,
		_w1411_,
		_w1412_
	);
	LUT3 #(
		.INIT('ha8)
	) name1195 (
		\datai[31]_pad ,
		_w266_,
		_w407_,
		_w1413_
	);
	LUT3 #(
		.INIT('ha8)
	) name1196 (
		\datai[30]_pad ,
		_w266_,
		_w407_,
		_w1414_
	);
	LUT4 #(
		.INIT('h0008)
	) name1197 (
		_w804_,
		_w806_,
		_w1267_,
		_w1414_,
		_w1415_
	);
	LUT3 #(
		.INIT('h82)
	) name1198 (
		_w601_,
		_w1413_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h8)
	) name1199 (
		_w525_,
		_w1413_,
		_w1417_
	);
	LUT4 #(
		.INIT('h0200)
	) name1200 (
		_w394_,
		_w624_,
		_w631_,
		_w813_,
		_w1418_
	);
	LUT4 #(
		.INIT('h000b)
	) name1201 (
		_w734_,
		_w737_,
		_w820_,
		_w1262_,
		_w1419_
	);
	LUT2 #(
		.INIT('h2)
	) name1202 (
		_w404_,
		_w1264_,
		_w1420_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w299_,
		_w1420_,
		_w1421_
	);
	LUT4 #(
		.INIT('h4055)
	) name1204 (
		_w1417_,
		_w1418_,
		_w1419_,
		_w1421_,
		_w1422_
	);
	LUT4 #(
		.INIT('h1311)
	) name1205 (
		_w970_,
		_w1305_,
		_w1416_,
		_w1422_,
		_w1423_
	);
	LUT3 #(
		.INIT('hce)
	) name1206 (
		_w1410_,
		_w1412_,
		_w1423_,
		_w1424_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1207 (
		_w256_,
		_w258_,
		_w261_,
		_w628_,
		_w1425_
	);
	LUT2 #(
		.INIT('h9)
	) name1208 (
		_w627_,
		_w631_,
		_w1426_
	);
	LUT3 #(
		.INIT('hd0)
	) name1209 (
		_w746_,
		_w768_,
		_w770_,
		_w1427_
	);
	LUT2 #(
		.INIT('h8)
	) name1210 (
		_w744_,
		_w746_,
		_w1428_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1211 (
		_w1322_,
		_w1323_,
		_w1324_,
		_w1428_,
		_w1429_
	);
	LUT2 #(
		.INIT('h8)
	) name1212 (
		_w778_,
		_w783_,
		_w1430_
	);
	LUT2 #(
		.INIT('h8)
	) name1213 (
		_w749_,
		_w777_,
		_w1431_
	);
	LUT4 #(
		.INIT('h8000)
	) name1214 (
		_w749_,
		_w777_,
		_w778_,
		_w783_,
		_w1432_
	);
	LUT3 #(
		.INIT('hb0)
	) name1215 (
		_w773_,
		_w777_,
		_w786_,
		_w1433_
	);
	LUT3 #(
		.INIT('hd0)
	) name1216 (
		_w783_,
		_w787_,
		_w792_,
		_w1434_
	);
	LUT3 #(
		.INIT('hd0)
	) name1217 (
		_w1430_,
		_w1433_,
		_w1434_,
		_w1435_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1218 (
		_w1427_,
		_w1429_,
		_w1432_,
		_w1435_,
		_w1436_
	);
	LUT4 #(
		.INIT('h1331)
	) name1219 (
		_w262_,
		_w1425_,
		_w1426_,
		_w1436_,
		_w1437_
	);
	LUT4 #(
		.INIT('h3933)
	) name1220 (
		_w394_,
		_w624_,
		_w631_,
		_w813_,
		_w1438_
	);
	LUT4 #(
		.INIT('h2a08)
	) name1221 (
		_w262_,
		_w266_,
		_w640_,
		_w1438_,
		_w1439_
	);
	LUT3 #(
		.INIT('ha8)
	) name1222 (
		_w404_,
		_w1425_,
		_w1439_,
		_w1440_
	);
	LUT4 #(
		.INIT('h2822)
	) name1223 (
		_w262_,
		_w627_,
		_w635_,
		_w804_,
		_w1441_
	);
	LUT3 #(
		.INIT('ha8)
	) name1224 (
		_w601_,
		_w1425_,
		_w1441_,
		_w1442_
	);
	LUT4 #(
		.INIT('hf800)
	) name1225 (
		_w698_,
		_w699_,
		_w701_,
		_w1330_,
		_w1443_
	);
	LUT4 #(
		.INIT('h2000)
	) name1226 (
		_w505_,
		_w697_,
		_w699_,
		_w1330_,
		_w1444_
	);
	LUT3 #(
		.INIT('h02)
	) name1227 (
		_w1329_,
		_w1443_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h8)
	) name1228 (
		_w690_,
		_w707_,
		_w1446_
	);
	LUT3 #(
		.INIT('h80)
	) name1229 (
		_w690_,
		_w707_,
		_w1328_,
		_w1447_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1230 (
		_w1329_,
		_w1443_,
		_w1444_,
		_w1447_,
		_w1448_
	);
	LUT3 #(
		.INIT('h07)
	) name1231 (
		_w690_,
		_w712_,
		_w715_,
		_w1449_
	);
	LUT3 #(
		.INIT('hb0)
	) name1232 (
		_w1327_,
		_w1446_,
		_w1449_,
		_w1450_
	);
	LUT2 #(
		.INIT('h8)
	) name1233 (
		_w649_,
		_w659_,
		_w1451_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		_w673_,
		_w688_,
		_w1452_
	);
	LUT4 #(
		.INIT('h8000)
	) name1235 (
		_w649_,
		_w659_,
		_w673_,
		_w688_,
		_w1453_
	);
	LUT3 #(
		.INIT('h07)
	) name1236 (
		_w673_,
		_w718_,
		_w721_,
		_w1454_
	);
	LUT3 #(
		.INIT('h0d)
	) name1237 (
		_w649_,
		_w723_,
		_w729_,
		_w1455_
	);
	LUT3 #(
		.INIT('hd0)
	) name1238 (
		_w1451_,
		_w1454_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1239 (
		_w1448_,
		_w1450_,
		_w1453_,
		_w1456_,
		_w1457_
	);
	LUT4 #(
		.INIT('h0880)
	) name1240 (
		_w262_,
		_w518_,
		_w1426_,
		_w1457_,
		_w1458_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1241 (
		_w256_,
		_w258_,
		_w261_,
		_w518_,
		_w1459_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name1242 (
		_w524_,
		_w526_,
		_w628_,
		_w1459_,
		_w1460_
	);
	LUT3 #(
		.INIT('h40)
	) name1243 (
		_w521_,
		_w522_,
		_w627_,
		_w1461_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w1460_,
		_w1461_,
		_w1462_
	);
	LUT3 #(
		.INIT('h10)
	) name1245 (
		_w1442_,
		_w1458_,
		_w1462_,
		_w1463_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1246 (
		_w587_,
		_w1437_,
		_w1440_,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h8)
	) name1247 (
		_w252_,
		_w628_,
		_w1465_
	);
	LUT4 #(
		.INIT('haa08)
	) name1248 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1464_,
		_w1465_,
		_w1466_
	);
	LUT2 #(
		.INIT('h2)
	) name1249 (
		\reg3_reg[26]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1467_
	);
	LUT3 #(
		.INIT('h07)
	) name1250 (
		_w606_,
		_w628_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('hb)
	) name1251 (
		_w1466_,
		_w1468_,
		_w1469_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1252 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[19]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1470_
	);
	LUT2 #(
		.INIT('h8)
	) name1253 (
		\reg0_reg[19]/NET0131 ,
		_w252_,
		_w1471_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1254 (
		\reg0_reg[19]/NET0131 ,
		_w846_,
		_w917_,
		_w1066_,
		_w1472_
	);
	LUT2 #(
		.INIT('h2)
	) name1255 (
		_w587_,
		_w1472_,
		_w1473_
	);
	LUT4 #(
		.INIT('hc535)
	) name1256 (
		\reg0_reg[19]/NET0131 ,
		_w876_,
		_w917_,
		_w1066_,
		_w1474_
	);
	LUT2 #(
		.INIT('h2)
	) name1257 (
		_w525_,
		_w686_,
		_w1475_
	);
	LUT3 #(
		.INIT('h01)
	) name1258 (
		_w1074_,
		_w1077_,
		_w1475_,
		_w1476_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1259 (
		_w917_,
		_w1074_,
		_w1077_,
		_w1475_,
		_w1477_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1260 (
		\reg0_reg[19]/NET0131 ,
		_w923_,
		_w924_,
		_w926_,
		_w1478_
	);
	LUT4 #(
		.INIT('h0031)
	) name1261 (
		_w518_,
		_w1477_,
		_w1474_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('h1311)
	) name1262 (
		_w254_,
		_w1471_,
		_w1473_,
		_w1479_,
		_w1480_
	);
	LUT3 #(
		.INIT('hce)
	) name1263 (
		\state_reg[0]/NET0131 ,
		_w1470_,
		_w1480_,
		_w1481_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1264 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[20]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1482_
	);
	LUT2 #(
		.INIT('h8)
	) name1265 (
		\reg0_reg[20]/NET0131 ,
		_w252_,
		_w1483_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1266 (
		\reg0_reg[20]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1484_
	);
	LUT4 #(
		.INIT('hb040)
	) name1267 (
		_w710_,
		_w720_,
		_w917_,
		_w1390_,
		_w1485_
	);
	LUT3 #(
		.INIT('ha8)
	) name1268 (
		_w518_,
		_w1484_,
		_w1485_,
		_w1486_
	);
	LUT4 #(
		.INIT('hc808)
	) name1269 (
		\reg0_reg[20]/NET0131 ,
		_w404_,
		_w917_,
		_w1394_,
		_w1487_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1270 (
		\reg0_reg[20]/NET0131 ,
		_w776_,
		_w917_,
		_w1390_,
		_w1488_
	);
	LUT2 #(
		.INIT('h8)
	) name1271 (
		_w525_,
		_w667_,
		_w1489_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1272 (
		_w601_,
		_w917_,
		_w1398_,
		_w1489_,
		_w1490_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1273 (
		\reg0_reg[20]/NET0131 ,
		_w923_,
		_w924_,
		_w1154_,
		_w1491_
	);
	LUT2 #(
		.INIT('h1)
	) name1274 (
		_w1490_,
		_w1491_,
		_w1492_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1275 (
		_w587_,
		_w1488_,
		_w1487_,
		_w1492_,
		_w1493_
	);
	LUT4 #(
		.INIT('h1311)
	) name1276 (
		_w254_,
		_w1483_,
		_w1486_,
		_w1493_,
		_w1494_
	);
	LUT3 #(
		.INIT('hce)
	) name1277 (
		\state_reg[0]/NET0131 ,
		_w1482_,
		_w1494_,
		_w1495_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1278 (
		\reg0_reg[29]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1496_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1279 (
		\reg0_reg[29]/NET0131 ,
		_w404_,
		_w917_,
		_w1265_,
		_w1497_
	);
	LUT4 #(
		.INIT('h8288)
	) name1280 (
		_w917_,
		_w1270_,
		_w1298_,
		_w1301_,
		_w1498_
	);
	LUT3 #(
		.INIT('ha8)
	) name1281 (
		_w587_,
		_w1496_,
		_w1498_,
		_w1499_
	);
	LUT4 #(
		.INIT('hc808)
	) name1282 (
		\reg0_reg[29]/NET0131 ,
		_w518_,
		_w917_,
		_w1287_,
		_w1500_
	);
	LUT4 #(
		.INIT('h8070)
	) name1283 (
		_w804_,
		_w806_,
		_w917_,
		_w1267_,
		_w1501_
	);
	LUT3 #(
		.INIT('h8a)
	) name1284 (
		\reg0_reg[29]/NET0131 ,
		_w923_,
		_w924_,
		_w1502_
	);
	LUT2 #(
		.INIT('h8)
	) name1285 (
		_w917_,
		_w1306_,
		_w1503_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w1502_,
		_w1503_,
		_w1504_
	);
	LUT4 #(
		.INIT('h5700)
	) name1287 (
		_w601_,
		_w1496_,
		_w1501_,
		_w1504_,
		_w1505_
	);
	LUT4 #(
		.INIT('h0100)
	) name1288 (
		_w1497_,
		_w1500_,
		_w1499_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h8)
	) name1289 (
		\reg0_reg[29]/NET0131 ,
		_w252_,
		_w1507_
	);
	LUT4 #(
		.INIT('haa08)
	) name1290 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1506_,
		_w1507_,
		_w1508_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1291 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[29]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1509_
	);
	LUT2 #(
		.INIT('he)
	) name1292 (
		_w1508_,
		_w1509_,
		_w1510_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1293 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[12]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1511_
	);
	LUT2 #(
		.INIT('h8)
	) name1294 (
		\reg1_reg[12]/NET0131 ,
		_w252_,
		_w1512_
	);
	LUT4 #(
		.INIT('haa02)
	) name1295 (
		\reg1_reg[12]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1513_
	);
	LUT4 #(
		.INIT('hd020)
	) name1296 (
		_w695_,
		_w706_,
		_w946_,
		_w1046_,
		_w1514_
	);
	LUT4 #(
		.INIT('hc535)
	) name1297 (
		\reg1_reg[12]/NET0131 ,
		_w423_,
		_w946_,
		_w1027_,
		_w1515_
	);
	LUT3 #(
		.INIT('ha2)
	) name1298 (
		\reg1_reg[12]/NET0131 ,
		_w924_,
		_w959_,
		_w1516_
	);
	LUT2 #(
		.INIT('h4)
	) name1299 (
		_w423_,
		_w525_,
		_w1517_
	);
	LUT2 #(
		.INIT('h8)
	) name1300 (
		_w946_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h1)
	) name1301 (
		_w1516_,
		_w1518_,
		_w1519_
	);
	LUT3 #(
		.INIT('hd0)
	) name1302 (
		_w601_,
		_w1515_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h5700)
	) name1303 (
		_w518_,
		_w1513_,
		_w1514_,
		_w1520_,
		_w1521_
	);
	LUT4 #(
		.INIT('h20d0)
	) name1304 (
		_w755_,
		_w766_,
		_w946_,
		_w1046_,
		_w1522_
	);
	LUT3 #(
		.INIT('ha8)
	) name1305 (
		_w587_,
		_w1513_,
		_w1522_,
		_w1523_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1306 (
		\reg1_reg[12]/NET0131 ,
		_w946_,
		_w1056_,
		_w1057_,
		_w1524_
	);
	LUT2 #(
		.INIT('h2)
	) name1307 (
		_w404_,
		_w1524_,
		_w1525_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1308 (
		_w254_,
		_w1523_,
		_w1525_,
		_w1521_,
		_w1526_
	);
	LUT4 #(
		.INIT('heeec)
	) name1309 (
		\state_reg[0]/NET0131 ,
		_w1511_,
		_w1512_,
		_w1526_,
		_w1527_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1310 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[19]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1528_
	);
	LUT2 #(
		.INIT('h8)
	) name1311 (
		\reg1_reg[19]/NET0131 ,
		_w252_,
		_w1529_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1312 (
		\reg1_reg[19]/NET0131 ,
		_w846_,
		_w946_,
		_w1066_,
		_w1530_
	);
	LUT2 #(
		.INIT('h2)
	) name1313 (
		_w587_,
		_w1530_,
		_w1531_
	);
	LUT4 #(
		.INIT('hc535)
	) name1314 (
		\reg1_reg[19]/NET0131 ,
		_w876_,
		_w946_,
		_w1066_,
		_w1532_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1315 (
		_w946_,
		_w1074_,
		_w1077_,
		_w1475_,
		_w1533_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1316 (
		\reg1_reg[19]/NET0131 ,
		_w924_,
		_w949_,
		_w950_,
		_w1534_
	);
	LUT4 #(
		.INIT('h0031)
	) name1317 (
		_w518_,
		_w1533_,
		_w1532_,
		_w1534_,
		_w1535_
	);
	LUT4 #(
		.INIT('h1311)
	) name1318 (
		_w254_,
		_w1529_,
		_w1531_,
		_w1535_,
		_w1536_
	);
	LUT3 #(
		.INIT('hce)
	) name1319 (
		\state_reg[0]/NET0131 ,
		_w1528_,
		_w1536_,
		_w1537_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1320 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[20]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1538_
	);
	LUT2 #(
		.INIT('h8)
	) name1321 (
		\reg1_reg[20]/NET0131 ,
		_w252_,
		_w1539_
	);
	LUT4 #(
		.INIT('haa02)
	) name1322 (
		\reg1_reg[20]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1540_
	);
	LUT4 #(
		.INIT('hb040)
	) name1323 (
		_w710_,
		_w720_,
		_w946_,
		_w1390_,
		_w1541_
	);
	LUT3 #(
		.INIT('ha8)
	) name1324 (
		_w518_,
		_w1540_,
		_w1541_,
		_w1542_
	);
	LUT4 #(
		.INIT('hc808)
	) name1325 (
		\reg1_reg[20]/NET0131 ,
		_w404_,
		_w946_,
		_w1394_,
		_w1543_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1326 (
		\reg1_reg[20]/NET0131 ,
		_w776_,
		_w946_,
		_w1390_,
		_w1544_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1327 (
		_w601_,
		_w946_,
		_w1398_,
		_w1489_,
		_w1545_
	);
	LUT3 #(
		.INIT('ha2)
	) name1328 (
		\reg1_reg[20]/NET0131 ,
		_w924_,
		_w949_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		_w1545_,
		_w1546_,
		_w1547_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1330 (
		_w587_,
		_w1544_,
		_w1543_,
		_w1547_,
		_w1548_
	);
	LUT4 #(
		.INIT('h1311)
	) name1331 (
		_w254_,
		_w1539_,
		_w1542_,
		_w1548_,
		_w1549_
	);
	LUT3 #(
		.INIT('hce)
	) name1332 (
		\state_reg[0]/NET0131 ,
		_w1538_,
		_w1549_,
		_w1550_
	);
	LUT4 #(
		.INIT('haa02)
	) name1333 (
		\reg1_reg[26]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1551_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1334 (
		\reg1_reg[26]/NET0131 ,
		_w946_,
		_w1426_,
		_w1436_,
		_w1552_
	);
	LUT4 #(
		.INIT('h7020)
	) name1335 (
		_w266_,
		_w640_,
		_w946_,
		_w1438_,
		_w1553_
	);
	LUT3 #(
		.INIT('ha8)
	) name1336 (
		_w404_,
		_w1551_,
		_w1553_,
		_w1554_
	);
	LUT4 #(
		.INIT('h2822)
	) name1337 (
		_w601_,
		_w627_,
		_w635_,
		_w804_,
		_w1555_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		_w525_,
		_w627_,
		_w1556_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1339 (
		_w518_,
		_w1426_,
		_w1457_,
		_w1556_,
		_w1557_
	);
	LUT4 #(
		.INIT('h0002)
	) name1340 (
		_w924_,
		_w959_,
		_w960_,
		_w1220_,
		_w1558_
	);
	LUT2 #(
		.INIT('h2)
	) name1341 (
		\reg1_reg[26]/NET0131 ,
		_w1558_,
		_w1559_
	);
	LUT4 #(
		.INIT('h0075)
	) name1342 (
		_w946_,
		_w1555_,
		_w1557_,
		_w1559_,
		_w1560_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1343 (
		_w587_,
		_w1552_,
		_w1554_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h8)
	) name1344 (
		\reg1_reg[26]/NET0131 ,
		_w252_,
		_w1562_
	);
	LUT4 #(
		.INIT('haa08)
	) name1345 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1561_,
		_w1562_,
		_w1563_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1346 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[26]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1564_
	);
	LUT2 #(
		.INIT('he)
	) name1347 (
		_w1563_,
		_w1564_,
		_w1565_
	);
	LUT4 #(
		.INIT('haa02)
	) name1348 (
		\reg1_reg[29]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1566_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1349 (
		\reg1_reg[29]/NET0131 ,
		_w404_,
		_w946_,
		_w1265_,
		_w1567_
	);
	LUT4 #(
		.INIT('h8288)
	) name1350 (
		_w946_,
		_w1270_,
		_w1298_,
		_w1301_,
		_w1568_
	);
	LUT3 #(
		.INIT('ha8)
	) name1351 (
		_w587_,
		_w1566_,
		_w1568_,
		_w1569_
	);
	LUT4 #(
		.INIT('hc808)
	) name1352 (
		\reg1_reg[29]/NET0131 ,
		_w518_,
		_w946_,
		_w1287_,
		_w1570_
	);
	LUT4 #(
		.INIT('h8070)
	) name1353 (
		_w804_,
		_w806_,
		_w946_,
		_w1267_,
		_w1571_
	);
	LUT3 #(
		.INIT('ha2)
	) name1354 (
		\reg1_reg[29]/NET0131 ,
		_w924_,
		_w959_,
		_w1572_
	);
	LUT2 #(
		.INIT('h8)
	) name1355 (
		_w946_,
		_w1306_,
		_w1573_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		_w1572_,
		_w1573_,
		_w1574_
	);
	LUT4 #(
		.INIT('h5700)
	) name1357 (
		_w601_,
		_w1566_,
		_w1571_,
		_w1574_,
		_w1575_
	);
	LUT4 #(
		.INIT('h0100)
	) name1358 (
		_w1567_,
		_w1570_,
		_w1569_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h8)
	) name1359 (
		\reg1_reg[29]/NET0131 ,
		_w252_,
		_w1577_
	);
	LUT4 #(
		.INIT('haa08)
	) name1360 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1576_,
		_w1577_,
		_w1578_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1361 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[29]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1579_
	);
	LUT2 #(
		.INIT('he)
	) name1362 (
		_w1578_,
		_w1579_,
		_w1580_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1363 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[12]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1581_
	);
	LUT2 #(
		.INIT('h8)
	) name1364 (
		\reg2_reg[12]/NET0131 ,
		_w252_,
		_w1582_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1365 (
		\reg2_reg[12]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1583_
	);
	LUT4 #(
		.INIT('hd020)
	) name1366 (
		_w695_,
		_w706_,
		_w970_,
		_w1046_,
		_w1584_
	);
	LUT4 #(
		.INIT('hc535)
	) name1367 (
		\reg2_reg[12]/NET0131 ,
		_w423_,
		_w970_,
		_w1027_,
		_w1585_
	);
	LUT3 #(
		.INIT('ha8)
	) name1368 (
		\reg2_reg[12]/NET0131 ,
		_w524_,
		_w976_,
		_w1586_
	);
	LUT2 #(
		.INIT('h8)
	) name1369 (
		_w520_,
		_w340_,
		_w1587_
	);
	LUT3 #(
		.INIT('h07)
	) name1370 (
		_w970_,
		_w1517_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h4)
	) name1371 (
		_w1586_,
		_w1588_,
		_w1589_
	);
	LUT3 #(
		.INIT('hd0)
	) name1372 (
		_w601_,
		_w1585_,
		_w1589_,
		_w1590_
	);
	LUT4 #(
		.INIT('h5700)
	) name1373 (
		_w518_,
		_w1583_,
		_w1584_,
		_w1590_,
		_w1591_
	);
	LUT4 #(
		.INIT('h20d0)
	) name1374 (
		_w755_,
		_w766_,
		_w970_,
		_w1046_,
		_w1592_
	);
	LUT3 #(
		.INIT('ha8)
	) name1375 (
		_w587_,
		_w1583_,
		_w1592_,
		_w1593_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1376 (
		\reg2_reg[12]/NET0131 ,
		_w970_,
		_w1056_,
		_w1057_,
		_w1594_
	);
	LUT2 #(
		.INIT('h2)
	) name1377 (
		_w404_,
		_w1594_,
		_w1595_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1378 (
		_w254_,
		_w1593_,
		_w1595_,
		_w1591_,
		_w1596_
	);
	LUT4 #(
		.INIT('heeec)
	) name1379 (
		\state_reg[0]/NET0131 ,
		_w1581_,
		_w1582_,
		_w1596_,
		_w1597_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1380 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[19]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1598_
	);
	LUT2 #(
		.INIT('h8)
	) name1381 (
		\reg2_reg[19]/NET0131 ,
		_w252_,
		_w1599_
	);
	LUT3 #(
		.INIT('h82)
	) name1382 (
		_w587_,
		_w846_,
		_w1066_,
		_w1600_
	);
	LUT3 #(
		.INIT('h28)
	) name1383 (
		_w518_,
		_w876_,
		_w1066_,
		_w1601_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1384 (
		_w970_,
		_w1476_,
		_w1601_,
		_w1600_,
		_w1602_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		_w520_,
		_w680_,
		_w1603_
	);
	LUT4 #(
		.INIT('h6662)
	) name1386 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w1604_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1387 (
		_w256_,
		_w258_,
		_w261_,
		_w1604_,
		_w1605_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1388 (
		\reg2_reg[19]/NET0131 ,
		_w524_,
		_w1237_,
		_w1605_,
		_w1606_
	);
	LUT2 #(
		.INIT('h1)
	) name1389 (
		_w1603_,
		_w1606_,
		_w1607_
	);
	LUT4 #(
		.INIT('h1311)
	) name1390 (
		_w254_,
		_w1599_,
		_w1602_,
		_w1607_,
		_w1608_
	);
	LUT3 #(
		.INIT('hce)
	) name1391 (
		\state_reg[0]/NET0131 ,
		_w1598_,
		_w1608_,
		_w1609_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1392 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[20]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1610_
	);
	LUT2 #(
		.INIT('h8)
	) name1393 (
		\reg2_reg[20]/NET0131 ,
		_w252_,
		_w1611_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1394 (
		\reg2_reg[20]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1612_
	);
	LUT4 #(
		.INIT('hb040)
	) name1395 (
		_w710_,
		_w720_,
		_w970_,
		_w1390_,
		_w1613_
	);
	LUT3 #(
		.INIT('ha8)
	) name1396 (
		_w518_,
		_w1612_,
		_w1613_,
		_w1614_
	);
	LUT4 #(
		.INIT('hc808)
	) name1397 (
		\reg2_reg[20]/NET0131 ,
		_w404_,
		_w970_,
		_w1394_,
		_w1615_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1398 (
		\reg2_reg[20]/NET0131 ,
		_w776_,
		_w970_,
		_w1390_,
		_w1616_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1399 (
		_w601_,
		_w970_,
		_w1398_,
		_w1489_,
		_w1617_
	);
	LUT2 #(
		.INIT('h8)
	) name1400 (
		_w520_,
		_w668_,
		_w1618_
	);
	LUT4 #(
		.INIT('h0057)
	) name1401 (
		\reg2_reg[20]/NET0131 ,
		_w524_,
		_w1237_,
		_w1618_,
		_w1619_
	);
	LUT2 #(
		.INIT('h4)
	) name1402 (
		_w1617_,
		_w1619_,
		_w1620_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1403 (
		_w587_,
		_w1616_,
		_w1615_,
		_w1620_,
		_w1621_
	);
	LUT4 #(
		.INIT('h1311)
	) name1404 (
		_w254_,
		_w1611_,
		_w1614_,
		_w1621_,
		_w1622_
	);
	LUT3 #(
		.INIT('hce)
	) name1405 (
		\state_reg[0]/NET0131 ,
		_w1610_,
		_w1622_,
		_w1623_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1406 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[12]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1624_
	);
	LUT2 #(
		.INIT('h8)
	) name1407 (
		\reg0_reg[12]/NET0131 ,
		_w252_,
		_w1625_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1408 (
		\reg0_reg[12]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1626_
	);
	LUT4 #(
		.INIT('h20d0)
	) name1409 (
		_w755_,
		_w766_,
		_w917_,
		_w1046_,
		_w1627_
	);
	LUT4 #(
		.INIT('hc535)
	) name1410 (
		\reg0_reg[12]/NET0131 ,
		_w423_,
		_w917_,
		_w1027_,
		_w1628_
	);
	LUT3 #(
		.INIT('h8a)
	) name1411 (
		\reg0_reg[12]/NET0131 ,
		_w923_,
		_w924_,
		_w1629_
	);
	LUT2 #(
		.INIT('h8)
	) name1412 (
		_w917_,
		_w1517_,
		_w1630_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		_w1629_,
		_w1630_,
		_w1631_
	);
	LUT3 #(
		.INIT('hd0)
	) name1414 (
		_w601_,
		_w1628_,
		_w1631_,
		_w1632_
	);
	LUT4 #(
		.INIT('h5700)
	) name1415 (
		_w587_,
		_w1626_,
		_w1627_,
		_w1632_,
		_w1633_
	);
	LUT4 #(
		.INIT('hd020)
	) name1416 (
		_w695_,
		_w706_,
		_w917_,
		_w1046_,
		_w1634_
	);
	LUT3 #(
		.INIT('ha8)
	) name1417 (
		_w518_,
		_w1626_,
		_w1634_,
		_w1635_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1418 (
		\reg0_reg[12]/NET0131 ,
		_w917_,
		_w1056_,
		_w1057_,
		_w1636_
	);
	LUT2 #(
		.INIT('h2)
	) name1419 (
		_w404_,
		_w1636_,
		_w1637_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1420 (
		_w254_,
		_w1635_,
		_w1637_,
		_w1633_,
		_w1638_
	);
	LUT4 #(
		.INIT('heeec)
	) name1421 (
		\state_reg[0]/NET0131 ,
		_w1624_,
		_w1625_,
		_w1638_,
		_w1639_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1422 (
		_w256_,
		_w258_,
		_w261_,
		_w387_,
		_w1640_
	);
	LUT4 #(
		.INIT('h10ef)
	) name1423 (
		_w389_,
		_w388_,
		_w390_,
		_w678_,
		_w1641_
	);
	LUT4 #(
		.INIT('h08a2)
	) name1424 (
		_w262_,
		_w1427_,
		_w1429_,
		_w1641_,
		_w1642_
	);
	LUT3 #(
		.INIT('ha8)
	) name1425 (
		_w587_,
		_w1640_,
		_w1642_,
		_w1643_
	);
	LUT4 #(
		.INIT('h5510)
	) name1426 (
		_w266_,
		_w394_,
		_w684_,
		_w898_,
		_w1644_
	);
	LUT4 #(
		.INIT('h0200)
	) name1427 (
		_w266_,
		_w382_,
		_w381_,
		_w383_,
		_w1645_
	);
	LUT4 #(
		.INIT('h3331)
	) name1428 (
		_w262_,
		_w1640_,
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT4 #(
		.INIT('h8070)
	) name1429 (
		_w596_,
		_w598_,
		_w601_,
		_w678_,
		_w1647_
	);
	LUT4 #(
		.INIT('h8a20)
	) name1430 (
		_w518_,
		_w1448_,
		_w1450_,
		_w1641_,
		_w1648_
	);
	LUT3 #(
		.INIT('h40)
	) name1431 (
		_w521_,
		_w522_,
		_w678_,
		_w1649_
	);
	LUT4 #(
		.INIT('h6e7d)
	) name1432 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w1650_
	);
	LUT4 #(
		.INIT('h001f)
	) name1433 (
		_w256_,
		_w258_,
		_w261_,
		_w1650_,
		_w1651_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1434 (
		_w387_,
		_w524_,
		_w526_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w1649_,
		_w1652_,
		_w1653_
	);
	LUT4 #(
		.INIT('h5700)
	) name1436 (
		_w262_,
		_w1647_,
		_w1648_,
		_w1653_,
		_w1654_
	);
	LUT3 #(
		.INIT('hd0)
	) name1437 (
		_w404_,
		_w1646_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h8)
	) name1438 (
		_w252_,
		_w387_,
		_w1656_
	);
	LUT4 #(
		.INIT('h0075)
	) name1439 (
		_w254_,
		_w1643_,
		_w1655_,
		_w1656_,
		_w1657_
	);
	LUT4 #(
		.INIT('h4800)
	) name1440 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w387_,
		_w1658_
	);
	LUT2 #(
		.INIT('h2)
	) name1441 (
		\reg3_reg[18]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1659_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		_w1658_,
		_w1659_,
		_w1660_
	);
	LUT3 #(
		.INIT('h2f)
	) name1443 (
		\state_reg[0]/NET0131 ,
		_w1657_,
		_w1660_,
		_w1661_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1444 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[25]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1662_
	);
	LUT2 #(
		.INIT('h8)
	) name1445 (
		\reg2_reg[25]/NET0131 ,
		_w252_,
		_w1663_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1446 (
		\reg2_reg[25]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1664_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name1447 (
		_w631_,
		_w640_,
		_w647_,
		_w899_,
		_w1665_
	);
	LUT4 #(
		.INIT('h2070)
	) name1448 (
		_w266_,
		_w647_,
		_w970_,
		_w1665_,
		_w1666_
	);
	LUT3 #(
		.INIT('ha8)
	) name1449 (
		_w404_,
		_w1664_,
		_w1666_,
		_w1667_
	);
	LUT4 #(
		.INIT('h5655)
	) name1450 (
		_w635_,
		_w638_,
		_w637_,
		_w639_,
		_w1668_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1451 (
		_w437_,
		_w452_,
		_w459_,
		_w1274_,
		_w1669_
	);
	LUT4 #(
		.INIT('h0070)
	) name1452 (
		_w513_,
		_w1275_,
		_w1276_,
		_w1669_,
		_w1670_
	);
	LUT4 #(
		.INIT('hc34b)
	) name1453 (
		_w1279_,
		_w1283_,
		_w1668_,
		_w1670_,
		_w1671_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1454 (
		\reg2_reg[25]/NET0131 ,
		_w518_,
		_w970_,
		_w1671_,
		_w1672_
	);
	LUT4 #(
		.INIT('ha200)
	) name1455 (
		_w555_,
		_w566_,
		_w584_,
		_w1291_,
		_w1673_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1456 (
		_w537_,
		_w540_,
		_w551_,
		_w1290_,
		_w1674_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1457 (
		_w1292_,
		_w1294_,
		_w1674_,
		_w1673_,
		_w1675_
	);
	LUT4 #(
		.INIT('h0a82)
	) name1458 (
		_w970_,
		_w1300_,
		_w1668_,
		_w1675_,
		_w1676_
	);
	LUT4 #(
		.INIT('h3c55)
	) name1459 (
		\reg2_reg[25]/NET0131 ,
		_w635_,
		_w804_,
		_w970_,
		_w1677_
	);
	LUT3 #(
		.INIT('ha8)
	) name1460 (
		\reg2_reg[25]/NET0131 ,
		_w524_,
		_w976_,
		_w1678_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		_w520_,
		_w636_,
		_w1679_
	);
	LUT2 #(
		.INIT('h8)
	) name1462 (
		_w525_,
		_w635_,
		_w1680_
	);
	LUT3 #(
		.INIT('h13)
	) name1463 (
		_w970_,
		_w1679_,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h4)
	) name1464 (
		_w1678_,
		_w1681_,
		_w1682_
	);
	LUT3 #(
		.INIT('hd0)
	) name1465 (
		_w601_,
		_w1677_,
		_w1682_,
		_w1683_
	);
	LUT4 #(
		.INIT('h5700)
	) name1466 (
		_w587_,
		_w1664_,
		_w1676_,
		_w1683_,
		_w1684_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1467 (
		_w254_,
		_w1667_,
		_w1672_,
		_w1684_,
		_w1685_
	);
	LUT4 #(
		.INIT('heeec)
	) name1468 (
		\state_reg[0]/NET0131 ,
		_w1662_,
		_w1663_,
		_w1685_,
		_w1686_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1469 (
		_w256_,
		_w258_,
		_w261_,
		_w654_,
		_w1687_
	);
	LUT2 #(
		.INIT('h9)
	) name1470 (
		_w652_,
		_w657_,
		_w1688_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1471 (
		_w1327_,
		_w1328_,
		_w1331_,
		_w1446_,
		_w1689_
	);
	LUT4 #(
		.INIT('h50d0)
	) name1472 (
		_w1452_,
		_w1449_,
		_w1454_,
		_w1689_,
		_w1690_
	);
	LUT4 #(
		.INIT('h3113)
	) name1473 (
		_w262_,
		_w1687_,
		_w1688_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('hb0)
	) name1474 (
		_w1427_,
		_w1431_,
		_w1433_,
		_w1692_
	);
	LUT4 #(
		.INIT('h87f0)
	) name1475 (
		_w1429_,
		_w1431_,
		_w1688_,
		_w1692_,
		_w1693_
	);
	LUT4 #(
		.INIT('h40c8)
	) name1476 (
		_w262_,
		_w587_,
		_w654_,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h2)
	) name1477 (
		_w266_,
		_w665_,
		_w1695_
	);
	LUT3 #(
		.INIT('h2a)
	) name1478 (
		_w615_,
		_w809_,
		_w1070_,
		_w1696_
	);
	LUT2 #(
		.INIT('h1)
	) name1479 (
		_w266_,
		_w899_,
		_w1697_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1480 (
		_w404_,
		_w1695_,
		_w1696_,
		_w1697_,
		_w1698_
	);
	LUT3 #(
		.INIT('h8a)
	) name1481 (
		_w652_,
		_w660_,
		_w1397_,
		_w1699_
	);
	LUT2 #(
		.INIT('h2)
	) name1482 (
		_w601_,
		_w1134_,
		_w1700_
	);
	LUT2 #(
		.INIT('h4)
	) name1483 (
		_w1699_,
		_w1700_,
		_w1701_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name1484 (
		_w524_,
		_w526_,
		_w654_,
		_w1078_,
		_w1702_
	);
	LUT3 #(
		.INIT('h40)
	) name1485 (
		_w521_,
		_w522_,
		_w652_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT4 #(
		.INIT('h5700)
	) name1487 (
		_w262_,
		_w1698_,
		_w1701_,
		_w1704_,
		_w1705_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1488 (
		_w518_,
		_w1691_,
		_w1694_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('h8)
	) name1489 (
		_w252_,
		_w654_,
		_w1707_
	);
	LUT4 #(
		.INIT('haa08)
	) name1490 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1706_,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h2)
	) name1491 (
		\reg3_reg[22]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1709_
	);
	LUT3 #(
		.INIT('h07)
	) name1492 (
		_w606_,
		_w654_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('hb)
	) name1493 (
		_w1708_,
		_w1710_,
		_w1711_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1494 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[30]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1712_
	);
	LUT2 #(
		.INIT('h8)
	) name1495 (
		\reg2_reg[30]/NET0131 ,
		_w252_,
		_w1713_
	);
	LUT4 #(
		.INIT('h08f7)
	) name1496 (
		_w804_,
		_w806_,
		_w1267_,
		_w1414_,
		_w1714_
	);
	LUT4 #(
		.INIT('h5455)
	) name1497 (
		\reg2_reg[30]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1715_
	);
	LUT2 #(
		.INIT('h2)
	) name1498 (
		_w601_,
		_w1715_,
		_w1716_
	);
	LUT3 #(
		.INIT('hd0)
	) name1499 (
		_w970_,
		_w1714_,
		_w1716_,
		_w1717_
	);
	LUT2 #(
		.INIT('h8)
	) name1500 (
		_w525_,
		_w1414_,
		_w1718_
	);
	LUT4 #(
		.INIT('h008f)
	) name1501 (
		_w1418_,
		_w1419_,
		_w1421_,
		_w1718_,
		_w1719_
	);
	LUT3 #(
		.INIT('h02)
	) name1502 (
		_w401_,
		_w398_,
		_w399_,
		_w1720_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1503 (
		_w256_,
		_w258_,
		_w261_,
		_w1720_,
		_w1721_
	);
	LUT4 #(
		.INIT('h0507)
	) name1504 (
		\reg2_reg[30]/NET0131 ,
		_w524_,
		_w1305_,
		_w1721_,
		_w1722_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1505 (
		_w970_,
		_w1719_,
		_w1717_,
		_w1722_,
		_w1723_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1506 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1713_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('he)
	) name1507 (
		_w1712_,
		_w1724_,
		_w1725_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1508 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[16]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1726_
	);
	LUT2 #(
		.INIT('h8)
	) name1509 (
		\reg0_reg[16]/NET0131 ,
		_w252_,
		_w1727_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1510 (
		\reg0_reg[16]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1728_
	);
	LUT4 #(
		.INIT('hd11d)
	) name1511 (
		\reg0_reg[16]/NET0131 ,
		_w917_,
		_w1347_,
		_w1348_,
		_w1729_
	);
	LUT2 #(
		.INIT('h2)
	) name1512 (
		_w587_,
		_w1729_,
		_w1730_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1513 (
		\reg0_reg[16]/NET0131 ,
		_w917_,
		_w1347_,
		_w1351_,
		_w1731_
	);
	LUT4 #(
		.INIT('h7020)
	) name1514 (
		_w266_,
		_w378_,
		_w917_,
		_w1353_,
		_w1732_
	);
	LUT3 #(
		.INIT('ha8)
	) name1515 (
		_w404_,
		_w1728_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('h4)
	) name1516 (
		_w446_,
		_w525_,
		_w1734_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1517 (
		_w601_,
		_w917_,
		_w1356_,
		_w1734_,
		_w1735_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1518 (
		\reg0_reg[16]/NET0131 ,
		_w923_,
		_w924_,
		_w1154_,
		_w1736_
	);
	LUT2 #(
		.INIT('h1)
	) name1519 (
		_w1735_,
		_w1736_,
		_w1737_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1520 (
		_w518_,
		_w1731_,
		_w1733_,
		_w1737_,
		_w1738_
	);
	LUT4 #(
		.INIT('h1311)
	) name1521 (
		_w254_,
		_w1727_,
		_w1730_,
		_w1738_,
		_w1739_
	);
	LUT3 #(
		.INIT('hce)
	) name1522 (
		\state_reg[0]/NET0131 ,
		_w1726_,
		_w1739_,
		_w1740_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1523 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[7]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1741_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		\reg2_reg[7]/NET0131 ,
		_w252_,
		_w1742_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1525 (
		\reg2_reg[7]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1743_
	);
	LUT4 #(
		.INIT('hc808)
	) name1526 (
		\reg2_reg[7]/NET0131 ,
		_w404_,
		_w970_,
		_w1371_,
		_w1744_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1527 (
		\reg2_reg[7]/NET0131 ,
		_w518_,
		_w970_,
		_w1374_,
		_w1745_
	);
	LUT4 #(
		.INIT('h20d0)
	) name1528 (
		_w562_,
		_w837_,
		_w970_,
		_w1373_,
		_w1746_
	);
	LUT2 #(
		.INIT('h4)
	) name1529 (
		_w467_,
		_w525_,
		_w1747_
	);
	LUT4 #(
		.INIT('h009f)
	) name1530 (
		_w467_,
		_w592_,
		_w601_,
		_w1747_,
		_w1748_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1531 (
		\reg2_reg[7]/NET0131 ,
		_w524_,
		_w976_,
		_w991_,
		_w1749_
	);
	LUT2 #(
		.INIT('h8)
	) name1532 (
		_w520_,
		_w324_,
		_w1750_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		_w1749_,
		_w1750_,
		_w1751_
	);
	LUT3 #(
		.INIT('hd0)
	) name1534 (
		_w970_,
		_w1748_,
		_w1751_,
		_w1752_
	);
	LUT4 #(
		.INIT('h5700)
	) name1535 (
		_w587_,
		_w1743_,
		_w1746_,
		_w1752_,
		_w1753_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1536 (
		_w254_,
		_w1744_,
		_w1745_,
		_w1753_,
		_w1754_
	);
	LUT4 #(
		.INIT('heeec)
	) name1537 (
		\state_reg[0]/NET0131 ,
		_w1741_,
		_w1742_,
		_w1754_,
		_w1755_
	);
	LUT4 #(
		.INIT('hd11d)
	) name1538 (
		\reg0_reg[22]/NET0131 ,
		_w917_,
		_w1688_,
		_w1690_,
		_w1756_
	);
	LUT2 #(
		.INIT('h2)
	) name1539 (
		_w518_,
		_w1756_,
		_w1757_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1540 (
		\reg0_reg[22]/NET0131 ,
		_w587_,
		_w917_,
		_w1693_,
		_w1758_
	);
	LUT2 #(
		.INIT('h8)
	) name1541 (
		_w525_,
		_w652_,
		_w1759_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1542 (
		_w917_,
		_w1698_,
		_w1701_,
		_w1759_,
		_w1760_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1543 (
		\reg0_reg[22]/NET0131 ,
		_w923_,
		_w924_,
		_w926_,
		_w1761_
	);
	LUT3 #(
		.INIT('h01)
	) name1544 (
		_w1758_,
		_w1760_,
		_w1761_,
		_w1762_
	);
	LUT2 #(
		.INIT('h8)
	) name1545 (
		\reg0_reg[22]/NET0131 ,
		_w252_,
		_w1763_
	);
	LUT4 #(
		.INIT('h0075)
	) name1546 (
		_w254_,
		_w1757_,
		_w1762_,
		_w1763_,
		_w1764_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1547 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[22]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1765_
	);
	LUT3 #(
		.INIT('hf2)
	) name1548 (
		\state_reg[0]/NET0131 ,
		_w1764_,
		_w1765_,
		_w1766_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1549 (
		\reg0_reg[26]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1767_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1550 (
		\reg0_reg[26]/NET0131 ,
		_w917_,
		_w1426_,
		_w1436_,
		_w1768_
	);
	LUT4 #(
		.INIT('h7020)
	) name1551 (
		_w266_,
		_w640_,
		_w917_,
		_w1438_,
		_w1769_
	);
	LUT3 #(
		.INIT('ha8)
	) name1552 (
		_w404_,
		_w1767_,
		_w1769_,
		_w1770_
	);
	LUT4 #(
		.INIT('h4e5d)
	) name1553 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w1771_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1554 (
		_w256_,
		_w258_,
		_w261_,
		_w1771_,
		_w1772_
	);
	LUT3 #(
		.INIT('ha2)
	) name1555 (
		\reg0_reg[26]/NET0131 ,
		_w924_,
		_w1772_,
		_w1773_
	);
	LUT4 #(
		.INIT('h0075)
	) name1556 (
		_w917_,
		_w1555_,
		_w1557_,
		_w1773_,
		_w1774_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1557 (
		_w587_,
		_w1768_,
		_w1770_,
		_w1774_,
		_w1775_
	);
	LUT2 #(
		.INIT('h8)
	) name1558 (
		\reg0_reg[26]/NET0131 ,
		_w252_,
		_w1776_
	);
	LUT4 #(
		.INIT('haa08)
	) name1559 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1775_,
		_w1776_,
		_w1777_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1560 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[26]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1778_
	);
	LUT2 #(
		.INIT('he)
	) name1561 (
		_w1777_,
		_w1778_,
		_w1779_
	);
	LUT2 #(
		.INIT('h8)
	) name1562 (
		_w601_,
		_w1714_,
		_w1780_
	);
	LUT2 #(
		.INIT('h8)
	) name1563 (
		_w917_,
		_w1410_,
		_w1781_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1564 (
		\reg0_reg[30]/NET0131 ,
		_w917_,
		_w924_,
		_w1410_,
		_w1782_
	);
	LUT4 #(
		.INIT('hffd0)
	) name1565 (
		_w1719_,
		_w1780_,
		_w1781_,
		_w1782_,
		_w1783_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1566 (
		\reg0_reg[31]/NET0131 ,
		_w917_,
		_w924_,
		_w1410_,
		_w1784_
	);
	LUT4 #(
		.INIT('hffb0)
	) name1567 (
		_w1416_,
		_w1422_,
		_w1781_,
		_w1784_,
		_w1785_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1568 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[7]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1786_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		\reg0_reg[7]/NET0131 ,
		_w252_,
		_w1787_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1570 (
		\reg0_reg[7]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1788_
	);
	LUT4 #(
		.INIT('hc808)
	) name1571 (
		\reg0_reg[7]/NET0131 ,
		_w404_,
		_w917_,
		_w1371_,
		_w1789_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1572 (
		\reg0_reg[7]/NET0131 ,
		_w518_,
		_w917_,
		_w1374_,
		_w1790_
	);
	LUT4 #(
		.INIT('h20d0)
	) name1573 (
		_w562_,
		_w837_,
		_w917_,
		_w1373_,
		_w1791_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1574 (
		\reg0_reg[7]/NET0131 ,
		_w923_,
		_w924_,
		_w1154_,
		_w1792_
	);
	LUT3 #(
		.INIT('h0d)
	) name1575 (
		_w917_,
		_w1748_,
		_w1792_,
		_w1793_
	);
	LUT4 #(
		.INIT('h5700)
	) name1576 (
		_w587_,
		_w1788_,
		_w1791_,
		_w1793_,
		_w1794_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1577 (
		_w254_,
		_w1789_,
		_w1790_,
		_w1794_,
		_w1795_
	);
	LUT4 #(
		.INIT('heeec)
	) name1578 (
		\state_reg[0]/NET0131 ,
		_w1786_,
		_w1787_,
		_w1795_,
		_w1796_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1579 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[8]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1797_
	);
	LUT2 #(
		.INIT('h8)
	) name1580 (
		\reg0_reg[8]/NET0131 ,
		_w252_,
		_w1798_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1581 (
		\reg0_reg[8]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1799_
	);
	LUT3 #(
		.INIT('h2a)
	) name1582 (
		_w266_,
		_w323_,
		_w325_,
		_w1800_
	);
	LUT3 #(
		.INIT('h8c)
	) name1583 (
		_w331_,
		_w335_,
		_w1369_,
		_w1801_
	);
	LUT2 #(
		.INIT('h1)
	) name1584 (
		_w266_,
		_w339_,
		_w1802_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1585 (
		_w917_,
		_w1800_,
		_w1801_,
		_w1802_,
		_w1803_
	);
	LUT3 #(
		.INIT('ha8)
	) name1586 (
		_w404_,
		_w1799_,
		_w1803_,
		_w1804_
	);
	LUT3 #(
		.INIT('h87)
	) name1587 (
		_w328_,
		_w330_,
		_w470_,
		_w1805_
	);
	LUT4 #(
		.INIT('h8f70)
	) name1588 (
		_w756_,
		_w760_,
		_w763_,
		_w1805_,
		_w1806_
	);
	LUT4 #(
		.INIT('hc808)
	) name1589 (
		\reg0_reg[8]/NET0131 ,
		_w587_,
		_w917_,
		_w1806_,
		_w1807_
	);
	LUT4 #(
		.INIT('h8f70)
	) name1590 (
		_w696_,
		_w700_,
		_w703_,
		_w1805_,
		_w1808_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1591 (
		\reg0_reg[8]/NET0131 ,
		_w518_,
		_w917_,
		_w1808_,
		_w1809_
	);
	LUT4 #(
		.INIT('h6c00)
	) name1592 (
		_w467_,
		_w470_,
		_w592_,
		_w917_,
		_w1810_
	);
	LUT3 #(
		.INIT('h8a)
	) name1593 (
		\reg0_reg[8]/NET0131 ,
		_w923_,
		_w924_,
		_w1811_
	);
	LUT2 #(
		.INIT('h4)
	) name1594 (
		_w470_,
		_w525_,
		_w1812_
	);
	LUT2 #(
		.INIT('h8)
	) name1595 (
		_w917_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h1)
	) name1596 (
		_w1811_,
		_w1813_,
		_w1814_
	);
	LUT4 #(
		.INIT('h5700)
	) name1597 (
		_w601_,
		_w1799_,
		_w1810_,
		_w1814_,
		_w1815_
	);
	LUT3 #(
		.INIT('h10)
	) name1598 (
		_w1809_,
		_w1807_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h1311)
	) name1599 (
		_w254_,
		_w1798_,
		_w1804_,
		_w1816_,
		_w1817_
	);
	LUT3 #(
		.INIT('hce)
	) name1600 (
		\state_reg[0]/NET0131 ,
		_w1797_,
		_w1817_,
		_w1818_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1601 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[11]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1602 (
		\reg1_reg[11]/NET0131 ,
		_w252_,
		_w1820_
	);
	LUT4 #(
		.INIT('haa02)
	) name1603 (
		\reg1_reg[11]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1821_
	);
	LUT4 #(
		.INIT('hb040)
	) name1604 (
		_w865_,
		_w866_,
		_w946_,
		_w1024_,
		_w1822_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1605 (
		_w418_,
		_w946_,
		_w1026_,
		_w1027_,
		_w1823_
	);
	LUT3 #(
		.INIT('ha2)
	) name1606 (
		\reg1_reg[11]/NET0131 ,
		_w924_,
		_w959_,
		_w1824_
	);
	LUT2 #(
		.INIT('h4)
	) name1607 (
		_w418_,
		_w525_,
		_w1825_
	);
	LUT2 #(
		.INIT('h8)
	) name1608 (
		_w946_,
		_w1825_,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name1609 (
		_w1824_,
		_w1826_,
		_w1827_
	);
	LUT4 #(
		.INIT('h5700)
	) name1610 (
		_w601_,
		_w1821_,
		_w1823_,
		_w1827_,
		_w1828_
	);
	LUT4 #(
		.INIT('h5700)
	) name1611 (
		_w518_,
		_w1821_,
		_w1822_,
		_w1828_,
		_w1829_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1612 (
		\reg1_reg[11]/NET0131 ,
		_w946_,
		_w1034_,
		_w1035_,
		_w1830_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1613 (
		\reg1_reg[11]/NET0131 ,
		_w840_,
		_w946_,
		_w1024_,
		_w1831_
	);
	LUT4 #(
		.INIT('hf531)
	) name1614 (
		_w404_,
		_w587_,
		_w1830_,
		_w1831_,
		_w1832_
	);
	LUT4 #(
		.INIT('h3111)
	) name1615 (
		_w254_,
		_w1820_,
		_w1829_,
		_w1832_,
		_w1833_
	);
	LUT3 #(
		.INIT('hce)
	) name1616 (
		\state_reg[0]/NET0131 ,
		_w1819_,
		_w1833_,
		_w1834_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1617 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[14]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1835_
	);
	LUT2 #(
		.INIT('h8)
	) name1618 (
		\reg1_reg[14]/NET0131 ,
		_w252_,
		_w1836_
	);
	LUT4 #(
		.INIT('hc808)
	) name1619 (
		\reg1_reg[14]/NET0131 ,
		_w404_,
		_w946_,
		_w1317_,
		_w1837_
	);
	LUT4 #(
		.INIT('hc808)
	) name1620 (
		\reg1_reg[14]/NET0131 ,
		_w587_,
		_w946_,
		_w1325_,
		_w1838_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1621 (
		\reg1_reg[14]/NET0131 ,
		_w518_,
		_w946_,
		_w1332_,
		_w1839_
	);
	LUT3 #(
		.INIT('ha2)
	) name1622 (
		\reg1_reg[14]/NET0131 ,
		_w924_,
		_w949_,
		_w1840_
	);
	LUT2 #(
		.INIT('h4)
	) name1623 (
		_w439_,
		_w525_,
		_w1841_
	);
	LUT4 #(
		.INIT('h009f)
	) name1624 (
		_w439_,
		_w596_,
		_w601_,
		_w1841_,
		_w1842_
	);
	LUT3 #(
		.INIT('h31)
	) name1625 (
		_w946_,
		_w1840_,
		_w1842_,
		_w1843_
	);
	LUT4 #(
		.INIT('h0100)
	) name1626 (
		_w1837_,
		_w1839_,
		_w1838_,
		_w1843_,
		_w1844_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1627 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1836_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('he)
	) name1628 (
		_w1835_,
		_w1845_,
		_w1846_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1629 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[16]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1847_
	);
	LUT2 #(
		.INIT('h8)
	) name1630 (
		\reg1_reg[16]/NET0131 ,
		_w252_,
		_w1848_
	);
	LUT4 #(
		.INIT('haa02)
	) name1631 (
		\reg1_reg[16]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1849_
	);
	LUT4 #(
		.INIT('hd11d)
	) name1632 (
		\reg1_reg[16]/NET0131 ,
		_w946_,
		_w1347_,
		_w1348_,
		_w1850_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		_w587_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1634 (
		\reg1_reg[16]/NET0131 ,
		_w946_,
		_w1347_,
		_w1351_,
		_w1852_
	);
	LUT4 #(
		.INIT('h7020)
	) name1635 (
		_w266_,
		_w378_,
		_w946_,
		_w1353_,
		_w1853_
	);
	LUT3 #(
		.INIT('ha8)
	) name1636 (
		_w404_,
		_w1849_,
		_w1853_,
		_w1854_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1637 (
		_w601_,
		_w946_,
		_w1356_,
		_w1734_,
		_w1855_
	);
	LUT3 #(
		.INIT('ha2)
	) name1638 (
		\reg1_reg[16]/NET0131 ,
		_w924_,
		_w949_,
		_w1856_
	);
	LUT2 #(
		.INIT('h1)
	) name1639 (
		_w1855_,
		_w1856_,
		_w1857_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1640 (
		_w518_,
		_w1852_,
		_w1854_,
		_w1857_,
		_w1858_
	);
	LUT4 #(
		.INIT('h1311)
	) name1641 (
		_w254_,
		_w1848_,
		_w1851_,
		_w1858_,
		_w1859_
	);
	LUT3 #(
		.INIT('hce)
	) name1642 (
		\state_reg[0]/NET0131 ,
		_w1847_,
		_w1859_,
		_w1860_
	);
	LUT4 #(
		.INIT('hd11d)
	) name1643 (
		\reg1_reg[22]/NET0131 ,
		_w946_,
		_w1688_,
		_w1690_,
		_w1861_
	);
	LUT2 #(
		.INIT('h2)
	) name1644 (
		_w518_,
		_w1861_,
		_w1862_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1645 (
		\reg1_reg[22]/NET0131 ,
		_w587_,
		_w946_,
		_w1693_,
		_w1863_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1646 (
		_w946_,
		_w1698_,
		_w1701_,
		_w1759_,
		_w1864_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1647 (
		\reg1_reg[22]/NET0131 ,
		_w924_,
		_w949_,
		_w950_,
		_w1865_
	);
	LUT3 #(
		.INIT('h01)
	) name1648 (
		_w1863_,
		_w1864_,
		_w1865_,
		_w1866_
	);
	LUT2 #(
		.INIT('h8)
	) name1649 (
		\reg1_reg[22]/NET0131 ,
		_w252_,
		_w1867_
	);
	LUT4 #(
		.INIT('h0075)
	) name1650 (
		_w254_,
		_w1862_,
		_w1866_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1651 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[22]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1869_
	);
	LUT3 #(
		.INIT('hf2)
	) name1652 (
		\state_reg[0]/NET0131 ,
		_w1868_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h8)
	) name1653 (
		_w946_,
		_w1410_,
		_w1871_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1654 (
		\reg1_reg[31]/NET0131 ,
		_w924_,
		_w946_,
		_w1410_,
		_w1872_
	);
	LUT4 #(
		.INIT('hffb0)
	) name1655 (
		_w1416_,
		_w1422_,
		_w1871_,
		_w1872_,
		_w1873_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1656 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[30]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1874_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1657 (
		_w256_,
		_w258_,
		_w261_,
		_w924_,
		_w1875_
	);
	LUT2 #(
		.INIT('h2)
	) name1658 (
		\reg1_reg[30]/NET0131 ,
		_w1875_,
		_w1876_
	);
	LUT4 #(
		.INIT('h005d)
	) name1659 (
		_w946_,
		_w1719_,
		_w1780_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		\reg1_reg[30]/NET0131 ,
		_w252_,
		_w1878_
	);
	LUT4 #(
		.INIT('haa08)
	) name1661 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1877_,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('he)
	) name1662 (
		_w1874_,
		_w1879_,
		_w1880_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1663 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[7]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1881_
	);
	LUT2 #(
		.INIT('h8)
	) name1664 (
		\reg1_reg[7]/NET0131 ,
		_w252_,
		_w1882_
	);
	LUT4 #(
		.INIT('haa02)
	) name1665 (
		\reg1_reg[7]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1883_
	);
	LUT4 #(
		.INIT('hc808)
	) name1666 (
		\reg1_reg[7]/NET0131 ,
		_w404_,
		_w946_,
		_w1371_,
		_w1884_
	);
	LUT4 #(
		.INIT('h20d0)
	) name1667 (
		_w562_,
		_w837_,
		_w946_,
		_w1373_,
		_w1885_
	);
	LUT3 #(
		.INIT('ha8)
	) name1668 (
		_w587_,
		_w1883_,
		_w1885_,
		_w1886_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1669 (
		\reg1_reg[7]/NET0131 ,
		_w518_,
		_w946_,
		_w1374_,
		_w1887_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1670 (
		\reg1_reg[7]/NET0131 ,
		_w924_,
		_w959_,
		_w960_,
		_w1888_
	);
	LUT3 #(
		.INIT('h0d)
	) name1671 (
		_w946_,
		_w1748_,
		_w1888_,
		_w1889_
	);
	LUT4 #(
		.INIT('h0100)
	) name1672 (
		_w1884_,
		_w1887_,
		_w1886_,
		_w1889_,
		_w1890_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1673 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1882_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('he)
	) name1674 (
		_w1881_,
		_w1891_,
		_w1892_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1675 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[11]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1893_
	);
	LUT2 #(
		.INIT('h8)
	) name1676 (
		\reg0_reg[11]/NET0131 ,
		_w252_,
		_w1894_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1677 (
		\reg0_reg[11]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1895_
	);
	LUT4 #(
		.INIT('hb040)
	) name1678 (
		_w865_,
		_w866_,
		_w917_,
		_w1024_,
		_w1896_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1679 (
		_w418_,
		_w917_,
		_w1026_,
		_w1027_,
		_w1897_
	);
	LUT3 #(
		.INIT('h8a)
	) name1680 (
		\reg0_reg[11]/NET0131 ,
		_w923_,
		_w924_,
		_w1898_
	);
	LUT2 #(
		.INIT('h8)
	) name1681 (
		_w917_,
		_w1825_,
		_w1899_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		_w1898_,
		_w1899_,
		_w1900_
	);
	LUT4 #(
		.INIT('h5700)
	) name1683 (
		_w601_,
		_w1895_,
		_w1897_,
		_w1900_,
		_w1901_
	);
	LUT4 #(
		.INIT('h5700)
	) name1684 (
		_w518_,
		_w1895_,
		_w1896_,
		_w1901_,
		_w1902_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1685 (
		\reg0_reg[11]/NET0131 ,
		_w917_,
		_w1034_,
		_w1035_,
		_w1903_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1686 (
		\reg0_reg[11]/NET0131 ,
		_w840_,
		_w917_,
		_w1024_,
		_w1904_
	);
	LUT4 #(
		.INIT('hf531)
	) name1687 (
		_w404_,
		_w587_,
		_w1903_,
		_w1904_,
		_w1905_
	);
	LUT4 #(
		.INIT('h3111)
	) name1688 (
		_w254_,
		_w1894_,
		_w1902_,
		_w1905_,
		_w1906_
	);
	LUT3 #(
		.INIT('hce)
	) name1689 (
		\state_reg[0]/NET0131 ,
		_w1893_,
		_w1906_,
		_w1907_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1690 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[14]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1908_
	);
	LUT2 #(
		.INIT('h8)
	) name1691 (
		\reg2_reg[14]/NET0131 ,
		_w252_,
		_w1909_
	);
	LUT4 #(
		.INIT('hc808)
	) name1692 (
		\reg2_reg[14]/NET0131 ,
		_w404_,
		_w970_,
		_w1317_,
		_w1910_
	);
	LUT4 #(
		.INIT('hc808)
	) name1693 (
		\reg2_reg[14]/NET0131 ,
		_w587_,
		_w970_,
		_w1325_,
		_w1911_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1694 (
		\reg2_reg[14]/NET0131 ,
		_w518_,
		_w970_,
		_w1332_,
		_w1912_
	);
	LUT2 #(
		.INIT('h8)
	) name1695 (
		_w520_,
		_w363_,
		_w1913_
	);
	LUT4 #(
		.INIT('h0057)
	) name1696 (
		\reg2_reg[14]/NET0131 ,
		_w524_,
		_w1237_,
		_w1913_,
		_w1914_
	);
	LUT3 #(
		.INIT('hd0)
	) name1697 (
		_w970_,
		_w1842_,
		_w1914_,
		_w1915_
	);
	LUT4 #(
		.INIT('h0100)
	) name1698 (
		_w1910_,
		_w1912_,
		_w1911_,
		_w1915_,
		_w1916_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1699 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1909_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('he)
	) name1700 (
		_w1908_,
		_w1917_,
		_w1918_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1701 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[16]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1919_
	);
	LUT2 #(
		.INIT('h8)
	) name1702 (
		\reg2_reg[16]/NET0131 ,
		_w252_,
		_w1920_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1703 (
		\reg2_reg[16]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1921_
	);
	LUT4 #(
		.INIT('hd11d)
	) name1704 (
		\reg2_reg[16]/NET0131 ,
		_w970_,
		_w1347_,
		_w1348_,
		_w1922_
	);
	LUT2 #(
		.INIT('h2)
	) name1705 (
		_w587_,
		_w1922_,
		_w1923_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1706 (
		\reg2_reg[16]/NET0131 ,
		_w970_,
		_w1347_,
		_w1351_,
		_w1924_
	);
	LUT4 #(
		.INIT('h7020)
	) name1707 (
		_w266_,
		_w378_,
		_w970_,
		_w1353_,
		_w1925_
	);
	LUT3 #(
		.INIT('ha8)
	) name1708 (
		_w404_,
		_w1921_,
		_w1925_,
		_w1926_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1709 (
		_w601_,
		_w970_,
		_w1356_,
		_w1734_,
		_w1927_
	);
	LUT2 #(
		.INIT('h8)
	) name1710 (
		_w520_,
		_w358_,
		_w1928_
	);
	LUT4 #(
		.INIT('h0057)
	) name1711 (
		\reg2_reg[16]/NET0131 ,
		_w524_,
		_w1237_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h4)
	) name1712 (
		_w1927_,
		_w1929_,
		_w1930_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1713 (
		_w518_,
		_w1924_,
		_w1926_,
		_w1930_,
		_w1931_
	);
	LUT4 #(
		.INIT('h1311)
	) name1714 (
		_w254_,
		_w1920_,
		_w1923_,
		_w1931_,
		_w1932_
	);
	LUT3 #(
		.INIT('hce)
	) name1715 (
		\state_reg[0]/NET0131 ,
		_w1919_,
		_w1932_,
		_w1933_
	);
	LUT4 #(
		.INIT('hd11d)
	) name1716 (
		\reg2_reg[22]/NET0131 ,
		_w970_,
		_w1688_,
		_w1690_,
		_w1934_
	);
	LUT2 #(
		.INIT('h2)
	) name1717 (
		_w518_,
		_w1934_,
		_w1935_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1718 (
		\reg2_reg[22]/NET0131 ,
		_w587_,
		_w970_,
		_w1693_,
		_w1936_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1719 (
		_w970_,
		_w1698_,
		_w1701_,
		_w1759_,
		_w1937_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		_w520_,
		_w654_,
		_w1938_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1721 (
		\reg2_reg[22]/NET0131 ,
		_w524_,
		_w990_,
		_w1237_,
		_w1939_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		_w1938_,
		_w1939_,
		_w1940_
	);
	LUT3 #(
		.INIT('h10)
	) name1723 (
		_w1936_,
		_w1937_,
		_w1940_,
		_w1941_
	);
	LUT2 #(
		.INIT('h8)
	) name1724 (
		\reg2_reg[22]/NET0131 ,
		_w252_,
		_w1942_
	);
	LUT4 #(
		.INIT('h0075)
	) name1725 (
		_w254_,
		_w1935_,
		_w1941_,
		_w1942_,
		_w1943_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1726 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[22]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1944_
	);
	LUT3 #(
		.INIT('hf2)
	) name1727 (
		\state_reg[0]/NET0131 ,
		_w1943_,
		_w1944_,
		_w1945_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1728 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[14]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1946_
	);
	LUT2 #(
		.INIT('h8)
	) name1729 (
		\reg0_reg[14]/NET0131 ,
		_w252_,
		_w1947_
	);
	LUT4 #(
		.INIT('hc808)
	) name1730 (
		\reg0_reg[14]/NET0131 ,
		_w404_,
		_w917_,
		_w1317_,
		_w1948_
	);
	LUT4 #(
		.INIT('hc808)
	) name1731 (
		\reg0_reg[14]/NET0131 ,
		_w587_,
		_w917_,
		_w1325_,
		_w1949_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1732 (
		\reg0_reg[14]/NET0131 ,
		_w518_,
		_w917_,
		_w1332_,
		_w1950_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1733 (
		\reg0_reg[14]/NET0131 ,
		_w923_,
		_w924_,
		_w1154_,
		_w1951_
	);
	LUT3 #(
		.INIT('h0d)
	) name1734 (
		_w917_,
		_w1842_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h0100)
	) name1735 (
		_w1948_,
		_w1950_,
		_w1949_,
		_w1952_,
		_w1953_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1736 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w1947_,
		_w1953_,
		_w1954_
	);
	LUT2 #(
		.INIT('he)
	) name1737 (
		_w1946_,
		_w1954_,
		_w1955_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1738 (
		\IR_reg[23]/NET0131 ,
		\reg3_reg[1]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1956_
	);
	LUT2 #(
		.INIT('h8)
	) name1739 (
		\reg3_reg[1]/NET0131 ,
		_w252_,
		_w1957_
	);
	LUT2 #(
		.INIT('h6)
	) name1740 (
		_w491_,
		_w493_,
		_w1958_
	);
	LUT3 #(
		.INIT('h60)
	) name1741 (
		_w491_,
		_w493_,
		_w601_,
		_w1959_
	);
	LUT4 #(
		.INIT('h5556)
	) name1742 (
		_w276_,
		_w280_,
		_w284_,
		_w299_,
		_w1960_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1743 (
		_w266_,
		_w282_,
		_w283_,
		_w404_,
		_w1961_
	);
	LUT3 #(
		.INIT('he0)
	) name1744 (
		_w266_,
		_w1960_,
		_w1961_,
		_w1962_
	);
	LUT3 #(
		.INIT('h87)
	) name1745 (
		_w278_,
		_w279_,
		_w491_,
		_w1963_
	);
	LUT3 #(
		.INIT('h84)
	) name1746 (
		_w494_,
		_w518_,
		_w1963_,
		_w1964_
	);
	LUT3 #(
		.INIT('h84)
	) name1747 (
		_w570_,
		_w587_,
		_w1963_,
		_w1965_
	);
	LUT2 #(
		.INIT('h1)
	) name1748 (
		_w1964_,
		_w1965_,
		_w1966_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1749 (
		_w262_,
		_w1959_,
		_w1962_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('h001f)
	) name1750 (
		_w256_,
		_w258_,
		_w261_,
		_w522_,
		_w1968_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1751 (
		\reg3_reg[1]/NET0131 ,
		_w524_,
		_w526_,
		_w1968_,
		_w1969_
	);
	LUT3 #(
		.INIT('h04)
	) name1752 (
		_w521_,
		_w522_,
		_w491_,
		_w1970_
	);
	LUT2 #(
		.INIT('h1)
	) name1753 (
		_w1969_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('h1311)
	) name1754 (
		_w254_,
		_w1957_,
		_w1967_,
		_w1971_,
		_w1972_
	);
	LUT3 #(
		.INIT('hce)
	) name1755 (
		\state_reg[0]/NET0131 ,
		_w1956_,
		_w1972_,
		_w1973_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1756 (
		\IR_reg[23]/NET0131 ,
		\reg3_reg[2]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w1974_
	);
	LUT2 #(
		.INIT('h8)
	) name1757 (
		\reg3_reg[2]/NET0131 ,
		_w252_,
		_w1975_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1758 (
		\reg3_reg[2]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w1976_
	);
	LUT3 #(
		.INIT('h80)
	) name1759 (
		_w266_,
		_w278_,
		_w279_,
		_w1977_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1760 (
		_w266_,
		_w301_,
		_w304_,
		_w1977_,
		_w1978_
	);
	LUT4 #(
		.INIT('he020)
	) name1761 (
		\reg3_reg[2]/NET0131 ,
		_w262_,
		_w404_,
		_w1978_,
		_w1979_
	);
	LUT3 #(
		.INIT('h87)
	) name1762 (
		_w273_,
		_w275_,
		_w497_,
		_w1980_
	);
	LUT4 #(
		.INIT('hf100)
	) name1763 (
		_w492_,
		_w494_,
		_w495_,
		_w1980_,
		_w1981_
	);
	LUT4 #(
		.INIT('h000e)
	) name1764 (
		_w492_,
		_w494_,
		_w495_,
		_w1980_,
		_w1982_
	);
	LUT3 #(
		.INIT('h02)
	) name1765 (
		_w518_,
		_w1982_,
		_w1981_,
		_w1983_
	);
	LUT4 #(
		.INIT('h7800)
	) name1766 (
		_w491_,
		_w493_,
		_w497_,
		_w601_,
		_w1984_
	);
	LUT4 #(
		.INIT('h0b07)
	) name1767 (
		_w571_,
		_w587_,
		_w1984_,
		_w1980_,
		_w1985_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1768 (
		_w256_,
		_w258_,
		_w261_,
		_w497_,
		_w1986_
	);
	LUT3 #(
		.INIT('ha8)
	) name1769 (
		_w525_,
		_w1976_,
		_w1986_,
		_w1987_
	);
	LUT2 #(
		.INIT('h2)
	) name1770 (
		_w520_,
		_w497_,
		_w1988_
	);
	LUT3 #(
		.INIT('h01)
	) name1771 (
		_w398_,
		_w399_,
		_w403_,
		_w1989_
	);
	LUT4 #(
		.INIT('h6664)
	) name1772 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w1990_
	);
	LUT4 #(
		.INIT('h001f)
	) name1773 (
		_w256_,
		_w258_,
		_w261_,
		_w1990_,
		_w1991_
	);
	LUT4 #(
		.INIT('h0507)
	) name1774 (
		\reg3_reg[2]/NET0131 ,
		_w524_,
		_w1988_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h4)
	) name1775 (
		_w1987_,
		_w1992_,
		_w1993_
	);
	LUT4 #(
		.INIT('h7500)
	) name1776 (
		_w262_,
		_w1983_,
		_w1985_,
		_w1993_,
		_w1994_
	);
	LUT4 #(
		.INIT('h1311)
	) name1777 (
		_w254_,
		_w1975_,
		_w1979_,
		_w1994_,
		_w1995_
	);
	LUT3 #(
		.INIT('hce)
	) name1778 (
		\state_reg[0]/NET0131 ,
		_w1974_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h8)
	) name1779 (
		_w252_,
		_w313_,
		_w1997_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1780 (
		_w256_,
		_w258_,
		_w261_,
		_w313_,
		_w1998_
	);
	LUT4 #(
		.INIT('h807f)
	) name1781 (
		_w301_,
		_w311_,
		_w322_,
		_w326_,
		_w1999_
	);
	LUT4 #(
		.INIT('h2a08)
	) name1782 (
		_w262_,
		_w266_,
		_w320_,
		_w1999_,
		_w2000_
	);
	LUT3 #(
		.INIT('ha8)
	) name1783 (
		_w404_,
		_w1998_,
		_w2000_,
		_w2001_
	);
	LUT3 #(
		.INIT('h78)
	) name1784 (
		_w312_,
		_w314_,
		_w475_,
		_w2002_
	);
	LUT4 #(
		.INIT('h208a)
	) name1785 (
		_w262_,
		_w760_,
		_w761_,
		_w2002_,
		_w2003_
	);
	LUT3 #(
		.INIT('ha8)
	) name1786 (
		_w587_,
		_w1998_,
		_w2003_,
		_w2004_
	);
	LUT4 #(
		.INIT('ha802)
	) name1787 (
		_w262_,
		_w700_,
		_w701_,
		_w2002_,
		_w2005_
	);
	LUT4 #(
		.INIT('h2800)
	) name1788 (
		_w262_,
		_w475_,
		_w591_,
		_w601_,
		_w2006_
	);
	LUT3 #(
		.INIT('ha8)
	) name1789 (
		_w313_,
		_w524_,
		_w906_,
		_w2007_
	);
	LUT3 #(
		.INIT('h04)
	) name1790 (
		_w521_,
		_w522_,
		_w475_,
		_w2008_
	);
	LUT2 #(
		.INIT('h1)
	) name1791 (
		_w2007_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h4)
	) name1792 (
		_w2006_,
		_w2009_,
		_w2010_
	);
	LUT4 #(
		.INIT('h5700)
	) name1793 (
		_w518_,
		_w1998_,
		_w2005_,
		_w2010_,
		_w2011_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1794 (
		_w254_,
		_w2001_,
		_w2004_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h2)
	) name1795 (
		\reg3_reg[6]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2013_
	);
	LUT4 #(
		.INIT('h4800)
	) name1796 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w313_,
		_w2014_
	);
	LUT2 #(
		.INIT('h1)
	) name1797 (
		_w2013_,
		_w2014_,
		_w2015_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1798 (
		\state_reg[0]/NET0131 ,
		_w1997_,
		_w2012_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h8)
	) name1799 (
		_w252_,
		_w329_,
		_w2017_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1800 (
		_w256_,
		_w258_,
		_w261_,
		_w329_,
		_w2018_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1801 (
		_w262_,
		_w1800_,
		_w1801_,
		_w1802_,
		_w2019_
	);
	LUT3 #(
		.INIT('ha8)
	) name1802 (
		_w404_,
		_w2018_,
		_w2019_,
		_w2020_
	);
	LUT4 #(
		.INIT('he040)
	) name1803 (
		_w262_,
		_w329_,
		_w587_,
		_w1806_,
		_w2021_
	);
	LUT4 #(
		.INIT('h40e0)
	) name1804 (
		_w262_,
		_w329_,
		_w518_,
		_w1808_,
		_w2022_
	);
	LUT4 #(
		.INIT('h28a0)
	) name1805 (
		_w262_,
		_w467_,
		_w470_,
		_w592_,
		_w2023_
	);
	LUT3 #(
		.INIT('h04)
	) name1806 (
		_w521_,
		_w522_,
		_w470_,
		_w2024_
	);
	LUT3 #(
		.INIT('ha8)
	) name1807 (
		_w329_,
		_w524_,
		_w526_,
		_w2025_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w2024_,
		_w2025_,
		_w2026_
	);
	LUT4 #(
		.INIT('h5700)
	) name1809 (
		_w601_,
		_w2018_,
		_w2023_,
		_w2026_,
		_w2027_
	);
	LUT3 #(
		.INIT('h10)
	) name1810 (
		_w2022_,
		_w2021_,
		_w2027_,
		_w2028_
	);
	LUT4 #(
		.INIT('h1311)
	) name1811 (
		_w254_,
		_w2017_,
		_w2020_,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h2)
	) name1812 (
		\reg3_reg[8]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2030_
	);
	LUT4 #(
		.INIT('h4800)
	) name1813 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w329_,
		_w2031_
	);
	LUT2 #(
		.INIT('h1)
	) name1814 (
		_w2030_,
		_w2031_,
		_w2032_
	);
	LUT3 #(
		.INIT('h2f)
	) name1815 (
		\state_reg[0]/NET0131 ,
		_w2029_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h8)
	) name1816 (
		_w252_,
		_w333_,
		_w2034_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1817 (
		_w256_,
		_w258_,
		_w261_,
		_w333_,
		_w2035_
	);
	LUT3 #(
		.INIT('h80)
	) name1818 (
		_w266_,
		_w328_,
		_w330_,
		_w2036_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1819 (
		_w266_,
		_w339_,
		_w353_,
		_w2036_,
		_w2037_
	);
	LUT4 #(
		.INIT('he040)
	) name1820 (
		_w262_,
		_w333_,
		_w404_,
		_w2037_,
		_w2038_
	);
	LUT3 #(
		.INIT('h87)
	) name1821 (
		_w332_,
		_w334_,
		_w431_,
		_w2039_
	);
	LUT4 #(
		.INIT('hd52a)
	) name1822 (
		_w486_,
		_w509_,
		_w512_,
		_w2039_,
		_w2040_
	);
	LUT4 #(
		.INIT('h40e0)
	) name1823 (
		_w262_,
		_w333_,
		_w518_,
		_w2040_,
		_w2041_
	);
	LUT4 #(
		.INIT('ha208)
	) name1824 (
		_w262_,
		_w566_,
		_w584_,
		_w2039_,
		_w2042_
	);
	LUT3 #(
		.INIT('ha8)
	) name1825 (
		_w587_,
		_w2035_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1826 (
		_w431_,
		_w467_,
		_w470_,
		_w592_,
		_w2044_
	);
	LUT4 #(
		.INIT('he040)
	) name1827 (
		_w262_,
		_w333_,
		_w601_,
		_w2044_,
		_w2045_
	);
	LUT3 #(
		.INIT('h04)
	) name1828 (
		_w521_,
		_w522_,
		_w431_,
		_w2046_
	);
	LUT3 #(
		.INIT('ha8)
	) name1829 (
		_w333_,
		_w524_,
		_w526_,
		_w2047_
	);
	LUT2 #(
		.INIT('h1)
	) name1830 (
		_w2046_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h4)
	) name1831 (
		_w2045_,
		_w2048_,
		_w2049_
	);
	LUT4 #(
		.INIT('h0100)
	) name1832 (
		_w2038_,
		_w2043_,
		_w2041_,
		_w2049_,
		_w2050_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1833 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2034_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h2)
	) name1834 (
		\reg3_reg[9]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2052_
	);
	LUT4 #(
		.INIT('h4800)
	) name1835 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w333_,
		_w2053_
	);
	LUT2 #(
		.INIT('h1)
	) name1836 (
		_w2052_,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('hb)
	) name1837 (
		_w2051_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h8)
	) name1838 (
		_w252_,
		_w636_,
		_w2056_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1839 (
		_w256_,
		_w258_,
		_w261_,
		_w636_,
		_w2057_
	);
	LUT4 #(
		.INIT('h082a)
	) name1840 (
		_w262_,
		_w266_,
		_w647_,
		_w1665_,
		_w2058_
	);
	LUT3 #(
		.INIT('ha8)
	) name1841 (
		_w404_,
		_w2057_,
		_w2058_,
		_w2059_
	);
	LUT4 #(
		.INIT('h0a82)
	) name1842 (
		_w262_,
		_w1300_,
		_w1668_,
		_w1675_,
		_w2060_
	);
	LUT3 #(
		.INIT('ha8)
	) name1843 (
		_w587_,
		_w2057_,
		_w2060_,
		_w2061_
	);
	LUT4 #(
		.INIT('h40c8)
	) name1844 (
		_w262_,
		_w518_,
		_w636_,
		_w1671_,
		_w2062_
	);
	LUT4 #(
		.INIT('h007d)
	) name1845 (
		_w262_,
		_w635_,
		_w804_,
		_w2057_,
		_w2063_
	);
	LUT3 #(
		.INIT('h40)
	) name1846 (
		_w521_,
		_w522_,
		_w635_,
		_w2064_
	);
	LUT3 #(
		.INIT('he0)
	) name1847 (
		_w524_,
		_w526_,
		_w636_,
		_w2065_
	);
	LUT2 #(
		.INIT('h1)
	) name1848 (
		_w2064_,
		_w2065_,
		_w2066_
	);
	LUT3 #(
		.INIT('hd0)
	) name1849 (
		_w601_,
		_w2063_,
		_w2066_,
		_w2067_
	);
	LUT4 #(
		.INIT('h0100)
	) name1850 (
		_w2062_,
		_w2059_,
		_w2061_,
		_w2067_,
		_w2068_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1851 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2056_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h2)
	) name1852 (
		\reg3_reg[25]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2070_
	);
	LUT3 #(
		.INIT('h07)
	) name1853 (
		_w606_,
		_w636_,
		_w2070_,
		_w2071_
	);
	LUT2 #(
		.INIT('hb)
	) name1854 (
		_w2069_,
		_w2071_,
		_w2072_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1855 (
		\reg2_reg[3]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2073_
	);
	LUT3 #(
		.INIT('h2a)
	) name1856 (
		_w266_,
		_w273_,
		_w275_,
		_w2074_
	);
	LUT4 #(
		.INIT('h0451)
	) name1857 (
		_w266_,
		_w301_,
		_w304_,
		_w309_,
		_w2075_
	);
	LUT4 #(
		.INIT('h111d)
	) name1858 (
		\reg2_reg[3]/NET0131 ,
		_w970_,
		_w2074_,
		_w2075_,
		_w2076_
	);
	LUT3 #(
		.INIT('h78)
	) name1859 (
		_w302_,
		_w303_,
		_w502_,
		_w2077_
	);
	LUT4 #(
		.INIT('he010)
	) name1860 (
		_w572_,
		_w574_,
		_w970_,
		_w2077_,
		_w2078_
	);
	LUT3 #(
		.INIT('ha8)
	) name1861 (
		_w587_,
		_w2073_,
		_w2078_,
		_w2079_
	);
	LUT4 #(
		.INIT('h10e0)
	) name1862 (
		_w499_,
		_w504_,
		_w970_,
		_w2077_,
		_w2080_
	);
	LUT2 #(
		.INIT('h4)
	) name1863 (
		_w502_,
		_w525_,
		_w2081_
	);
	LUT4 #(
		.INIT('h009f)
	) name1864 (
		_w502_,
		_w589_,
		_w601_,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h4)
	) name1865 (
		\reg3_reg[3]/NET0131 ,
		_w520_,
		_w2083_
	);
	LUT4 #(
		.INIT('h0057)
	) name1866 (
		\reg2_reg[3]/NET0131 ,
		_w524_,
		_w1237_,
		_w2083_,
		_w2084_
	);
	LUT3 #(
		.INIT('hd0)
	) name1867 (
		_w970_,
		_w2082_,
		_w2084_,
		_w2085_
	);
	LUT4 #(
		.INIT('h5700)
	) name1868 (
		_w518_,
		_w2073_,
		_w2080_,
		_w2085_,
		_w2086_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1869 (
		_w404_,
		_w2076_,
		_w2079_,
		_w2086_,
		_w2087_
	);
	LUT2 #(
		.INIT('h8)
	) name1870 (
		\reg2_reg[3]/NET0131 ,
		_w252_,
		_w2088_
	);
	LUT4 #(
		.INIT('haa08)
	) name1871 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2087_,
		_w2088_,
		_w2089_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1872 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[3]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2090_
	);
	LUT2 #(
		.INIT('he)
	) name1873 (
		_w2089_,
		_w2090_,
		_w2091_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1874 (
		\reg0_reg[18]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2092_
	);
	LUT4 #(
		.INIT('h08a2)
	) name1875 (
		_w917_,
		_w1427_,
		_w1429_,
		_w1641_,
		_w2093_
	);
	LUT3 #(
		.INIT('ha8)
	) name1876 (
		_w587_,
		_w2092_,
		_w2093_,
		_w2094_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1877 (
		\reg0_reg[18]/NET0131 ,
		_w917_,
		_w1644_,
		_w1645_,
		_w2095_
	);
	LUT2 #(
		.INIT('h8)
	) name1878 (
		_w525_,
		_w678_,
		_w2096_
	);
	LUT3 #(
		.INIT('h01)
	) name1879 (
		_w1647_,
		_w1648_,
		_w2096_,
		_w2097_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1880 (
		_w917_,
		_w1647_,
		_w1648_,
		_w2096_,
		_w2098_
	);
	LUT3 #(
		.INIT('ha2)
	) name1881 (
		\reg0_reg[18]/NET0131 ,
		_w924_,
		_w1772_,
		_w2099_
	);
	LUT4 #(
		.INIT('h0031)
	) name1882 (
		_w404_,
		_w2098_,
		_w2095_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h8)
	) name1883 (
		\reg0_reg[18]/NET0131 ,
		_w252_,
		_w2101_
	);
	LUT4 #(
		.INIT('h0075)
	) name1884 (
		_w254_,
		_w2094_,
		_w2100_,
		_w2101_,
		_w2102_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1885 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[18]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2103_
	);
	LUT3 #(
		.INIT('hf2)
	) name1886 (
		\state_reg[0]/NET0131 ,
		_w2102_,
		_w2103_,
		_w2104_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1887 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[25]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2105_
	);
	LUT2 #(
		.INIT('h8)
	) name1888 (
		\reg0_reg[25]/NET0131 ,
		_w252_,
		_w2106_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1889 (
		\reg0_reg[25]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2107_
	);
	LUT4 #(
		.INIT('h2070)
	) name1890 (
		_w266_,
		_w647_,
		_w917_,
		_w1665_,
		_w2108_
	);
	LUT3 #(
		.INIT('ha8)
	) name1891 (
		_w404_,
		_w2107_,
		_w2108_,
		_w2109_
	);
	LUT4 #(
		.INIT('h0a82)
	) name1892 (
		_w917_,
		_w1300_,
		_w1668_,
		_w1675_,
		_w2110_
	);
	LUT3 #(
		.INIT('ha8)
	) name1893 (
		_w587_,
		_w2107_,
		_w2110_,
		_w2111_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1894 (
		\reg0_reg[25]/NET0131 ,
		_w518_,
		_w917_,
		_w1671_,
		_w2112_
	);
	LUT4 #(
		.INIT('h3c55)
	) name1895 (
		\reg0_reg[25]/NET0131 ,
		_w635_,
		_w804_,
		_w917_,
		_w2113_
	);
	LUT3 #(
		.INIT('h8a)
	) name1896 (
		\reg0_reg[25]/NET0131 ,
		_w923_,
		_w924_,
		_w2114_
	);
	LUT2 #(
		.INIT('h8)
	) name1897 (
		_w917_,
		_w1680_,
		_w2115_
	);
	LUT2 #(
		.INIT('h1)
	) name1898 (
		_w2114_,
		_w2115_,
		_w2116_
	);
	LUT3 #(
		.INIT('hd0)
	) name1899 (
		_w601_,
		_w2113_,
		_w2116_,
		_w2117_
	);
	LUT4 #(
		.INIT('h0100)
	) name1900 (
		_w2112_,
		_w2109_,
		_w2111_,
		_w2117_,
		_w2118_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1901 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2106_,
		_w2118_,
		_w2119_
	);
	LUT2 #(
		.INIT('he)
	) name1902 (
		_w2105_,
		_w2119_,
		_w2120_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1903 (
		\reg0_reg[3]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2121_
	);
	LUT4 #(
		.INIT('h111d)
	) name1904 (
		\reg0_reg[3]/NET0131 ,
		_w917_,
		_w2074_,
		_w2075_,
		_w2122_
	);
	LUT4 #(
		.INIT('he010)
	) name1905 (
		_w572_,
		_w574_,
		_w917_,
		_w2077_,
		_w2123_
	);
	LUT3 #(
		.INIT('ha8)
	) name1906 (
		_w587_,
		_w2121_,
		_w2123_,
		_w2124_
	);
	LUT4 #(
		.INIT('h10e0)
	) name1907 (
		_w499_,
		_w504_,
		_w518_,
		_w2077_,
		_w2125_
	);
	LUT3 #(
		.INIT('ha2)
	) name1908 (
		\reg0_reg[3]/NET0131 ,
		_w924_,
		_w1772_,
		_w2126_
	);
	LUT4 #(
		.INIT('h005d)
	) name1909 (
		_w917_,
		_w2082_,
		_w2125_,
		_w2126_,
		_w2127_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1910 (
		_w404_,
		_w2122_,
		_w2124_,
		_w2127_,
		_w2128_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		\reg0_reg[3]/NET0131 ,
		_w252_,
		_w2129_
	);
	LUT4 #(
		.INIT('haa08)
	) name1912 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2128_,
		_w2129_,
		_w2130_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1913 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[3]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2131_
	);
	LUT2 #(
		.INIT('he)
	) name1914 (
		_w2130_,
		_w2131_,
		_w2132_
	);
	LUT4 #(
		.INIT('h5014)
	) name1915 (
		_w266_,
		_w339_,
		_w348_,
		_w353_,
		_w2133_
	);
	LUT3 #(
		.INIT('h80)
	) name1916 (
		_w266_,
		_w332_,
		_w334_,
		_w2134_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1917 (
		\reg1_reg[10]/NET0131 ,
		_w946_,
		_w2133_,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h2)
	) name1918 (
		_w404_,
		_w2135_,
		_w2136_
	);
	LUT3 #(
		.INIT('h78)
	) name1919 (
		_w350_,
		_w352_,
		_w427_,
		_w2137_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1920 (
		\reg1_reg[10]/NET0131 ,
		_w946_,
		_w1322_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h2)
	) name1921 (
		_w587_,
		_w2138_,
		_w2139_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1922 (
		_w427_,
		_w467_,
		_w592_,
		_w593_,
		_w2140_
	);
	LUT2 #(
		.INIT('h4)
	) name1923 (
		_w427_,
		_w525_,
		_w2141_
	);
	LUT3 #(
		.INIT('h07)
	) name1924 (
		_w601_,
		_w2140_,
		_w2141_,
		_w2142_
	);
	LUT4 #(
		.INIT('hd700)
	) name1925 (
		_w518_,
		_w1445_,
		_w2137_,
		_w2142_,
		_w2143_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1926 (
		\reg1_reg[10]/NET0131 ,
		_w924_,
		_w949_,
		_w1220_,
		_w2144_
	);
	LUT3 #(
		.INIT('h0d)
	) name1927 (
		_w946_,
		_w2143_,
		_w2144_,
		_w2145_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1928 (
		_w254_,
		_w2136_,
		_w2139_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h8)
	) name1929 (
		\reg1_reg[10]/NET0131 ,
		_w252_,
		_w2147_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1930 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[10]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2148_
	);
	LUT4 #(
		.INIT('hffa8)
	) name1931 (
		\state_reg[0]/NET0131 ,
		_w2146_,
		_w2147_,
		_w2148_,
		_w2149_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1932 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[25]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2150_
	);
	LUT2 #(
		.INIT('h8)
	) name1933 (
		\reg1_reg[25]/NET0131 ,
		_w252_,
		_w2151_
	);
	LUT4 #(
		.INIT('haa02)
	) name1934 (
		\reg1_reg[25]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2152_
	);
	LUT4 #(
		.INIT('h2070)
	) name1935 (
		_w266_,
		_w647_,
		_w946_,
		_w1665_,
		_w2153_
	);
	LUT3 #(
		.INIT('ha8)
	) name1936 (
		_w404_,
		_w2152_,
		_w2153_,
		_w2154_
	);
	LUT4 #(
		.INIT('h0a82)
	) name1937 (
		_w946_,
		_w1300_,
		_w1668_,
		_w1675_,
		_w2155_
	);
	LUT3 #(
		.INIT('ha8)
	) name1938 (
		_w587_,
		_w2152_,
		_w2155_,
		_w2156_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1939 (
		\reg1_reg[25]/NET0131 ,
		_w518_,
		_w946_,
		_w1671_,
		_w2157_
	);
	LUT4 #(
		.INIT('h3c55)
	) name1940 (
		\reg1_reg[25]/NET0131 ,
		_w635_,
		_w804_,
		_w946_,
		_w2158_
	);
	LUT3 #(
		.INIT('ha2)
	) name1941 (
		\reg1_reg[25]/NET0131 ,
		_w924_,
		_w959_,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1942 (
		_w946_,
		_w1680_,
		_w2160_
	);
	LUT2 #(
		.INIT('h1)
	) name1943 (
		_w2159_,
		_w2160_,
		_w2161_
	);
	LUT3 #(
		.INIT('hd0)
	) name1944 (
		_w601_,
		_w2158_,
		_w2161_,
		_w2162_
	);
	LUT4 #(
		.INIT('h0100)
	) name1945 (
		_w2157_,
		_w2154_,
		_w2156_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1946 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2151_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('he)
	) name1947 (
		_w2150_,
		_w2164_,
		_w2165_
	);
	LUT4 #(
		.INIT('haa02)
	) name1948 (
		\reg1_reg[3]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2166_
	);
	LUT4 #(
		.INIT('h111d)
	) name1949 (
		\reg1_reg[3]/NET0131 ,
		_w946_,
		_w2074_,
		_w2075_,
		_w2167_
	);
	LUT4 #(
		.INIT('he010)
	) name1950 (
		_w572_,
		_w574_,
		_w946_,
		_w2077_,
		_w2168_
	);
	LUT3 #(
		.INIT('ha8)
	) name1951 (
		_w587_,
		_w2166_,
		_w2168_,
		_w2169_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1952 (
		\reg1_reg[3]/NET0131 ,
		_w924_,
		_w949_,
		_w1220_,
		_w2170_
	);
	LUT4 #(
		.INIT('h005d)
	) name1953 (
		_w946_,
		_w2082_,
		_w2125_,
		_w2170_,
		_w2171_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1954 (
		_w404_,
		_w2167_,
		_w2169_,
		_w2171_,
		_w2172_
	);
	LUT2 #(
		.INIT('h8)
	) name1955 (
		\reg1_reg[3]/NET0131 ,
		_w252_,
		_w2173_
	);
	LUT4 #(
		.INIT('haa08)
	) name1956 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2172_,
		_w2173_,
		_w2174_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1957 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[3]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2175_
	);
	LUT2 #(
		.INIT('he)
	) name1958 (
		_w2174_,
		_w2175_,
		_w2176_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1959 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[10]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2177_
	);
	LUT2 #(
		.INIT('h8)
	) name1960 (
		\reg2_reg[10]/NET0131 ,
		_w252_,
		_w2178_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1961 (
		\reg2_reg[10]/NET0131 ,
		_w970_,
		_w2133_,
		_w2134_,
		_w2179_
	);
	LUT2 #(
		.INIT('h2)
	) name1962 (
		_w404_,
		_w2179_,
		_w2180_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1963 (
		\reg2_reg[10]/NET0131 ,
		_w970_,
		_w1322_,
		_w2137_,
		_w2181_
	);
	LUT2 #(
		.INIT('h2)
	) name1964 (
		_w587_,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('h8)
	) name1965 (
		_w520_,
		_w351_,
		_w2183_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1966 (
		_w256_,
		_w258_,
		_w261_,
		_w1650_,
		_w2184_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1967 (
		\reg2_reg[10]/NET0131 ,
		_w524_,
		_w976_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h1)
	) name1968 (
		_w2183_,
		_w2185_,
		_w2186_
	);
	LUT3 #(
		.INIT('hd0)
	) name1969 (
		_w970_,
		_w2143_,
		_w2186_,
		_w2187_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1970 (
		_w254_,
		_w2180_,
		_w2182_,
		_w2187_,
		_w2188_
	);
	LUT4 #(
		.INIT('heeec)
	) name1971 (
		\state_reg[0]/NET0131 ,
		_w2177_,
		_w2178_,
		_w2188_,
		_w2189_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1972 (
		\reg0_reg[10]/NET0131 ,
		_w917_,
		_w2133_,
		_w2134_,
		_w2190_
	);
	LUT2 #(
		.INIT('h2)
	) name1973 (
		_w404_,
		_w2190_,
		_w2191_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1974 (
		\reg0_reg[10]/NET0131 ,
		_w917_,
		_w1322_,
		_w2137_,
		_w2192_
	);
	LUT2 #(
		.INIT('h2)
	) name1975 (
		_w587_,
		_w2192_,
		_w2193_
	);
	LUT3 #(
		.INIT('ha2)
	) name1976 (
		\reg0_reg[10]/NET0131 ,
		_w924_,
		_w1772_,
		_w2194_
	);
	LUT3 #(
		.INIT('h0d)
	) name1977 (
		_w917_,
		_w2143_,
		_w2194_,
		_w2195_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1978 (
		_w254_,
		_w2191_,
		_w2193_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		\reg0_reg[10]/NET0131 ,
		_w252_,
		_w2197_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1980 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[10]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2198_
	);
	LUT4 #(
		.INIT('hffa8)
	) name1981 (
		\state_reg[0]/NET0131 ,
		_w2196_,
		_w2197_,
		_w2198_,
		_w2199_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name1982 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[18]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2200_
	);
	LUT2 #(
		.INIT('h8)
	) name1983 (
		\reg2_reg[18]/NET0131 ,
		_w252_,
		_w2201_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1984 (
		\reg2_reg[18]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2202_
	);
	LUT4 #(
		.INIT('h08a2)
	) name1985 (
		_w970_,
		_w1427_,
		_w1429_,
		_w1641_,
		_w2203_
	);
	LUT3 #(
		.INIT('ha8)
	) name1986 (
		_w587_,
		_w2202_,
		_w2203_,
		_w2204_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1987 (
		\reg2_reg[18]/NET0131 ,
		_w970_,
		_w1644_,
		_w1645_,
		_w2205_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1988 (
		_w970_,
		_w1647_,
		_w1648_,
		_w2096_,
		_w2206_
	);
	LUT2 #(
		.INIT('h8)
	) name1989 (
		_w520_,
		_w387_,
		_w2207_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1990 (
		\reg2_reg[18]/NET0131 ,
		_w524_,
		_w976_,
		_w2184_,
		_w2208_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		_w2207_,
		_w2208_,
		_w2209_
	);
	LUT4 #(
		.INIT('h3100)
	) name1992 (
		_w404_,
		_w2206_,
		_w2205_,
		_w2209_,
		_w2210_
	);
	LUT4 #(
		.INIT('h1311)
	) name1993 (
		_w254_,
		_w2201_,
		_w2204_,
		_w2210_,
		_w2211_
	);
	LUT3 #(
		.INIT('hce)
	) name1994 (
		\state_reg[0]/NET0131 ,
		_w2200_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h8)
	) name1995 (
		_w252_,
		_w306_,
		_w2213_
	);
	LUT3 #(
		.INIT('h87)
	) name1996 (
		_w307_,
		_w308_,
		_w488_,
		_w2214_
	);
	LUT4 #(
		.INIT('h000d)
	) name1997 (
		_w505_,
		_w697_,
		_w698_,
		_w2214_,
		_w2215_
	);
	LUT4 #(
		.INIT('hf200)
	) name1998 (
		_w505_,
		_w697_,
		_w698_,
		_w2214_,
		_w2216_
	);
	LUT3 #(
		.INIT('h02)
	) name1999 (
		_w518_,
		_w2216_,
		_w2215_,
		_w2217_
	);
	LUT3 #(
		.INIT('h60)
	) name2000 (
		_w488_,
		_w590_,
		_w601_,
		_w2218_
	);
	LUT4 #(
		.INIT('h0d07)
	) name2001 (
		_w587_,
		_w758_,
		_w2218_,
		_w2214_,
		_w2219_
	);
	LUT3 #(
		.INIT('h8a)
	) name2002 (
		_w262_,
		_w2217_,
		_w2219_,
		_w2220_
	);
	LUT4 #(
		.INIT('h1540)
	) name2003 (
		_w266_,
		_w301_,
		_w311_,
		_w320_,
		_w2221_
	);
	LUT3 #(
		.INIT('h80)
	) name2004 (
		_w266_,
		_w302_,
		_w303_,
		_w2222_
	);
	LUT4 #(
		.INIT('h001f)
	) name2005 (
		_w256_,
		_w258_,
		_w261_,
		_w306_,
		_w2223_
	);
	LUT2 #(
		.INIT('h2)
	) name2006 (
		_w404_,
		_w2223_,
		_w2224_
	);
	LUT4 #(
		.INIT('h5700)
	) name2007 (
		_w262_,
		_w2221_,
		_w2222_,
		_w2224_,
		_w2225_
	);
	LUT3 #(
		.INIT('h04)
	) name2008 (
		_w521_,
		_w522_,
		_w488_,
		_w2226_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2009 (
		_w256_,
		_w258_,
		_w261_,
		_w517_,
		_w2227_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2010 (
		_w306_,
		_w524_,
		_w906_,
		_w2227_,
		_w2228_
	);
	LUT2 #(
		.INIT('h1)
	) name2011 (
		_w2226_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h4)
	) name2012 (
		_w2225_,
		_w2229_,
		_w2230_
	);
	LUT4 #(
		.INIT('h1311)
	) name2013 (
		_w254_,
		_w2213_,
		_w2220_,
		_w2230_,
		_w2231_
	);
	LUT3 #(
		.INIT('h6c)
	) name2014 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2232_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2015 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2232_,
		_w2233_
	);
	LUT3 #(
		.INIT('hf2)
	) name2016 (
		\state_reg[0]/NET0131 ,
		_w2231_,
		_w2233_,
		_w2234_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2017 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[6]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name2018 (
		\reg2_reg[6]/NET0131 ,
		_w252_,
		_w2236_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2019 (
		\reg2_reg[6]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2237_
	);
	LUT4 #(
		.INIT('h7020)
	) name2020 (
		_w266_,
		_w320_,
		_w970_,
		_w1999_,
		_w2238_
	);
	LUT3 #(
		.INIT('ha8)
	) name2021 (
		_w404_,
		_w2237_,
		_w2238_,
		_w2239_
	);
	LUT4 #(
		.INIT('h40b0)
	) name2022 (
		_w760_,
		_w761_,
		_w970_,
		_w2002_,
		_w2240_
	);
	LUT3 #(
		.INIT('ha8)
	) name2023 (
		_w587_,
		_w2237_,
		_w2240_,
		_w2241_
	);
	LUT4 #(
		.INIT('he010)
	) name2024 (
		_w700_,
		_w701_,
		_w970_,
		_w2002_,
		_w2242_
	);
	LUT2 #(
		.INIT('h4)
	) name2025 (
		_w475_,
		_w525_,
		_w2243_
	);
	LUT4 #(
		.INIT('h009f)
	) name2026 (
		_w475_,
		_w591_,
		_w601_,
		_w2243_,
		_w2244_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2027 (
		\reg2_reg[6]/NET0131 ,
		_w524_,
		_w976_,
		_w991_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name2028 (
		_w520_,
		_w313_,
		_w2246_
	);
	LUT2 #(
		.INIT('h1)
	) name2029 (
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT3 #(
		.INIT('hd0)
	) name2030 (
		_w970_,
		_w2244_,
		_w2247_,
		_w2248_
	);
	LUT4 #(
		.INIT('h5700)
	) name2031 (
		_w518_,
		_w2237_,
		_w2242_,
		_w2248_,
		_w2249_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2032 (
		_w254_,
		_w2239_,
		_w2241_,
		_w2249_,
		_w2250_
	);
	LUT4 #(
		.INIT('heeec)
	) name2033 (
		\state_reg[0]/NET0131 ,
		_w2235_,
		_w2236_,
		_w2250_,
		_w2251_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2034 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[8]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2252_
	);
	LUT2 #(
		.INIT('h8)
	) name2035 (
		\reg2_reg[8]/NET0131 ,
		_w252_,
		_w2253_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2036 (
		\reg2_reg[8]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2254_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2037 (
		_w970_,
		_w1800_,
		_w1801_,
		_w1802_,
		_w2255_
	);
	LUT3 #(
		.INIT('ha8)
	) name2038 (
		_w404_,
		_w2254_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('hc808)
	) name2039 (
		\reg2_reg[8]/NET0131 ,
		_w587_,
		_w970_,
		_w1806_,
		_w2257_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2040 (
		\reg2_reg[8]/NET0131 ,
		_w518_,
		_w970_,
		_w1808_,
		_w2258_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2041 (
		_w467_,
		_w470_,
		_w592_,
		_w970_,
		_w2259_
	);
	LUT3 #(
		.INIT('ha8)
	) name2042 (
		\reg2_reg[8]/NET0131 ,
		_w524_,
		_w976_,
		_w2260_
	);
	LUT2 #(
		.INIT('h8)
	) name2043 (
		_w520_,
		_w329_,
		_w2261_
	);
	LUT3 #(
		.INIT('h07)
	) name2044 (
		_w970_,
		_w1812_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h4)
	) name2045 (
		_w2260_,
		_w2262_,
		_w2263_
	);
	LUT4 #(
		.INIT('h5700)
	) name2046 (
		_w601_,
		_w2254_,
		_w2259_,
		_w2263_,
		_w2264_
	);
	LUT3 #(
		.INIT('h10)
	) name2047 (
		_w2258_,
		_w2257_,
		_w2264_,
		_w2265_
	);
	LUT4 #(
		.INIT('h1311)
	) name2048 (
		_w254_,
		_w2253_,
		_w2256_,
		_w2265_,
		_w2266_
	);
	LUT3 #(
		.INIT('hce)
	) name2049 (
		\state_reg[0]/NET0131 ,
		_w2252_,
		_w2266_,
		_w2267_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2050 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[17]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2268_
	);
	LUT2 #(
		.INIT('h8)
	) name2051 (
		\reg0_reg[17]/NET0131 ,
		_w252_,
		_w2269_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2052 (
		\reg0_reg[17]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2270_
	);
	LUT4 #(
		.INIT('hfc55)
	) name2053 (
		\reg0_reg[17]/NET0131 ,
		_w395_,
		_w396_,
		_w917_,
		_w2271_
	);
	LUT2 #(
		.INIT('h2)
	) name2054 (
		_w404_,
		_w2271_,
		_w2272_
	);
	LUT4 #(
		.INIT('h30a0)
	) name2055 (
		\reg0_reg[17]/NET0131 ,
		_w514_,
		_w518_,
		_w917_,
		_w2273_
	);
	LUT2 #(
		.INIT('h8)
	) name2056 (
		_w411_,
		_w525_,
		_w2274_
	);
	LUT2 #(
		.INIT('h8)
	) name2057 (
		_w917_,
		_w2274_,
		_w2275_
	);
	LUT3 #(
		.INIT('h8a)
	) name2058 (
		\reg0_reg[17]/NET0131 ,
		_w923_,
		_w924_,
		_w2276_
	);
	LUT2 #(
		.INIT('h1)
	) name2059 (
		_w2275_,
		_w2276_,
		_w2277_
	);
	LUT4 #(
		.INIT('h5900)
	) name2060 (
		_w414_,
		_w552_,
		_w585_,
		_w917_,
		_w2278_
	);
	LUT3 #(
		.INIT('ha8)
	) name2061 (
		_w587_,
		_w2270_,
		_w2278_,
		_w2279_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2062 (
		_w411_,
		_w597_,
		_w599_,
		_w917_,
		_w2280_
	);
	LUT3 #(
		.INIT('ha8)
	) name2063 (
		_w601_,
		_w2270_,
		_w2280_,
		_w2281_
	);
	LUT4 #(
		.INIT('h0100)
	) name2064 (
		_w2273_,
		_w2279_,
		_w2281_,
		_w2277_,
		_w2282_
	);
	LUT4 #(
		.INIT('h1311)
	) name2065 (
		_w254_,
		_w2269_,
		_w2272_,
		_w2282_,
		_w2283_
	);
	LUT3 #(
		.INIT('hce)
	) name2066 (
		\state_reg[0]/NET0131 ,
		_w2268_,
		_w2283_,
		_w2284_
	);
	LUT2 #(
		.INIT('h4)
	) name2067 (
		_w491_,
		_w525_,
		_w2285_
	);
	LUT4 #(
		.INIT('h0010)
	) name2068 (
		_w1959_,
		_w1962_,
		_w1966_,
		_w2285_,
		_w2286_
	);
	LUT4 #(
		.INIT('hf7e2)
	) name2069 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w2287_
	);
	LUT4 #(
		.INIT('h4066)
	) name2070 (
		_w401_,
		_w398_,
		_w403_,
		_w400_,
		_w2288_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2071 (
		_w256_,
		_w258_,
		_w261_,
		_w2288_,
		_w2289_
	);
	LUT2 #(
		.INIT('h2)
	) name2072 (
		_w1410_,
		_w2289_,
		_w2290_
	);
	LUT3 #(
		.INIT('h2a)
	) name2073 (
		\reg0_reg[1]/NET0131 ,
		_w1155_,
		_w2290_,
		_w2291_
	);
	LUT3 #(
		.INIT('hf2)
	) name2074 (
		_w1781_,
		_w2286_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2075 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[21]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2293_
	);
	LUT2 #(
		.INIT('h8)
	) name2076 (
		\reg0_reg[21]/NET0131 ,
		_w252_,
		_w2294_
	);
	LUT4 #(
		.INIT('h999f)
	) name2077 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w2295_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2078 (
		_w256_,
		_w258_,
		_w261_,
		_w2295_,
		_w2296_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2079 (
		\reg0_reg[21]/NET0131 ,
		_w923_,
		_w924_,
		_w2296_,
		_w2297_
	);
	LUT2 #(
		.INIT('h8)
	) name2080 (
		_w525_,
		_w660_,
		_w2298_
	);
	LUT3 #(
		.INIT('h82)
	) name2081 (
		_w601_,
		_w660_,
		_w1397_,
		_w2299_
	);
	LUT2 #(
		.INIT('h9)
	) name2082 (
		_w660_,
		_w665_,
		_w2300_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2083 (
		_w1289_,
		_w1291_,
		_w1293_,
		_w2300_,
		_w2301_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2084 (
		_w1289_,
		_w1291_,
		_w1293_,
		_w2300_,
		_w2302_
	);
	LUT3 #(
		.INIT('h02)
	) name2085 (
		_w587_,
		_w2302_,
		_w2301_,
		_w2303_
	);
	LUT3 #(
		.INIT('h28)
	) name2086 (
		_w518_,
		_w1278_,
		_w2300_,
		_w2304_
	);
	LUT4 #(
		.INIT('h0001)
	) name2087 (
		_w2298_,
		_w2303_,
		_w2304_,
		_w2299_,
		_w2305_
	);
	LUT4 #(
		.INIT('h4144)
	) name2088 (
		_w266_,
		_w657_,
		_w665_,
		_w1070_,
		_w2306_
	);
	LUT2 #(
		.INIT('h8)
	) name2089 (
		_w266_,
		_w671_,
		_w2307_
	);
	LUT3 #(
		.INIT('h02)
	) name2090 (
		_w404_,
		_w2306_,
		_w2307_,
		_w2308_
	);
	LUT4 #(
		.INIT('h1131)
	) name2091 (
		_w917_,
		_w2297_,
		_w2305_,
		_w2308_,
		_w2309_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2092 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2294_,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('he)
	) name2093 (
		_w2293_,
		_w2310_,
		_w2311_
	);
	LUT4 #(
		.INIT('h0040)
	) name2094 (
		_w923_,
		_w924_,
		_w1410_,
		_w2296_,
		_w2312_
	);
	LUT2 #(
		.INIT('h2)
	) name2095 (
		\reg0_reg[2]/NET0131 ,
		_w2312_,
		_w2313_
	);
	LUT2 #(
		.INIT('h4)
	) name2096 (
		_w497_,
		_w525_,
		_w2314_
	);
	LUT3 #(
		.INIT('h04)
	) name2097 (
		_w1983_,
		_w1985_,
		_w2314_,
		_w2315_
	);
	LUT2 #(
		.INIT('h8)
	) name2098 (
		_w404_,
		_w1978_,
		_w2316_
	);
	LUT4 #(
		.INIT('h8808)
	) name2099 (
		_w917_,
		_w1410_,
		_w2315_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('he)
	) name2100 (
		_w2313_,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('h2)
	) name2101 (
		\reg0_reg[4]/NET0131 ,
		_w2312_,
		_w2319_
	);
	LUT3 #(
		.INIT('h02)
	) name2102 (
		_w404_,
		_w2221_,
		_w2222_,
		_w2320_
	);
	LUT2 #(
		.INIT('h4)
	) name2103 (
		_w488_,
		_w525_,
		_w2321_
	);
	LUT4 #(
		.INIT('h0004)
	) name2104 (
		_w2217_,
		_w2219_,
		_w2321_,
		_w2320_,
		_w2322_
	);
	LUT4 #(
		.INIT('hf0f8)
	) name2105 (
		_w917_,
		_w1410_,
		_w2319_,
		_w2322_,
		_w2323_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2106 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[5]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2324_
	);
	LUT2 #(
		.INIT('h8)
	) name2107 (
		\reg0_reg[5]/NET0131 ,
		_w252_,
		_w2325_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2108 (
		\reg0_reg[5]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2326_
	);
	LUT3 #(
		.INIT('h2a)
	) name2109 (
		_w266_,
		_w307_,
		_w308_,
		_w2327_
	);
	LUT4 #(
		.INIT('hf070)
	) name2110 (
		_w301_,
		_w311_,
		_w315_,
		_w320_,
		_w2328_
	);
	LUT4 #(
		.INIT('h1555)
	) name2111 (
		_w266_,
		_w301_,
		_w311_,
		_w322_,
		_w2329_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2112 (
		_w917_,
		_w2327_,
		_w2328_,
		_w2329_,
		_w2330_
	);
	LUT3 #(
		.INIT('ha8)
	) name2113 (
		_w404_,
		_w2326_,
		_w2330_,
		_w2331_
	);
	LUT3 #(
		.INIT('h87)
	) name2114 (
		_w318_,
		_w319_,
		_w479_,
		_w2332_
	);
	LUT4 #(
		.INIT('hc535)
	) name2115 (
		\reg0_reg[5]/NET0131 ,
		_w509_,
		_w917_,
		_w2332_,
		_w2333_
	);
	LUT4 #(
		.INIT('hf40b)
	) name2116 (
		_w572_,
		_w577_,
		_w580_,
		_w2332_,
		_w2334_
	);
	LUT4 #(
		.INIT('hc808)
	) name2117 (
		\reg0_reg[5]/NET0131 ,
		_w587_,
		_w917_,
		_w2334_,
		_w2335_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2118 (
		\reg0_reg[5]/NET0131 ,
		_w923_,
		_w924_,
		_w1154_,
		_w2336_
	);
	LUT2 #(
		.INIT('h4)
	) name2119 (
		_w479_,
		_w525_,
		_w2337_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2120 (
		_w479_,
		_w488_,
		_w590_,
		_w601_,
		_w2338_
	);
	LUT4 #(
		.INIT('h1113)
	) name2121 (
		_w917_,
		_w2336_,
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT4 #(
		.INIT('h3100)
	) name2122 (
		_w518_,
		_w2335_,
		_w2333_,
		_w2339_,
		_w2340_
	);
	LUT4 #(
		.INIT('h1311)
	) name2123 (
		_w254_,
		_w2325_,
		_w2331_,
		_w2340_,
		_w2341_
	);
	LUT3 #(
		.INIT('hce)
	) name2124 (
		\state_reg[0]/NET0131 ,
		_w2324_,
		_w2341_,
		_w2342_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2125 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[6]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2343_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		\reg0_reg[6]/NET0131 ,
		_w252_,
		_w2344_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2127 (
		\reg0_reg[6]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2345_
	);
	LUT4 #(
		.INIT('h7020)
	) name2128 (
		_w266_,
		_w320_,
		_w917_,
		_w1999_,
		_w2346_
	);
	LUT3 #(
		.INIT('ha8)
	) name2129 (
		_w404_,
		_w2345_,
		_w2346_,
		_w2347_
	);
	LUT4 #(
		.INIT('h40b0)
	) name2130 (
		_w760_,
		_w761_,
		_w917_,
		_w2002_,
		_w2348_
	);
	LUT3 #(
		.INIT('ha8)
	) name2131 (
		_w587_,
		_w2345_,
		_w2348_,
		_w2349_
	);
	LUT4 #(
		.INIT('he010)
	) name2132 (
		_w700_,
		_w701_,
		_w917_,
		_w2002_,
		_w2350_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2133 (
		\reg0_reg[6]/NET0131 ,
		_w923_,
		_w924_,
		_w1154_,
		_w2351_
	);
	LUT3 #(
		.INIT('h0d)
	) name2134 (
		_w917_,
		_w2244_,
		_w2351_,
		_w2352_
	);
	LUT4 #(
		.INIT('h5700)
	) name2135 (
		_w518_,
		_w2345_,
		_w2350_,
		_w2352_,
		_w2353_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2136 (
		_w254_,
		_w2347_,
		_w2349_,
		_w2353_,
		_w2354_
	);
	LUT4 #(
		.INIT('heeec)
	) name2137 (
		\state_reg[0]/NET0131 ,
		_w2343_,
		_w2344_,
		_w2354_,
		_w2355_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2138 (
		\IR_reg[23]/NET0131 ,
		\reg0_reg[9]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2356_
	);
	LUT2 #(
		.INIT('h8)
	) name2139 (
		\reg0_reg[9]/NET0131 ,
		_w252_,
		_w2357_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2140 (
		\reg0_reg[9]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2358_
	);
	LUT4 #(
		.INIT('hc808)
	) name2141 (
		\reg0_reg[9]/NET0131 ,
		_w404_,
		_w917_,
		_w2037_,
		_w2359_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2142 (
		\reg0_reg[9]/NET0131 ,
		_w518_,
		_w917_,
		_w2040_,
		_w2360_
	);
	LUT4 #(
		.INIT('hd020)
	) name2143 (
		_w566_,
		_w584_,
		_w917_,
		_w2039_,
		_w2361_
	);
	LUT3 #(
		.INIT('ha8)
	) name2144 (
		_w587_,
		_w2358_,
		_w2361_,
		_w2362_
	);
	LUT4 #(
		.INIT('hc808)
	) name2145 (
		\reg0_reg[9]/NET0131 ,
		_w601_,
		_w917_,
		_w2044_,
		_w2363_
	);
	LUT2 #(
		.INIT('h4)
	) name2146 (
		_w431_,
		_w525_,
		_w2364_
	);
	LUT2 #(
		.INIT('h8)
	) name2147 (
		_w917_,
		_w2364_,
		_w2365_
	);
	LUT3 #(
		.INIT('h8a)
	) name2148 (
		\reg0_reg[9]/NET0131 ,
		_w923_,
		_w924_,
		_w2366_
	);
	LUT2 #(
		.INIT('h1)
	) name2149 (
		_w2365_,
		_w2366_,
		_w2367_
	);
	LUT2 #(
		.INIT('h4)
	) name2150 (
		_w2363_,
		_w2367_,
		_w2368_
	);
	LUT4 #(
		.INIT('h0100)
	) name2151 (
		_w2359_,
		_w2362_,
		_w2360_,
		_w2368_,
		_w2369_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2152 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2357_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('he)
	) name2153 (
		_w2356_,
		_w2370_,
		_w2371_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2154 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[17]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2372_
	);
	LUT2 #(
		.INIT('h8)
	) name2155 (
		\reg1_reg[17]/NET0131 ,
		_w252_,
		_w2373_
	);
	LUT4 #(
		.INIT('haa02)
	) name2156 (
		\reg1_reg[17]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2374_
	);
	LUT4 #(
		.INIT('hfc55)
	) name2157 (
		\reg1_reg[17]/NET0131 ,
		_w395_,
		_w396_,
		_w946_,
		_w2375_
	);
	LUT2 #(
		.INIT('h2)
	) name2158 (
		_w404_,
		_w2375_,
		_w2376_
	);
	LUT4 #(
		.INIT('h30a0)
	) name2159 (
		\reg1_reg[17]/NET0131 ,
		_w514_,
		_w518_,
		_w946_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		_w946_,
		_w2274_,
		_w2378_
	);
	LUT3 #(
		.INIT('ha2)
	) name2161 (
		\reg1_reg[17]/NET0131 ,
		_w924_,
		_w959_,
		_w2379_
	);
	LUT2 #(
		.INIT('h1)
	) name2162 (
		_w2378_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('h5900)
	) name2163 (
		_w414_,
		_w552_,
		_w585_,
		_w946_,
		_w2381_
	);
	LUT3 #(
		.INIT('ha8)
	) name2164 (
		_w587_,
		_w2374_,
		_w2381_,
		_w2382_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2165 (
		_w411_,
		_w597_,
		_w599_,
		_w946_,
		_w2383_
	);
	LUT3 #(
		.INIT('ha8)
	) name2166 (
		_w601_,
		_w2374_,
		_w2383_,
		_w2384_
	);
	LUT4 #(
		.INIT('h0100)
	) name2167 (
		_w2377_,
		_w2382_,
		_w2384_,
		_w2380_,
		_w2385_
	);
	LUT4 #(
		.INIT('h1311)
	) name2168 (
		_w254_,
		_w2373_,
		_w2376_,
		_w2385_,
		_w2386_
	);
	LUT3 #(
		.INIT('hce)
	) name2169 (
		\state_reg[0]/NET0131 ,
		_w2372_,
		_w2386_,
		_w2387_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2170 (
		_w256_,
		_w258_,
		_w261_,
		_w2288_,
		_w2388_
	);
	LUT4 #(
		.INIT('h0020)
	) name2171 (
		_w924_,
		_w949_,
		_w1410_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h2)
	) name2172 (
		\reg1_reg[1]/NET0131 ,
		_w2389_,
		_w2390_
	);
	LUT3 #(
		.INIT('hf2)
	) name2173 (
		_w1871_,
		_w2286_,
		_w2390_,
		_w2391_
	);
	LUT4 #(
		.INIT('hf100)
	) name2174 (
		_w256_,
		_w258_,
		_w261_,
		_w2295_,
		_w2392_
	);
	LUT4 #(
		.INIT('h0020)
	) name2175 (
		_w924_,
		_w959_,
		_w1410_,
		_w2392_,
		_w2393_
	);
	LUT2 #(
		.INIT('h2)
	) name2176 (
		\reg1_reg[2]/NET0131 ,
		_w2393_,
		_w2394_
	);
	LUT4 #(
		.INIT('h8808)
	) name2177 (
		_w946_,
		_w1410_,
		_w2315_,
		_w2316_,
		_w2395_
	);
	LUT2 #(
		.INIT('he)
	) name2178 (
		_w2394_,
		_w2395_,
		_w2396_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2179 (
		_w256_,
		_w258_,
		_w261_,
		_w1604_,
		_w2397_
	);
	LUT2 #(
		.INIT('h2)
	) name2180 (
		_w1410_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('h2a)
	) name2181 (
		\reg1_reg[4]/NET0131 ,
		_w961_,
		_w2398_,
		_w2399_
	);
	LUT4 #(
		.INIT('hff08)
	) name2182 (
		_w946_,
		_w1410_,
		_w2322_,
		_w2399_,
		_w2400_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2183 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[5]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2401_
	);
	LUT2 #(
		.INIT('h8)
	) name2184 (
		\reg1_reg[5]/NET0131 ,
		_w252_,
		_w2402_
	);
	LUT4 #(
		.INIT('haa02)
	) name2185 (
		\reg1_reg[5]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2403_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2186 (
		_w946_,
		_w2327_,
		_w2328_,
		_w2329_,
		_w2404_
	);
	LUT3 #(
		.INIT('ha8)
	) name2187 (
		_w404_,
		_w2403_,
		_w2404_,
		_w2405_
	);
	LUT4 #(
		.INIT('hc535)
	) name2188 (
		\reg1_reg[5]/NET0131 ,
		_w509_,
		_w946_,
		_w2332_,
		_w2406_
	);
	LUT4 #(
		.INIT('hc808)
	) name2189 (
		\reg1_reg[5]/NET0131 ,
		_w587_,
		_w946_,
		_w2334_,
		_w2407_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2190 (
		\reg1_reg[5]/NET0131 ,
		_w924_,
		_w959_,
		_w960_,
		_w2408_
	);
	LUT4 #(
		.INIT('h0057)
	) name2191 (
		_w946_,
		_w2337_,
		_w2338_,
		_w2408_,
		_w2409_
	);
	LUT4 #(
		.INIT('h3100)
	) name2192 (
		_w518_,
		_w2407_,
		_w2406_,
		_w2409_,
		_w2410_
	);
	LUT4 #(
		.INIT('h1311)
	) name2193 (
		_w254_,
		_w2402_,
		_w2405_,
		_w2410_,
		_w2411_
	);
	LUT3 #(
		.INIT('hce)
	) name2194 (
		\state_reg[0]/NET0131 ,
		_w2401_,
		_w2411_,
		_w2412_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2195 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[6]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2413_
	);
	LUT2 #(
		.INIT('h8)
	) name2196 (
		\reg1_reg[6]/NET0131 ,
		_w252_,
		_w2414_
	);
	LUT4 #(
		.INIT('haa02)
	) name2197 (
		\reg1_reg[6]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2415_
	);
	LUT4 #(
		.INIT('h7020)
	) name2198 (
		_w266_,
		_w320_,
		_w946_,
		_w1999_,
		_w2416_
	);
	LUT3 #(
		.INIT('ha8)
	) name2199 (
		_w404_,
		_w2415_,
		_w2416_,
		_w2417_
	);
	LUT4 #(
		.INIT('h40b0)
	) name2200 (
		_w760_,
		_w761_,
		_w946_,
		_w2002_,
		_w2418_
	);
	LUT3 #(
		.INIT('ha8)
	) name2201 (
		_w587_,
		_w2415_,
		_w2418_,
		_w2419_
	);
	LUT4 #(
		.INIT('he010)
	) name2202 (
		_w700_,
		_w701_,
		_w946_,
		_w2002_,
		_w2420_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2203 (
		\reg1_reg[6]/NET0131 ,
		_w924_,
		_w959_,
		_w960_,
		_w2421_
	);
	LUT3 #(
		.INIT('h0d)
	) name2204 (
		_w946_,
		_w2244_,
		_w2421_,
		_w2422_
	);
	LUT4 #(
		.INIT('h5700)
	) name2205 (
		_w518_,
		_w2415_,
		_w2420_,
		_w2422_,
		_w2423_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2206 (
		_w254_,
		_w2417_,
		_w2419_,
		_w2423_,
		_w2424_
	);
	LUT4 #(
		.INIT('heeec)
	) name2207 (
		\state_reg[0]/NET0131 ,
		_w2413_,
		_w2414_,
		_w2424_,
		_w2425_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2208 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[8]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2426_
	);
	LUT2 #(
		.INIT('h8)
	) name2209 (
		\reg1_reg[8]/NET0131 ,
		_w252_,
		_w2427_
	);
	LUT4 #(
		.INIT('haa02)
	) name2210 (
		\reg1_reg[8]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2428_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2211 (
		_w946_,
		_w1800_,
		_w1801_,
		_w1802_,
		_w2429_
	);
	LUT3 #(
		.INIT('ha8)
	) name2212 (
		_w404_,
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT4 #(
		.INIT('hc808)
	) name2213 (
		\reg1_reg[8]/NET0131 ,
		_w587_,
		_w946_,
		_w1806_,
		_w2431_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2214 (
		\reg1_reg[8]/NET0131 ,
		_w518_,
		_w946_,
		_w1808_,
		_w2432_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2215 (
		_w467_,
		_w470_,
		_w592_,
		_w946_,
		_w2433_
	);
	LUT2 #(
		.INIT('h8)
	) name2216 (
		_w946_,
		_w1812_,
		_w2434_
	);
	LUT3 #(
		.INIT('ha2)
	) name2217 (
		\reg1_reg[8]/NET0131 ,
		_w924_,
		_w959_,
		_w2435_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		_w2434_,
		_w2435_,
		_w2436_
	);
	LUT4 #(
		.INIT('h5700)
	) name2219 (
		_w601_,
		_w2428_,
		_w2433_,
		_w2436_,
		_w2437_
	);
	LUT3 #(
		.INIT('h10)
	) name2220 (
		_w2432_,
		_w2431_,
		_w2437_,
		_w2438_
	);
	LUT4 #(
		.INIT('h1311)
	) name2221 (
		_w254_,
		_w2427_,
		_w2430_,
		_w2438_,
		_w2439_
	);
	LUT3 #(
		.INIT('hce)
	) name2222 (
		\state_reg[0]/NET0131 ,
		_w2426_,
		_w2439_,
		_w2440_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2223 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[9]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2441_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		\reg1_reg[9]/NET0131 ,
		_w252_,
		_w2442_
	);
	LUT4 #(
		.INIT('haa02)
	) name2225 (
		\reg1_reg[9]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2443_
	);
	LUT4 #(
		.INIT('hc808)
	) name2226 (
		\reg1_reg[9]/NET0131 ,
		_w404_,
		_w946_,
		_w2037_,
		_w2444_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2227 (
		\reg1_reg[9]/NET0131 ,
		_w518_,
		_w946_,
		_w2040_,
		_w2445_
	);
	LUT4 #(
		.INIT('hd020)
	) name2228 (
		_w566_,
		_w584_,
		_w946_,
		_w2039_,
		_w2446_
	);
	LUT3 #(
		.INIT('ha8)
	) name2229 (
		_w587_,
		_w2443_,
		_w2446_,
		_w2447_
	);
	LUT4 #(
		.INIT('hc808)
	) name2230 (
		\reg1_reg[9]/NET0131 ,
		_w601_,
		_w946_,
		_w2044_,
		_w2448_
	);
	LUT2 #(
		.INIT('h8)
	) name2231 (
		_w946_,
		_w2364_,
		_w2449_
	);
	LUT3 #(
		.INIT('ha2)
	) name2232 (
		\reg1_reg[9]/NET0131 ,
		_w924_,
		_w959_,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		_w2449_,
		_w2450_,
		_w2451_
	);
	LUT2 #(
		.INIT('h4)
	) name2234 (
		_w2448_,
		_w2451_,
		_w2452_
	);
	LUT4 #(
		.INIT('h0100)
	) name2235 (
		_w2444_,
		_w2447_,
		_w2445_,
		_w2452_,
		_w2453_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2236 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2442_,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('he)
	) name2237 (
		_w2441_,
		_w2454_,
		_w2455_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2238 (
		\IR_reg[23]/NET0131 ,
		\reg3_reg[0]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2456_
	);
	LUT2 #(
		.INIT('h8)
	) name2239 (
		\reg3_reg[0]/NET0131 ,
		_w252_,
		_w2457_
	);
	LUT2 #(
		.INIT('h4)
	) name2240 (
		_w493_,
		_w905_,
		_w2458_
	);
	LUT4 #(
		.INIT('h1114)
	) name2241 (
		_w266_,
		_w280_,
		_w284_,
		_w299_,
		_w2459_
	);
	LUT3 #(
		.INIT('h70)
	) name2242 (
		_w282_,
		_w283_,
		_w493_,
		_w2460_
	);
	LUT3 #(
		.INIT('h87)
	) name2243 (
		_w282_,
		_w283_,
		_w493_,
		_w2461_
	);
	LUT4 #(
		.INIT('h7800)
	) name2244 (
		_w282_,
		_w283_,
		_w493_,
		_w517_,
		_w2462_
	);
	LUT4 #(
		.INIT('h0013)
	) name2245 (
		_w404_,
		_w2458_,
		_w2459_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h2)
	) name2246 (
		_w520_,
		_w493_,
		_w2464_
	);
	LUT4 #(
		.INIT('h0057)
	) name2247 (
		\reg3_reg[0]/NET0131 ,
		_w521_,
		_w524_,
		_w2464_,
		_w2465_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2248 (
		_w254_,
		_w262_,
		_w2463_,
		_w2465_,
		_w2466_
	);
	LUT4 #(
		.INIT('heeec)
	) name2249 (
		\state_reg[0]/NET0131 ,
		_w2456_,
		_w2457_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h8)
	) name2250 (
		_w252_,
		_w662_,
		_w2468_
	);
	LUT4 #(
		.INIT('h001f)
	) name2251 (
		_w256_,
		_w258_,
		_w261_,
		_w662_,
		_w2469_
	);
	LUT2 #(
		.INIT('h2)
	) name2252 (
		_w404_,
		_w2469_,
		_w2470_
	);
	LUT4 #(
		.INIT('h5700)
	) name2253 (
		_w262_,
		_w2306_,
		_w2307_,
		_w2470_,
		_w2471_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2254 (
		_w262_,
		_w2303_,
		_w2304_,
		_w2299_,
		_w2472_
	);
	LUT3 #(
		.INIT('h40)
	) name2255 (
		_w521_,
		_w522_,
		_w660_,
		_w2473_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name2256 (
		_w524_,
		_w526_,
		_w662_,
		_w1991_,
		_w2474_
	);
	LUT2 #(
		.INIT('h1)
	) name2257 (
		_w2473_,
		_w2474_,
		_w2475_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2258 (
		_w254_,
		_w2472_,
		_w2471_,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h2)
	) name2259 (
		\reg3_reg[21]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2477_
	);
	LUT3 #(
		.INIT('h07)
	) name2260 (
		_w606_,
		_w662_,
		_w2477_,
		_w2478_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2261 (
		\state_reg[0]/NET0131 ,
		_w2468_,
		_w2476_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2262 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[4]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2480_
	);
	LUT2 #(
		.INIT('h8)
	) name2263 (
		\reg2_reg[4]/NET0131 ,
		_w252_,
		_w2481_
	);
	LUT2 #(
		.INIT('h8)
	) name2264 (
		_w520_,
		_w306_,
		_w2482_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2265 (
		_w256_,
		_w258_,
		_w261_,
		_w2287_,
		_w2483_
	);
	LUT4 #(
		.INIT('h0001)
	) name2266 (
		_w524_,
		_w976_,
		_w2184_,
		_w2483_,
		_w2484_
	);
	LUT3 #(
		.INIT('h31)
	) name2267 (
		\reg2_reg[4]/NET0131 ,
		_w2482_,
		_w2484_,
		_w2485_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2268 (
		_w254_,
		_w970_,
		_w2322_,
		_w2485_,
		_w2486_
	);
	LUT4 #(
		.INIT('heeec)
	) name2269 (
		\state_reg[0]/NET0131 ,
		_w2480_,
		_w2481_,
		_w2486_,
		_w2487_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2270 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[5]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2488_
	);
	LUT2 #(
		.INIT('h8)
	) name2271 (
		\reg2_reg[5]/NET0131 ,
		_w252_,
		_w2489_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2272 (
		\reg2_reg[5]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2490_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2273 (
		_w970_,
		_w2327_,
		_w2328_,
		_w2329_,
		_w2491_
	);
	LUT3 #(
		.INIT('ha8)
	) name2274 (
		_w404_,
		_w2490_,
		_w2491_,
		_w2492_
	);
	LUT4 #(
		.INIT('hc535)
	) name2275 (
		\reg2_reg[5]/NET0131 ,
		_w509_,
		_w970_,
		_w2332_,
		_w2493_
	);
	LUT4 #(
		.INIT('hc808)
	) name2276 (
		\reg2_reg[5]/NET0131 ,
		_w587_,
		_w970_,
		_w2334_,
		_w2494_
	);
	LUT3 #(
		.INIT('ha8)
	) name2277 (
		_w970_,
		_w2337_,
		_w2338_,
		_w2495_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2278 (
		\reg2_reg[5]/NET0131 ,
		_w524_,
		_w976_,
		_w991_,
		_w2496_
	);
	LUT2 #(
		.INIT('h8)
	) name2279 (
		_w520_,
		_w317_,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name2280 (
		_w2496_,
		_w2497_,
		_w2498_
	);
	LUT2 #(
		.INIT('h4)
	) name2281 (
		_w2495_,
		_w2498_,
		_w2499_
	);
	LUT4 #(
		.INIT('h3100)
	) name2282 (
		_w518_,
		_w2494_,
		_w2493_,
		_w2499_,
		_w2500_
	);
	LUT4 #(
		.INIT('h1311)
	) name2283 (
		_w254_,
		_w2489_,
		_w2492_,
		_w2500_,
		_w2501_
	);
	LUT3 #(
		.INIT('hce)
	) name2284 (
		\state_reg[0]/NET0131 ,
		_w2488_,
		_w2501_,
		_w2502_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2285 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[9]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2503_
	);
	LUT2 #(
		.INIT('h8)
	) name2286 (
		\reg2_reg[9]/NET0131 ,
		_w252_,
		_w2504_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2287 (
		\reg2_reg[9]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2505_
	);
	LUT4 #(
		.INIT('hc808)
	) name2288 (
		\reg2_reg[9]/NET0131 ,
		_w404_,
		_w970_,
		_w2037_,
		_w2506_
	);
	LUT4 #(
		.INIT('hd020)
	) name2289 (
		_w566_,
		_w584_,
		_w970_,
		_w2039_,
		_w2507_
	);
	LUT3 #(
		.INIT('ha8)
	) name2290 (
		_w587_,
		_w2505_,
		_w2507_,
		_w2508_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2291 (
		\reg2_reg[9]/NET0131 ,
		_w518_,
		_w970_,
		_w2040_,
		_w2509_
	);
	LUT4 #(
		.INIT('hc808)
	) name2292 (
		\reg2_reg[9]/NET0131 ,
		_w601_,
		_w970_,
		_w2044_,
		_w2510_
	);
	LUT3 #(
		.INIT('ha8)
	) name2293 (
		\reg2_reg[9]/NET0131 ,
		_w524_,
		_w976_,
		_w2511_
	);
	LUT2 #(
		.INIT('h8)
	) name2294 (
		_w520_,
		_w333_,
		_w2512_
	);
	LUT3 #(
		.INIT('h07)
	) name2295 (
		_w970_,
		_w2364_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('h4)
	) name2296 (
		_w2511_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h4)
	) name2297 (
		_w2510_,
		_w2514_,
		_w2515_
	);
	LUT4 #(
		.INIT('h0100)
	) name2298 (
		_w2506_,
		_w2509_,
		_w2508_,
		_w2515_,
		_w2516_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2299 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2504_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('he)
	) name2300 (
		_w2503_,
		_w2517_,
		_w2518_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2301 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[21]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2519_
	);
	LUT2 #(
		.INIT('h8)
	) name2302 (
		\reg1_reg[21]/NET0131 ,
		_w252_,
		_w2520_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2303 (
		\reg1_reg[21]/NET0131 ,
		_w924_,
		_w959_,
		_w2392_,
		_w2521_
	);
	LUT4 #(
		.INIT('h005d)
	) name2304 (
		_w946_,
		_w2305_,
		_w2308_,
		_w2521_,
		_w2522_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2305 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2520_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('he)
	) name2306 (
		_w2519_,
		_w2523_,
		_w2524_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2307 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[1]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2525_
	);
	LUT2 #(
		.INIT('h8)
	) name2308 (
		\reg2_reg[1]/NET0131 ,
		_w252_,
		_w2526_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2309 (
		_w970_,
		_w1962_,
		_w1966_,
		_w2285_,
		_w2527_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2310 (
		\reg2_reg[1]/NET0131 ,
		_w524_,
		_w976_,
		_w1605_,
		_w2528_
	);
	LUT2 #(
		.INIT('h8)
	) name2311 (
		\reg3_reg[1]/NET0131 ,
		_w520_,
		_w2529_
	);
	LUT4 #(
		.INIT('hc808)
	) name2312 (
		\reg2_reg[1]/NET0131 ,
		_w601_,
		_w970_,
		_w1958_,
		_w2530_
	);
	LUT3 #(
		.INIT('h01)
	) name2313 (
		_w2529_,
		_w2528_,
		_w2530_,
		_w2531_
	);
	LUT4 #(
		.INIT('h1311)
	) name2314 (
		_w254_,
		_w2526_,
		_w2527_,
		_w2531_,
		_w2532_
	);
	LUT3 #(
		.INIT('hce)
	) name2315 (
		\state_reg[0]/NET0131 ,
		_w2525_,
		_w2532_,
		_w2533_
	);
	LUT4 #(
		.INIT('h0020)
	) name2316 (
		_w924_,
		_w949_,
		_w1410_,
		_w2397_,
		_w2534_
	);
	LUT2 #(
		.INIT('h2)
	) name2317 (
		\reg1_reg[0]/NET0131 ,
		_w2534_,
		_w2535_
	);
	LUT3 #(
		.INIT('hf2)
	) name2318 (
		_w1871_,
		_w2463_,
		_w2535_,
		_w2536_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2319 (
		\IR_reg[23]/NET0131 ,
		\reg1_reg[13]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2537_
	);
	LUT2 #(
		.INIT('h8)
	) name2320 (
		\reg1_reg[13]/NET0131 ,
		_w252_,
		_w2538_
	);
	LUT2 #(
		.INIT('h4)
	) name2321 (
		_w442_,
		_w525_,
		_w2539_
	);
	LUT3 #(
		.INIT('h78)
	) name2322 (
		_w370_,
		_w371_,
		_w442_,
		_w2540_
	);
	LUT3 #(
		.INIT('h82)
	) name2323 (
		_w587_,
		_w1289_,
		_w2540_,
		_w2541_
	);
	LUT4 #(
		.INIT('h8a20)
	) name2324 (
		_w518_,
		_w1271_,
		_w1273_,
		_w2540_,
		_w2542_
	);
	LUT3 #(
		.INIT('h13)
	) name2325 (
		_w423_,
		_w442_,
		_w1027_,
		_w2543_
	);
	LUT2 #(
		.INIT('h4)
	) name2326 (
		_w596_,
		_w601_,
		_w2544_
	);
	LUT2 #(
		.INIT('h4)
	) name2327 (
		_w2543_,
		_w2544_,
		_w2545_
	);
	LUT4 #(
		.INIT('h0001)
	) name2328 (
		_w2539_,
		_w2542_,
		_w2541_,
		_w2545_,
		_w2546_
	);
	LUT4 #(
		.INIT('h08f7)
	) name2329 (
		_w339_,
		_w356_,
		_w372_,
		_w367_,
		_w2547_
	);
	LUT4 #(
		.INIT('h80d0)
	) name2330 (
		_w266_,
		_w343_,
		_w946_,
		_w2547_,
		_w2548_
	);
	LUT4 #(
		.INIT('h5501)
	) name2331 (
		\reg1_reg[13]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2549_
	);
	LUT2 #(
		.INIT('h2)
	) name2332 (
		_w404_,
		_w2549_,
		_w2550_
	);
	LUT4 #(
		.INIT('h4644)
	) name2333 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w2551_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2334 (
		_w256_,
		_w258_,
		_w261_,
		_w2551_,
		_w2552_
	);
	LUT3 #(
		.INIT('ha2)
	) name2335 (
		\reg1_reg[13]/NET0131 ,
		_w924_,
		_w2552_,
		_w2553_
	);
	LUT3 #(
		.INIT('h0b)
	) name2336 (
		_w2548_,
		_w2550_,
		_w2553_,
		_w2554_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2337 (
		_w254_,
		_w946_,
		_w2546_,
		_w2554_,
		_w2555_
	);
	LUT4 #(
		.INIT('heeec)
	) name2338 (
		\state_reg[0]/NET0131 ,
		_w2537_,
		_w2538_,
		_w2555_,
		_w2556_
	);
	LUT3 #(
		.INIT('ha2)
	) name2339 (
		_w404_,
		_w917_,
		_w2459_,
		_w2557_
	);
	LUT4 #(
		.INIT('h1540)
	) name2340 (
		_w515_,
		_w282_,
		_w283_,
		_w493_,
		_w2558_
	);
	LUT4 #(
		.INIT('hb9bb)
	) name2341 (
		_w401_,
		_w398_,
		_w399_,
		_w403_,
		_w2559_
	);
	LUT3 #(
		.INIT('hd0)
	) name2342 (
		_w917_,
		_w2558_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name2343 (
		\reg0_reg[0]/NET0131 ,
		_w924_,
		_w2561_
	);
	LUT4 #(
		.INIT('h8088)
	) name2344 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w493_,
		_w905_,
		_w2562_
	);
	LUT2 #(
		.INIT('h4)
	) name2345 (
		_w2561_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h4)
	) name2346 (
		_w2560_,
		_w2563_,
		_w2564_
	);
	LUT3 #(
		.INIT('h15)
	) name2347 (
		\reg0_reg[0]/NET0131 ,
		_w917_,
		_w1410_,
		_w2565_
	);
	LUT3 #(
		.INIT('h0b)
	) name2348 (
		_w2557_,
		_w2564_,
		_w2565_,
		_w2566_
	);
	LUT4 #(
		.INIT('h0100)
	) name2349 (
		_w524_,
		_w990_,
		_w1237_,
		_w1410_,
		_w2567_
	);
	LUT2 #(
		.INIT('h2)
	) name2350 (
		\reg2_reg[0]/NET0131 ,
		_w2567_,
		_w2568_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name2351 (
		_w404_,
		_w970_,
		_w2458_,
		_w2459_,
		_w2569_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		\reg3_reg[0]/NET0131 ,
		_w520_,
		_w2570_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2353 (
		\reg2_reg[0]/NET0131 ,
		_w517_,
		_w970_,
		_w2461_,
		_w2571_
	);
	LUT2 #(
		.INIT('h1)
	) name2354 (
		_w2570_,
		_w2571_,
		_w2572_
	);
	LUT4 #(
		.INIT('hecee)
	) name2355 (
		_w1410_,
		_w2568_,
		_w2569_,
		_w2572_,
		_w2573_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2356 (
		\IR_reg[23]/NET0131 ,
		\reg2_reg[13]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2574_
	);
	LUT2 #(
		.INIT('h8)
	) name2357 (
		\reg2_reg[13]/NET0131 ,
		_w252_,
		_w2575_
	);
	LUT4 #(
		.INIT('h7020)
	) name2358 (
		_w266_,
		_w343_,
		_w404_,
		_w2547_,
		_w2576_
	);
	LUT4 #(
		.INIT('h0001)
	) name2359 (
		_w2542_,
		_w2541_,
		_w2545_,
		_w2576_,
		_w2577_
	);
	LUT2 #(
		.INIT('h8)
	) name2360 (
		_w520_,
		_w369_,
		_w2578_
	);
	LUT4 #(
		.INIT('h0001)
	) name2361 (
		_w524_,
		_w976_,
		_w991_,
		_w1605_,
		_w2579_
	);
	LUT3 #(
		.INIT('h31)
	) name2362 (
		\reg2_reg[13]/NET0131 ,
		_w2578_,
		_w2579_,
		_w2580_
	);
	LUT4 #(
		.INIT('h7500)
	) name2363 (
		_w970_,
		_w2539_,
		_w2577_,
		_w2580_,
		_w2581_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2364 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w2575_,
		_w2581_,
		_w2582_
	);
	LUT2 #(
		.INIT('he)
	) name2365 (
		_w2574_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h2)
	) name2366 (
		\reg0_reg[13]/NET0131 ,
		_w2312_,
		_w2584_
	);
	LUT4 #(
		.INIT('hff8a)
	) name2367 (
		_w1781_,
		_w2539_,
		_w2577_,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h1)
	) name2368 (
		\reg3_reg[2]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2586_
	);
	LUT2 #(
		.INIT('h2)
	) name2369 (
		_w266_,
		_w407_,
		_w2587_
	);
	LUT2 #(
		.INIT('h8)
	) name2370 (
		\IR_reg[0]/NET0131 ,
		\reg1_reg[0]/NET0131 ,
		_w2588_
	);
	LUT2 #(
		.INIT('h6)
	) name2371 (
		\IR_reg[0]/NET0131 ,
		\reg1_reg[0]/NET0131 ,
		_w2589_
	);
	LUT2 #(
		.INIT('h8)
	) name2372 (
		_w266_,
		_w407_,
		_w2590_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		\IR_reg[0]/NET0131 ,
		\reg2_reg[0]/NET0131 ,
		_w2591_
	);
	LUT2 #(
		.INIT('h6)
	) name2374 (
		\IR_reg[0]/NET0131 ,
		\reg2_reg[0]/NET0131 ,
		_w2592_
	);
	LUT4 #(
		.INIT('h57df)
	) name2375 (
		_w266_,
		_w407_,
		_w2589_,
		_w2592_,
		_w2593_
	);
	LUT4 #(
		.INIT('h8882)
	) name2376 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[28]/NET0131 ,
		_w238_,
		_w265_,
		_w2594_
	);
	LUT3 #(
		.INIT('h08)
	) name2377 (
		_w241_,
		_w250_,
		_w2594_,
		_w2595_
	);
	LUT3 #(
		.INIT('h15)
	) name2378 (
		\addr[2]_pad ,
		_w241_,
		_w250_,
		_w2596_
	);
	LUT4 #(
		.INIT('h153f)
	) name2379 (
		_w516_,
		_w2593_,
		_w2595_,
		_w2596_,
		_w2597_
	);
	LUT4 #(
		.INIT('h0900)
	) name2380 (
		\IR_reg[23]/NET0131 ,
		_w236_,
		_w401_,
		_w398_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		_w252_,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h9)
	) name2382 (
		\reg2_reg[2]/NET0131 ,
		_w496_,
		_w2600_
	);
	LUT3 #(
		.INIT('he8)
	) name2383 (
		\reg2_reg[1]/NET0131 ,
		_w490_,
		_w2591_,
		_w2601_
	);
	LUT2 #(
		.INIT('h6)
	) name2384 (
		_w2600_,
		_w2601_,
		_w2602_
	);
	LUT4 #(
		.INIT('h73fb)
	) name2385 (
		_w266_,
		_w407_,
		_w496_,
		_w2602_,
		_w2603_
	);
	LUT2 #(
		.INIT('h9)
	) name2386 (
		\reg1_reg[2]/NET0131 ,
		_w496_,
		_w2604_
	);
	LUT3 #(
		.INIT('he8)
	) name2387 (
		\reg1_reg[1]/NET0131 ,
		_w490_,
		_w2588_,
		_w2605_
	);
	LUT2 #(
		.INIT('h6)
	) name2388 (
		_w2604_,
		_w2605_,
		_w2606_
	);
	LUT4 #(
		.INIT('hf1fd)
	) name2389 (
		\addr[2]_pad ,
		_w266_,
		_w407_,
		_w2606_,
		_w2607_
	);
	LUT4 #(
		.INIT('h1000)
	) name2390 (
		_w252_,
		_w2598_,
		_w2603_,
		_w2607_,
		_w2608_
	);
	LUT4 #(
		.INIT('haa02)
	) name2391 (
		\state_reg[0]/NET0131 ,
		_w237_,
		_w2597_,
		_w2608_,
		_w2609_
	);
	LUT2 #(
		.INIT('h1)
	) name2392 (
		_w2586_,
		_w2609_,
		_w2610_
	);
	LUT3 #(
		.INIT('h15)
	) name2393 (
		\addr[4]_pad ,
		_w241_,
		_w250_,
		_w2611_
	);
	LUT4 #(
		.INIT('h153f)
	) name2394 (
		_w516_,
		_w2593_,
		_w2595_,
		_w2611_,
		_w2612_
	);
	LUT4 #(
		.INIT('h3c96)
	) name2395 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		\reg2_reg[4]/NET0131 ,
		_w227_,
		_w2613_
	);
	LUT3 #(
		.INIT('h12)
	) name2396 (
		\IR_reg[3]/NET0131 ,
		\reg2_reg[3]/NET0131 ,
		_w500_,
		_w2614_
	);
	LUT3 #(
		.INIT('h84)
	) name2397 (
		\IR_reg[3]/NET0131 ,
		\reg2_reg[3]/NET0131 ,
		_w500_,
		_w2615_
	);
	LUT4 #(
		.INIT('h004d)
	) name2398 (
		\reg2_reg[2]/NET0131 ,
		_w496_,
		_w2601_,
		_w2615_,
		_w2616_
	);
	LUT3 #(
		.INIT('h02)
	) name2399 (
		_w2613_,
		_w2614_,
		_w2616_,
		_w2617_
	);
	LUT3 #(
		.INIT('h54)
	) name2400 (
		_w2613_,
		_w2614_,
		_w2616_,
		_w2618_
	);
	LUT4 #(
		.INIT('h0008)
	) name2401 (
		_w266_,
		_w407_,
		_w2618_,
		_w2617_,
		_w2619_
	);
	LUT4 #(
		.INIT('h3c96)
	) name2402 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		\reg1_reg[4]/NET0131 ,
		_w227_,
		_w2620_
	);
	LUT3 #(
		.INIT('h12)
	) name2403 (
		\IR_reg[3]/NET0131 ,
		\reg1_reg[3]/NET0131 ,
		_w500_,
		_w2621_
	);
	LUT3 #(
		.INIT('h84)
	) name2404 (
		\IR_reg[3]/NET0131 ,
		\reg1_reg[3]/NET0131 ,
		_w500_,
		_w2622_
	);
	LUT4 #(
		.INIT('h004d)
	) name2405 (
		\reg1_reg[2]/NET0131 ,
		_w496_,
		_w2605_,
		_w2622_,
		_w2623_
	);
	LUT3 #(
		.INIT('h02)
	) name2406 (
		_w2620_,
		_w2621_,
		_w2623_,
		_w2624_
	);
	LUT3 #(
		.INIT('h54)
	) name2407 (
		_w2620_,
		_w2621_,
		_w2623_,
		_w2625_
	);
	LUT4 #(
		.INIT('h0002)
	) name2408 (
		_w266_,
		_w407_,
		_w2625_,
		_w2624_,
		_w2626_
	);
	LUT4 #(
		.INIT('hfdcd)
	) name2409 (
		\addr[4]_pad ,
		_w266_,
		_w407_,
		_w487_,
		_w2627_
	);
	LUT3 #(
		.INIT('h10)
	) name2410 (
		_w2626_,
		_w2619_,
		_w2627_,
		_w2628_
	);
	LUT4 #(
		.INIT('h32fa)
	) name2411 (
		_w237_,
		_w2599_,
		_w2612_,
		_w2628_,
		_w2629_
	);
	LUT3 #(
		.INIT('he2)
	) name2412 (
		\reg3_reg[4]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2629_,
		_w2630_
	);
	LUT3 #(
		.INIT('h10)
	) name2413 (
		\addr[12]_pad ,
		_w401_,
		_w398_,
		_w2631_
	);
	LUT4 #(
		.INIT('h3313)
	) name2414 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2631_,
		_w2632_
	);
	LUT4 #(
		.INIT('h4448)
	) name2415 (
		\IR_reg[12]/NET0131 ,
		\reg1_reg[12]/NET0131 ,
		_w420_,
		_w421_,
		_w2633_
	);
	LUT4 #(
		.INIT('h2221)
	) name2416 (
		\IR_reg[12]/NET0131 ,
		\reg1_reg[12]/NET0131 ,
		_w420_,
		_w421_,
		_w2634_
	);
	LUT4 #(
		.INIT('h9996)
	) name2417 (
		\IR_reg[12]/NET0131 ,
		\reg1_reg[12]/NET0131 ,
		_w420_,
		_w421_,
		_w2635_
	);
	LUT2 #(
		.INIT('h8)
	) name2418 (
		\reg1_reg[11]/NET0131 ,
		_w417_,
		_w2636_
	);
	LUT2 #(
		.INIT('h1)
	) name2419 (
		\reg1_reg[10]/NET0131 ,
		_w426_,
		_w2637_
	);
	LUT4 #(
		.INIT('h0309)
	) name2420 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		\reg1_reg[9]/NET0131 ,
		_w415_,
		_w2638_
	);
	LUT3 #(
		.INIT('h84)
	) name2421 (
		\IR_reg[7]/NET0131 ,
		\reg1_reg[7]/NET0131 ,
		_w465_,
		_w2639_
	);
	LUT3 #(
		.INIT('h12)
	) name2422 (
		\IR_reg[6]/NET0131 ,
		\reg1_reg[6]/NET0131 ,
		_w473_,
		_w2640_
	);
	LUT3 #(
		.INIT('h84)
	) name2423 (
		\IR_reg[6]/NET0131 ,
		\reg1_reg[6]/NET0131 ,
		_w473_,
		_w2641_
	);
	LUT4 #(
		.INIT('h222b)
	) name2424 (
		\reg1_reg[4]/NET0131 ,
		_w487_,
		_w2621_,
		_w2623_,
		_w2642_
	);
	LUT4 #(
		.INIT('h0107)
	) name2425 (
		\reg1_reg[5]/NET0131 ,
		_w478_,
		_w2641_,
		_w2642_,
		_w2643_
	);
	LUT3 #(
		.INIT('h21)
	) name2426 (
		\IR_reg[8]/NET0131 ,
		\reg1_reg[8]/NET0131 ,
		_w420_,
		_w2644_
	);
	LUT3 #(
		.INIT('h12)
	) name2427 (
		\IR_reg[7]/NET0131 ,
		\reg1_reg[7]/NET0131 ,
		_w465_,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name2428 (
		_w2644_,
		_w2645_,
		_w2646_
	);
	LUT4 #(
		.INIT('hab00)
	) name2429 (
		_w2639_,
		_w2640_,
		_w2643_,
		_w2646_,
		_w2647_
	);
	LUT4 #(
		.INIT('hc060)
	) name2430 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		\reg1_reg[9]/NET0131 ,
		_w415_,
		_w2648_
	);
	LUT3 #(
		.INIT('h48)
	) name2431 (
		\IR_reg[8]/NET0131 ,
		\reg1_reg[8]/NET0131 ,
		_w420_,
		_w2649_
	);
	LUT2 #(
		.INIT('h1)
	) name2432 (
		_w2648_,
		_w2649_,
		_w2650_
	);
	LUT3 #(
		.INIT('h45)
	) name2433 (
		_w2638_,
		_w2647_,
		_w2650_,
		_w2651_
	);
	LUT2 #(
		.INIT('h8)
	) name2434 (
		\reg1_reg[10]/NET0131 ,
		_w426_,
		_w2652_
	);
	LUT4 #(
		.INIT('h00ba)
	) name2435 (
		_w2638_,
		_w2647_,
		_w2650_,
		_w2652_,
		_w2653_
	);
	LUT4 #(
		.INIT('h888e)
	) name2436 (
		\reg1_reg[11]/NET0131 ,
		_w417_,
		_w2637_,
		_w2653_,
		_w2654_
	);
	LUT3 #(
		.INIT('h28)
	) name2437 (
		_w2587_,
		_w2635_,
		_w2654_,
		_w2655_
	);
	LUT4 #(
		.INIT('h4448)
	) name2438 (
		\IR_reg[12]/NET0131 ,
		\reg2_reg[12]/NET0131 ,
		_w420_,
		_w421_,
		_w2656_
	);
	LUT4 #(
		.INIT('h2221)
	) name2439 (
		\IR_reg[12]/NET0131 ,
		\reg2_reg[12]/NET0131 ,
		_w420_,
		_w421_,
		_w2657_
	);
	LUT4 #(
		.INIT('h9996)
	) name2440 (
		\IR_reg[12]/NET0131 ,
		\reg2_reg[12]/NET0131 ,
		_w420_,
		_w421_,
		_w2658_
	);
	LUT2 #(
		.INIT('h8)
	) name2441 (
		\reg2_reg[11]/NET0131 ,
		_w417_,
		_w2659_
	);
	LUT4 #(
		.INIT('he8c0)
	) name2442 (
		\reg2_reg[10]/NET0131 ,
		\reg2_reg[11]/NET0131 ,
		_w417_,
		_w426_,
		_w2660_
	);
	LUT2 #(
		.INIT('h1)
	) name2443 (
		\reg2_reg[10]/NET0131 ,
		_w426_,
		_w2661_
	);
	LUT4 #(
		.INIT('hfca8)
	) name2444 (
		\reg2_reg[10]/NET0131 ,
		\reg2_reg[11]/NET0131 ,
		_w417_,
		_w426_,
		_w2662_
	);
	LUT4 #(
		.INIT('h0309)
	) name2445 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		\reg2_reg[9]/NET0131 ,
		_w415_,
		_w2663_
	);
	LUT3 #(
		.INIT('h21)
	) name2446 (
		\IR_reg[8]/NET0131 ,
		\reg2_reg[8]/NET0131 ,
		_w420_,
		_w2664_
	);
	LUT3 #(
		.INIT('h12)
	) name2447 (
		\IR_reg[7]/NET0131 ,
		\reg2_reg[7]/NET0131 ,
		_w465_,
		_w2665_
	);
	LUT3 #(
		.INIT('h84)
	) name2448 (
		\IR_reg[7]/NET0131 ,
		\reg2_reg[7]/NET0131 ,
		_w465_,
		_w2666_
	);
	LUT3 #(
		.INIT('h12)
	) name2449 (
		\IR_reg[6]/NET0131 ,
		\reg2_reg[6]/NET0131 ,
		_w473_,
		_w2667_
	);
	LUT3 #(
		.INIT('h84)
	) name2450 (
		\IR_reg[6]/NET0131 ,
		\reg2_reg[6]/NET0131 ,
		_w473_,
		_w2668_
	);
	LUT4 #(
		.INIT('h222b)
	) name2451 (
		\reg2_reg[4]/NET0131 ,
		_w487_,
		_w2614_,
		_w2616_,
		_w2669_
	);
	LUT4 #(
		.INIT('h0107)
	) name2452 (
		\reg2_reg[5]/NET0131 ,
		_w478_,
		_w2668_,
		_w2669_,
		_w2670_
	);
	LUT4 #(
		.INIT('h888e)
	) name2453 (
		\reg2_reg[7]/NET0131 ,
		_w466_,
		_w2667_,
		_w2670_,
		_w2671_
	);
	LUT3 #(
		.INIT('h48)
	) name2454 (
		\IR_reg[8]/NET0131 ,
		\reg2_reg[8]/NET0131 ,
		_w420_,
		_w2672_
	);
	LUT4 #(
		.INIT('hc060)
	) name2455 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		\reg2_reg[9]/NET0131 ,
		_w415_,
		_w2673_
	);
	LUT2 #(
		.INIT('h1)
	) name2456 (
		_w2672_,
		_w2673_,
		_w2674_
	);
	LUT4 #(
		.INIT('h1055)
	) name2457 (
		_w2663_,
		_w2664_,
		_w2671_,
		_w2674_,
		_w2675_
	);
	LUT3 #(
		.INIT('h15)
	) name2458 (
		_w2660_,
		_w2662_,
		_w2675_,
		_w2676_
	);
	LUT3 #(
		.INIT('h40)
	) name2459 (
		_w266_,
		_w407_,
		_w422_,
		_w2677_
	);
	LUT4 #(
		.INIT('h070f)
	) name2460 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w408_,
		_w516_,
		_w2678_
	);
	LUT3 #(
		.INIT('h31)
	) name2461 (
		\addr[12]_pad ,
		_w2677_,
		_w2678_,
		_w2679_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2462 (
		_w2590_,
		_w2658_,
		_w2676_,
		_w2679_,
		_w2680_
	);
	LUT4 #(
		.INIT('hbabb)
	) name2463 (
		_w1062_,
		_w2632_,
		_w2655_,
		_w2680_,
		_w2681_
	);
	LUT3 #(
		.INIT('h10)
	) name2464 (
		\addr[13]_pad ,
		_w401_,
		_w398_,
		_w2682_
	);
	LUT4 #(
		.INIT('h3313)
	) name2465 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2682_,
		_w2683_
	);
	LUT4 #(
		.INIT('hfca8)
	) name2466 (
		\reg1_reg[10]/NET0131 ,
		\reg1_reg[11]/NET0131 ,
		_w417_,
		_w426_,
		_w2684_
	);
	LUT3 #(
		.INIT('h07)
	) name2467 (
		\reg1_reg[11]/NET0131 ,
		_w417_,
		_w2633_,
		_w2685_
	);
	LUT4 #(
		.INIT('h1055)
	) name2468 (
		_w2634_,
		_w2653_,
		_w2684_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h1)
	) name2469 (
		\reg1_reg[13]/NET0131 ,
		_w441_,
		_w2687_
	);
	LUT4 #(
		.INIT('h9060)
	) name2470 (
		\reg1_reg[13]/NET0131 ,
		_w441_,
		_w2587_,
		_w2686_,
		_w2688_
	);
	LUT2 #(
		.INIT('h6)
	) name2471 (
		\reg2_reg[13]/NET0131 ,
		_w441_,
		_w2689_
	);
	LUT2 #(
		.INIT('h1)
	) name2472 (
		_w2664_,
		_w2665_,
		_w2690_
	);
	LUT3 #(
		.INIT('h17)
	) name2473 (
		\reg2_reg[8]/NET0131 ,
		_w469_,
		_w2666_,
		_w2691_
	);
	LUT4 #(
		.INIT('hef00)
	) name2474 (
		_w2667_,
		_w2670_,
		_w2690_,
		_w2691_,
		_w2692_
	);
	LUT3 #(
		.INIT('h07)
	) name2475 (
		\reg2_reg[10]/NET0131 ,
		_w426_,
		_w2673_,
		_w2693_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2476 (
		_w2662_,
		_w2663_,
		_w2692_,
		_w2693_,
		_w2694_
	);
	LUT3 #(
		.INIT('h07)
	) name2477 (
		\reg2_reg[11]/NET0131 ,
		_w417_,
		_w2656_,
		_w2695_
	);
	LUT3 #(
		.INIT('h45)
	) name2478 (
		_w2657_,
		_w2694_,
		_w2695_,
		_w2696_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name2479 (
		\addr[13]_pad ,
		_w266_,
		_w407_,
		_w441_,
		_w2697_
	);
	LUT4 #(
		.INIT('hd700)
	) name2480 (
		_w2590_,
		_w2689_,
		_w2696_,
		_w2697_,
		_w2698_
	);
	LUT4 #(
		.INIT('h8000)
	) name2481 (
		\addr[13]_pad ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w516_,
		_w2699_
	);
	LUT2 #(
		.INIT('h2)
	) name2482 (
		\reg3_reg[13]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2700_
	);
	LUT2 #(
		.INIT('h1)
	) name2483 (
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT4 #(
		.INIT('h45ff)
	) name2484 (
		_w2683_,
		_w2688_,
		_w2698_,
		_w2701_,
		_w2702_
	);
	LUT3 #(
		.INIT('h10)
	) name2485 (
		\addr[14]_pad ,
		_w401_,
		_w398_,
		_w2703_
	);
	LUT4 #(
		.INIT('h3313)
	) name2486 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h2)
	) name2487 (
		\reg1_reg[14]/NET0131 ,
		_w438_,
		_w2705_
	);
	LUT2 #(
		.INIT('h4)
	) name2488 (
		\reg1_reg[14]/NET0131 ,
		_w438_,
		_w2706_
	);
	LUT2 #(
		.INIT('h9)
	) name2489 (
		\reg1_reg[14]/NET0131 ,
		_w438_,
		_w2707_
	);
	LUT3 #(
		.INIT('h07)
	) name2490 (
		\reg1_reg[13]/NET0131 ,
		_w441_,
		_w2633_,
		_w2708_
	);
	LUT4 #(
		.INIT('h040f)
	) name2491 (
		_w2634_,
		_w2654_,
		_w2687_,
		_w2708_,
		_w2709_
	);
	LUT3 #(
		.INIT('h28)
	) name2492 (
		_w2587_,
		_w2707_,
		_w2709_,
		_w2710_
	);
	LUT2 #(
		.INIT('h2)
	) name2493 (
		\reg2_reg[14]/NET0131 ,
		_w438_,
		_w2711_
	);
	LUT2 #(
		.INIT('h4)
	) name2494 (
		\reg2_reg[14]/NET0131 ,
		_w438_,
		_w2712_
	);
	LUT2 #(
		.INIT('h9)
	) name2495 (
		\reg2_reg[14]/NET0131 ,
		_w438_,
		_w2713_
	);
	LUT3 #(
		.INIT('h0e)
	) name2496 (
		\reg2_reg[13]/NET0131 ,
		_w441_,
		_w2657_,
		_w2714_
	);
	LUT4 #(
		.INIT('hea00)
	) name2497 (
		_w2660_,
		_w2662_,
		_w2675_,
		_w2714_,
		_w2715_
	);
	LUT3 #(
		.INIT('h17)
	) name2498 (
		\reg2_reg[13]/NET0131 ,
		_w441_,
		_w2656_,
		_w2716_
	);
	LUT4 #(
		.INIT('h2822)
	) name2499 (
		_w2590_,
		_w2713_,
		_w2715_,
		_w2716_,
		_w2717_
	);
	LUT3 #(
		.INIT('h04)
	) name2500 (
		_w266_,
		_w407_,
		_w438_,
		_w2718_
	);
	LUT3 #(
		.INIT('h0d)
	) name2501 (
		\addr[14]_pad ,
		_w2678_,
		_w2718_,
		_w2719_
	);
	LUT2 #(
		.INIT('h4)
	) name2502 (
		_w2717_,
		_w2719_,
		_w2720_
	);
	LUT4 #(
		.INIT('hbabb)
	) name2503 (
		_w1341_,
		_w2704_,
		_w2710_,
		_w2720_,
		_w2721_
	);
	LUT3 #(
		.INIT('h10)
	) name2504 (
		\addr[15]_pad ,
		_w401_,
		_w398_,
		_w2722_
	);
	LUT4 #(
		.INIT('h3313)
	) name2505 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2722_,
		_w2723_
	);
	LUT3 #(
		.INIT('h84)
	) name2506 (
		\IR_reg[15]/NET0131 ,
		\reg1_reg[15]/NET0131 ,
		_w447_,
		_w2724_
	);
	LUT3 #(
		.INIT('h12)
	) name2507 (
		\IR_reg[15]/NET0131 ,
		\reg1_reg[15]/NET0131 ,
		_w447_,
		_w2725_
	);
	LUT3 #(
		.INIT('h69)
	) name2508 (
		\IR_reg[15]/NET0131 ,
		\reg1_reg[15]/NET0131 ,
		_w447_,
		_w2726_
	);
	LUT4 #(
		.INIT('h51f3)
	) name2509 (
		\reg1_reg[13]/NET0131 ,
		\reg1_reg[14]/NET0131 ,
		_w438_,
		_w441_,
		_w2727_
	);
	LUT4 #(
		.INIT('h020f)
	) name2510 (
		_w2686_,
		_w2687_,
		_w2706_,
		_w2727_,
		_w2728_
	);
	LUT3 #(
		.INIT('h84)
	) name2511 (
		\IR_reg[15]/NET0131 ,
		\reg2_reg[15]/NET0131 ,
		_w447_,
		_w2729_
	);
	LUT3 #(
		.INIT('h12)
	) name2512 (
		\IR_reg[15]/NET0131 ,
		\reg2_reg[15]/NET0131 ,
		_w447_,
		_w2730_
	);
	LUT3 #(
		.INIT('h69)
	) name2513 (
		\IR_reg[15]/NET0131 ,
		\reg2_reg[15]/NET0131 ,
		_w447_,
		_w2731_
	);
	LUT2 #(
		.INIT('h4)
	) name2514 (
		_w2712_,
		_w2714_,
		_w2732_
	);
	LUT4 #(
		.INIT('h71f3)
	) name2515 (
		\reg2_reg[13]/NET0131 ,
		\reg2_reg[14]/NET0131 ,
		_w438_,
		_w441_,
		_w2733_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2516 (
		_w2694_,
		_w2695_,
		_w2732_,
		_w2733_,
		_w2734_
	);
	LUT3 #(
		.INIT('h40)
	) name2517 (
		_w266_,
		_w407_,
		_w448_,
		_w2735_
	);
	LUT3 #(
		.INIT('h0d)
	) name2518 (
		\addr[15]_pad ,
		_w2678_,
		_w2735_,
		_w2736_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2519 (
		_w2590_,
		_w2731_,
		_w2734_,
		_w2736_,
		_w2737_
	);
	LUT4 #(
		.INIT('hd700)
	) name2520 (
		_w2587_,
		_w2726_,
		_w2728_,
		_w2737_,
		_w2738_
	);
	LUT3 #(
		.INIT('hab)
	) name2521 (
		_w1019_,
		_w2723_,
		_w2738_,
		_w2739_
	);
	LUT3 #(
		.INIT('h10)
	) name2522 (
		\addr[17]_pad ,
		_w401_,
		_w398_,
		_w2740_
	);
	LUT4 #(
		.INIT('h3313)
	) name2523 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2740_,
		_w2741_
	);
	LUT4 #(
		.INIT('h4448)
	) name2524 (
		\IR_reg[17]/NET0131 ,
		\reg1_reg[17]/NET0131 ,
		_w238_,
		_w409_,
		_w2742_
	);
	LUT4 #(
		.INIT('h2221)
	) name2525 (
		\IR_reg[17]/NET0131 ,
		\reg1_reg[17]/NET0131 ,
		_w238_,
		_w409_,
		_w2743_
	);
	LUT4 #(
		.INIT('h9996)
	) name2526 (
		\IR_reg[17]/NET0131 ,
		\reg1_reg[17]/NET0131 ,
		_w238_,
		_w409_,
		_w2744_
	);
	LUT4 #(
		.INIT('h0509)
	) name2527 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[16]/NET0131 ,
		_w233_,
		_w2745_
	);
	LUT4 #(
		.INIT('ha060)
	) name2528 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[16]/NET0131 ,
		_w233_,
		_w2746_
	);
	LUT2 #(
		.INIT('h1)
	) name2529 (
		_w2724_,
		_w2746_,
		_w2747_
	);
	LUT4 #(
		.INIT('h040f)
	) name2530 (
		_w2725_,
		_w2728_,
		_w2745_,
		_w2747_,
		_w2748_
	);
	LUT4 #(
		.INIT('h4448)
	) name2531 (
		\IR_reg[17]/NET0131 ,
		\reg2_reg[17]/NET0131 ,
		_w238_,
		_w409_,
		_w2749_
	);
	LUT4 #(
		.INIT('h2221)
	) name2532 (
		\IR_reg[17]/NET0131 ,
		\reg2_reg[17]/NET0131 ,
		_w238_,
		_w409_,
		_w2750_
	);
	LUT4 #(
		.INIT('h9996)
	) name2533 (
		\IR_reg[17]/NET0131 ,
		\reg2_reg[17]/NET0131 ,
		_w238_,
		_w409_,
		_w2751_
	);
	LUT4 #(
		.INIT('h0509)
	) name2534 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[16]/NET0131 ,
		_w233_,
		_w2752_
	);
	LUT4 #(
		.INIT('ha060)
	) name2535 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[16]/NET0131 ,
		_w233_,
		_w2753_
	);
	LUT2 #(
		.INIT('h1)
	) name2536 (
		_w2729_,
		_w2753_,
		_w2754_
	);
	LUT4 #(
		.INIT('h010f)
	) name2537 (
		_w2730_,
		_w2734_,
		_w2752_,
		_w2754_,
		_w2755_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name2538 (
		\addr[17]_pad ,
		_w266_,
		_w407_,
		_w410_,
		_w2756_
	);
	LUT4 #(
		.INIT('hd700)
	) name2539 (
		_w2590_,
		_w2751_,
		_w2755_,
		_w2756_,
		_w2757_
	);
	LUT4 #(
		.INIT('hd700)
	) name2540 (
		_w2587_,
		_w2744_,
		_w2748_,
		_w2757_,
		_w2758_
	);
	LUT4 #(
		.INIT('h8000)
	) name2541 (
		\addr[17]_pad ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w516_,
		_w2759_
	);
	LUT2 #(
		.INIT('h1)
	) name2542 (
		_w605_,
		_w2759_,
		_w2760_
	);
	LUT3 #(
		.INIT('h1f)
	) name2543 (
		_w2741_,
		_w2758_,
		_w2760_,
		_w2761_
	);
	LUT3 #(
		.INIT('h10)
	) name2544 (
		\addr[18]_pad ,
		_w401_,
		_w398_,
		_w2762_
	);
	LUT4 #(
		.INIT('h3313)
	) name2545 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2762_,
		_w2763_
	);
	LUT4 #(
		.INIT('h4448)
	) name2546 (
		\IR_reg[18]/NET0131 ,
		\reg1_reg[18]/NET0131 ,
		_w238_,
		_w676_,
		_w2764_
	);
	LUT4 #(
		.INIT('h2221)
	) name2547 (
		\IR_reg[18]/NET0131 ,
		\reg1_reg[18]/NET0131 ,
		_w238_,
		_w676_,
		_w2765_
	);
	LUT4 #(
		.INIT('h9996)
	) name2548 (
		\IR_reg[18]/NET0131 ,
		\reg1_reg[18]/NET0131 ,
		_w238_,
		_w676_,
		_w2766_
	);
	LUT2 #(
		.INIT('h1)
	) name2549 (
		_w2705_,
		_w2724_,
		_w2767_
	);
	LUT4 #(
		.INIT('h040f)
	) name2550 (
		_w2706_,
		_w2709_,
		_w2725_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h1)
	) name2551 (
		_w2742_,
		_w2746_,
		_w2769_
	);
	LUT4 #(
		.INIT('h1055)
	) name2552 (
		_w2743_,
		_w2745_,
		_w2768_,
		_w2769_,
		_w2770_
	);
	LUT3 #(
		.INIT('h28)
	) name2553 (
		_w2587_,
		_w2766_,
		_w2770_,
		_w2771_
	);
	LUT4 #(
		.INIT('h4448)
	) name2554 (
		\IR_reg[18]/NET0131 ,
		\reg2_reg[18]/NET0131 ,
		_w238_,
		_w676_,
		_w2772_
	);
	LUT4 #(
		.INIT('h2221)
	) name2555 (
		\IR_reg[18]/NET0131 ,
		\reg2_reg[18]/NET0131 ,
		_w238_,
		_w676_,
		_w2773_
	);
	LUT4 #(
		.INIT('h9996)
	) name2556 (
		\IR_reg[18]/NET0131 ,
		\reg2_reg[18]/NET0131 ,
		_w238_,
		_w676_,
		_w2774_
	);
	LUT2 #(
		.INIT('h1)
	) name2557 (
		_w2711_,
		_w2729_,
		_w2775_
	);
	LUT4 #(
		.INIT('hba00)
	) name2558 (
		_w2712_,
		_w2715_,
		_w2716_,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('h1)
	) name2559 (
		_w2749_,
		_w2753_,
		_w2777_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2560 (
		_w2730_,
		_w2752_,
		_w2776_,
		_w2777_,
		_w2778_
	);
	LUT4 #(
		.INIT('ha082)
	) name2561 (
		_w2590_,
		_w2750_,
		_w2774_,
		_w2778_,
		_w2779_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name2562 (
		\addr[18]_pad ,
		_w266_,
		_w407_,
		_w677_,
		_w2780_
	);
	LUT2 #(
		.INIT('h4)
	) name2563 (
		_w2779_,
		_w2780_,
		_w2781_
	);
	LUT4 #(
		.INIT('h8000)
	) name2564 (
		\addr[18]_pad ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w516_,
		_w2782_
	);
	LUT2 #(
		.INIT('h1)
	) name2565 (
		_w1659_,
		_w2782_,
		_w2783_
	);
	LUT4 #(
		.INIT('h45ff)
	) name2566 (
		_w2763_,
		_w2771_,
		_w2781_,
		_w2783_,
		_w2784_
	);
	LUT3 #(
		.INIT('h10)
	) name2567 (
		\addr[19]_pad ,
		_w401_,
		_w398_,
		_w2785_
	);
	LUT4 #(
		.INIT('h3313)
	) name2568 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2785_,
		_w2786_
	);
	LUT2 #(
		.INIT('h1)
	) name2569 (
		_w2743_,
		_w2765_,
		_w2787_
	);
	LUT4 #(
		.INIT('h010f)
	) name2570 (
		_w2742_,
		_w2748_,
		_w2764_,
		_w2787_,
		_w2788_
	);
	LUT4 #(
		.INIT('h9996)
	) name2571 (
		\IR_reg[19]/NET0131 ,
		\reg1_reg[19]/NET0131 ,
		_w238_,
		_w402_,
		_w2789_
	);
	LUT3 #(
		.INIT('h82)
	) name2572 (
		_w2587_,
		_w2788_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h1)
	) name2573 (
		_w2749_,
		_w2772_,
		_w2791_
	);
	LUT4 #(
		.INIT('h040f)
	) name2574 (
		_w2750_,
		_w2755_,
		_w2773_,
		_w2791_,
		_w2792_
	);
	LUT4 #(
		.INIT('h9060)
	) name2575 (
		\reg2_reg[19]/NET0131 ,
		_w403_,
		_w2590_,
		_w2792_,
		_w2793_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2576 (
		\addr[19]_pad ,
		_w403_,
		_w266_,
		_w407_,
		_w2794_
	);
	LUT2 #(
		.INIT('h4)
	) name2577 (
		_w2793_,
		_w2794_,
		_w2795_
	);
	LUT4 #(
		.INIT('h8000)
	) name2578 (
		\addr[19]_pad ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w516_,
		_w2796_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w1087_,
		_w2796_,
		_w2797_
	);
	LUT4 #(
		.INIT('h45ff)
	) name2580 (
		_w2786_,
		_w2790_,
		_w2795_,
		_w2797_,
		_w2798_
	);
	LUT2 #(
		.INIT('h2)
	) name2581 (
		\reg3_reg[1]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2799_
	);
	LUT3 #(
		.INIT('h10)
	) name2582 (
		\addr[1]_pad ,
		_w401_,
		_w398_,
		_w2800_
	);
	LUT4 #(
		.INIT('h3313)
	) name2583 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2800_,
		_w2801_
	);
	LUT4 #(
		.INIT('h936c)
	) name2584 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[1]/NET0131 ,
		_w2802_
	);
	LUT2 #(
		.INIT('h6)
	) name2585 (
		_w2591_,
		_w2802_,
		_w2803_
	);
	LUT3 #(
		.INIT('h80)
	) name2586 (
		_w266_,
		_w407_,
		_w2803_,
		_w2804_
	);
	LUT4 #(
		.INIT('h936c)
	) name2587 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[1]/NET0131 ,
		_w2805_
	);
	LUT2 #(
		.INIT('h6)
	) name2588 (
		_w2588_,
		_w2805_,
		_w2806_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name2589 (
		_w266_,
		_w407_,
		_w490_,
		_w2806_,
		_w2807_
	);
	LUT2 #(
		.INIT('h4)
	) name2590 (
		_w2804_,
		_w2807_,
		_w2808_
	);
	LUT4 #(
		.INIT('h020f)
	) name2591 (
		\addr[1]_pad ,
		_w2678_,
		_w2801_,
		_w2808_,
		_w2809_
	);
	LUT2 #(
		.INIT('he)
	) name2592 (
		_w2799_,
		_w2809_,
		_w2810_
	);
	LUT2 #(
		.INIT('h2)
	) name2593 (
		\reg3_reg[3]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2811_
	);
	LUT3 #(
		.INIT('h10)
	) name2594 (
		\addr[3]_pad ,
		_w401_,
		_w398_,
		_w2812_
	);
	LUT4 #(
		.INIT('h3313)
	) name2595 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2812_,
		_w2813_
	);
	LUT3 #(
		.INIT('h69)
	) name2596 (
		\IR_reg[3]/NET0131 ,
		\reg1_reg[3]/NET0131 ,
		_w500_,
		_w2814_
	);
	LUT4 #(
		.INIT('h4db2)
	) name2597 (
		\reg1_reg[2]/NET0131 ,
		_w496_,
		_w2605_,
		_w2814_,
		_w2815_
	);
	LUT3 #(
		.INIT('h20)
	) name2598 (
		_w266_,
		_w407_,
		_w2815_,
		_w2816_
	);
	LUT3 #(
		.INIT('h69)
	) name2599 (
		\IR_reg[3]/NET0131 ,
		\reg2_reg[3]/NET0131 ,
		_w500_,
		_w2817_
	);
	LUT4 #(
		.INIT('h4db2)
	) name2600 (
		\reg2_reg[2]/NET0131 ,
		_w496_,
		_w2601_,
		_w2817_,
		_w2818_
	);
	LUT4 #(
		.INIT('h37bf)
	) name2601 (
		_w266_,
		_w407_,
		_w501_,
		_w2818_,
		_w2819_
	);
	LUT2 #(
		.INIT('h4)
	) name2602 (
		_w2816_,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('h020f)
	) name2603 (
		\addr[3]_pad ,
		_w2678_,
		_w2813_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('he)
	) name2604 (
		_w2811_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h6)
	) name2605 (
		\reg2_reg[5]/NET0131 ,
		_w478_,
		_w2823_
	);
	LUT4 #(
		.INIT('h0880)
	) name2606 (
		_w266_,
		_w407_,
		_w2669_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h6)
	) name2607 (
		\reg1_reg[5]/NET0131 ,
		_w478_,
		_w2825_
	);
	LUT4 #(
		.INIT('h0220)
	) name2608 (
		_w266_,
		_w407_,
		_w2642_,
		_w2825_,
		_w2826_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name2609 (
		\addr[5]_pad ,
		_w266_,
		_w407_,
		_w478_,
		_w2827_
	);
	LUT3 #(
		.INIT('h10)
	) name2610 (
		_w2826_,
		_w2824_,
		_w2827_,
		_w2828_
	);
	LUT3 #(
		.INIT('h02)
	) name2611 (
		\state_reg[0]/NET0131 ,
		_w252_,
		_w2598_,
		_w2829_
	);
	LUT4 #(
		.INIT('h8000)
	) name2612 (
		\addr[5]_pad ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w516_,
		_w2830_
	);
	LUT2 #(
		.INIT('h2)
	) name2613 (
		\reg3_reg[5]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2831_
	);
	LUT4 #(
		.INIT('hefee)
	) name2614 (
		_w2830_,
		_w2831_,
		_w2828_,
		_w2829_,
		_w2832_
	);
	LUT3 #(
		.INIT('h10)
	) name2615 (
		\addr[6]_pad ,
		_w401_,
		_w398_,
		_w2833_
	);
	LUT4 #(
		.INIT('h3313)
	) name2616 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2833_,
		_w2834_
	);
	LUT3 #(
		.INIT('h40)
	) name2617 (
		_w266_,
		_w407_,
		_w474_,
		_w2835_
	);
	LUT3 #(
		.INIT('h0d)
	) name2618 (
		\addr[6]_pad ,
		_w2678_,
		_w2835_,
		_w2836_
	);
	LUT3 #(
		.INIT('h69)
	) name2619 (
		\IR_reg[6]/NET0131 ,
		\reg1_reg[6]/NET0131 ,
		_w473_,
		_w2837_
	);
	LUT4 #(
		.INIT('he800)
	) name2620 (
		\reg1_reg[5]/NET0131 ,
		_w478_,
		_w2642_,
		_w2837_,
		_w2838_
	);
	LUT4 #(
		.INIT('h0017)
	) name2621 (
		\reg1_reg[5]/NET0131 ,
		_w478_,
		_w2642_,
		_w2837_,
		_w2839_
	);
	LUT3 #(
		.INIT('h02)
	) name2622 (
		_w2587_,
		_w2839_,
		_w2838_,
		_w2840_
	);
	LUT3 #(
		.INIT('h69)
	) name2623 (
		\IR_reg[6]/NET0131 ,
		\reg2_reg[6]/NET0131 ,
		_w473_,
		_w2841_
	);
	LUT4 #(
		.INIT('he800)
	) name2624 (
		\reg2_reg[5]/NET0131 ,
		_w478_,
		_w2669_,
		_w2841_,
		_w2842_
	);
	LUT4 #(
		.INIT('h0017)
	) name2625 (
		\reg2_reg[5]/NET0131 ,
		_w478_,
		_w2669_,
		_w2841_,
		_w2843_
	);
	LUT3 #(
		.INIT('h02)
	) name2626 (
		_w2590_,
		_w2843_,
		_w2842_,
		_w2844_
	);
	LUT2 #(
		.INIT('h1)
	) name2627 (
		_w2840_,
		_w2844_,
		_w2845_
	);
	LUT4 #(
		.INIT('habbb)
	) name2628 (
		_w2013_,
		_w2834_,
		_w2836_,
		_w2845_,
		_w2846_
	);
	LUT3 #(
		.INIT('h10)
	) name2629 (
		\addr[7]_pad ,
		_w401_,
		_w398_,
		_w2847_
	);
	LUT4 #(
		.INIT('h3313)
	) name2630 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2847_,
		_w2848_
	);
	LUT3 #(
		.INIT('h69)
	) name2631 (
		\IR_reg[7]/NET0131 ,
		\reg1_reg[7]/NET0131 ,
		_w465_,
		_w2849_
	);
	LUT4 #(
		.INIT('ha802)
	) name2632 (
		_w2587_,
		_w2640_,
		_w2643_,
		_w2849_,
		_w2850_
	);
	LUT3 #(
		.INIT('h69)
	) name2633 (
		\IR_reg[7]/NET0131 ,
		\reg2_reg[7]/NET0131 ,
		_w465_,
		_w2851_
	);
	LUT4 #(
		.INIT('ha802)
	) name2634 (
		_w2590_,
		_w2667_,
		_w2670_,
		_w2851_,
		_w2852_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name2635 (
		\addr[7]_pad ,
		_w266_,
		_w407_,
		_w466_,
		_w2853_
	);
	LUT4 #(
		.INIT('h5455)
	) name2636 (
		_w2848_,
		_w2852_,
		_w2850_,
		_w2853_,
		_w2854_
	);
	LUT4 #(
		.INIT('h8000)
	) name2637 (
		\addr[7]_pad ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w516_,
		_w2855_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		_w1384_,
		_w2855_,
		_w2856_
	);
	LUT2 #(
		.INIT('hb)
	) name2639 (
		_w2854_,
		_w2856_,
		_w2857_
	);
	LUT3 #(
		.INIT('h10)
	) name2640 (
		\addr[8]_pad ,
		_w401_,
		_w398_,
		_w2858_
	);
	LUT4 #(
		.INIT('h3313)
	) name2641 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('h888e)
	) name2642 (
		\reg1_reg[7]/NET0131 ,
		_w466_,
		_w2640_,
		_w2643_,
		_w2860_
	);
	LUT3 #(
		.INIT('h96)
	) name2643 (
		\IR_reg[8]/NET0131 ,
		\reg1_reg[8]/NET0131 ,
		_w420_,
		_w2861_
	);
	LUT3 #(
		.INIT('h28)
	) name2644 (
		_w2587_,
		_w2860_,
		_w2861_,
		_w2862_
	);
	LUT3 #(
		.INIT('h96)
	) name2645 (
		\IR_reg[8]/NET0131 ,
		\reg2_reg[8]/NET0131 ,
		_w420_,
		_w2863_
	);
	LUT3 #(
		.INIT('h28)
	) name2646 (
		_w2590_,
		_w2671_,
		_w2863_,
		_w2864_
	);
	LUT3 #(
		.INIT('h40)
	) name2647 (
		_w266_,
		_w407_,
		_w469_,
		_w2865_
	);
	LUT3 #(
		.INIT('h0d)
	) name2648 (
		\addr[8]_pad ,
		_w2678_,
		_w2865_,
		_w2866_
	);
	LUT4 #(
		.INIT('h5455)
	) name2649 (
		_w2859_,
		_w2864_,
		_w2862_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('he)
	) name2650 (
		_w2030_,
		_w2867_,
		_w2868_
	);
	LUT3 #(
		.INIT('h10)
	) name2651 (
		\addr[9]_pad ,
		_w401_,
		_w398_,
		_w2869_
	);
	LUT4 #(
		.INIT('h3313)
	) name2652 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2869_,
		_w2870_
	);
	LUT4 #(
		.INIT('h3c96)
	) name2653 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		\reg1_reg[9]/NET0131 ,
		_w415_,
		_w2871_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2654 (
		_w2587_,
		_w2647_,
		_w2649_,
		_w2871_,
		_w2872_
	);
	LUT4 #(
		.INIT('h3c96)
	) name2655 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		\reg2_reg[9]/NET0131 ,
		_w415_,
		_w2873_
	);
	LUT3 #(
		.INIT('h82)
	) name2656 (
		_w2590_,
		_w2692_,
		_w2873_,
		_w2874_
	);
	LUT3 #(
		.INIT('h04)
	) name2657 (
		_w266_,
		_w407_,
		_w430_,
		_w2875_
	);
	LUT3 #(
		.INIT('h0d)
	) name2658 (
		\addr[9]_pad ,
		_w2678_,
		_w2875_,
		_w2876_
	);
	LUT4 #(
		.INIT('h5455)
	) name2659 (
		_w2870_,
		_w2872_,
		_w2874_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('he)
	) name2660 (
		_w2052_,
		_w2877_,
		_w2878_
	);
	LUT3 #(
		.INIT('h10)
	) name2661 (
		\addr[11]_pad ,
		_w401_,
		_w398_,
		_w2879_
	);
	LUT4 #(
		.INIT('h3313)
	) name2662 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2879_,
		_w2880_
	);
	LUT3 #(
		.INIT('h10)
	) name2663 (
		_w2636_,
		_w2653_,
		_w2684_,
		_w2881_
	);
	LUT2 #(
		.INIT('h6)
	) name2664 (
		\reg1_reg[11]/NET0131 ,
		_w417_,
		_w2882_
	);
	LUT4 #(
		.INIT('haa02)
	) name2665 (
		_w2587_,
		_w2637_,
		_w2653_,
		_w2882_,
		_w2883_
	);
	LUT2 #(
		.INIT('h4)
	) name2666 (
		_w2881_,
		_w2883_,
		_w2884_
	);
	LUT2 #(
		.INIT('h4)
	) name2667 (
		_w2659_,
		_w2694_,
		_w2885_
	);
	LUT2 #(
		.INIT('h6)
	) name2668 (
		\reg2_reg[11]/NET0131 ,
		_w417_,
		_w2886_
	);
	LUT4 #(
		.INIT('h0155)
	) name2669 (
		_w2661_,
		_w2663_,
		_w2692_,
		_w2693_,
		_w2887_
	);
	LUT3 #(
		.INIT('ha8)
	) name2670 (
		_w2590_,
		_w2886_,
		_w2887_,
		_w2888_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name2671 (
		\addr[11]_pad ,
		_w266_,
		_w407_,
		_w417_,
		_w2889_
	);
	LUT3 #(
		.INIT('hb0)
	) name2672 (
		_w2885_,
		_w2888_,
		_w2889_,
		_w2890_
	);
	LUT4 #(
		.INIT('h8000)
	) name2673 (
		\addr[11]_pad ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w516_,
		_w2891_
	);
	LUT2 #(
		.INIT('h1)
	) name2674 (
		_w1040_,
		_w2891_,
		_w2892_
	);
	LUT4 #(
		.INIT('h45ff)
	) name2675 (
		_w2880_,
		_w2884_,
		_w2890_,
		_w2892_,
		_w2893_
	);
	LUT4 #(
		.INIT('h5557)
	) name2676 (
		\state_reg[0]/NET0131 ,
		_w252_,
		_w408_,
		_w2598_,
		_w2894_
	);
	LUT2 #(
		.INIT('h2)
	) name2677 (
		\reg3_reg[0]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2895_
	);
	LUT3 #(
		.INIT('h10)
	) name2678 (
		\addr[0]_pad ,
		_w401_,
		_w398_,
		_w2896_
	);
	LUT4 #(
		.INIT('h3313)
	) name2679 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h8)
	) name2680 (
		_w407_,
		_w2594_,
		_w2898_
	);
	LUT2 #(
		.INIT('h2)
	) name2681 (
		_w2593_,
		_w2898_,
		_w2899_
	);
	LUT4 #(
		.INIT('h020f)
	) name2682 (
		\addr[0]_pad ,
		_w2678_,
		_w2897_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('he)
	) name2683 (
		_w2895_,
		_w2900_,
		_w2901_
	);
	LUT2 #(
		.INIT('h2)
	) name2684 (
		\reg3_reg[10]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2902_
	);
	LUT3 #(
		.INIT('h10)
	) name2685 (
		\addr[10]_pad ,
		_w401_,
		_w398_,
		_w2903_
	);
	LUT4 #(
		.INIT('h3313)
	) name2686 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h6)
	) name2687 (
		\reg2_reg[10]/NET0131 ,
		_w426_,
		_w2905_
	);
	LUT3 #(
		.INIT('h28)
	) name2688 (
		_w2590_,
		_w2675_,
		_w2905_,
		_w2906_
	);
	LUT2 #(
		.INIT('h6)
	) name2689 (
		\reg1_reg[10]/NET0131 ,
		_w426_,
		_w2907_
	);
	LUT3 #(
		.INIT('h40)
	) name2690 (
		_w266_,
		_w407_,
		_w426_,
		_w2908_
	);
	LUT3 #(
		.INIT('h0d)
	) name2691 (
		\addr[10]_pad ,
		_w2678_,
		_w2908_,
		_w2909_
	);
	LUT4 #(
		.INIT('hd700)
	) name2692 (
		_w2587_,
		_w2651_,
		_w2907_,
		_w2909_,
		_w2910_
	);
	LUT4 #(
		.INIT('hbabb)
	) name2693 (
		_w2902_,
		_w2904_,
		_w2906_,
		_w2910_,
		_w2911_
	);
	LUT3 #(
		.INIT('h10)
	) name2694 (
		\addr[16]_pad ,
		_w401_,
		_w398_,
		_w2912_
	);
	LUT4 #(
		.INIT('h3313)
	) name2695 (
		\state_reg[0]/NET0131 ,
		_w606_,
		_w254_,
		_w2912_,
		_w2913_
	);
	LUT4 #(
		.INIT('h5a96)
	) name2696 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[16]/NET0131 ,
		_w233_,
		_w2914_
	);
	LUT3 #(
		.INIT('h28)
	) name2697 (
		_w2587_,
		_w2768_,
		_w2914_,
		_w2915_
	);
	LUT4 #(
		.INIT('h5a96)
	) name2698 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[16]/NET0131 ,
		_w233_,
		_w2916_
	);
	LUT4 #(
		.INIT('ha802)
	) name2699 (
		_w2590_,
		_w2730_,
		_w2776_,
		_w2916_,
		_w2917_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name2700 (
		\addr[16]_pad ,
		_w266_,
		_w407_,
		_w445_,
		_w2918_
	);
	LUT2 #(
		.INIT('h4)
	) name2701 (
		_w2917_,
		_w2918_,
		_w2919_
	);
	LUT4 #(
		.INIT('h8000)
	) name2702 (
		\addr[16]_pad ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w516_,
		_w2920_
	);
	LUT2 #(
		.INIT('h1)
	) name2703 (
		_w1364_,
		_w2920_,
		_w2921_
	);
	LUT4 #(
		.INIT('h45ff)
	) name2704 (
		_w2913_,
		_w2915_,
		_w2919_,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h8)
	) name2705 (
		\state_reg[0]/NET0131 ,
		_w252_,
		_w2923_
	);
	LUT3 #(
		.INIT('h2a)
	) name2706 (
		\datao[15]_pad ,
		_w241_,
		_w250_,
		_w2924_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2707 (
		_w251_,
		_w376_,
		_w375_,
		_w377_,
		_w2925_
	);
	LUT2 #(
		.INIT('he)
	) name2708 (
		_w2924_,
		_w2925_,
		_w2926_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2709 (
		\datao[28]_pad ,
		_w251_,
		_w734_,
		_w737_,
		_w2927_
	);
	LUT4 #(
		.INIT('h2eee)
	) name2710 (
		\datao[8]_pad ,
		_w251_,
		_w328_,
		_w330_,
		_w2928_
	);
	LUT4 #(
		.INIT('h4448)
	) name2711 (
		\IR_reg[27]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w248_,
		_w406_,
		_w2929_
	);
	LUT2 #(
		.INIT('h2)
	) name2712 (
		\datai[27]_pad ,
		\state_reg[0]/NET0131 ,
		_w2930_
	);
	LUT2 #(
		.INIT('he)
	) name2713 (
		_w2929_,
		_w2930_,
		_w2931_
	);
	LUT4 #(
		.INIT('h4448)
	) name2714 (
		\IR_reg[30]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w244_,
		_w271_,
		_w2932_
	);
	LUT2 #(
		.INIT('h2)
	) name2715 (
		\datai[30]_pad ,
		\state_reg[0]/NET0131 ,
		_w2933_
	);
	LUT2 #(
		.INIT('he)
	) name2716 (
		_w2932_,
		_w2933_,
		_w2934_
	);
	LUT4 #(
		.INIT('h4448)
	) name2717 (
		\IR_reg[28]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w238_,
		_w265_,
		_w2935_
	);
	LUT2 #(
		.INIT('h2)
	) name2718 (
		\datai[28]_pad ,
		\state_reg[0]/NET0131 ,
		_w2936_
	);
	LUT2 #(
		.INIT('he)
	) name2719 (
		_w2935_,
		_w2936_,
		_w2937_
	);
	LUT4 #(
		.INIT('ha060)
	) name2720 (
		\IR_reg[29]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w268_,
		_w2938_
	);
	LUT2 #(
		.INIT('h2)
	) name2721 (
		\datai[29]_pad ,
		\state_reg[0]/NET0131 ,
		_w2939_
	);
	LUT2 #(
		.INIT('he)
	) name2722 (
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT3 #(
		.INIT('h10)
	) name2723 (
		\IR_reg[29]/NET0131 ,
		\IR_reg[30]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w2941_
	);
	LUT4 #(
		.INIT('he222)
	) name2724 (
		\datai[31]_pad ,
		\state_reg[0]/NET0131 ,
		_w268_,
		_w2941_,
		_w2942_
	);
	LUT4 #(
		.INIT('hac5c)
	) name2725 (
		\IR_reg[15]/NET0131 ,
		\datai[15]_pad ,
		\state_reg[0]/NET0131 ,
		_w447_,
		_w2943_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2726 (
		\IR_reg[23]/NET0131 ,
		\datai[23]_pad ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w2944_
	);
	LUT4 #(
		.INIT('h4448)
	) name2727 (
		\IR_reg[24]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w238_,
		_w240_,
		_w2945_
	);
	LUT2 #(
		.INIT('h2)
	) name2728 (
		\datai[24]_pad ,
		\state_reg[0]/NET0131 ,
		_w2946_
	);
	LUT2 #(
		.INIT('he)
	) name2729 (
		_w2945_,
		_w2946_,
		_w2947_
	);
	LUT4 #(
		.INIT('h8884)
	) name2730 (
		\IR_reg[17]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w238_,
		_w409_,
		_w2948_
	);
	LUT2 #(
		.INIT('h1)
	) name2731 (
		\datai[17]_pad ,
		\state_reg[0]/NET0131 ,
		_w2949_
	);
	LUT2 #(
		.INIT('h1)
	) name2732 (
		_w2948_,
		_w2949_,
		_w2950_
	);
	LUT3 #(
		.INIT('h2e)
	) name2733 (
		\datai[22]_pad ,
		\state_reg[0]/NET0131 ,
		_w401_,
		_w2951_
	);
	LUT4 #(
		.INIT('h4448)
	) name2734 (
		\IR_reg[19]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w238_,
		_w402_,
		_w2952_
	);
	LUT2 #(
		.INIT('h2)
	) name2735 (
		\datai[19]_pad ,
		\state_reg[0]/NET0131 ,
		_w2953_
	);
	LUT2 #(
		.INIT('he)
	) name2736 (
		_w2952_,
		_w2953_,
		_w2954_
	);
	LUT2 #(
		.INIT('h1)
	) name2737 (
		\datai[16]_pad ,
		\state_reg[0]/NET0131 ,
		_w2955_
	);
	LUT4 #(
		.INIT('h5090)
	) name2738 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w233_,
		_w2956_
	);
	LUT2 #(
		.INIT('h1)
	) name2739 (
		_w2955_,
		_w2956_,
		_w2957_
	);
	LUT3 #(
		.INIT('he2)
	) name2740 (
		\datai[21]_pad ,
		\state_reg[0]/NET0131 ,
		_w398_,
		_w2958_
	);
	LUT2 #(
		.INIT('h1)
	) name2741 (
		\datai[20]_pad ,
		\state_reg[0]/NET0131 ,
		_w2959_
	);
	LUT4 #(
		.INIT('h5090)
	) name2742 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w235_,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name2743 (
		_w2959_,
		_w2960_,
		_w2961_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2744 (
		\IR_reg[26]/NET0131 ,
		\datai[26]_pad ,
		\state_reg[0]/NET0131 ,
		_w244_,
		_w2962_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2745 (
		\IR_reg[25]/NET0131 ,
		\datai[25]_pad ,
		\state_reg[0]/NET0131 ,
		_w248_,
		_w2963_
	);
	LUT3 #(
		.INIT('he2)
	) name2746 (
		\datai[11]_pad ,
		\state_reg[0]/NET0131 ,
		_w417_,
		_w2964_
	);
	LUT3 #(
		.INIT('he2)
	) name2747 (
		\datai[13]_pad ,
		\state_reg[0]/NET0131 ,
		_w441_,
		_w2965_
	);
	LUT3 #(
		.INIT('h2e)
	) name2748 (
		\datai[14]_pad ,
		\state_reg[0]/NET0131 ,
		_w438_,
		_w2966_
	);
	LUT4 #(
		.INIT('h4448)
	) name2749 (
		\IR_reg[12]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w420_,
		_w421_,
		_w2967_
	);
	LUT2 #(
		.INIT('h2)
	) name2750 (
		\datai[12]_pad ,
		\state_reg[0]/NET0131 ,
		_w2968_
	);
	LUT2 #(
		.INIT('he)
	) name2751 (
		_w2967_,
		_w2968_,
		_w2969_
	);
	LUT4 #(
		.INIT('h8884)
	) name2752 (
		\IR_reg[18]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w238_,
		_w676_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name2753 (
		\datai[18]_pad ,
		\state_reg[0]/NET0131 ,
		_w2971_
	);
	LUT2 #(
		.INIT('h1)
	) name2754 (
		_w2970_,
		_w2971_,
		_w2972_
	);
	LUT4 #(
		.INIT('hc060)
	) name2755 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w415_,
		_w2973_
	);
	LUT2 #(
		.INIT('h2)
	) name2756 (
		\datai[9]_pad ,
		\state_reg[0]/NET0131 ,
		_w2974_
	);
	LUT2 #(
		.INIT('he)
	) name2757 (
		_w2973_,
		_w2974_,
		_w2975_
	);
	LUT4 #(
		.INIT('hac5c)
	) name2758 (
		\IR_reg[7]/NET0131 ,
		\datai[7]_pad ,
		\state_reg[0]/NET0131 ,
		_w465_,
		_w2976_
	);
	LUT3 #(
		.INIT('he2)
	) name2759 (
		\datai[10]_pad ,
		\state_reg[0]/NET0131 ,
		_w426_,
		_w2977_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2760 (
		\IR_reg[8]/NET0131 ,
		\datai[8]_pad ,
		\state_reg[0]/NET0131 ,
		_w420_,
		_w2978_
	);
	LUT4 #(
		.INIT('hac5c)
	) name2761 (
		\IR_reg[6]/NET0131 ,
		\datai[6]_pad ,
		\state_reg[0]/NET0131 ,
		_w473_,
		_w2979_
	);
	LUT4 #(
		.INIT('hc060)
	) name2762 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w227_,
		_w2980_
	);
	LUT2 #(
		.INIT('h2)
	) name2763 (
		\datai[4]_pad ,
		\state_reg[0]/NET0131 ,
		_w2981_
	);
	LUT2 #(
		.INIT('he)
	) name2764 (
		_w2980_,
		_w2981_,
		_w2982_
	);
	LUT3 #(
		.INIT('he2)
	) name2765 (
		\datai[5]_pad ,
		\state_reg[0]/NET0131 ,
		_w478_,
		_w2983_
	);
	LUT4 #(
		.INIT('hac5c)
	) name2766 (
		\IR_reg[3]/NET0131 ,
		\datai[3]_pad ,
		\state_reg[0]/NET0131 ,
		_w500_,
		_w2984_
	);
	LUT3 #(
		.INIT('h2e)
	) name2767 (
		\datai[2]_pad ,
		\state_reg[0]/NET0131 ,
		_w496_,
		_w2985_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2768 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2986_
	);
	LUT2 #(
		.INIT('h2)
	) name2769 (
		\datai[1]_pad ,
		\state_reg[0]/NET0131 ,
		_w2987_
	);
	LUT2 #(
		.INIT('he)
	) name2770 (
		_w2986_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('haa2a)
	) name2771 (
		\reg2_reg[24]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w524_,
		_w2989_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2772 (
		\reg2_reg[24]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w2990_
	);
	LUT4 #(
		.INIT('h0c84)
	) name2773 (
		_w788_,
		_w970_,
		_w1092_,
		_w1095_,
		_w2991_
	);
	LUT3 #(
		.INIT('ha8)
	) name2774 (
		_w587_,
		_w2990_,
		_w2991_,
		_w2992_
	);
	LUT4 #(
		.INIT('h8288)
	) name2775 (
		_w970_,
		_w1092_,
		_w1100_,
		_w1103_,
		_w2993_
	);
	LUT3 #(
		.INIT('ha8)
	) name2776 (
		_w518_,
		_w2990_,
		_w2993_,
		_w2994_
	);
	LUT4 #(
		.INIT('h111d)
	) name2777 (
		\reg2_reg[24]/NET0131 ,
		_w970_,
		_w1106_,
		_w1107_,
		_w2995_
	);
	LUT4 #(
		.INIT('h9500)
	) name2778 (
		_w643_,
		_w799_,
		_w802_,
		_w970_,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name2779 (
		_w520_,
		_w644_,
		_w2997_
	);
	LUT4 #(
		.INIT('h1000)
	) name2780 (
		_w256_,
		_w258_,
		_w261_,
		_w643_,
		_w2998_
	);
	LUT4 #(
		.INIT('h1113)
	) name2781 (
		_w525_,
		_w2997_,
		_w2990_,
		_w2998_,
		_w2999_
	);
	LUT4 #(
		.INIT('h5700)
	) name2782 (
		_w601_,
		_w2990_,
		_w2996_,
		_w2999_,
		_w3000_
	);
	LUT3 #(
		.INIT('hd0)
	) name2783 (
		_w404_,
		_w2995_,
		_w3000_,
		_w3001_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2784 (
		_w1410_,
		_w2992_,
		_w2994_,
		_w3001_,
		_w3002_
	);
	LUT2 #(
		.INIT('he)
	) name2785 (
		_w2989_,
		_w3002_,
		_w3003_
	);
	LUT4 #(
		.INIT('h0155)
	) name2786 (
		\reg3_reg[3]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w3004_
	);
	LUT4 #(
		.INIT('h222e)
	) name2787 (
		\reg3_reg[3]/NET0131 ,
		_w262_,
		_w2074_,
		_w2075_,
		_w3005_
	);
	LUT4 #(
		.INIT('ha802)
	) name2788 (
		_w262_,
		_w572_,
		_w574_,
		_w2077_,
		_w3006_
	);
	LUT3 #(
		.INIT('ha8)
	) name2789 (
		_w587_,
		_w3004_,
		_w3006_,
		_w3007_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2790 (
		_w262_,
		_w499_,
		_w504_,
		_w2077_,
		_w3008_
	);
	LUT2 #(
		.INIT('h2)
	) name2791 (
		_w520_,
		_w502_,
		_w3009_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2792 (
		\reg3_reg[3]/NET0131 ,
		_w524_,
		_w906_,
		_w3009_,
		_w3010_
	);
	LUT3 #(
		.INIT('hd0)
	) name2793 (
		_w262_,
		_w2082_,
		_w3010_,
		_w3011_
	);
	LUT4 #(
		.INIT('h5700)
	) name2794 (
		_w518_,
		_w3004_,
		_w3008_,
		_w3011_,
		_w3012_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2795 (
		_w404_,
		_w3005_,
		_w3007_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h4)
	) name2796 (
		\reg3_reg[3]/NET0131 ,
		_w252_,
		_w3014_
	);
	LUT4 #(
		.INIT('haa08)
	) name2797 (
		\state_reg[0]/NET0131 ,
		_w254_,
		_w3013_,
		_w3014_,
		_w3015_
	);
	LUT4 #(
		.INIT('he3d3)
	) name2798 (
		\IR_reg[23]/NET0131 ,
		\reg3_reg[3]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w3016_
	);
	LUT2 #(
		.INIT('hb)
	) name2799 (
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT4 #(
		.INIT('haa2a)
	) name2800 (
		\reg2_reg[11]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w524_,
		_w3018_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2801 (
		\reg2_reg[11]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w3019_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2802 (
		\reg2_reg[11]/NET0131 ,
		_w970_,
		_w1034_,
		_w1035_,
		_w3020_
	);
	LUT4 #(
		.INIT('h00c8)
	) name2803 (
		_w418_,
		_w970_,
		_w1026_,
		_w1027_,
		_w3021_
	);
	LUT2 #(
		.INIT('h8)
	) name2804 (
		_w520_,
		_w346_,
		_w3022_
	);
	LUT4 #(
		.INIT('h0010)
	) name2805 (
		_w256_,
		_w258_,
		_w261_,
		_w418_,
		_w3023_
	);
	LUT4 #(
		.INIT('h1113)
	) name2806 (
		_w525_,
		_w3022_,
		_w3019_,
		_w3023_,
		_w3024_
	);
	LUT4 #(
		.INIT('h5700)
	) name2807 (
		_w601_,
		_w3019_,
		_w3021_,
		_w3024_,
		_w3025_
	);
	LUT3 #(
		.INIT('hd0)
	) name2808 (
		_w404_,
		_w3020_,
		_w3025_,
		_w3026_
	);
	LUT4 #(
		.INIT('hb040)
	) name2809 (
		_w865_,
		_w866_,
		_w970_,
		_w1024_,
		_w3027_
	);
	LUT3 #(
		.INIT('ha8)
	) name2810 (
		_w518_,
		_w3019_,
		_w3027_,
		_w3028_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2811 (
		\reg2_reg[11]/NET0131 ,
		_w840_,
		_w970_,
		_w1024_,
		_w3029_
	);
	LUT2 #(
		.INIT('h2)
	) name2812 (
		_w587_,
		_w3029_,
		_w3030_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2813 (
		_w1410_,
		_w3028_,
		_w3030_,
		_w3026_,
		_w3031_
	);
	LUT2 #(
		.INIT('he)
	) name2814 (
		_w3018_,
		_w3031_,
		_w3032_
	);
	LUT2 #(
		.INIT('h8)
	) name2815 (
		_w252_,
		_w369_,
		_w3033_
	);
	LUT3 #(
		.INIT('h04)
	) name2816 (
		_w521_,
		_w522_,
		_w442_,
		_w3034_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2817 (
		_w369_,
		_w524_,
		_w526_,
		_w1968_,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name2818 (
		_w3034_,
		_w3035_,
		_w3036_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2819 (
		_w254_,
		_w262_,
		_w2577_,
		_w3036_,
		_w3037_
	);
	LUT4 #(
		.INIT('h4800)
	) name2820 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w369_,
		_w3038_
	);
	LUT2 #(
		.INIT('h1)
	) name2821 (
		_w2700_,
		_w3038_,
		_w3039_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2822 (
		\state_reg[0]/NET0131 ,
		_w3033_,
		_w3037_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h8)
	) name2823 (
		_w252_,
		_w351_,
		_w3041_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2824 (
		_w256_,
		_w258_,
		_w261_,
		_w351_,
		_w3042_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2825 (
		_w262_,
		_w2133_,
		_w2134_,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h2)
	) name2826 (
		_w404_,
		_w3043_,
		_w3044_
	);
	LUT4 #(
		.INIT('h007d)
	) name2827 (
		_w262_,
		_w1322_,
		_w2137_,
		_w3042_,
		_w3045_
	);
	LUT2 #(
		.INIT('h2)
	) name2828 (
		_w587_,
		_w3045_,
		_w3046_
	);
	LUT4 #(
		.INIT('he040)
	) name2829 (
		_w262_,
		_w351_,
		_w601_,
		_w2140_,
		_w3047_
	);
	LUT4 #(
		.INIT('h0880)
	) name2830 (
		_w262_,
		_w518_,
		_w1445_,
		_w2137_,
		_w3048_
	);
	LUT3 #(
		.INIT('h04)
	) name2831 (
		_w521_,
		_w522_,
		_w427_,
		_w3049_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2832 (
		_w351_,
		_w524_,
		_w526_,
		_w1459_,
		_w3050_
	);
	LUT2 #(
		.INIT('h1)
	) name2833 (
		_w3049_,
		_w3050_,
		_w3051_
	);
	LUT3 #(
		.INIT('h10)
	) name2834 (
		_w3047_,
		_w3048_,
		_w3051_,
		_w3052_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2835 (
		_w254_,
		_w3044_,
		_w3046_,
		_w3052_,
		_w3053_
	);
	LUT4 #(
		.INIT('h4800)
	) name2836 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w351_,
		_w3054_
	);
	LUT2 #(
		.INIT('h1)
	) name2837 (
		_w2902_,
		_w3054_,
		_w3055_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2838 (
		\state_reg[0]/NET0131 ,
		_w3041_,
		_w3053_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h8)
	) name2839 (
		_w252_,
		_w317_,
		_w3057_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2840 (
		_w256_,
		_w258_,
		_w261_,
		_w317_,
		_w3058_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2841 (
		_w262_,
		_w2327_,
		_w2328_,
		_w2329_,
		_w3059_
	);
	LUT3 #(
		.INIT('ha8)
	) name2842 (
		_w404_,
		_w3058_,
		_w3059_,
		_w3060_
	);
	LUT4 #(
		.INIT('he040)
	) name2843 (
		_w262_,
		_w317_,
		_w587_,
		_w2334_,
		_w3061_
	);
	LUT4 #(
		.INIT('h00d7)
	) name2844 (
		_w262_,
		_w509_,
		_w2332_,
		_w3058_,
		_w3062_
	);
	LUT3 #(
		.INIT('ha8)
	) name2845 (
		_w317_,
		_w524_,
		_w906_,
		_w3063_
	);
	LUT3 #(
		.INIT('h04)
	) name2846 (
		_w521_,
		_w522_,
		_w479_,
		_w3064_
	);
	LUT4 #(
		.INIT('h0007)
	) name2847 (
		_w262_,
		_w2338_,
		_w3063_,
		_w3064_,
		_w3065_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2848 (
		_w518_,
		_w3062_,
		_w3061_,
		_w3065_,
		_w3066_
	);
	LUT4 #(
		.INIT('h1311)
	) name2849 (
		_w254_,
		_w3057_,
		_w3060_,
		_w3066_,
		_w3067_
	);
	LUT4 #(
		.INIT('h4800)
	) name2850 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w236_,
		_w317_,
		_w3068_
	);
	LUT2 #(
		.INIT('h1)
	) name2851 (
		_w2831_,
		_w3068_,
		_w3069_
	);
	LUT3 #(
		.INIT('h2f)
	) name2852 (
		\state_reg[0]/NET0131 ,
		_w3067_,
		_w3069_,
		_w3070_
	);
	LUT4 #(
		.INIT('haa2a)
	) name2853 (
		\reg2_reg[17]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w524_,
		_w3071_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2854 (
		\reg2_reg[17]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w3072_
	);
	LUT4 #(
		.INIT('hfc55)
	) name2855 (
		\reg2_reg[17]/NET0131 ,
		_w395_,
		_w396_,
		_w970_,
		_w3073_
	);
	LUT2 #(
		.INIT('h2)
	) name2856 (
		_w404_,
		_w3073_,
		_w3074_
	);
	LUT4 #(
		.INIT('h30a0)
	) name2857 (
		\reg2_reg[17]/NET0131 ,
		_w514_,
		_w518_,
		_w970_,
		_w3075_
	);
	LUT2 #(
		.INIT('h8)
	) name2858 (
		_w224_,
		_w520_,
		_w3076_
	);
	LUT4 #(
		.INIT('h1000)
	) name2859 (
		_w256_,
		_w258_,
		_w261_,
		_w411_,
		_w3077_
	);
	LUT4 #(
		.INIT('h1113)
	) name2860 (
		_w525_,
		_w3076_,
		_w3072_,
		_w3077_,
		_w3078_
	);
	LUT4 #(
		.INIT('h5900)
	) name2861 (
		_w414_,
		_w552_,
		_w585_,
		_w970_,
		_w3079_
	);
	LUT3 #(
		.INIT('ha8)
	) name2862 (
		_w587_,
		_w3072_,
		_w3079_,
		_w3080_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2863 (
		_w411_,
		_w597_,
		_w599_,
		_w970_,
		_w3081_
	);
	LUT3 #(
		.INIT('ha8)
	) name2864 (
		_w601_,
		_w3072_,
		_w3081_,
		_w3082_
	);
	LUT4 #(
		.INIT('h0100)
	) name2865 (
		_w3075_,
		_w3080_,
		_w3082_,
		_w3078_,
		_w3083_
	);
	LUT4 #(
		.INIT('hecee)
	) name2866 (
		_w1410_,
		_w3071_,
		_w3074_,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('haa2a)
	) name2867 (
		\reg2_reg[2]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w524_,
		_w3085_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2868 (
		\reg2_reg[2]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w3086_
	);
	LUT4 #(
		.INIT('hc808)
	) name2869 (
		\reg2_reg[2]/NET0131 ,
		_w404_,
		_w970_,
		_w1978_,
		_w3087_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2870 (
		_w970_,
		_w1983_,
		_w1985_,
		_w2314_,
		_w3088_
	);
	LUT2 #(
		.INIT('h8)
	) name2871 (
		\reg3_reg[2]/NET0131 ,
		_w520_,
		_w3089_
	);
	LUT3 #(
		.INIT('h51)
	) name2872 (
		_w3089_,
		_w3086_,
		_w2551_,
		_w3090_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2873 (
		_w1410_,
		_w3087_,
		_w3088_,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('he)
	) name2874 (
		_w3085_,
		_w3091_,
		_w3092_
	);
	LUT4 #(
		.INIT('haa2a)
	) name2875 (
		\reg2_reg[21]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w524_,
		_w3093_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2876 (
		\reg2_reg[21]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w3094_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2877 (
		\reg2_reg[21]/NET0131 ,
		_w970_,
		_w2306_,
		_w2307_,
		_w3095_
	);
	LUT2 #(
		.INIT('h2)
	) name2878 (
		_w404_,
		_w3095_,
		_w3096_
	);
	LUT2 #(
		.INIT('h8)
	) name2879 (
		_w520_,
		_w662_,
		_w3097_
	);
	LUT3 #(
		.INIT('h23)
	) name2880 (
		_w2551_,
		_w3097_,
		_w3094_,
		_w3098_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2881 (
		_w970_,
		_w2305_,
		_w3096_,
		_w3098_,
		_w3099_
	);
	LUT3 #(
		.INIT('hce)
	) name2882 (
		_w1410_,
		_w3093_,
		_w3099_,
		_w3100_
	);
	LUT4 #(
		.INIT('haa2a)
	) name2883 (
		\reg2_reg[26]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w254_,
		_w524_,
		_w3101_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2884 (
		\reg2_reg[26]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w3102_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2885 (
		\reg2_reg[26]/NET0131 ,
		_w970_,
		_w1426_,
		_w1436_,
		_w3103_
	);
	LUT4 #(
		.INIT('h7020)
	) name2886 (
		_w266_,
		_w640_,
		_w970_,
		_w1438_,
		_w3104_
	);
	LUT3 #(
		.INIT('ha8)
	) name2887 (
		_w404_,
		_w3102_,
		_w3104_,
		_w3105_
	);
	LUT4 #(
		.INIT('h6500)
	) name2888 (
		_w627_,
		_w635_,
		_w804_,
		_w970_,
		_w3106_
	);
	LUT3 #(
		.INIT('ha8)
	) name2889 (
		_w601_,
		_w3102_,
		_w3106_,
		_w3107_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2890 (
		\reg2_reg[26]/NET0131 ,
		_w970_,
		_w1426_,
		_w1457_,
		_w3108_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		_w520_,
		_w628_,
		_w3109_
	);
	LUT4 #(
		.INIT('h1000)
	) name2892 (
		_w256_,
		_w258_,
		_w261_,
		_w627_,
		_w3110_
	);
	LUT4 #(
		.INIT('h1113)
	) name2893 (
		_w525_,
		_w3109_,
		_w3102_,
		_w3110_,
		_w3111_
	);
	LUT4 #(
		.INIT('h3100)
	) name2894 (
		_w518_,
		_w3107_,
		_w3108_,
		_w3111_,
		_w3112_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2895 (
		_w587_,
		_w3103_,
		_w3105_,
		_w3112_,
		_w3113_
	);
	LUT3 #(
		.INIT('hce)
	) name2896 (
		_w1410_,
		_w3101_,
		_w3113_,
		_w3114_
	);
	LUT4 #(
		.INIT('haa02)
	) name2897 (
		\reg1_reg[18]/NET0131 ,
		_w256_,
		_w258_,
		_w261_,
		_w3115_
	);
	LUT4 #(
		.INIT('h2d00)
	) name2898 (
		_w1427_,
		_w1429_,
		_w1641_,
		_w1871_,
		_w3116_
	);
	LUT3 #(
		.INIT('ha8)
	) name2899 (
		_w587_,
		_w3115_,
		_w3116_,
		_w3117_
	);
	LUT3 #(
		.INIT('h02)
	) name2900 (
		_w404_,
		_w1644_,
		_w1645_,
		_w3118_
	);
	LUT3 #(
		.INIT('h2a)
	) name2901 (
		\reg1_reg[18]/NET0131 ,
		_w1221_,
		_w1410_,
		_w3119_
	);
	LUT4 #(
		.INIT('h005d)
	) name2902 (
		_w1871_,
		_w2097_,
		_w3118_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('hb)
	) name2903 (
		_w3117_,
		_w3120_,
		_w3121_
	);
	LUT4 #(
		.INIT('h7000)
	) name2904 (
		_w241_,
		_w250_,
		_w266_,
		_w407_,
		_w3122_
	);
	LUT4 #(
		.INIT('ha888)
	) name2905 (
		\state_reg[0]/NET0131 ,
		_w237_,
		_w404_,
		_w3122_,
		_w3123_
	);
	LUT2 #(
		.INIT('h2)
	) name2906 (
		\B_reg/NET0131 ,
		_w3123_,
		_w3124_
	);
	LUT4 #(
		.INIT('h0705)
	) name2907 (
		_w634_,
		_w649_,
		_w725_,
		_w889_,
		_w3125_
	);
	LUT4 #(
		.INIT('h0705)
	) name2908 (
		_w659_,
		_w673_,
		_w722_,
		_w886_,
		_w3126_
	);
	LUT4 #(
		.INIT('h2302)
	) name2909 (
		_w335_,
		_w429_,
		_w431_,
		_w471_,
		_w3127_
	);
	LUT3 #(
		.INIT('h51)
	) name2910 (
		_w435_,
		_w692_,
		_w3127_,
		_w3128_
	);
	LUT4 #(
		.INIT('h008e)
	) name2911 (
		_w372_,
		_w424_,
		_w442_,
		_w453_,
		_w3129_
	);
	LUT3 #(
		.INIT('h51)
	) name2912 (
		_w457_,
		_w707_,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h1)
	) name2913 (
		_w3128_,
		_w3130_,
		_w3131_
	);
	LUT3 #(
		.INIT('ha8)
	) name2914 (
		_w713_,
		_w3128_,
		_w3130_,
		_w3132_
	);
	LUT4 #(
		.INIT('h020b)
	) name2915 (
		_w280_,
		_w491_,
		_w498_,
		_w2460_,
		_w3133_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2916 (
		_w505_,
		_w508_,
		_w699_,
		_w3133_,
		_w3134_
	);
	LUT4 #(
		.INIT('h0001)
	) name2917 (
		_w429_,
		_w432_,
		_w434_,
		_w435_,
		_w3135_
	);
	LUT3 #(
		.INIT('h01)
	) name2918 (
		_w457_,
		_w483_,
		_w484_,
		_w3136_
	);
	LUT3 #(
		.INIT('h80)
	) name2919 (
		_w455_,
		_w3135_,
		_w3136_,
		_w3137_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2920 (
		_w481_,
		_w696_,
		_w3134_,
		_w3137_,
		_w3138_
	);
	LUT4 #(
		.INIT('h000b)
	) name2921 (
		_w361_,
		_w446_,
		_w714_,
		_w717_,
		_w3139_
	);
	LUT3 #(
		.INIT('h8a)
	) name2922 (
		_w688_,
		_w690_,
		_w872_,
		_w3140_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2923 (
		_w3132_,
		_w3138_,
		_w3139_,
		_w3140_,
		_w3141_
	);
	LUT3 #(
		.INIT('h40)
	) name2924 (
		_w722_,
		_w884_,
		_w886_,
		_w3142_
	);
	LUT2 #(
		.INIT('h8)
	) name2925 (
		_w726_,
		_w728_,
		_w3143_
	);
	LUT4 #(
		.INIT('hba00)
	) name2926 (
		_w3126_,
		_w3141_,
		_w3142_,
		_w3143_,
		_w3144_
	);
	LUT4 #(
		.INIT('h00ba)
	) name2927 (
		_w733_,
		_w734_,
		_w737_,
		_w1269_,
		_w3145_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2928 (
		_w296_,
		_w1260_,
		_w1261_,
		_w1414_,
		_w3146_
	);
	LUT4 #(
		.INIT('h1000)
	) name2929 (
		_w296_,
		_w297_,
		_w298_,
		_w1413_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name2930 (
		_w3146_,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h8)
	) name2931 (
		_w3145_,
		_w3148_,
		_w3149_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2932 (
		_w296_,
		_w297_,
		_w298_,
		_w1413_,
		_w3150_
	);
	LUT4 #(
		.INIT('h1000)
	) name2933 (
		_w296_,
		_w1260_,
		_w1261_,
		_w1414_,
		_w3151_
	);
	LUT2 #(
		.INIT('h1)
	) name2934 (
		_w3150_,
		_w3151_,
		_w3152_
	);
	LUT4 #(
		.INIT('h00df)
	) name2935 (
		_w733_,
		_w734_,
		_w737_,
		_w1268_,
		_w3153_
	);
	LUT2 #(
		.INIT('h1)
	) name2936 (
		_w1269_,
		_w3146_,
		_w3154_
	);
	LUT4 #(
		.INIT('h1303)
	) name2937 (
		_w3153_,
		_w3147_,
		_w3152_,
		_w3154_,
		_w3155_
	);
	LUT4 #(
		.INIT('h001f)
	) name2938 (
		_w3125_,
		_w3144_,
		_w3149_,
		_w3155_,
		_w3156_
	);
	LUT3 #(
		.INIT('h84)
	) name2939 (
		_w403_,
		_w400_,
		_w3156_,
		_w3157_
	);
	LUT3 #(
		.INIT('hc8)
	) name2940 (
		_w299_,
		_w1413_,
		_w3146_,
		_w3158_
	);
	LUT2 #(
		.INIT('h1)
	) name2941 (
		_w1268_,
		_w3145_,
		_w3159_
	);
	LUT2 #(
		.INIT('h8)
	) name2942 (
		_w675_,
		_w691_,
		_w3160_
	);
	LUT4 #(
		.INIT('hccc8)
	) name2943 (
		_w477_,
		_w696_,
		_w700_,
		_w701_,
		_w3161_
	);
	LUT2 #(
		.INIT('h1)
	) name2944 (
		_w484_,
		_w1101_,
		_w3162_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2945 (
		_w713_,
		_w3131_,
		_w3161_,
		_w3162_,
		_w3163_
	);
	LUT4 #(
		.INIT('h002a)
	) name2946 (
		_w650_,
		_w719_,
		_w724_,
		_w3126_,
		_w3164_
	);
	LUT2 #(
		.INIT('h1)
	) name2947 (
		_w730_,
		_w3164_,
		_w3165_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2948 (
		_w3153_,
		_w3160_,
		_w3163_,
		_w3165_,
		_w3166_
	);
	LUT4 #(
		.INIT('h001f)
	) name2949 (
		_w299_,
		_w1262_,
		_w1414_,
		_w3150_,
		_w3167_
	);
	LUT4 #(
		.INIT('h0155)
	) name2950 (
		_w3158_,
		_w3159_,
		_w3166_,
		_w3167_,
		_w3168_
	);
	LUT4 #(
		.INIT('h2818)
	) name2951 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w235_,
		_w3169_
	);
	LUT3 #(
		.INIT('h60)
	) name2952 (
		_w403_,
		_w3168_,
		_w3169_,
		_w3170_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name2953 (
		_w1268_,
		_w3145_,
		_w3148_,
		_w3151_,
		_w3171_
	);
	LUT2 #(
		.INIT('h1)
	) name2954 (
		_w3150_,
		_w3171_,
		_w3172_
	);
	LUT2 #(
		.INIT('h8)
	) name2955 (
		_w3153_,
		_w3152_,
		_w3173_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2956 (
		_w1351_,
		_w3160_,
		_w3165_,
		_w3173_,
		_w3174_
	);
	LUT3 #(
		.INIT('h02)
	) name2957 (
		_w1989_,
		_w3172_,
		_w3174_,
		_w3175_
	);
	LUT3 #(
		.INIT('h10)
	) name2958 (
		_w398_,
		_w399_,
		_w403_,
		_w3176_
	);
	LUT2 #(
		.INIT('h2)
	) name2959 (
		\B_reg/NET0131 ,
		_w401_,
		_w3177_
	);
	LUT4 #(
		.INIT('h1428)
	) name2960 (
		_w615_,
		_w643_,
		_w647_,
		_w651_,
		_w3178_
	);
	LUT4 #(
		.INIT('h0990)
	) name2961 (
		_w361_,
		_w446_,
		_w667_,
		_w671_,
		_w3179_
	);
	LUT2 #(
		.INIT('h8)
	) name2962 (
		_w3178_,
		_w3179_,
		_w3180_
	);
	LUT4 #(
		.INIT('h4000)
	) name2963 (
		_w1373_,
		_w1805_,
		_w1963_,
		_w1980_,
		_w3181_
	);
	LUT3 #(
		.INIT('h01)
	) name2964 (
		_w414_,
		_w1024_,
		_w1046_,
		_w3182_
	);
	LUT4 #(
		.INIT('h0080)
	) name2965 (
		_w2214_,
		_w2332_,
		_w2461_,
		_w2540_,
		_w3183_
	);
	LUT4 #(
		.INIT('h0004)
	) name2966 (
		_w2002_,
		_w2039_,
		_w2077_,
		_w2137_,
		_w3184_
	);
	LUT4 #(
		.INIT('h8000)
	) name2967 (
		_w3183_,
		_w3184_,
		_w3181_,
		_w3182_,
		_w3185_
	);
	LUT3 #(
		.INIT('h06)
	) name2968 (
		_w652_,
		_w657_,
		_w1668_,
		_w3186_
	);
	LUT3 #(
		.INIT('h10)
	) name2969 (
		_w861_,
		_w2300_,
		_w3186_,
		_w3187_
	);
	LUT3 #(
		.INIT('h80)
	) name2970 (
		_w3180_,
		_w3185_,
		_w3187_,
		_w3188_
	);
	LUT3 #(
		.INIT('h01)
	) name2971 (
		_w1641_,
		_w3146_,
		_w3147_,
		_w3189_
	);
	LUT4 #(
		.INIT('h1000)
	) name2972 (
		_w1006_,
		_w1066_,
		_w1270_,
		_w1319_,
		_w3190_
	);
	LUT4 #(
		.INIT('h4000)
	) name2973 (
		_w1426_,
		_w3152_,
		_w3189_,
		_w3190_,
		_w3191_
	);
	LUT2 #(
		.INIT('h4)
	) name2974 (
		_w741_,
		_w3191_,
		_w3192_
	);
	LUT4 #(
		.INIT('h8242)
	) name2975 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w235_,
		_w3193_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2976 (
		_w403_,
		_w3188_,
		_w3192_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h1)
	) name2977 (
		_w3177_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2978 (
		_w3172_,
		_w3174_,
		_w3176_,
		_w3195_,
		_w3196_
	);
	LUT2 #(
		.INIT('h4)
	) name2979 (
		_w3175_,
		_w3196_,
		_w3197_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2980 (
		_w606_,
		_w3170_,
		_w3157_,
		_w3197_,
		_w3198_
	);
	LUT2 #(
		.INIT('he)
	) name2981 (
		_w3124_,
		_w3198_,
		_w3199_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g22/_0_  = _w609_ ;
	assign \g32_dup/_0_  = _w616_ ;
	assign \g35904/_0_  = _w833_ ;
	assign \g35905/_0_  = _w916_ ;
	assign \g35906/_0_  = _w933_ ;
	assign \g35907/_0_  = _w945_ ;
	assign \g35908/_0_  = _w956_ ;
	assign \g35909/_0_  = _w969_ ;
	assign \g35910/_0_  = _w986_ ;
	assign \g35911/_0_  = _w999_ ;
	assign \g35932/_0_  = _w1021_ ;
	assign \g35955/_0_  = _w1043_ ;
	assign \g35956/_0_  = _w1064_ ;
	assign \g35957/_0_  = _w1089_ ;
	assign \g35962/_0_  = _w1118_ ;
	assign \g35967/_0_  = _w1144_ ;
	assign \g35968/_0_  = _w1160_ ;
	assign \g35971/_0_  = _w1174_ ;
	assign \g35972/_0_  = _w1192_ ;
	assign \g35973/_0_  = _w1204_ ;
	assign \g35974/_0_  = _w1216_ ;
	assign \g35975/_0_  = _w1228_ ;
	assign \g35976/_0_  = _w1242_ ;
	assign \g35977/_0_  = _w1255_ ;
	assign \g35978/_0_  = _w1313_ ;
	assign \g36015/_0_  = _w1344_ ;
	assign \g36016/_0_  = _w1366_ ;
	assign \g36018/_0_  = _w1387_ ;
	assign \g36022/_0_  = _w1408_ ;
	assign \g36023/_0_  = _w1424_ ;
	assign \g36025/_0_  = _w1469_ ;
	assign \g36029/_0_  = _w1481_ ;
	assign \g36030/_0_  = _w1495_ ;
	assign \g36031/_0_  = _w1510_ ;
	assign \g36032/_0_  = _w1527_ ;
	assign \g36033/_0_  = _w1537_ ;
	assign \g36034/_0_  = _w1550_ ;
	assign \g36035/_0_  = _w1565_ ;
	assign \g36036/_0_  = _w1580_ ;
	assign \g36038/_0_  = _w1597_ ;
	assign \g36039/_0_  = _w1609_ ;
	assign \g36040/_0_  = _w1623_ ;
	assign \g36041/_0_  = _w1639_ ;
	assign \g36073/_0_  = _w1661_ ;
	assign \g36087/_0_  = _w1686_ ;
	assign \g36091/_0_  = _w1711_ ;
	assign \g36092/_0_  = _w1725_ ;
	assign \g36093/_0_  = _w1740_ ;
	assign \g36094/_0_  = _w1755_ ;
	assign \g36096/_0_  = _w1766_ ;
	assign \g36097/_0_  = _w1779_ ;
	assign \g36098/_0_  = _w1783_ ;
	assign \g36099/_0_  = _w1785_ ;
	assign \g36100/_0_  = _w1796_ ;
	assign \g36101/_0_  = _w1818_ ;
	assign \g36102/_0_  = _w1834_ ;
	assign \g36103/_0_  = _w1846_ ;
	assign \g36104/_0_  = _w1860_ ;
	assign \g36105/_0_  = _w1870_ ;
	assign \g36106/_0_  = _w1873_ ;
	assign \g36107/_0_  = _w1880_ ;
	assign \g36108/_0_  = _w1892_ ;
	assign \g36109/_0_  = _w1907_ ;
	assign \g36110/_0_  = _w1918_ ;
	assign \g36111/_0_  = _w1933_ ;
	assign \g36112/_0_  = _w1945_ ;
	assign \g36113/_0_  = _w1955_ ;
	assign \g36165/_0_  = _w1973_ ;
	assign \g36169/_0_  = _w1996_ ;
	assign \g36170/_0_  = _w2016_ ;
	assign \g36171/_0_  = _w2033_ ;
	assign \g36172/_0_  = _w2055_ ;
	assign \g36198/_0_  = _w2072_ ;
	assign \g36199/_0_  = _w2091_ ;
	assign \g36200/_0_  = _w2104_ ;
	assign \g36201/_0_  = _w2120_ ;
	assign \g36202/_0_  = _w2132_ ;
	assign \g36203/_0_  = _w2149_ ;
	assign \g36205/_0_  = _w2165_ ;
	assign \g36206/_0_  = _w2176_ ;
	assign \g36207/_0_  = _w2189_ ;
	assign \g36208/_0_  = _w2199_ ;
	assign \g36209/_0_  = _w2212_ ;
	assign \g36240/_0_  = _w2234_ ;
	assign \g36281/_0_  = _w2251_ ;
	assign \g36282/_0_  = _w2267_ ;
	assign \g36283/_0_  = _w2284_ ;
	assign \g36284/_0_  = _w2292_ ;
	assign \g36285/_0_  = _w2311_ ;
	assign \g36286/_0_  = _w2318_ ;
	assign \g36287/_0_  = _w2323_ ;
	assign \g36288/_0_  = _w2342_ ;
	assign \g36289/_0_  = _w2355_ ;
	assign \g36290/_0_  = _w2371_ ;
	assign \g36291/_0_  = _w2387_ ;
	assign \g36292/_0_  = _w2391_ ;
	assign \g36293/_0_  = _w2396_ ;
	assign \g36294/_0_  = _w2400_ ;
	assign \g36295/_0_  = _w2412_ ;
	assign \g36296/_0_  = _w2425_ ;
	assign \g36297/_0_  = _w2440_ ;
	assign \g36298/_0_  = _w2455_ ;
	assign \g36330/_0_  = _w2467_ ;
	assign \g36385/_0_  = _w2479_ ;
	assign \g36390/_0_  = _w2487_ ;
	assign \g36391/_0_  = _w2502_ ;
	assign \g36392/_0_  = _w2518_ ;
	assign \g36393/_0_  = _w2524_ ;
	assign \g36394/_0_  = _w2533_ ;
	assign \g36470/_0_  = _w2536_ ;
	assign \g36471/_0_  = _w2556_ ;
	assign \g36472/_0_  = _w2566_ ;
	assign \g36473/_0_  = _w2573_ ;
	assign \g36474/_0_  = _w2583_ ;
	assign \g36475/_0_  = _w2585_ ;
	assign \g38/_0_  = _w368_ ;
	assign \g38399/_0_  = _w2610_ ;
	assign \g38400/_0_  = _w2630_ ;
	assign \g39639/_0_  = _w2681_ ;
	assign \g39641/_0_  = _w2702_ ;
	assign \g39644/_0_  = _w2721_ ;
	assign \g39647/_0_  = _w2739_ ;
	assign \g39648/_0_  = _w2761_ ;
	assign \g39650/_0_  = _w2784_ ;
	assign \g39654/_0_  = _w2798_ ;
	assign \g39658/_0_  = _w2810_ ;
	assign \g39660/_0_  = _w2822_ ;
	assign \g39662/_0_  = _w2832_ ;
	assign \g39663/_0_  = _w2846_ ;
	assign \g39665/_0_  = _w2857_ ;
	assign \g39666/_0_  = _w2868_ ;
	assign \g39667/_0_  = _w2878_ ;
	assign \g39730/_0_  = _w2893_ ;
	assign \g39796/_0_  = _w2894_ ;
	assign \g39930/_0_  = _w2901_ ;
	assign \g39931/_0_  = _w2911_ ;
	assign \g39932/_0_  = _w2922_ ;
	assign \g40045/_0_  = _w259_ ;
	assign \g40150/u3_syn_4  = _w1410_ ;
	assign \g40608/_0_  = _w261_ ;
	assign \g41017/u3_syn_4  = _w2923_ ;
	assign \g42159/_0_  = _w2926_ ;
	assign \g42169/_0_  = _w2927_ ;
	assign \g42174/_0_  = _w2928_ ;
	assign \g42483/_0_  = _w821_ ;
	assign \g42736/_0_  = _w310_ ;
	assign \g42746/_0_  = _w373_ ;
	assign \g42755/_0_  = _w305_ ;
	assign \g42767/_0_  = _w281_ ;
	assign \g42776/_0_  = _w327_ ;
	assign \g42871_dup/_1_  = _w666_ ;
	assign \g42908/_0_  = _w648_ ;
	assign \g42938/_0_  = _w354_ ;
	assign \g42969/_0_  = _w344_ ;
	assign \g43022/_0_  = _w672_ ;
	assign \g44035/_1__syn_2  = _w931_ ;
	assign \g44227/_3_  = _w2931_ ;
	assign \g44260/_3_  = _w2934_ ;
	assign \g44261/_3_  = _w2937_ ;
	assign \g44262/_3_  = _w2940_ ;
	assign \g44311/_3_  = _w2942_ ;
	assign \g44378/_3_  = _w2943_ ;
	assign \g44379/_3_  = _w2944_ ;
	assign \g44383/_3_  = _w2947_ ;
	assign \g44384/_3_  = _w2950_ ;
	assign \g44385/_3_  = _w2951_ ;
	assign \g44386/_3_  = _w2954_ ;
	assign \g44390/_3_  = _w2957_ ;
	assign \g44391/_3_  = _w2958_ ;
	assign \g44492/_3_  = _w2961_ ;
	assign \g44493/_3_  = _w2962_ ;
	assign \g44494/_3_  = _w2963_ ;
	assign \g44495/_3_  = _w2964_ ;
	assign \g44496/_3_  = _w2965_ ;
	assign \g44497/_3_  = _w2966_ ;
	assign \g44498/_3_  = _w2969_ ;
	assign \g44499/_3_  = _w2972_ ;
	assign \g44575/_3_  = _w2975_ ;
	assign \g44589/_3_  = _w2976_ ;
	assign \g44596/_3_  = _w2977_ ;
	assign \g44615/_3_  = _w2978_ ;
	assign \g44795/_3_  = _w2979_ ;
	assign \g44803/_3_  = _w2982_ ;
	assign \g44804/_3_  = _w2983_ ;
	assign \g44888/_3_  = _w2984_ ;
	assign \g44889/_3_  = _w2985_ ;
	assign \g45004/_3_  = _w2988_ ;
	assign \g46129/_0_  = _w285_ ;
	assign \g46133/_0_  = _w300_ ;
	assign \g46265/_2_  = _w321_ ;
	assign \g46313/_0_  = _w3003_ ;
	assign \g46372/_0_  = _w3017_ ;
	assign \g46377/_0_  = _w3032_ ;
	assign \g46399/_0_  = _w3040_ ;
	assign \g46405/_0_  = _w3056_ ;
	assign \g46427/_0_  = _w3070_ ;
	assign \g46461/_0_  = _w3084_ ;
	assign \g46526/_0_  = _w3092_ ;
	assign \g46576/_0_  = _w362_ ;
	assign \g46608/_0_  = _w277_ ;
	assign \g46697/_0_  = _w658_ ;
	assign \g46778/_0_  = _w316_ ;
	assign \g47007/_0_  = _w336_ ;
	assign \g47023/_0_  = _w3100_ ;
	assign \g47077/_1_  = _w392_ ;
	assign \g47097/_0_  = _w685_ ;
	assign \g47109/_1_  = _w632_ ;
	assign \g47142_dup/_1_  = _w349_ ;
	assign \g47256/_0_  = _w625_ ;
	assign \g47328/_0_  = _w3114_ ;
	assign \g47373/_0_  = _w3121_ ;
	assign \g47465/_0_  = _w1263_ ;
	assign \g47518/_0_  = _w3199_ ;
	assign \g47556/_1_  = _w641_ ;
	assign \g56/_0_  = _w385_ ;
	assign \state_reg[0]/NET0131_syn_2  = _w218_ ;
endmodule;