module top (\101GAT(25)_pad , \106GAT(26)_pad , \111GAT(27)_pad , \116GAT(28)_pad , \121GAT(29)_pad , \126GAT(30)_pad , \130GAT(31)_pad , \135GAT(32)_pad , \138GAT(33)_pad , \13GAT(2)_pad , \143GAT(34)_pad , \146GAT(35)_pad , \149GAT(36)_pad , \152GAT(37)_pad , \153GAT(38)_pad , \156GAT(39)_pad , \159GAT(40)_pad , \165GAT(41)_pad , \171GAT(42)_pad , \177GAT(43)_pad , \17GAT(3)_pad , \183GAT(44)_pad , \189GAT(45)_pad , \195GAT(46)_pad , \1GAT(0)_pad , \201GAT(47)_pad , \207GAT(48)_pad , \210GAT(49)_pad , \219GAT(50)_pad , \228GAT(51)_pad , \237GAT(52)_pad , \246GAT(53)_pad , \255GAT(54)_pad , \259GAT(55)_pad , \260GAT(56)_pad , \261GAT(57)_pad , \267GAT(58)_pad , \268GAT(59)_pad , \26GAT(4)_pad , \29GAT(5)_pad , \36GAT(6)_pad , \42GAT(7)_pad , \51GAT(8)_pad , \55GAT(9)_pad , \59GAT(10)_pad , \68GAT(11)_pad , \72GAT(12)_pad , \73GAT(13)_pad , \74GAT(14)_pad , \75GAT(15)_pad , \80GAT(16)_pad , \85GAT(17)_pad , \86GAT(18)_pad , \87GAT(19)_pad , \88GAT(20)_pad , \89GAT(21)_pad , \8GAT(1)_pad , \90GAT(22)_pad , \91GAT(23)_pad , \96GAT(24)_pad , \273GAT(103) , \388GAT(133)_pad , \389GAT(132)_pad , \391GAT(124)_pad , \393GAT(165) , \418GAT(168)_pad , \419GAT(164)_pad , \420GAT(158)_pad , \421GAT(162)_pad , \422GAT(161)_pad , \423GAT(155)_pad , \446GAT(183)_pad , \448GAT(179)_pad , \449GAT(176)_pad , \450GAT(173)_pad , \767GAT(349)_pad , \768GAT(334)_pad , \811GAT(378) , \837GAT(396) , \838GAT(395) , \839GAT(394) , \854GAT(419) , \866GAT(426)_pad , \867GAT(432) , \868GAT(431) , \869GAT(430) );
	input \101GAT(25)_pad  ;
	input \106GAT(26)_pad  ;
	input \111GAT(27)_pad  ;
	input \116GAT(28)_pad  ;
	input \121GAT(29)_pad  ;
	input \126GAT(30)_pad  ;
	input \130GAT(31)_pad  ;
	input \135GAT(32)_pad  ;
	input \138GAT(33)_pad  ;
	input \13GAT(2)_pad  ;
	input \143GAT(34)_pad  ;
	input \146GAT(35)_pad  ;
	input \149GAT(36)_pad  ;
	input \152GAT(37)_pad  ;
	input \153GAT(38)_pad  ;
	input \156GAT(39)_pad  ;
	input \159GAT(40)_pad  ;
	input \165GAT(41)_pad  ;
	input \171GAT(42)_pad  ;
	input \177GAT(43)_pad  ;
	input \17GAT(3)_pad  ;
	input \183GAT(44)_pad  ;
	input \189GAT(45)_pad  ;
	input \195GAT(46)_pad  ;
	input \1GAT(0)_pad  ;
	input \201GAT(47)_pad  ;
	input \207GAT(48)_pad  ;
	input \210GAT(49)_pad  ;
	input \219GAT(50)_pad  ;
	input \228GAT(51)_pad  ;
	input \237GAT(52)_pad  ;
	input \246GAT(53)_pad  ;
	input \255GAT(54)_pad  ;
	input \259GAT(55)_pad  ;
	input \260GAT(56)_pad  ;
	input \261GAT(57)_pad  ;
	input \267GAT(58)_pad  ;
	input \268GAT(59)_pad  ;
	input \26GAT(4)_pad  ;
	input \29GAT(5)_pad  ;
	input \36GAT(6)_pad  ;
	input \42GAT(7)_pad  ;
	input \51GAT(8)_pad  ;
	input \55GAT(9)_pad  ;
	input \59GAT(10)_pad  ;
	input \68GAT(11)_pad  ;
	input \72GAT(12)_pad  ;
	input \73GAT(13)_pad  ;
	input \74GAT(14)_pad  ;
	input \75GAT(15)_pad  ;
	input \80GAT(16)_pad  ;
	input \85GAT(17)_pad  ;
	input \86GAT(18)_pad  ;
	input \87GAT(19)_pad  ;
	input \88GAT(20)_pad  ;
	input \89GAT(21)_pad  ;
	input \8GAT(1)_pad  ;
	input \90GAT(22)_pad  ;
	input \91GAT(23)_pad  ;
	input \96GAT(24)_pad  ;
	output \273GAT(103)  ;
	output \388GAT(133)_pad  ;
	output \389GAT(132)_pad  ;
	output \391GAT(124)_pad  ;
	output \393GAT(165)  ;
	output \418GAT(168)_pad  ;
	output \419GAT(164)_pad  ;
	output \420GAT(158)_pad  ;
	output \421GAT(162)_pad  ;
	output \422GAT(161)_pad  ;
	output \423GAT(155)_pad  ;
	output \446GAT(183)_pad  ;
	output \448GAT(179)_pad  ;
	output \449GAT(176)_pad  ;
	output \450GAT(173)_pad  ;
	output \767GAT(349)_pad  ;
	output \768GAT(334)_pad  ;
	output \811GAT(378)  ;
	output \837GAT(396)  ;
	output \838GAT(395)  ;
	output \839GAT(394)  ;
	output \854GAT(419)  ;
	output \866GAT(426)_pad  ;
	output \867GAT(432)  ;
	output \868GAT(431)  ;
	output \869GAT(430)  ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\29GAT(5)_pad ,
		\36GAT(6)_pad ,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\42GAT(7)_pad ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\29GAT(5)_pad ,
		\75GAT(15)_pad ,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\42GAT(7)_pad ,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\80GAT(16)_pad ,
		_w61_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\85GAT(17)_pad ,
		\86GAT(18)_pad ,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\1GAT(0)_pad ,
		\26GAT(4)_pad ,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\51GAT(8)_pad ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\13GAT(2)_pad ,
		\17GAT(3)_pad ,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\1GAT(0)_pad ,
		\8GAT(1)_pad ,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w69_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w67_,
		_w69_,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		_w62_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\59GAT(10)_pad ,
		\75GAT(15)_pad ,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\80GAT(16)_pad ,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\36GAT(6)_pad ,
		\59GAT(10)_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\80GAT(16)_pad ,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\42GAT(7)_pad ,
		_w76_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\87GAT(19)_pad ,
		\88GAT(20)_pad ,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\90GAT(22)_pad ,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w62_,
		_w72_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\13GAT(2)_pad ,
		\55GAT(9)_pad ,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w70_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\29GAT(5)_pad ,
		\68GAT(11)_pad ,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\59GAT(10)_pad ,
		\68GAT(11)_pad ,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w83_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\74GAT(14)_pad ,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\89GAT(21)_pad ,
		_w79_,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\111GAT(27)_pad ,
		\91GAT(23)_pad ,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		\111GAT(27)_pad ,
		\91GAT(23)_pad ,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w90_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\126GAT(30)_pad ,
		\96GAT(24)_pad ,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\126GAT(30)_pad ,
		\96GAT(24)_pad ,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w93_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		_w92_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w92_,
		_w95_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\101GAT(25)_pad ,
		\121GAT(29)_pad ,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\101GAT(25)_pad ,
		\121GAT(29)_pad ,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w99_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		\116GAT(28)_pad ,
		\135GAT(32)_pad ,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		\116GAT(28)_pad ,
		\135GAT(32)_pad ,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w102_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w101_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w101_,
		_w104_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		\106GAT(26)_pad ,
		\130GAT(31)_pad ,
		_w108_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\106GAT(26)_pad ,
		\130GAT(31)_pad ,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w108_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		_w107_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w107_,
		_w110_,
		_w112_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w111_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w98_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w98_,
		_w113_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w114_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\171GAT(42)_pad ,
		\177GAT(43)_pad ,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\171GAT(42)_pad ,
		\177GAT(43)_pad ,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w117_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\130GAT(31)_pad ,
		\183GAT(44)_pad ,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\130GAT(31)_pad ,
		\183GAT(44)_pad ,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		_w119_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		_w119_,
		_w122_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\159GAT(40)_pad ,
		\195GAT(46)_pad ,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\159GAT(40)_pad ,
		\195GAT(46)_pad ,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w126_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\189GAT(45)_pad ,
		\207GAT(48)_pad ,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		\189GAT(45)_pad ,
		\207GAT(48)_pad ,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w128_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w128_,
		_w131_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		\165GAT(41)_pad ,
		\201GAT(47)_pad ,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		\165GAT(41)_pad ,
		\201GAT(47)_pad ,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w135_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		_w134_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		_w134_,
		_w137_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w138_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w125_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w125_,
		_w140_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w141_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\42GAT(7)_pad ,
		\72GAT(12)_pad ,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\73GAT(13)_pad ,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w87_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		\201GAT(47)_pad ,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\17GAT(3)_pad ,
		\51GAT(8)_pad ,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\42GAT(7)_pad ,
		_w74_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w70_,
		_w148_,
		_w150_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w149_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\156GAT(39)_pad ,
		\59GAT(10)_pad ,
		_w152_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\17GAT(3)_pad ,
		\42GAT(7)_pad ,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		\17GAT(3)_pad ,
		\42GAT(7)_pad ,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w68_,
		_w152_,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w155_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w151_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\126GAT(30)_pad ,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\55GAT(9)_pad ,
		_w68_,
		_w160_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		\268GAT(59)_pad ,
		\80GAT(16)_pad ,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w63_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w160_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w67_,
		_w148_,
		_w164_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w152_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\1GAT(0)_pad ,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		\153GAT(38)_pad ,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w163_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w159_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		\201GAT(47)_pad ,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\201GAT(47)_pad ,
		_w169_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w170_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		\261GAT(57)_pad ,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		\261GAT(57)_pad ,
		_w171_,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w170_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\219GAT(50)_pad ,
		_w173_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		_w175_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\228GAT(51)_pad ,
		_w172_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\201GAT(47)_pad ,
		\237GAT(52)_pad ,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		\246GAT(53)_pad ,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w169_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		\121GAT(29)_pad ,
		\210GAT(49)_pad ,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\255GAT(54)_pad ,
		\267GAT(58)_pad ,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		_w147_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w181_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		_w178_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		_w177_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\183GAT(44)_pad ,
		_w146_,
		_w189_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		\111GAT(27)_pad ,
		_w158_,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		\143GAT(34)_pad ,
		_w166_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w163_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w190_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\183GAT(44)_pad ,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		\183GAT(44)_pad ,
		_w193_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		\121GAT(29)_pad ,
		_w158_,
		_w197_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		\149GAT(36)_pad ,
		_w166_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w163_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		_w197_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\195GAT(46)_pad ,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w170_,
		_w174_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w201_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		\195GAT(46)_pad ,
		_w200_,
		_w204_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		\116GAT(28)_pad ,
		_w158_,
		_w205_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\146GAT(35)_pad ,
		_w166_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w163_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		_w205_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		\189GAT(45)_pad ,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w204_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w203_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		\189GAT(45)_pad ,
		_w208_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w211_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w196_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h2)
	) name154 (
		_w196_,
		_w213_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\219GAT(50)_pad ,
		_w214_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\183GAT(44)_pad ,
		\237GAT(52)_pad ,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\246GAT(53)_pad ,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		_w193_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\106GAT(26)_pad ,
		\210GAT(49)_pad ,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\228GAT(51)_pad ,
		_w196_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w189_,
		_w221_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		_w220_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w222_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h4)
	) name165 (
		_w217_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w209_,
		_w212_,
		_w227_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		\228GAT(51)_pad ,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w202_,
		_w204_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w201_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		_w227_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		_w227_,
		_w230_,
		_w232_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\219GAT(50)_pad ,
		_w231_,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\189GAT(45)_pad ,
		\237GAT(52)_pad ,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		\246GAT(53)_pad ,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w208_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		\111GAT(27)_pad ,
		\210GAT(49)_pad ,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\189GAT(45)_pad ,
		_w146_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		\255GAT(54)_pad ,
		\259GAT(55)_pad ,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w238_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		_w239_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w237_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w228_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		_w234_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w201_,
		_w204_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		\228GAT(51)_pad ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		_w202_,
		_w246_,
		_w248_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		_w202_,
		_w246_,
		_w249_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		\219GAT(50)_pad ,
		_w248_,
		_w250_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w249_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		\116GAT(28)_pad ,
		\210GAT(49)_pad ,
		_w252_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\195GAT(46)_pad ,
		_w146_,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		\195GAT(46)_pad ,
		\237GAT(52)_pad ,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		\246GAT(53)_pad ,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w200_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\255GAT(54)_pad ,
		\260GAT(56)_pad ,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w252_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w253_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w256_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		_w247_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w251_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		\106GAT(26)_pad ,
		_w158_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		_w152_,
		_w160_,
		_w264_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		\153GAT(38)_pad ,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\138GAT(33)_pad ,
		\152GAT(37)_pad ,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w162_,
		_w164_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w266_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w265_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		_w263_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		\177GAT(43)_pad ,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		\177GAT(43)_pad ,
		_w270_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\228GAT(51)_pad ,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w194_,
		_w215_,
		_w275_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		_w273_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		_w273_,
		_w275_,
		_w277_
	);
	LUT2 #(
		.INIT('h2)
	) name217 (
		\219GAT(50)_pad ,
		_w276_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\177GAT(43)_pad ,
		\237GAT(52)_pad ,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		\246GAT(53)_pad ,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w270_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		\177GAT(43)_pad ,
		_w146_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\101GAT(25)_pad ,
		\210GAT(49)_pad ,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w283_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w282_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w274_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w279_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		\91GAT(23)_pad ,
		_w158_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		\138GAT(33)_pad ,
		\8GAT(1)_pad ,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		\143GAT(34)_pad ,
		_w264_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w267_,
		_w290_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		_w291_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w289_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		\159GAT(40)_pad ,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		\159GAT(40)_pad ,
		_w294_,
		_w296_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		\101GAT(25)_pad ,
		_w158_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		\138GAT(33)_pad ,
		\17GAT(3)_pad ,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\149GAT(36)_pad ,
		_w264_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w267_,
		_w298_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		_w297_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h2)
	) name242 (
		\171GAT(42)_pad ,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w272_,
		_w275_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w271_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h4)
	) name245 (
		_w303_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		\171GAT(42)_pad ,
		_w302_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		\96GAT(24)_pad ,
		_w158_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		\138GAT(33)_pad ,
		\51GAT(8)_pad ,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		\146GAT(35)_pad ,
		_w264_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w267_,
		_w309_,
		_w311_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		_w310_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w308_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h4)
	) name253 (
		\165GAT(41)_pad ,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		_w307_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name255 (
		_w306_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		\165GAT(41)_pad ,
		_w313_,
		_w317_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w316_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w296_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w295_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w295_,
		_w296_,
		_w321_
	);
	LUT2 #(
		.INIT('h4)
	) name261 (
		_w318_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		_w318_,
		_w321_,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\219GAT(50)_pad ,
		_w322_,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w323_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\228GAT(51)_pad ,
		_w321_,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		\159GAT(40)_pad ,
		\237GAT(52)_pad ,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		\246GAT(53)_pad ,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w294_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		\159GAT(40)_pad ,
		_w146_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		\210GAT(49)_pad ,
		\268GAT(59)_pad ,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w330_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		_w329_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w326_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h4)
	) name274 (
		_w325_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\165GAT(41)_pad ,
		_w146_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w314_,
		_w317_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w305_,
		_w307_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w303_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h4)
	) name279 (
		_w337_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		_w337_,
		_w339_,
		_w341_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		\219GAT(50)_pad ,
		_w340_,
		_w342_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w341_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		\165GAT(41)_pad ,
		\237GAT(52)_pad ,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		\246GAT(53)_pad ,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w313_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		\210GAT(49)_pad ,
		\91GAT(23)_pad ,
		_w347_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\228GAT(51)_pad ,
		_w337_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w336_,
		_w347_,
		_w349_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w346_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		_w348_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		_w343_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w303_,
		_w307_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		\228GAT(51)_pad ,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		_w305_,
		_w353_,
		_w355_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		_w305_,
		_w353_,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		\219GAT(50)_pad ,
		_w355_,
		_w357_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w356_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		\171GAT(42)_pad ,
		\237GAT(52)_pad ,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		\246GAT(53)_pad ,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w302_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		\171GAT(42)_pad ,
		_w146_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		\210GAT(49)_pad ,
		\96GAT(24)_pad ,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w362_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name304 (
		_w361_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w354_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		_w358_,
		_w366_,
		_w367_
	);
	assign \273GAT(103)  = _w62_ ;
	assign \388GAT(133)_pad  = _w64_ ;
	assign \389GAT(132)_pad  = _w65_ ;
	assign \391GAT(124)_pad  = _w66_ ;
	assign \393GAT(165)  = _w68_ ;
	assign \418GAT(168)_pad  = _w71_ ;
	assign \419GAT(164)_pad  = _w73_ ;
	assign \420GAT(158)_pad  = _w75_ ;
	assign \421GAT(162)_pad  = _w77_ ;
	assign \422GAT(161)_pad  = _w78_ ;
	assign \423GAT(155)_pad  = _w80_ ;
	assign \446GAT(183)_pad  = _w81_ ;
	assign \448GAT(179)_pad  = _w85_ ;
	assign \449GAT(176)_pad  = _w88_ ;
	assign \450GAT(173)_pad  = _w89_ ;
	assign \767GAT(349)_pad  = _w116_ ;
	assign \768GAT(334)_pad  = _w143_ ;
	assign \811GAT(378)  = _w188_ ;
	assign \837GAT(396)  = _w226_ ;
	assign \838GAT(395)  = _w245_ ;
	assign \839GAT(394)  = _w262_ ;
	assign \854GAT(419)  = _w288_ ;
	assign \866GAT(426)_pad  = _w320_ ;
	assign \867GAT(432)  = _w335_ ;
	assign \868GAT(431)  = _w352_ ;
	assign \869GAT(430)  = _w367_ ;
endmodule;