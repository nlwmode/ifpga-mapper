module top (\1(0)_pad , \107(12)_pad , \116(13)_pad , \124(14)_pad , \125(15)_pad , \128(16)_pad , \13(1)_pad , \132(17)_pad , \137(18)_pad , \143(19)_pad , \150(20)_pad , \159(21)_pad , \169(22)_pad , \1698(48)_pad , \179(23)_pad , \190(24)_pad , \20(2)_pad , \200(25)_pad , \213(26)_pad , \222(27)_pad , \223(28)_pad , \226(29)_pad , \232(30)_pad , \238(31)_pad , \244(32)_pad , \250(33)_pad , \257(34)_pad , \264(35)_pad , \270(36)_pad , \274(37)_pad , \283(38)_pad , \2897(49)_pad , \294(39)_pad , \303(40)_pad , \311(41)_pad , \317(42)_pad , \322(43)_pad , \326(44)_pad , \329(45)_pad , \33(3)_pad , \330(46)_pad , \343(47)_pad , \41(4)_pad , \45(5)_pad , \50(6)_pad , \58(7)_pad , \68(8)_pad , \77(9)_pad , \87(10)_pad , \97(11)_pad , \2690(1611) , \2709(1587) , \353(405)_pad , \355(399)_pad , \358(1161)_pad , \361(940)_pad , \364(1484)_pad , \367(1585)_pad , \369(1321)_pad , \372(1243)_pad , \381(1626)_pad , \384(1553)_pad , \387(1616)_pad , \390(1603)_pad , \393(1605)_pad , \396(1504)_pad , \399(1428)_pad , \402(1718)_pad , \404(1714) , \407(1657)_pad , \409(1670)_pad , \605(1186) );
	input \1(0)_pad  ;
	input \107(12)_pad  ;
	input \116(13)_pad  ;
	input \124(14)_pad  ;
	input \125(15)_pad  ;
	input \128(16)_pad  ;
	input \13(1)_pad  ;
	input \132(17)_pad  ;
	input \137(18)_pad  ;
	input \143(19)_pad  ;
	input \150(20)_pad  ;
	input \159(21)_pad  ;
	input \169(22)_pad  ;
	input \1698(48)_pad  ;
	input \179(23)_pad  ;
	input \190(24)_pad  ;
	input \20(2)_pad  ;
	input \200(25)_pad  ;
	input \213(26)_pad  ;
	input \222(27)_pad  ;
	input \223(28)_pad  ;
	input \226(29)_pad  ;
	input \232(30)_pad  ;
	input \238(31)_pad  ;
	input \244(32)_pad  ;
	input \250(33)_pad  ;
	input \257(34)_pad  ;
	input \264(35)_pad  ;
	input \270(36)_pad  ;
	input \274(37)_pad  ;
	input \283(38)_pad  ;
	input \2897(49)_pad  ;
	input \294(39)_pad  ;
	input \303(40)_pad  ;
	input \311(41)_pad  ;
	input \317(42)_pad  ;
	input \322(43)_pad  ;
	input \326(44)_pad  ;
	input \329(45)_pad  ;
	input \33(3)_pad  ;
	input \330(46)_pad  ;
	input \343(47)_pad  ;
	input \41(4)_pad  ;
	input \45(5)_pad  ;
	input \50(6)_pad  ;
	input \58(7)_pad  ;
	input \68(8)_pad  ;
	input \77(9)_pad  ;
	input \87(10)_pad  ;
	input \97(11)_pad  ;
	output \2690(1611)  ;
	output \2709(1587)  ;
	output \353(405)_pad  ;
	output \355(399)_pad  ;
	output \358(1161)_pad  ;
	output \361(940)_pad  ;
	output \364(1484)_pad  ;
	output \367(1585)_pad  ;
	output \369(1321)_pad  ;
	output \372(1243)_pad  ;
	output \381(1626)_pad  ;
	output \384(1553)_pad  ;
	output \387(1616)_pad  ;
	output \390(1603)_pad  ;
	output \393(1605)_pad  ;
	output \396(1504)_pad  ;
	output \399(1428)_pad  ;
	output \402(1718)_pad  ;
	output \404(1714)  ;
	output \407(1657)_pad  ;
	output \409(1670)_pad  ;
	output \605(1186)  ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	LUT4 #(
		.INIT('h0400)
	) name0 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\213(26)_pad ,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\343(47)_pad ,
		_w52_,
		_w53_
	);
	LUT4 #(
		.INIT('h1015)
	) name2 (
		\20(2)_pad ,
		\283(38)_pad ,
		\33(3)_pad ,
		\97(11)_pad ,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\1(0)_pad ,
		\20(2)_pad ,
		_w55_
	);
	LUT4 #(
		.INIT('h5777)
	) name4 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		\116(13)_pad ,
		\20(2)_pad ,
		_w57_
	);
	LUT3 #(
		.INIT('h01)
	) name6 (
		_w56_,
		_w57_,
		_w54_,
		_w58_
	);
	LUT4 #(
		.INIT('h1000)
	) name7 (
		\1(0)_pad ,
		\116(13)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		_w59_
	);
	LUT4 #(
		.INIT('h0237)
	) name8 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		_w60_
	);
	LUT3 #(
		.INIT('h07)
	) name9 (
		\116(13)_pad ,
		_w60_,
		_w59_,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		_w58_,
		_w61_,
		_w62_
	);
	LUT4 #(
		.INIT('h0888)
	) name11 (
		\1(0)_pad ,
		\13(1)_pad ,
		\33(3)_pad ,
		\41(4)_pad ,
		_w63_
	);
	LUT3 #(
		.INIT('h10)
	) name12 (
		\1(0)_pad ,
		\41(4)_pad ,
		\45(5)_pad ,
		_w64_
	);
	LUT3 #(
		.INIT('h20)
	) name13 (
		\274(37)_pad ,
		_w63_,
		_w64_,
		_w65_
	);
	LUT3 #(
		.INIT('h04)
	) name14 (
		\1698(48)_pad ,
		\257(34)_pad ,
		\33(3)_pad ,
		_w66_
	);
	LUT4 #(
		.INIT('h0f77)
	) name15 (
		\1698(48)_pad ,
		\264(35)_pad ,
		\303(40)_pad ,
		\33(3)_pad ,
		_w67_
	);
	LUT3 #(
		.INIT('h8a)
	) name16 (
		_w63_,
		_w66_,
		_w67_,
		_w68_
	);
	LUT3 #(
		.INIT('h02)
	) name17 (
		\270(36)_pad ,
		_w63_,
		_w64_,
		_w69_
	);
	LUT3 #(
		.INIT('h01)
	) name18 (
		_w65_,
		_w68_,
		_w69_,
		_w70_
	);
	LUT4 #(
		.INIT('haaa8)
	) name19 (
		\169(22)_pad ,
		_w65_,
		_w68_,
		_w69_,
		_w71_
	);
	LUT4 #(
		.INIT('h0002)
	) name20 (
		\179(23)_pad ,
		_w65_,
		_w68_,
		_w69_,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w71_,
		_w72_,
		_w73_
	);
	LUT3 #(
		.INIT('h54)
	) name22 (
		_w62_,
		_w71_,
		_w72_,
		_w74_
	);
	LUT4 #(
		.INIT('h0002)
	) name23 (
		\190(24)_pad ,
		_w65_,
		_w68_,
		_w69_,
		_w75_
	);
	LUT4 #(
		.INIT('haaa8)
	) name24 (
		\200(25)_pad ,
		_w65_,
		_w68_,
		_w69_,
		_w76_
	);
	LUT3 #(
		.INIT('h02)
	) name25 (
		_w62_,
		_w76_,
		_w75_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w74_,
		_w77_,
		_w78_
	);
	LUT3 #(
		.INIT('h08)
	) name27 (
		\1698(48)_pad ,
		\244(32)_pad ,
		\33(3)_pad ,
		_w79_
	);
	LUT4 #(
		.INIT('h55cf)
	) name28 (
		\116(13)_pad ,
		\1698(48)_pad ,
		\238(31)_pad ,
		\33(3)_pad ,
		_w80_
	);
	LUT3 #(
		.INIT('h8a)
	) name29 (
		_w63_,
		_w79_,
		_w80_,
		_w81_
	);
	LUT3 #(
		.INIT('h10)
	) name30 (
		\1(0)_pad ,
		\274(37)_pad ,
		\45(5)_pad ,
		_w82_
	);
	LUT3 #(
		.INIT('h23)
	) name31 (
		\1(0)_pad ,
		\250(33)_pad ,
		\45(5)_pad ,
		_w83_
	);
	LUT3 #(
		.INIT('h01)
	) name32 (
		_w63_,
		_w83_,
		_w82_,
		_w84_
	);
	LUT3 #(
		.INIT('h02)
	) name33 (
		\179(23)_pad ,
		_w81_,
		_w84_,
		_w85_
	);
	LUT4 #(
		.INIT('h5553)
	) name34 (
		\169(22)_pad ,
		\179(23)_pad ,
		_w81_,
		_w84_,
		_w86_
	);
	LUT4 #(
		.INIT('hccc8)
	) name35 (
		\107(12)_pad ,
		\20(2)_pad ,
		\87(10)_pad ,
		\97(11)_pad ,
		_w87_
	);
	LUT4 #(
		.INIT('h23ef)
	) name36 (
		\20(2)_pad ,
		\33(3)_pad ,
		\68(8)_pad ,
		\97(11)_pad ,
		_w88_
	);
	LUT3 #(
		.INIT('h45)
	) name37 (
		_w56_,
		_w87_,
		_w88_,
		_w89_
	);
	LUT4 #(
		.INIT('h0040)
	) name38 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\87(10)_pad ,
		_w90_
	);
	LUT3 #(
		.INIT('h13)
	) name39 (
		\87(10)_pad ,
		_w90_,
		_w60_,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		_w89_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w86_,
		_w92_,
		_w93_
	);
	LUT3 #(
		.INIT('ha8)
	) name42 (
		\200(25)_pad ,
		_w81_,
		_w84_,
		_w94_
	);
	LUT3 #(
		.INIT('h02)
	) name43 (
		\190(24)_pad ,
		_w81_,
		_w84_,
		_w95_
	);
	LUT3 #(
		.INIT('h02)
	) name44 (
		_w92_,
		_w95_,
		_w94_,
		_w96_
	);
	LUT4 #(
		.INIT('heee2)
	) name45 (
		_w86_,
		_w92_,
		_w95_,
		_w94_,
		_w97_
	);
	LUT3 #(
		.INIT('h04)
	) name46 (
		\1698(48)_pad ,
		\250(33)_pad ,
		\33(3)_pad ,
		_w98_
	);
	LUT4 #(
		.INIT('h0f77)
	) name47 (
		\1698(48)_pad ,
		\257(34)_pad ,
		\294(39)_pad ,
		\33(3)_pad ,
		_w99_
	);
	LUT3 #(
		.INIT('h8a)
	) name48 (
		_w63_,
		_w98_,
		_w99_,
		_w100_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name49 (
		\264(35)_pad ,
		\274(37)_pad ,
		_w63_,
		_w64_,
		_w101_
	);
	LUT3 #(
		.INIT('h8a)
	) name50 (
		\200(25)_pad ,
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\107(12)_pad ,
		_w60_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\13(1)_pad ,
		\33(3)_pad ,
		_w104_
	);
	LUT4 #(
		.INIT('h1f3f)
	) name53 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		_w105_
	);
	LUT4 #(
		.INIT('h2320)
	) name54 (
		\116(13)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		\87(10)_pad ,
		_w106_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name55 (
		\107(12)_pad ,
		_w56_,
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w103_,
		_w107_,
		_w108_
	);
	LUT3 #(
		.INIT('h20)
	) name57 (
		\190(24)_pad ,
		_w100_,
		_w101_,
		_w109_
	);
	LUT3 #(
		.INIT('h02)
	) name58 (
		_w108_,
		_w109_,
		_w102_,
		_w110_
	);
	LUT3 #(
		.INIT('h08)
	) name59 (
		\1698(48)_pad ,
		\250(33)_pad ,
		\33(3)_pad ,
		_w111_
	);
	LUT4 #(
		.INIT('h0fbb)
	) name60 (
		\1698(48)_pad ,
		\244(32)_pad ,
		\283(38)_pad ,
		\33(3)_pad ,
		_w112_
	);
	LUT3 #(
		.INIT('h8a)
	) name61 (
		_w63_,
		_w111_,
		_w112_,
		_w113_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name62 (
		\257(34)_pad ,
		\274(37)_pad ,
		_w63_,
		_w64_,
		_w114_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		_w113_,
		_w114_,
		_w115_
	);
	LUT3 #(
		.INIT('h8a)
	) name64 (
		\200(25)_pad ,
		_w113_,
		_w114_,
		_w116_
	);
	LUT3 #(
		.INIT('h20)
	) name65 (
		\190(24)_pad ,
		_w113_,
		_w114_,
		_w117_
	);
	LUT3 #(
		.INIT('h48)
	) name66 (
		\107(12)_pad ,
		\20(2)_pad ,
		\97(11)_pad ,
		_w118_
	);
	LUT4 #(
		.INIT('h1013)
	) name67 (
		\107(12)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		\77(9)_pad ,
		_w119_
	);
	LUT3 #(
		.INIT('h01)
	) name68 (
		_w56_,
		_w119_,
		_w118_,
		_w120_
	);
	LUT4 #(
		.INIT('h0040)
	) name69 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\97(11)_pad ,
		_w121_
	);
	LUT3 #(
		.INIT('h07)
	) name70 (
		\97(11)_pad ,
		_w60_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w120_,
		_w122_,
		_w123_
	);
	LUT3 #(
		.INIT('h04)
	) name72 (
		_w117_,
		_w123_,
		_w116_,
		_w124_
	);
	LUT3 #(
		.INIT('h10)
	) name73 (
		\179(23)_pad ,
		_w100_,
		_w101_,
		_w125_
	);
	LUT3 #(
		.INIT('h45)
	) name74 (
		\169(22)_pad ,
		_w100_,
		_w101_,
		_w126_
	);
	LUT3 #(
		.INIT('h01)
	) name75 (
		_w108_,
		_w126_,
		_w125_,
		_w127_
	);
	LUT3 #(
		.INIT('h10)
	) name76 (
		\179(23)_pad ,
		_w113_,
		_w114_,
		_w128_
	);
	LUT3 #(
		.INIT('h45)
	) name77 (
		\169(22)_pad ,
		_w113_,
		_w114_,
		_w129_
	);
	LUT3 #(
		.INIT('h01)
	) name78 (
		_w123_,
		_w129_,
		_w128_,
		_w130_
	);
	LUT4 #(
		.INIT('h0001)
	) name79 (
		_w127_,
		_w110_,
		_w124_,
		_w130_,
		_w131_
	);
	LUT3 #(
		.INIT('h80)
	) name80 (
		_w78_,
		_w97_,
		_w131_,
		_w132_
	);
	LUT4 #(
		.INIT('h1555)
	) name81 (
		_w53_,
		_w78_,
		_w97_,
		_w131_,
		_w133_
	);
	LUT3 #(
		.INIT('h54)
	) name82 (
		\179(23)_pad ,
		_w81_,
		_w84_,
		_w134_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name83 (
		_w100_,
		_w101_,
		_w113_,
		_w114_,
		_w135_
	);
	LUT3 #(
		.INIT('h40)
	) name84 (
		_w70_,
		_w134_,
		_w135_,
		_w136_
	);
	LUT4 #(
		.INIT('h0100)
	) name85 (
		_w68_,
		_w69_,
		_w100_,
		_w101_,
		_w137_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name86 (
		_w53_,
		_w85_,
		_w115_,
		_w137_,
		_w138_
	);
	LUT3 #(
		.INIT('h8a)
	) name87 (
		\330(46)_pad ,
		_w136_,
		_w138_,
		_w139_
	);
	LUT4 #(
		.INIT('h000e)
	) name88 (
		_w74_,
		_w127_,
		_w110_,
		_w124_,
		_w140_
	);
	LUT4 #(
		.INIT('h5501)
	) name89 (
		_w93_,
		_w140_,
		_w130_,
		_w96_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w53_,
		_w141_,
		_w142_
	);
	LUT4 #(
		.INIT('h04ee)
	) name91 (
		_w53_,
		_w141_,
		_w132_,
		_w139_,
		_w143_
	);
	LUT3 #(
		.INIT('h08)
	) name92 (
		\1698(48)_pad ,
		\232(30)_pad ,
		\33(3)_pad ,
		_w144_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name93 (
		\1698(48)_pad ,
		\226(29)_pad ,
		\33(3)_pad ,
		\97(11)_pad ,
		_w145_
	);
	LUT3 #(
		.INIT('h8a)
	) name94 (
		_w63_,
		_w144_,
		_w145_,
		_w146_
	);
	LUT3 #(
		.INIT('h54)
	) name95 (
		\1(0)_pad ,
		\41(4)_pad ,
		\45(5)_pad ,
		_w147_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name96 (
		\238(31)_pad ,
		\274(37)_pad ,
		_w63_,
		_w147_,
		_w148_
	);
	LUT3 #(
		.INIT('h10)
	) name97 (
		\179(23)_pad ,
		_w146_,
		_w148_,
		_w149_
	);
	LUT4 #(
		.INIT('h0727)
	) name98 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\68(8)_pad ,
		_w150_,
		_w151_
	);
	LUT4 #(
		.INIT('h5410)
	) name100 (
		\20(2)_pad ,
		\33(3)_pad ,
		\50(6)_pad ,
		\77(9)_pad ,
		_w152_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name101 (
		\68(8)_pad ,
		_w56_,
		_w105_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w151_,
		_w153_,
		_w154_
	);
	LUT3 #(
		.INIT('h45)
	) name103 (
		\169(22)_pad ,
		_w146_,
		_w148_,
		_w155_
	);
	LUT3 #(
		.INIT('h01)
	) name104 (
		_w154_,
		_w155_,
		_w149_,
		_w156_
	);
	LUT3 #(
		.INIT('h8a)
	) name105 (
		\200(25)_pad ,
		_w146_,
		_w148_,
		_w157_
	);
	LUT3 #(
		.INIT('h20)
	) name106 (
		\190(24)_pad ,
		_w146_,
		_w148_,
		_w158_
	);
	LUT3 #(
		.INIT('h02)
	) name107 (
		_w154_,
		_w158_,
		_w157_,
		_w159_
	);
	LUT3 #(
		.INIT('h08)
	) name108 (
		\1698(48)_pad ,
		\226(29)_pad ,
		\33(3)_pad ,
		_w160_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name109 (
		\1698(48)_pad ,
		\223(28)_pad ,
		\33(3)_pad ,
		\87(10)_pad ,
		_w161_
	);
	LUT3 #(
		.INIT('h8a)
	) name110 (
		_w63_,
		_w160_,
		_w161_,
		_w162_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name111 (
		\232(30)_pad ,
		\274(37)_pad ,
		_w63_,
		_w147_,
		_w163_
	);
	LUT3 #(
		.INIT('h10)
	) name112 (
		\179(23)_pad ,
		_w162_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\58(7)_pad ,
		_w150_,
		_w165_
	);
	LUT3 #(
		.INIT('h82)
	) name114 (
		\20(2)_pad ,
		\58(7)_pad ,
		\68(8)_pad ,
		_w166_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name115 (
		\159(21)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		\68(8)_pad ,
		_w167_
	);
	LUT4 #(
		.INIT('h0040)
	) name116 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\58(7)_pad ,
		_w168_
	);
	LUT4 #(
		.INIT('h00ba)
	) name117 (
		_w56_,
		_w166_,
		_w167_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w165_,
		_w169_,
		_w170_
	);
	LUT3 #(
		.INIT('h45)
	) name119 (
		\169(22)_pad ,
		_w162_,
		_w163_,
		_w171_
	);
	LUT3 #(
		.INIT('h01)
	) name120 (
		_w170_,
		_w171_,
		_w164_,
		_w172_
	);
	LUT3 #(
		.INIT('h8a)
	) name121 (
		\200(25)_pad ,
		_w162_,
		_w163_,
		_w173_
	);
	LUT3 #(
		.INIT('h20)
	) name122 (
		\190(24)_pad ,
		_w162_,
		_w163_,
		_w174_
	);
	LUT3 #(
		.INIT('h02)
	) name123 (
		_w170_,
		_w174_,
		_w173_,
		_w175_
	);
	LUT4 #(
		.INIT('h0001)
	) name124 (
		_w172_,
		_w156_,
		_w159_,
		_w175_,
		_w176_
	);
	LUT3 #(
		.INIT('h08)
	) name125 (
		\1698(48)_pad ,
		\238(31)_pad ,
		\33(3)_pad ,
		_w177_
	);
	LUT4 #(
		.INIT('h55cf)
	) name126 (
		\107(12)_pad ,
		\1698(48)_pad ,
		\232(30)_pad ,
		\33(3)_pad ,
		_w178_
	);
	LUT3 #(
		.INIT('h8a)
	) name127 (
		_w63_,
		_w177_,
		_w178_,
		_w179_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name128 (
		\244(32)_pad ,
		\274(37)_pad ,
		_w63_,
		_w147_,
		_w180_
	);
	LUT3 #(
		.INIT('h10)
	) name129 (
		\179(23)_pad ,
		_w179_,
		_w180_,
		_w181_
	);
	LUT4 #(
		.INIT('h0145)
	) name130 (
		\20(2)_pad ,
		\33(3)_pad ,
		\58(7)_pad ,
		\87(10)_pad ,
		_w182_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		\20(2)_pad ,
		\77(9)_pad ,
		_w183_
	);
	LUT3 #(
		.INIT('h01)
	) name132 (
		_w56_,
		_w183_,
		_w182_,
		_w184_
	);
	LUT4 #(
		.INIT('h0040)
	) name133 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\77(9)_pad ,
		_w185_
	);
	LUT3 #(
		.INIT('h07)
	) name134 (
		\77(9)_pad ,
		_w150_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w184_,
		_w186_,
		_w187_
	);
	LUT3 #(
		.INIT('h45)
	) name136 (
		\169(22)_pad ,
		_w179_,
		_w180_,
		_w188_
	);
	LUT3 #(
		.INIT('h01)
	) name137 (
		_w187_,
		_w188_,
		_w181_,
		_w189_
	);
	LUT3 #(
		.INIT('h20)
	) name138 (
		\190(24)_pad ,
		_w179_,
		_w180_,
		_w190_
	);
	LUT3 #(
		.INIT('h8a)
	) name139 (
		\200(25)_pad ,
		_w179_,
		_w180_,
		_w191_
	);
	LUT3 #(
		.INIT('h02)
	) name140 (
		_w187_,
		_w191_,
		_w190_,
		_w192_
	);
	LUT3 #(
		.INIT('h08)
	) name141 (
		\1698(48)_pad ,
		\223(28)_pad ,
		\33(3)_pad ,
		_w193_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name142 (
		\1698(48)_pad ,
		\222(27)_pad ,
		\33(3)_pad ,
		\77(9)_pad ,
		_w194_
	);
	LUT3 #(
		.INIT('h8a)
	) name143 (
		_w63_,
		_w193_,
		_w194_,
		_w195_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name144 (
		\226(29)_pad ,
		\274(37)_pad ,
		_w63_,
		_w147_,
		_w196_
	);
	LUT3 #(
		.INIT('h10)
	) name145 (
		\179(23)_pad ,
		_w195_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\50(6)_pad ,
		_w150_,
		_w198_
	);
	LUT4 #(
		.INIT('haaa8)
	) name147 (
		\20(2)_pad ,
		\50(6)_pad ,
		\58(7)_pad ,
		\68(8)_pad ,
		_w199_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name148 (
		\150(20)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		\58(7)_pad ,
		_w200_
	);
	LUT4 #(
		.INIT('h0040)
	) name149 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\50(6)_pad ,
		_w201_
	);
	LUT4 #(
		.INIT('h00ba)
	) name150 (
		_w56_,
		_w199_,
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		_w198_,
		_w202_,
		_w203_
	);
	LUT3 #(
		.INIT('h45)
	) name152 (
		\169(22)_pad ,
		_w195_,
		_w196_,
		_w204_
	);
	LUT3 #(
		.INIT('h01)
	) name153 (
		_w203_,
		_w204_,
		_w197_,
		_w205_
	);
	LUT3 #(
		.INIT('h8a)
	) name154 (
		\200(25)_pad ,
		_w195_,
		_w196_,
		_w206_
	);
	LUT3 #(
		.INIT('h20)
	) name155 (
		\190(24)_pad ,
		_w195_,
		_w196_,
		_w207_
	);
	LUT3 #(
		.INIT('h02)
	) name156 (
		_w203_,
		_w207_,
		_w206_,
		_w208_
	);
	LUT4 #(
		.INIT('h0001)
	) name157 (
		_w189_,
		_w192_,
		_w205_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w176_,
		_w209_,
		_w210_
	);
	LUT4 #(
		.INIT('h00ba)
	) name159 (
		_w156_,
		_w159_,
		_w189_,
		_w175_,
		_w211_
	);
	LUT4 #(
		.INIT('h3031)
	) name160 (
		_w172_,
		_w205_,
		_w208_,
		_w211_,
		_w212_
	);
	LUT3 #(
		.INIT('hb0)
	) name161 (
		_w143_,
		_w210_,
		_w212_,
		_w213_
	);
	LUT3 #(
		.INIT('h8a)
	) name162 (
		_w53_,
		_w151_,
		_w153_,
		_w214_
	);
	LUT3 #(
		.INIT('h01)
	) name163 (
		_w156_,
		_w159_,
		_w214_,
		_w215_
	);
	LUT4 #(
		.INIT('h5f52)
	) name164 (
		_w53_,
		_w154_,
		_w156_,
		_w159_,
		_w216_
	);
	LUT3 #(
		.INIT('h8a)
	) name165 (
		_w53_,
		_w184_,
		_w186_,
		_w217_
	);
	LUT3 #(
		.INIT('h01)
	) name166 (
		_w189_,
		_w217_,
		_w192_,
		_w218_
	);
	LUT4 #(
		.INIT('h5f52)
	) name167 (
		_w53_,
		_w187_,
		_w189_,
		_w192_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w219_,
		_w216_,
		_w220_
	);
	LUT4 #(
		.INIT('h04fb)
	) name169 (
		_w133_,
		_w139_,
		_w219_,
		_w216_,
		_w221_
	);
	LUT4 #(
		.INIT('h4544)
	) name170 (
		_w53_,
		_w189_,
		_w141_,
		_w218_,
		_w222_
	);
	LUT2 #(
		.INIT('h9)
	) name171 (
		_w221_,
		_w222_,
		_w223_
	);
	LUT4 #(
		.INIT('h8a88)
	) name172 (
		_w215_,
		_w189_,
		_w141_,
		_w218_,
		_w224_
	);
	LUT4 #(
		.INIT('h0001)
	) name173 (
		_w52_,
		_w170_,
		_w171_,
		_w164_,
		_w225_
	);
	LUT3 #(
		.INIT('h8a)
	) name174 (
		_w52_,
		_w165_,
		_w169_,
		_w226_
	);
	LUT4 #(
		.INIT('h3331)
	) name175 (
		_w170_,
		_w226_,
		_w174_,
		_w173_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w172_,
		_w227_,
		_w228_
	);
	LUT3 #(
		.INIT('h32)
	) name177 (
		_w172_,
		_w225_,
		_w227_,
		_w229_
	);
	LUT3 #(
		.INIT('h02)
	) name178 (
		_w229_,
		_w219_,
		_w216_,
		_w230_
	);
	LUT4 #(
		.INIT('hb4f0)
	) name179 (
		_w133_,
		_w139_,
		_w229_,
		_w220_,
		_w231_
	);
	LUT4 #(
		.INIT('h54ab)
	) name180 (
		_w53_,
		_w156_,
		_w224_,
		_w231_,
		_w232_
	);
	LUT3 #(
		.INIT('ha8)
	) name181 (
		_w213_,
		_w223_,
		_w232_,
		_w233_
	);
	LUT4 #(
		.INIT('h0054)
	) name182 (
		_w53_,
		_w156_,
		_w224_,
		_w228_,
		_w234_
	);
	LUT4 #(
		.INIT('h5f52)
	) name183 (
		_w52_,
		_w203_,
		_w205_,
		_w208_,
		_w235_
	);
	LUT4 #(
		.INIT('h6555)
	) name184 (
		_w235_,
		_w133_,
		_w139_,
		_w230_,
		_w236_
	);
	LUT3 #(
		.INIT('h20)
	) name185 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		_w237_
	);
	LUT4 #(
		.INIT('h0020)
	) name186 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\41(4)_pad ,
		_w238_
	);
	LUT4 #(
		.INIT('h1e00)
	) name187 (
		_w225_,
		_w234_,
		_w236_,
		_w238_,
		_w239_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name188 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\45(5)_pad ,
		_w240_
	);
	LUT4 #(
		.INIT('h001e)
	) name189 (
		_w225_,
		_w234_,
		_w236_,
		_w240_,
		_w241_
	);
	LUT4 #(
		.INIT('h8088)
	) name190 (
		\1(0)_pad ,
		\13(1)_pad ,
		\169(22)_pad ,
		\20(2)_pad ,
		_w242_
	);
	LUT3 #(
		.INIT('h08)
	) name191 (
		\179(23)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w243_
	);
	LUT4 #(
		.INIT('h0020)
	) name192 (
		\179(23)_pad ,
		\190(24)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		\87(10)_pad ,
		_w244_,
		_w245_
	);
	LUT4 #(
		.INIT('h8000)
	) name194 (
		\179(23)_pad ,
		\190(24)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w246_
	);
	LUT3 #(
		.INIT('h37)
	) name195 (
		\179(23)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w247_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		\190(24)_pad ,
		\20(2)_pad ,
		_w248_
	);
	LUT4 #(
		.INIT('h0f4f)
	) name197 (
		\179(23)_pad ,
		\190(24)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w249_
	);
	LUT4 #(
		.INIT('h135f)
	) name198 (
		\116(13)_pad ,
		\68(8)_pad ,
		_w246_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w245_,
		_w250_,
		_w251_
	);
	LUT3 #(
		.INIT('h40)
	) name200 (
		\179(23)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w252_
	);
	LUT4 #(
		.INIT('h1000)
	) name201 (
		\179(23)_pad ,
		\190(24)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w253_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		\33(3)_pad ,
		\41(4)_pad ,
		_w254_
	);
	LUT3 #(
		.INIT('h70)
	) name203 (
		\58(7)_pad ,
		_w253_,
		_w254_,
		_w255_
	);
	LUT4 #(
		.INIT('h0010)
	) name204 (
		\179(23)_pad ,
		\190(24)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w256_
	);
	LUT4 #(
		.INIT('h4000)
	) name205 (
		\179(23)_pad ,
		\190(24)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w257_
	);
	LUT4 #(
		.INIT('h135f)
	) name206 (
		\283(38)_pad ,
		\77(9)_pad ,
		_w256_,
		_w257_,
		_w258_
	);
	LUT4 #(
		.INIT('h2000)
	) name207 (
		\179(23)_pad ,
		\190(24)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w259_
	);
	LUT4 #(
		.INIT('h0080)
	) name208 (
		\179(23)_pad ,
		\190(24)_pad ,
		\20(2)_pad ,
		\200(25)_pad ,
		_w260_
	);
	LUT4 #(
		.INIT('h135f)
	) name209 (
		\107(12)_pad ,
		\97(11)_pad ,
		_w260_,
		_w259_,
		_w261_
	);
	LUT3 #(
		.INIT('h80)
	) name210 (
		_w255_,
		_w258_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		_w251_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name212 (
		\41(4)_pad ,
		\50(6)_pad ,
		_w264_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\159(21)_pad ,
		_w253_,
		_w265_
	);
	LUT4 #(
		.INIT('h135f)
	) name214 (
		\132(17)_pad ,
		\143(19)_pad ,
		_w259_,
		_w257_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		_w265_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		\33(3)_pad ,
		\41(4)_pad ,
		_w268_
	);
	LUT3 #(
		.INIT('h70)
	) name217 (
		\125(15)_pad ,
		_w246_,
		_w268_,
		_w269_
	);
	LUT4 #(
		.INIT('h153f)
	) name218 (
		\128(16)_pad ,
		\150(20)_pad ,
		_w249_,
		_w260_,
		_w270_
	);
	LUT4 #(
		.INIT('h135f)
	) name219 (
		\124(14)_pad ,
		\137(18)_pad ,
		_w256_,
		_w244_,
		_w271_
	);
	LUT3 #(
		.INIT('h80)
	) name220 (
		_w269_,
		_w270_,
		_w271_,
		_w272_
	);
	LUT3 #(
		.INIT('h15)
	) name221 (
		_w264_,
		_w267_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		_w240_,
		_w238_,
		_w274_
	);
	LUT3 #(
		.INIT('h01)
	) name223 (
		\50(6)_pad ,
		_w104_,
		_w242_,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		_w274_,
		_w275_,
		_w276_
	);
	LUT4 #(
		.INIT('h7500)
	) name225 (
		_w242_,
		_w263_,
		_w273_,
		_w276_,
		_w277_
	);
	LUT3 #(
		.INIT('h70)
	) name226 (
		_w104_,
		_w235_,
		_w277_,
		_w278_
	);
	LUT4 #(
		.INIT('h1011)
	) name227 (
		_w241_,
		_w278_,
		_w233_,
		_w239_,
		_w279_
	);
	LUT4 #(
		.INIT('hefee)
	) name228 (
		_w241_,
		_w278_,
		_w233_,
		_w239_,
		_w280_
	);
	LUT4 #(
		.INIT('h08a2)
	) name229 (
		_w238_,
		_w213_,
		_w223_,
		_w232_,
		_w281_
	);
	LUT4 #(
		.INIT('h4070)
	) name230 (
		_w52_,
		_w172_,
		_w104_,
		_w227_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		\159(21)_pad ,
		_w249_,
		_w283_
	);
	LUT4 #(
		.INIT('h135f)
	) name232 (
		\128(16)_pad ,
		\150(20)_pad ,
		_w246_,
		_w257_,
		_w284_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w283_,
		_w284_,
		_w285_
	);
	LUT3 #(
		.INIT('h13)
	) name234 (
		\137(18)_pad ,
		\33(3)_pad ,
		_w259_,
		_w286_
	);
	LUT4 #(
		.INIT('h135f)
	) name235 (
		\132(17)_pad ,
		\50(6)_pad ,
		_w260_,
		_w253_,
		_w287_
	);
	LUT4 #(
		.INIT('h135f)
	) name236 (
		\125(15)_pad ,
		\143(19)_pad ,
		_w256_,
		_w244_,
		_w288_
	);
	LUT3 #(
		.INIT('h80)
	) name237 (
		_w286_,
		_w287_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\283(38)_pad ,
		_w246_,
		_w290_
	);
	LUT4 #(
		.INIT('h153f)
	) name239 (
		\107(12)_pad ,
		\77(9)_pad ,
		_w249_,
		_w259_,
		_w291_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		_w290_,
		_w291_,
		_w292_
	);
	LUT3 #(
		.INIT('h2a)
	) name241 (
		\33(3)_pad ,
		\68(8)_pad ,
		_w253_,
		_w293_
	);
	LUT4 #(
		.INIT('h135f)
	) name242 (
		\294(39)_pad ,
		\87(10)_pad ,
		_w256_,
		_w257_,
		_w294_
	);
	LUT4 #(
		.INIT('h47ff)
	) name243 (
		\116(13)_pad ,
		\190(24)_pad ,
		\97(11)_pad ,
		_w243_,
		_w295_
	);
	LUT3 #(
		.INIT('h80)
	) name244 (
		_w293_,
		_w294_,
		_w295_,
		_w296_
	);
	LUT4 #(
		.INIT('h0777)
	) name245 (
		_w285_,
		_w289_,
		_w292_,
		_w296_,
		_w297_
	);
	LUT3 #(
		.INIT('h01)
	) name246 (
		\58(7)_pad ,
		_w104_,
		_w242_,
		_w298_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		_w274_,
		_w298_,
		_w299_
	);
	LUT3 #(
		.INIT('hd0)
	) name248 (
		_w242_,
		_w297_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		_w282_,
		_w300_,
		_w301_
	);
	LUT3 #(
		.INIT('h0e)
	) name250 (
		_w240_,
		_w232_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		_w281_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('hb)
	) name252 (
		_w281_,
		_w302_,
		_w304_
	);
	LUT4 #(
		.INIT('h0001)
	) name253 (
		\50(6)_pad ,
		\58(7)_pad ,
		\68(8)_pad ,
		\77(9)_pad ,
		_w305_
	);
	LUT3 #(
		.INIT('hc8)
	) name254 (
		\107(12)_pad ,
		\87(10)_pad ,
		\97(11)_pad ,
		_w306_
	);
	LUT3 #(
		.INIT('h37)
	) name255 (
		\107(12)_pad ,
		\87(10)_pad ,
		\97(11)_pad ,
		_w307_
	);
	LUT4 #(
		.INIT('h9669)
	) name256 (
		\250(33)_pad ,
		\257(34)_pad ,
		\264(35)_pad ,
		\270(36)_pad ,
		_w308_
	);
	LUT4 #(
		.INIT('h6996)
	) name257 (
		\226(29)_pad ,
		\232(30)_pad ,
		\238(31)_pad ,
		\244(32)_pad ,
		_w309_
	);
	LUT2 #(
		.INIT('h6)
	) name258 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT4 #(
		.INIT('h135f)
	) name259 (
		\107(12)_pad ,
		\116(13)_pad ,
		\264(35)_pad ,
		\270(36)_pad ,
		_w311_
	);
	LUT4 #(
		.INIT('h135f)
	) name260 (
		\238(31)_pad ,
		\257(34)_pad ,
		\68(8)_pad ,
		\97(11)_pad ,
		_w312_
	);
	LUT4 #(
		.INIT('h135f)
	) name261 (
		\226(29)_pad ,
		\232(30)_pad ,
		\50(6)_pad ,
		\58(7)_pad ,
		_w313_
	);
	LUT4 #(
		.INIT('h135f)
	) name262 (
		\244(32)_pad ,
		\250(33)_pad ,
		\77(9)_pad ,
		\87(10)_pad ,
		_w314_
	);
	LUT4 #(
		.INIT('h8000)
	) name263 (
		_w313_,
		_w314_,
		_w311_,
		_w312_,
		_w315_
	);
	LUT3 #(
		.INIT('ha8)
	) name264 (
		\50(6)_pad ,
		\58(7)_pad ,
		\68(8)_pad ,
		_w316_
	);
	LUT3 #(
		.INIT('h80)
	) name265 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		_w317_
	);
	LUT3 #(
		.INIT('ha8)
	) name266 (
		\250(33)_pad ,
		\257(34)_pad ,
		\264(35)_pad ,
		_w318_
	);
	LUT4 #(
		.INIT('h153f)
	) name267 (
		_w237_,
		_w316_,
		_w317_,
		_w318_,
		_w319_
	);
	LUT3 #(
		.INIT('he0)
	) name268 (
		_w55_,
		_w315_,
		_w319_,
		_w320_
	);
	LUT4 #(
		.INIT('h0001)
	) name269 (
		\107(12)_pad ,
		\116(13)_pad ,
		\87(10)_pad ,
		\97(11)_pad ,
		_w321_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name270 (
		\1(0)_pad ,
		_w238_,
		_w316_,
		_w321_,
		_w322_
	);
	LUT3 #(
		.INIT('h1f)
	) name271 (
		\1(0)_pad ,
		_w143_,
		_w322_,
		_w323_
	);
	LUT4 #(
		.INIT('h87af)
	) name272 (
		\50(6)_pad ,
		\58(7)_pad ,
		\68(8)_pad ,
		\77(9)_pad ,
		_w324_
	);
	LUT3 #(
		.INIT('h48)
	) name273 (
		\107(12)_pad ,
		\116(13)_pad ,
		\97(11)_pad ,
		_w325_
	);
	LUT4 #(
		.INIT('h72fa)
	) name274 (
		\13(1)_pad ,
		\20(2)_pad ,
		_w324_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		\1(0)_pad ,
		_w326_,
		_w327_
	);
	LUT4 #(
		.INIT('h0440)
	) name276 (
		_w133_,
		_w139_,
		_w230_,
		_w210_,
		_w328_
	);
	LUT3 #(
		.INIT('h1e)
	) name277 (
		_w225_,
		_w234_,
		_w328_,
		_w329_
	);
	LUT4 #(
		.INIT('hef00)
	) name278 (
		_w53_,
		_w141_,
		_w210_,
		_w212_,
		_w330_
	);
	LUT3 #(
		.INIT('ha2)
	) name279 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		_w331_
	);
	LUT4 #(
		.INIT('hbaab)
	) name280 (
		_w327_,
		_w331_,
		_w329_,
		_w330_,
		_w332_
	);
	LUT3 #(
		.INIT('h4f)
	) name281 (
		_w141_,
		_w210_,
		_w212_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w132_,
		_w210_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		\303(40)_pad ,
		_w256_,
		_w335_
	);
	LUT4 #(
		.INIT('h153f)
	) name284 (
		\116(13)_pad ,
		\283(38)_pad ,
		_w260_,
		_w259_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name285 (
		_w335_,
		_w336_,
		_w337_
	);
	LUT3 #(
		.INIT('h2a)
	) name286 (
		\33(3)_pad ,
		\87(10)_pad ,
		_w249_,
		_w338_
	);
	LUT4 #(
		.INIT('h1bff)
	) name287 (
		\190(24)_pad ,
		\77(9)_pad ,
		\97(11)_pad ,
		_w252_,
		_w339_
	);
	LUT4 #(
		.INIT('h153f)
	) name288 (
		\107(12)_pad ,
		\294(39)_pad ,
		_w246_,
		_w244_,
		_w340_
	);
	LUT3 #(
		.INIT('h80)
	) name289 (
		_w338_,
		_w339_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		\150(20)_pad ,
		_w244_,
		_w342_
	);
	LUT4 #(
		.INIT('h153f)
	) name291 (
		\143(19)_pad ,
		\50(6)_pad ,
		_w249_,
		_w259_,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name292 (
		_w342_,
		_w343_,
		_w344_
	);
	LUT3 #(
		.INIT('h15)
	) name293 (
		\33(3)_pad ,
		\58(7)_pad ,
		_w253_,
		_w345_
	);
	LUT4 #(
		.INIT('h135f)
	) name294 (
		\132(17)_pad ,
		\159(21)_pad ,
		_w246_,
		_w257_,
		_w346_
	);
	LUT4 #(
		.INIT('h153f)
	) name295 (
		\128(16)_pad ,
		\137(18)_pad ,
		_w260_,
		_w256_,
		_w347_
	);
	LUT3 #(
		.INIT('h80)
	) name296 (
		_w345_,
		_w346_,
		_w347_,
		_w348_
	);
	LUT4 #(
		.INIT('h0777)
	) name297 (
		_w337_,
		_w341_,
		_w344_,
		_w348_,
		_w349_
	);
	LUT3 #(
		.INIT('h01)
	) name298 (
		\68(8)_pad ,
		_w104_,
		_w242_,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		_w274_,
		_w350_,
		_w351_
	);
	LUT3 #(
		.INIT('hd0)
	) name300 (
		_w242_,
		_w349_,
		_w351_,
		_w352_
	);
	LUT3 #(
		.INIT('h70)
	) name301 (
		_w104_,
		_w216_,
		_w352_,
		_w353_
	);
	LUT4 #(
		.INIT('h00eb)
	) name302 (
		_w240_,
		_w221_,
		_w222_,
		_w353_,
		_w354_
	);
	LUT4 #(
		.INIT('h7d00)
	) name303 (
		_w238_,
		_w213_,
		_w223_,
		_w354_,
		_w355_
	);
	LUT4 #(
		.INIT('h82ff)
	) name304 (
		_w238_,
		_w213_,
		_w223_,
		_w354_,
		_w356_
	);
	LUT3 #(
		.INIT('h4b)
	) name305 (
		_w133_,
		_w139_,
		_w219_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\311(41)_pad ,
		_w256_,
		_w358_
	);
	LUT4 #(
		.INIT('h153f)
	) name307 (
		\283(38)_pad ,
		\294(39)_pad ,
		_w260_,
		_w259_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		_w358_,
		_w359_,
		_w360_
	);
	LUT3 #(
		.INIT('h2a)
	) name309 (
		\33(3)_pad ,
		\97(11)_pad ,
		_w249_,
		_w361_
	);
	LUT4 #(
		.INIT('h47ff)
	) name310 (
		\107(12)_pad ,
		\190(24)_pad ,
		\87(10)_pad ,
		_w252_,
		_w362_
	);
	LUT4 #(
		.INIT('h153f)
	) name311 (
		\116(13)_pad ,
		\303(40)_pad ,
		_w246_,
		_w244_,
		_w363_
	);
	LUT3 #(
		.INIT('h80)
	) name312 (
		_w361_,
		_w362_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		\159(21)_pad ,
		_w244_,
		_w365_
	);
	LUT4 #(
		.INIT('h153f)
	) name314 (
		\150(20)_pad ,
		\58(7)_pad ,
		_w249_,
		_w259_,
		_w366_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		_w365_,
		_w366_,
		_w367_
	);
	LUT3 #(
		.INIT('h15)
	) name316 (
		\33(3)_pad ,
		\68(8)_pad ,
		_w253_,
		_w368_
	);
	LUT4 #(
		.INIT('h135f)
	) name317 (
		\137(18)_pad ,
		\50(6)_pad ,
		_w246_,
		_w257_,
		_w369_
	);
	LUT4 #(
		.INIT('h153f)
	) name318 (
		\132(17)_pad ,
		\143(19)_pad ,
		_w260_,
		_w256_,
		_w370_
	);
	LUT3 #(
		.INIT('h80)
	) name319 (
		_w368_,
		_w369_,
		_w370_,
		_w371_
	);
	LUT4 #(
		.INIT('h0777)
	) name320 (
		_w360_,
		_w364_,
		_w367_,
		_w371_,
		_w372_
	);
	LUT3 #(
		.INIT('h01)
	) name321 (
		\77(9)_pad ,
		_w104_,
		_w242_,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		_w274_,
		_w373_,
		_w374_
	);
	LUT3 #(
		.INIT('hd0)
	) name323 (
		_w242_,
		_w372_,
		_w374_,
		_w375_
	);
	LUT3 #(
		.INIT('h70)
	) name324 (
		_w104_,
		_w219_,
		_w375_,
		_w376_
	);
	LUT4 #(
		.INIT('h00eb)
	) name325 (
		_w274_,
		_w142_,
		_w357_,
		_w376_,
		_w377_
	);
	LUT4 #(
		.INIT('hff14)
	) name326 (
		_w274_,
		_w142_,
		_w357_,
		_w376_,
		_w378_
	);
	LUT3 #(
		.INIT('h01)
	) name327 (
		\13(1)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		_w379_
	);
	LUT3 #(
		.INIT('h8a)
	) name328 (
		_w53_,
		_w89_,
		_w91_,
		_w380_
	);
	LUT3 #(
		.INIT('h02)
	) name329 (
		_w53_,
		_w86_,
		_w92_,
		_w381_
	);
	LUT3 #(
		.INIT('h0d)
	) name330 (
		_w97_,
		_w380_,
		_w381_,
		_w382_
	);
	LUT4 #(
		.INIT('h00c4)
	) name331 (
		_w97_,
		_w379_,
		_w380_,
		_w381_,
		_w383_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		\50(6)_pad ,
		_w244_,
		_w384_
	);
	LUT4 #(
		.INIT('h135f)
	) name333 (
		\150(20)_pad ,
		\58(7)_pad ,
		_w260_,
		_w257_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w384_,
		_w385_,
		_w386_
	);
	LUT3 #(
		.INIT('h15)
	) name335 (
		\33(3)_pad ,
		\68(8)_pad ,
		_w249_,
		_w387_
	);
	LUT4 #(
		.INIT('h135f)
	) name336 (
		\159(21)_pad ,
		\77(9)_pad ,
		_w259_,
		_w253_,
		_w388_
	);
	LUT4 #(
		.INIT('h153f)
	) name337 (
		\137(18)_pad ,
		\143(19)_pad ,
		_w246_,
		_w256_,
		_w389_
	);
	LUT3 #(
		.INIT('h80)
	) name338 (
		_w387_,
		_w388_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\107(12)_pad ,
		_w249_,
		_w391_
	);
	LUT4 #(
		.INIT('h153f)
	) name340 (
		\116(13)_pad ,
		\283(38)_pad ,
		_w244_,
		_w257_,
		_w392_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w391_,
		_w392_,
		_w393_
	);
	LUT3 #(
		.INIT('h4c)
	) name342 (
		\294(39)_pad ,
		\33(3)_pad ,
		_w259_,
		_w394_
	);
	LUT4 #(
		.INIT('h135f)
	) name343 (
		\311(41)_pad ,
		\97(11)_pad ,
		_w246_,
		_w253_,
		_w395_
	);
	LUT4 #(
		.INIT('h135f)
	) name344 (
		\303(40)_pad ,
		\317(42)_pad ,
		_w260_,
		_w256_,
		_w396_
	);
	LUT3 #(
		.INIT('h80)
	) name345 (
		_w394_,
		_w395_,
		_w396_,
		_w397_
	);
	LUT4 #(
		.INIT('h0777)
	) name346 (
		_w386_,
		_w390_,
		_w393_,
		_w397_,
		_w398_
	);
	LUT4 #(
		.INIT('h2000)
	) name347 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		_w399_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		_w308_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w242_,
		_w379_,
		_w401_
	);
	LUT4 #(
		.INIT('hdf00)
	) name350 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\87(10)_pad ,
		_w402_
	);
	LUT3 #(
		.INIT('h01)
	) name351 (
		_w242_,
		_w379_,
		_w402_,
		_w403_
	);
	LUT3 #(
		.INIT('h8a)
	) name352 (
		_w274_,
		_w400_,
		_w403_,
		_w404_
	);
	LUT3 #(
		.INIT('hd0)
	) name353 (
		_w242_,
		_w398_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		_w383_,
		_w405_,
		_w406_
	);
	LUT3 #(
		.INIT('h8a)
	) name355 (
		_w53_,
		_w58_,
		_w61_,
		_w407_
	);
	LUT4 #(
		.INIT('hccf1)
	) name356 (
		_w62_,
		_w73_,
		_w77_,
		_w407_,
		_w408_
	);
	LUT4 #(
		.INIT('h1110)
	) name357 (
		_w53_,
		_w62_,
		_w71_,
		_w72_,
		_w409_
	);
	LUT4 #(
		.INIT('h0001)
	) name358 (
		_w53_,
		_w108_,
		_w126_,
		_w125_,
		_w410_
	);
	LUT3 #(
		.INIT('h8a)
	) name359 (
		_w53_,
		_w103_,
		_w107_,
		_w411_
	);
	LUT4 #(
		.INIT('h00fd)
	) name360 (
		_w108_,
		_w109_,
		_w102_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w127_,
		_w412_,
		_w413_
	);
	LUT4 #(
		.INIT('h0407)
	) name362 (
		_w53_,
		_w127_,
		_w409_,
		_w412_,
		_w414_
	);
	LUT3 #(
		.INIT('h10)
	) name363 (
		_w127_,
		_w110_,
		_w409_,
		_w415_
	);
	LUT4 #(
		.INIT('hddd2)
	) name364 (
		\330(46)_pad ,
		_w408_,
		_w414_,
		_w415_,
		_w416_
	);
	LUT4 #(
		.INIT('h0001)
	) name365 (
		_w53_,
		_w123_,
		_w129_,
		_w128_,
		_w417_
	);
	LUT3 #(
		.INIT('h8a)
	) name366 (
		_w53_,
		_w120_,
		_w122_,
		_w418_
	);
	LUT4 #(
		.INIT('h00fb)
	) name367 (
		_w117_,
		_w123_,
		_w116_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w130_,
		_w419_,
		_w420_
	);
	LUT3 #(
		.INIT('h32)
	) name369 (
		_w130_,
		_w417_,
		_w419_,
		_w421_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name370 (
		\330(46)_pad ,
		_w408_,
		_w410_,
		_w413_,
		_w422_
	);
	LUT2 #(
		.INIT('hb)
	) name371 (
		_w415_,
		_w422_,
		_w423_
	);
	LUT3 #(
		.INIT('h96)
	) name372 (
		_w415_,
		_w421_,
		_w422_,
		_w424_
	);
	LUT4 #(
		.INIT('h222a)
	) name373 (
		_w238_,
		_w143_,
		_w416_,
		_w424_,
		_w425_
	);
	LUT4 #(
		.INIT('h3132)
	) name374 (
		_w415_,
		_w417_,
		_w420_,
		_w422_,
		_w426_
	);
	LUT2 #(
		.INIT('h6)
	) name375 (
		_w382_,
		_w426_,
		_w427_
	);
	LUT4 #(
		.INIT('h0233)
	) name376 (
		_w240_,
		_w406_,
		_w425_,
		_w427_,
		_w428_
	);
	LUT4 #(
		.INIT('hfdcc)
	) name377 (
		_w240_,
		_w406_,
		_w425_,
		_w427_,
		_w429_
	);
	LUT4 #(
		.INIT('h08a2)
	) name378 (
		_w238_,
		_w143_,
		_w416_,
		_w424_,
		_w430_
	);
	LUT4 #(
		.INIT('h1441)
	) name379 (
		_w240_,
		_w415_,
		_w421_,
		_w422_,
		_w431_
	);
	LUT4 #(
		.INIT('h4070)
	) name380 (
		_w53_,
		_w130_,
		_w379_,
		_w419_,
		_w432_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		\303(40)_pad ,
		_w259_,
		_w433_
	);
	LUT4 #(
		.INIT('h153f)
	) name382 (
		\311(41)_pad ,
		\317(42)_pad ,
		_w246_,
		_w260_,
		_w434_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		_w433_,
		_w434_,
		_w435_
	);
	LUT3 #(
		.INIT('h4c)
	) name384 (
		\116(13)_pad ,
		\33(3)_pad ,
		_w249_,
		_w436_
	);
	LUT4 #(
		.INIT('h153f)
	) name385 (
		\294(39)_pad ,
		\322(43)_pad ,
		_w256_,
		_w244_,
		_w437_
	);
	LUT4 #(
		.INIT('h1dff)
	) name386 (
		\107(12)_pad ,
		\190(24)_pad ,
		\283(38)_pad ,
		_w252_,
		_w438_
	);
	LUT3 #(
		.INIT('h80)
	) name387 (
		_w436_,
		_w437_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		\58(7)_pad ,
		_w244_,
		_w440_
	);
	LUT4 #(
		.INIT('h135f)
	) name389 (
		\159(21)_pad ,
		\68(8)_pad ,
		_w260_,
		_w257_,
		_w441_
	);
	LUT2 #(
		.INIT('h4)
	) name390 (
		_w440_,
		_w441_,
		_w442_
	);
	LUT3 #(
		.INIT('h15)
	) name391 (
		\33(3)_pad ,
		\77(9)_pad ,
		_w249_,
		_w443_
	);
	LUT4 #(
		.INIT('h135f)
	) name392 (
		\50(6)_pad ,
		\87(10)_pad ,
		_w259_,
		_w253_,
		_w444_
	);
	LUT4 #(
		.INIT('h153f)
	) name393 (
		\143(19)_pad ,
		\150(20)_pad ,
		_w246_,
		_w256_,
		_w445_
	);
	LUT3 #(
		.INIT('h80)
	) name394 (
		_w443_,
		_w444_,
		_w445_,
		_w446_
	);
	LUT4 #(
		.INIT('h0777)
	) name395 (
		_w435_,
		_w439_,
		_w442_,
		_w446_,
		_w447_
	);
	LUT4 #(
		.INIT('h6996)
	) name396 (
		\107(12)_pad ,
		\116(13)_pad ,
		\87(10)_pad ,
		\97(11)_pad ,
		_w448_
	);
	LUT2 #(
		.INIT('h2)
	) name397 (
		_w399_,
		_w448_,
		_w449_
	);
	LUT4 #(
		.INIT('hdf00)
	) name398 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\97(11)_pad ,
		_w450_
	);
	LUT3 #(
		.INIT('h01)
	) name399 (
		_w242_,
		_w379_,
		_w450_,
		_w451_
	);
	LUT3 #(
		.INIT('h8a)
	) name400 (
		_w274_,
		_w449_,
		_w451_,
		_w452_
	);
	LUT3 #(
		.INIT('hd0)
	) name401 (
		_w242_,
		_w447_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		_w432_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w431_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w430_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('hb)
	) name405 (
		_w430_,
		_w455_,
		_w457_
	);
	LUT4 #(
		.INIT('h4070)
	) name406 (
		_w53_,
		_w127_,
		_w379_,
		_w412_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		\159(21)_pad ,
		_w246_,
		_w459_
	);
	LUT4 #(
		.INIT('h153f)
	) name408 (
		\58(7)_pad ,
		\68(8)_pad ,
		_w244_,
		_w259_,
		_w460_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		_w459_,
		_w460_,
		_w461_
	);
	LUT3 #(
		.INIT('h15)
	) name410 (
		\33(3)_pad ,
		\77(9)_pad ,
		_w257_,
		_w462_
	);
	LUT4 #(
		.INIT('h135f)
	) name411 (
		\87(10)_pad ,
		\97(11)_pad ,
		_w249_,
		_w253_,
		_w463_
	);
	LUT4 #(
		.INIT('h153f)
	) name412 (
		\150(20)_pad ,
		\50(6)_pad ,
		_w260_,
		_w256_,
		_w464_
	);
	LUT3 #(
		.INIT('h80)
	) name413 (
		_w462_,
		_w463_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		\311(41)_pad ,
		_w259_,
		_w466_
	);
	LUT4 #(
		.INIT('h153f)
	) name415 (
		\294(39)_pad ,
		\322(43)_pad ,
		_w246_,
		_w257_,
		_w467_
	);
	LUT2 #(
		.INIT('h4)
	) name416 (
		_w466_,
		_w467_,
		_w468_
	);
	LUT3 #(
		.INIT('h4c)
	) name417 (
		\303(40)_pad ,
		\33(3)_pad ,
		_w244_,
		_w469_
	);
	LUT4 #(
		.INIT('h153f)
	) name418 (
		\116(13)_pad ,
		\317(42)_pad ,
		_w260_,
		_w253_,
		_w470_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name419 (
		\283(38)_pad ,
		\326(44)_pad ,
		_w247_,
		_w248_,
		_w471_
	);
	LUT3 #(
		.INIT('h80)
	) name420 (
		_w469_,
		_w470_,
		_w471_,
		_w472_
	);
	LUT4 #(
		.INIT('h0777)
	) name421 (
		_w461_,
		_w465_,
		_w468_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		\45(5)_pad ,
		_w309_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		\68(8)_pad ,
		\77(9)_pad ,
		_w475_
	);
	LUT3 #(
		.INIT('h10)
	) name424 (
		\45(5)_pad ,
		\50(6)_pad ,
		\58(7)_pad ,
		_w476_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name425 (
		_w321_,
		_w399_,
		_w475_,
		_w476_,
		_w477_
	);
	LUT4 #(
		.INIT('h3133)
	) name426 (
		\1(0)_pad ,
		\107(12)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		_w478_
	);
	LUT4 #(
		.INIT('h0020)
	) name427 (
		\1(0)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		\33(3)_pad ,
		_w479_
	);
	LUT3 #(
		.INIT('h23)
	) name428 (
		_w321_,
		_w478_,
		_w479_,
		_w480_
	);
	LUT4 #(
		.INIT('h20aa)
	) name429 (
		_w401_,
		_w474_,
		_w477_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		_w274_,
		_w481_,
		_w482_
	);
	LUT3 #(
		.INIT('hd0)
	) name431 (
		_w242_,
		_w473_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h4)
	) name432 (
		_w458_,
		_w483_,
		_w484_
	);
	LUT3 #(
		.INIT('h0e)
	) name433 (
		_w240_,
		_w416_,
		_w484_,
		_w485_
	);
	LUT4 #(
		.INIT('h7d00)
	) name434 (
		_w238_,
		_w143_,
		_w416_,
		_w485_,
		_w486_
	);
	LUT4 #(
		.INIT('h82ff)
	) name435 (
		_w238_,
		_w143_,
		_w416_,
		_w485_,
		_w487_
	);
	LUT3 #(
		.INIT('h21)
	) name436 (
		\330(46)_pad ,
		_w274_,
		_w408_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		\283(38)_pad ,
		_w253_,
		_w489_
	);
	LUT4 #(
		.INIT('h153f)
	) name438 (
		\303(40)_pad ,
		\326(44)_pad ,
		_w246_,
		_w257_,
		_w490_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w489_,
		_w490_,
		_w491_
	);
	LUT3 #(
		.INIT('h4c)
	) name440 (
		\322(43)_pad ,
		\33(3)_pad ,
		_w260_,
		_w492_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name441 (
		\294(39)_pad ,
		\329(45)_pad ,
		_w247_,
		_w248_,
		_w493_
	);
	LUT4 #(
		.INIT('h135f)
	) name442 (
		\311(41)_pad ,
		\317(42)_pad ,
		_w244_,
		_w259_,
		_w494_
	);
	LUT3 #(
		.INIT('h80)
	) name443 (
		_w492_,
		_w493_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		\50(6)_pad ,
		_w246_,
		_w496_
	);
	LUT4 #(
		.INIT('h27ff)
	) name445 (
		\190(24)_pad ,
		\58(7)_pad ,
		\77(9)_pad ,
		_w243_,
		_w497_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w496_,
		_w497_,
		_w498_
	);
	LUT3 #(
		.INIT('h15)
	) name447 (
		\33(3)_pad ,
		\87(10)_pad ,
		_w257_,
		_w499_
	);
	LUT4 #(
		.INIT('h153f)
	) name448 (
		\107(12)_pad ,
		\97(11)_pad ,
		_w249_,
		_w253_,
		_w500_
	);
	LUT4 #(
		.INIT('h135f)
	) name449 (
		\159(21)_pad ,
		\68(8)_pad ,
		_w256_,
		_w259_,
		_w501_
	);
	LUT3 #(
		.INIT('h80)
	) name450 (
		_w499_,
		_w500_,
		_w501_,
		_w502_
	);
	LUT4 #(
		.INIT('h0777)
	) name451 (
		_w491_,
		_w495_,
		_w498_,
		_w502_,
		_w503_
	);
	LUT4 #(
		.INIT('h9669)
	) name452 (
		\50(6)_pad ,
		\58(7)_pad ,
		\68(8)_pad ,
		\77(9)_pad ,
		_w504_
	);
	LUT4 #(
		.INIT('h10b0)
	) name453 (
		\45(5)_pad ,
		_w316_,
		_w399_,
		_w504_,
		_w505_
	);
	LUT4 #(
		.INIT('h3133)
	) name454 (
		\1(0)_pad ,
		\116(13)_pad ,
		\13(1)_pad ,
		\20(2)_pad ,
		_w506_
	);
	LUT3 #(
		.INIT('h0b)
	) name455 (
		_w306_,
		_w479_,
		_w506_,
		_w507_
	);
	LUT4 #(
		.INIT('h2a22)
	) name456 (
		_w274_,
		_w401_,
		_w505_,
		_w507_,
		_w508_
	);
	LUT3 #(
		.INIT('hd0)
	) name457 (
		_w242_,
		_w503_,
		_w508_,
		_w509_
	);
	LUT3 #(
		.INIT('h70)
	) name458 (
		_w379_,
		_w408_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w488_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('he)
	) name460 (
		_w488_,
		_w510_,
		_w512_
	);
	LUT2 #(
		.INIT('h9)
	) name461 (
		_w486_,
		_w511_,
		_w513_
	);
	LUT2 #(
		.INIT('h6)
	) name462 (
		_w428_,
		_w513_,
		_w514_
	);
	LUT3 #(
		.INIT('h96)
	) name463 (
		_w355_,
		_w377_,
		_w456_,
		_w515_
	);
	LUT2 #(
		.INIT('h6)
	) name464 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT4 #(
		.INIT('h6996)
	) name465 (
		_w279_,
		_w303_,
		_w514_,
		_w515_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		\213(26)_pad ,
		\343(47)_pad ,
		_w518_
	);
	LUT4 #(
		.INIT('haa3c)
	) name467 (
		\2897(49)_pad ,
		_w279_,
		_w303_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h6)
	) name468 (
		_w516_,
		_w519_,
		_w520_
	);
	LUT3 #(
		.INIT('h80)
	) name469 (
		_w377_,
		_w486_,
		_w511_,
		_w521_
	);
	LUT4 #(
		.INIT('h8000)
	) name470 (
		_w355_,
		_w428_,
		_w456_,
		_w521_,
		_w522_
	);
	LUT3 #(
		.INIT('h7f)
	) name471 (
		_w279_,
		_w303_,
		_w522_,
		_w523_
	);
	LUT3 #(
		.INIT('h80)
	) name472 (
		_w279_,
		_w303_,
		_w518_,
		_w524_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name473 (
		\213(26)_pad ,
		_w279_,
		_w303_,
		_w522_,
		_w525_
	);
	LUT2 #(
		.INIT('hb)
	) name474 (
		_w524_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h6)
	) name475 (
		_w448_,
		_w504_,
		_w527_
	);
	assign \2690(1611)  = _w280_ ;
	assign \2709(1587)  = _w304_ ;
	assign \353(405)_pad  = _w305_ ;
	assign \355(399)_pad  = _w307_ ;
	assign \358(1161)_pad  = _w310_ ;
	assign \361(940)_pad  = _w320_ ;
	assign \364(1484)_pad  = _w323_ ;
	assign \367(1585)_pad  = _w332_ ;
	assign \369(1321)_pad  = _w333_ ;
	assign \372(1243)_pad  = _w334_ ;
	assign \381(1626)_pad  = _w356_ ;
	assign \384(1553)_pad  = _w378_ ;
	assign \387(1616)_pad  = _w429_ ;
	assign \390(1603)_pad  = _w457_ ;
	assign \393(1605)_pad  = _w487_ ;
	assign \396(1504)_pad  = _w512_ ;
	assign \399(1428)_pad  = _w423_ ;
	assign \402(1718)_pad  = _w517_ ;
	assign \404(1714)  = _w520_ ;
	assign \407(1657)_pad  = _w523_ ;
	assign \409(1670)_pad  = _w526_ ;
	assign \605(1186)  = _w527_ ;
endmodule;