module top (\g102_pad , \g10_reg/NET0131 , \g11_reg/NET0131 , \g1293_pad , \g14_reg/NET0131 , \g15_reg/NET0131 , \g18_reg/NET0131 , \g197_reg/NET0131 , \g19_reg/NET0131 , \g1_reg/NET0131 , \g204_reg/NET0131 , \g205_reg/NET0131 , \g206_reg/NET0131 , \g207_reg/NET0131 , \g208_reg/NET0131 , \g209_reg/NET0131 , \g210_reg/NET0131 , \g211_reg/NET0131 , \g212_reg/NET0131 , \g218_reg/NET0131 , \g224_reg/NET0131 , \g230_reg/NET0131 , \g236_reg/NET0131 , \g242_reg/NET0131 , \g248_reg/NET0131 , \g24_reg/NET0131 , \g254_reg/NET0131 , \g25_reg/NET0131 , \g260_reg/NET0131 , \g266_reg/NET0131 , \g269_reg/NET0131 , \g276_reg/NET0131 , \g277_reg/NET0131 , \g278_reg/NET0131 , \g279_reg/NET0131 , \g280_reg/NET0131 , \g281_reg/NET0131 , \g282_reg/NET0131 , \g283_reg/NET0131 , \g28_reg/NET0131 , \g293_reg/NET0131 , \g297_reg/NET0131 , \g29_reg/NET0131 , \g2_reg/NET0131 , \g33_reg/NET0131 , \g3_reg/NET0131 , \g402_reg/NET0131 , \g406_reg/NET0131 , \g4099_pad , \g4100_pad , \g4101_pad , \g4102_pad , \g4103_pad , \g4104_pad , \g4105_pad , \g4108_pad , \g410_reg/NET0131 , \g4110_pad , \g4112_pad , \g414_reg/NET0131 , \g418_reg/NET0131 , \g422_reg/NET0131 , \g426_reg/NET0131 , \g430_reg/NET0131 , \g434_reg/NET0131 , \g437_reg/NET0131 , \g441_reg/NET0131 , \g4422_pad , \g445_reg/NET0131 , \g449_reg/NET0131 , \g453_reg/NET0131 , \g457_reg/NET0131 , \g461_reg/NET0131 , \g465_reg/NET0131 , \g471_reg/NET0131 , \g478_reg/NET0131 , \g486_reg/NET0131 , \g489_reg/NET0131 , \g48_reg/NET0131 , \g492_reg/NET0131 , \g496_reg/NET0131 , \g500_reg/NET0131 , \g504_reg/NET0131 , \g508_reg/NET0131 , \g512_reg/NET0131 , \g536_reg/NET0131 , \g541_reg/NET0131 , \g545_reg/NET0131 , \g548_reg/NET0131 , \g551_reg/NET0131 , \g554_reg/NET0131 , \g557_pad , \g558_pad , \g559_pad , \g560_pad , \g561_pad , \g562_pad , \g563_pad , \g567_pad , \g571_reg/NET0131 , \g574_reg/NET0131 , \g578_reg/NET0131 , \g582_reg/NET0131 , \g586_reg/NET0131 , \g590_reg/NET0131 , \g594_reg/NET0131 , \g598_reg/NET0131 , \g602_reg/NET0131 , \g606_reg/NET0131 , \g610_reg/NET0131 , \g613_reg/NET0131 , \g616_reg/NET0131 , \g619_reg/NET0131 , \g622_reg/NET0131 , \g625_reg/NET0131 , \g628_reg/NET0131 , \g631_reg/NET0131 , \g634_reg/NET0131 , \g638_reg/NET0131 , \g639_pad , \g642_reg/NET0131 , \g646_reg/NET0131 , \g650_reg/NET0131 , \g654_reg/NET0131 , \g662_reg/NET0131 , \g669_reg/NET0131 , \g672_reg/NET0131 , \g675_reg/NET0131 , \g676_reg/NET0131 , \g677_reg/NET0131 , \g678_reg/NET0131 , \g679_reg/NET0131 , \g680_reg/NET0131 , \g681_reg/NET0131 , \g682_reg/NET0131 , \g683_reg/NET0131 , \g684_reg/NET0131 , \g685_reg/NET0131 , \g687_reg/NET0131 , \g688_reg/NET0131 , \g689_reg/NET0131 , \g698_reg/NET0131 , \g6_reg/NET0131 , \g702_pad , \g7_reg/NET0131 , \g89_pad , \_al_n1 , \g10560/_0_ , \g10562/_1_ , \g10564/_1_ , \g10566/_1_ , \g10567/_0_ , \g10569/_1_ , \g10580/_0_ , \g10616/_2_ , \g10627/_2_ , \g10628/_0_ , \g10629/_2_ , \g10630/_2_ , \g10633/_2_ , \g10635/_2_ , \g10636/_2_ , \g10637/_2_ , \g10641/_0_ , \g10649/_0_ , \g10672/_0_ , \g10673/_0_ , \g10680/_0_ , \g10683/_0_ , \g10686/_0_ , \g10695/_0_ , \g10700/_0_ , \g10703/_0_ , \g10704/_0_ , \g10748/_0_ , \g10750/_2_ , \g10757/_0_ , \g10758/_0_ , \g10782/_0_ , \g10826/_0_ , \g10827/_0_ , \g10828/_1_ , \g10832/_2_ , \g10834/_2_ , \g10836/_0_ , \g10837/_1__syn_2 , \g10868/_0_ , \g10904/_0_ , \g10913/_0_ , \g10915/_0_ , \g10922/_0_ , \g10938/_0_ , \g10939/_0_ , \g10940/_0_ , \g10941/_0_ , \g10942/_0_ , \g10944/_2_ , \g10977/_0_ , \g10980/_0_ , \g11020/_0_ , \g11028/_0_ , \g11051/_0_ , \g11057/_0_ , \g11109/_0_ , \g11113/_2_ , \g11156/_0_ , \g11172/_3_ , \g11193/_0_ , \g11219/_0_ , \g11355/_0_ , \g11384/_0_ , \g11442/_0_ , \g11448/_0_ , \g11558/_0_ , \g11559/_0_ , \g11824/_1_ , \g11853/_0_ , \g11854/_0_ , \g11977/_0_ , \g11981/_0_ , \g2584_pad , \g4121_pad , \g4809_pad , \g5692_pad , \g6282_pad , \g6284_pad , \g6360_pad , \g6362_pad , \g6364_pad , \g6366_pad , \g6368_pad , \g6370_pad , \g6372_pad , \g6374_pad );
	input \g102_pad  ;
	input \g10_reg/NET0131  ;
	input \g11_reg/NET0131  ;
	input \g1293_pad  ;
	input \g14_reg/NET0131  ;
	input \g15_reg/NET0131  ;
	input \g18_reg/NET0131  ;
	input \g197_reg/NET0131  ;
	input \g19_reg/NET0131  ;
	input \g1_reg/NET0131  ;
	input \g204_reg/NET0131  ;
	input \g205_reg/NET0131  ;
	input \g206_reg/NET0131  ;
	input \g207_reg/NET0131  ;
	input \g208_reg/NET0131  ;
	input \g209_reg/NET0131  ;
	input \g210_reg/NET0131  ;
	input \g211_reg/NET0131  ;
	input \g212_reg/NET0131  ;
	input \g218_reg/NET0131  ;
	input \g224_reg/NET0131  ;
	input \g230_reg/NET0131  ;
	input \g236_reg/NET0131  ;
	input \g242_reg/NET0131  ;
	input \g248_reg/NET0131  ;
	input \g24_reg/NET0131  ;
	input \g254_reg/NET0131  ;
	input \g25_reg/NET0131  ;
	input \g260_reg/NET0131  ;
	input \g266_reg/NET0131  ;
	input \g269_reg/NET0131  ;
	input \g276_reg/NET0131  ;
	input \g277_reg/NET0131  ;
	input \g278_reg/NET0131  ;
	input \g279_reg/NET0131  ;
	input \g280_reg/NET0131  ;
	input \g281_reg/NET0131  ;
	input \g282_reg/NET0131  ;
	input \g283_reg/NET0131  ;
	input \g28_reg/NET0131  ;
	input \g293_reg/NET0131  ;
	input \g297_reg/NET0131  ;
	input \g29_reg/NET0131  ;
	input \g2_reg/NET0131  ;
	input \g33_reg/NET0131  ;
	input \g3_reg/NET0131  ;
	input \g402_reg/NET0131  ;
	input \g406_reg/NET0131  ;
	input \g4099_pad  ;
	input \g4100_pad  ;
	input \g4101_pad  ;
	input \g4102_pad  ;
	input \g4103_pad  ;
	input \g4104_pad  ;
	input \g4105_pad  ;
	input \g4108_pad  ;
	input \g410_reg/NET0131  ;
	input \g4110_pad  ;
	input \g4112_pad  ;
	input \g414_reg/NET0131  ;
	input \g418_reg/NET0131  ;
	input \g422_reg/NET0131  ;
	input \g426_reg/NET0131  ;
	input \g430_reg/NET0131  ;
	input \g434_reg/NET0131  ;
	input \g437_reg/NET0131  ;
	input \g441_reg/NET0131  ;
	input \g4422_pad  ;
	input \g445_reg/NET0131  ;
	input \g449_reg/NET0131  ;
	input \g453_reg/NET0131  ;
	input \g457_reg/NET0131  ;
	input \g461_reg/NET0131  ;
	input \g465_reg/NET0131  ;
	input \g471_reg/NET0131  ;
	input \g478_reg/NET0131  ;
	input \g486_reg/NET0131  ;
	input \g489_reg/NET0131  ;
	input \g48_reg/NET0131  ;
	input \g492_reg/NET0131  ;
	input \g496_reg/NET0131  ;
	input \g500_reg/NET0131  ;
	input \g504_reg/NET0131  ;
	input \g508_reg/NET0131  ;
	input \g512_reg/NET0131  ;
	input \g536_reg/NET0131  ;
	input \g541_reg/NET0131  ;
	input \g545_reg/NET0131  ;
	input \g548_reg/NET0131  ;
	input \g551_reg/NET0131  ;
	input \g554_reg/NET0131  ;
	input \g557_pad  ;
	input \g558_pad  ;
	input \g559_pad  ;
	input \g560_pad  ;
	input \g561_pad  ;
	input \g562_pad  ;
	input \g563_pad  ;
	input \g567_pad  ;
	input \g571_reg/NET0131  ;
	input \g574_reg/NET0131  ;
	input \g578_reg/NET0131  ;
	input \g582_reg/NET0131  ;
	input \g586_reg/NET0131  ;
	input \g590_reg/NET0131  ;
	input \g594_reg/NET0131  ;
	input \g598_reg/NET0131  ;
	input \g602_reg/NET0131  ;
	input \g606_reg/NET0131  ;
	input \g610_reg/NET0131  ;
	input \g613_reg/NET0131  ;
	input \g616_reg/NET0131  ;
	input \g619_reg/NET0131  ;
	input \g622_reg/NET0131  ;
	input \g625_reg/NET0131  ;
	input \g628_reg/NET0131  ;
	input \g631_reg/NET0131  ;
	input \g634_reg/NET0131  ;
	input \g638_reg/NET0131  ;
	input \g639_pad  ;
	input \g642_reg/NET0131  ;
	input \g646_reg/NET0131  ;
	input \g650_reg/NET0131  ;
	input \g654_reg/NET0131  ;
	input \g662_reg/NET0131  ;
	input \g669_reg/NET0131  ;
	input \g672_reg/NET0131  ;
	input \g675_reg/NET0131  ;
	input \g676_reg/NET0131  ;
	input \g677_reg/NET0131  ;
	input \g678_reg/NET0131  ;
	input \g679_reg/NET0131  ;
	input \g680_reg/NET0131  ;
	input \g681_reg/NET0131  ;
	input \g682_reg/NET0131  ;
	input \g683_reg/NET0131  ;
	input \g684_reg/NET0131  ;
	input \g685_reg/NET0131  ;
	input \g687_reg/NET0131  ;
	input \g688_reg/NET0131  ;
	input \g689_reg/NET0131  ;
	input \g698_reg/NET0131  ;
	input \g6_reg/NET0131  ;
	input \g702_pad  ;
	input \g7_reg/NET0131  ;
	input \g89_pad  ;
	output \_al_n1  ;
	output \g10560/_0_  ;
	output \g10562/_1_  ;
	output \g10564/_1_  ;
	output \g10566/_1_  ;
	output \g10567/_0_  ;
	output \g10569/_1_  ;
	output \g10580/_0_  ;
	output \g10616/_2_  ;
	output \g10627/_2_  ;
	output \g10628/_0_  ;
	output \g10629/_2_  ;
	output \g10630/_2_  ;
	output \g10633/_2_  ;
	output \g10635/_2_  ;
	output \g10636/_2_  ;
	output \g10637/_2_  ;
	output \g10641/_0_  ;
	output \g10649/_0_  ;
	output \g10672/_0_  ;
	output \g10673/_0_  ;
	output \g10680/_0_  ;
	output \g10683/_0_  ;
	output \g10686/_0_  ;
	output \g10695/_0_  ;
	output \g10700/_0_  ;
	output \g10703/_0_  ;
	output \g10704/_0_  ;
	output \g10748/_0_  ;
	output \g10750/_2_  ;
	output \g10757/_0_  ;
	output \g10758/_0_  ;
	output \g10782/_0_  ;
	output \g10826/_0_  ;
	output \g10827/_0_  ;
	output \g10828/_1_  ;
	output \g10832/_2_  ;
	output \g10834/_2_  ;
	output \g10836/_0_  ;
	output \g10837/_1__syn_2  ;
	output \g10868/_0_  ;
	output \g10904/_0_  ;
	output \g10913/_0_  ;
	output \g10915/_0_  ;
	output \g10922/_0_  ;
	output \g10938/_0_  ;
	output \g10939/_0_  ;
	output \g10940/_0_  ;
	output \g10941/_0_  ;
	output \g10942/_0_  ;
	output \g10944/_2_  ;
	output \g10977/_0_  ;
	output \g10980/_0_  ;
	output \g11020/_0_  ;
	output \g11028/_0_  ;
	output \g11051/_0_  ;
	output \g11057/_0_  ;
	output \g11109/_0_  ;
	output \g11113/_2_  ;
	output \g11156/_0_  ;
	output \g11172/_3_  ;
	output \g11193/_0_  ;
	output \g11219/_0_  ;
	output \g11355/_0_  ;
	output \g11384/_0_  ;
	output \g11442/_0_  ;
	output \g11448/_0_  ;
	output \g11558/_0_  ;
	output \g11559/_0_  ;
	output \g11824/_1_  ;
	output \g11853/_0_  ;
	output \g11854/_0_  ;
	output \g11977/_0_  ;
	output \g11981/_0_  ;
	output \g2584_pad  ;
	output \g4121_pad  ;
	output \g4809_pad  ;
	output \g5692_pad  ;
	output \g6282_pad  ;
	output \g6284_pad  ;
	output \g6360_pad  ;
	output \g6362_pad  ;
	output \g6364_pad  ;
	output \g6366_pad  ;
	output \g6368_pad  ;
	output \g6370_pad  ;
	output \g6372_pad  ;
	output \g6374_pad  ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w262_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w164_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w165_ ;
	wire _w263_ ;
	wire _w136_ ;
	wire _w393_ ;
	wire _w195_ ;
	wire _w180_ ;
	wire _w153_ ;
	wire _w163_ ;
	wire _w261_ ;
	wire _w134_ ;
	wire _w391_ ;
	wire _w193_ ;
	wire _w160_ ;
	wire _w152_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w32_ ;
	wire _w289_ ;
	wire _w159_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w62_ ;
	wire _w319_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w194_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w392_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\g266_reg/NET0131 ,
		_w32_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\g4112_pad ,
		_w62_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\g677_reg/NET0131 ,
		_w134_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\g678_reg/NET0131 ,
		_w136_
	);
	LUT3 #(
		.INIT('h80)
	) name4 (
		\g602_reg/NET0131 ,
		\g610_reg/NET0131 ,
		\g613_reg/NET0131 ,
		_w152_
	);
	LUT4 #(
		.INIT('h8000)
	) name5 (
		\g602_reg/NET0131 ,
		\g610_reg/NET0131 ,
		\g613_reg/NET0131 ,
		\g616_reg/NET0131 ,
		_w153_
	);
	LUT3 #(
		.INIT('h80)
	) name6 (
		\g619_reg/NET0131 ,
		\g622_reg/NET0131 ,
		_w153_,
		_w154_
	);
	LUT4 #(
		.INIT('h8000)
	) name7 (
		\g619_reg/NET0131 ,
		\g622_reg/NET0131 ,
		\g625_reg/NET0131 ,
		_w153_,
		_w155_
	);
	LUT4 #(
		.INIT('h8000)
	) name8 (
		\g578_reg/NET0131 ,
		\g628_reg/NET0131 ,
		\g631_reg/NET0131 ,
		_w155_,
		_w156_
	);
	LUT4 #(
		.INIT('h8000)
	) name9 (
		\g574_reg/NET0131 ,
		\g582_reg/NET0131 ,
		\g586_reg/NET0131 ,
		_w156_,
		_w157_
	);
	LUT4 #(
		.INIT('h70f0)
	) name10 (
		\g590_reg/NET0131 ,
		\g594_reg/NET0131 ,
		\g639_pad ,
		_w157_,
		_w158_
	);
	LUT4 #(
		.INIT('hdfaf)
	) name11 (
		\g590_reg/NET0131 ,
		\g594_reg/NET0131 ,
		\g639_pad ,
		_w157_,
		_w159_
	);
	LUT2 #(
		.INIT('h6)
	) name12 (
		\g582_reg/NET0131 ,
		_w156_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w158_,
		_w160_,
		_w161_
	);
	LUT3 #(
		.INIT('h6c)
	) name14 (
		\g582_reg/NET0131 ,
		\g586_reg/NET0131 ,
		_w156_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w158_,
		_w162_,
		_w163_
	);
	LUT4 #(
		.INIT('h60c0)
	) name16 (
		\g590_reg/NET0131 ,
		\g594_reg/NET0131 ,
		\g639_pad ,
		_w157_,
		_w164_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name17 (
		\g574_reg/NET0131 ,
		\g582_reg/NET0131 ,
		\g586_reg/NET0131 ,
		_w156_,
		_w165_
	);
	LUT2 #(
		.INIT('hd)
	) name18 (
		_w158_,
		_w165_,
		_w166_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name19 (
		\g578_reg/NET0131 ,
		\g628_reg/NET0131 ,
		\g631_reg/NET0131 ,
		_w155_,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w158_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h9)
	) name21 (
		\g19_reg/NET0131 ,
		\g25_reg/NET0131 ,
		_w169_
	);
	LUT3 #(
		.INIT('h96)
	) name22 (
		\g33_reg/NET0131 ,
		\g3_reg/NET0131 ,
		\g7_reg/NET0131 ,
		_w170_
	);
	LUT3 #(
		.INIT('h69)
	) name23 (
		\g11_reg/NET0131 ,
		\g15_reg/NET0131 ,
		\g29_reg/NET0131 ,
		_w171_
	);
	LUT3 #(
		.INIT('h69)
	) name24 (
		_w169_,
		_w170_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\g1293_pad ,
		\g702_pad ,
		_w173_
	);
	LUT3 #(
		.INIT('h40)
	) name26 (
		\g266_reg/NET0131 ,
		\g4110_pad ,
		\g662_reg/NET0131 ,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w173_,
		_w174_,
		_w175_
	);
	LUT4 #(
		.INIT('h2000)
	) name28 (
		\g676_reg/NET0131 ,
		\g698_reg/NET0131 ,
		_w173_,
		_w174_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\g688_reg/NET0131 ,
		\g689_reg/NET0131 ,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w176_,
		_w177_,
		_w178_
	);
	LUT3 #(
		.INIT('h40)
	) name31 (
		\g687_reg/NET0131 ,
		_w176_,
		_w177_,
		_w179_
	);
	LUT4 #(
		.INIT('h8000)
	) name32 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		\g206_reg/NET0131 ,
		\g207_reg/NET0131 ,
		_w180_
	);
	LUT3 #(
		.INIT('h80)
	) name33 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w182_
	);
	LUT2 #(
		.INIT('h9)
	) name35 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w183_
	);
	LUT4 #(
		.INIT('h4206)
	) name36 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g471_reg/NET0131 ,
		_w180_,
		_w184_
	);
	LUT4 #(
		.INIT('h0213)
	) name37 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		\g679_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w185_
	);
	LUT4 #(
		.INIT('h084c)
	) name38 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		\g677_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w186_
	);
	LUT3 #(
		.INIT('ha8)
	) name39 (
		\g206_reg/NET0131 ,
		_w185_,
		_w186_,
		_w187_
	);
	LUT4 #(
		.INIT('h0213)
	) name40 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		\g683_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w188_
	);
	LUT4 #(
		.INIT('h084c)
	) name41 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		\g681_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w189_
	);
	LUT3 #(
		.INIT('h54)
	) name42 (
		\g206_reg/NET0131 ,
		_w188_,
		_w189_,
		_w190_
	);
	LUT4 #(
		.INIT('h8884)
	) name43 (
		\g471_reg/NET0131 ,
		_w183_,
		_w187_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\g210_reg/NET0131 ,
		\g211_reg/NET0131 ,
		_w192_
	);
	LUT4 #(
		.INIT('ha800)
	) name45 (
		_w181_,
		_w184_,
		_w191_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		\g210_reg/NET0131 ,
		\g211_reg/NET0131 ,
		_w194_
	);
	LUT4 #(
		.INIT('h8000)
	) name47 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w180_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\g210_reg/NET0131 ,
		\g211_reg/NET0131 ,
		_w196_
	);
	LUT4 #(
		.INIT('h8000)
	) name49 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w180_,
		_w196_,
		_w197_
	);
	LUT3 #(
		.INIT('h01)
	) name50 (
		\g210_reg/NET0131 ,
		\g211_reg/NET0131 ,
		\g471_reg/NET0131 ,
		_w198_
	);
	LUT4 #(
		.INIT('hd900)
	) name51 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w180_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w197_,
		_w199_,
		_w200_
	);
	LUT3 #(
		.INIT('h70)
	) name53 (
		_w191_,
		_w195_,
		_w200_,
		_w201_
	);
	LUT3 #(
		.INIT('h20)
	) name54 (
		\g211_reg/NET0131 ,
		_w193_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w191_,
		_w195_,
		_w203_
	);
	LUT4 #(
		.INIT('h7f00)
	) name56 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w180_,
		_w192_,
		_w204_
	);
	LUT3 #(
		.INIT('h70)
	) name57 (
		\g208_reg/NET0131 ,
		_w180_,
		_w194_,
		_w205_
	);
	LUT4 #(
		.INIT('h131f)
	) name58 (
		_w184_,
		_w191_,
		_w204_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		_w203_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('hb)
	) name60 (
		_w202_,
		_w207_,
		_w208_
	);
	LUT4 #(
		.INIT('h1b11)
	) name61 (
		\g197_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w202_,
		_w207_,
		_w209_
	);
	LUT4 #(
		.INIT('he4ee)
	) name62 (
		\g197_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w202_,
		_w207_,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		_w179_,
		_w209_,
		_w211_
	);
	LUT3 #(
		.INIT('h80)
	) name64 (
		\g687_reg/NET0131 ,
		_w176_,
		_w177_,
		_w212_
	);
	LUT4 #(
		.INIT('h8000)
	) name65 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		\g278_reg/NET0131 ,
		\g279_reg/NET0131 ,
		_w213_
	);
	LUT3 #(
		.INIT('h80)
	) name66 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w215_
	);
	LUT2 #(
		.INIT('h9)
	) name68 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w216_
	);
	LUT4 #(
		.INIT('h0213)
	) name69 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		\g679_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w217_
	);
	LUT4 #(
		.INIT('h084c)
	) name70 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		\g677_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w218_
	);
	LUT3 #(
		.INIT('ha8)
	) name71 (
		\g278_reg/NET0131 ,
		_w217_,
		_w218_,
		_w219_
	);
	LUT4 #(
		.INIT('h0213)
	) name72 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		\g683_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w220_
	);
	LUT4 #(
		.INIT('h084c)
	) name73 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		\g681_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w221_
	);
	LUT3 #(
		.INIT('h54)
	) name74 (
		\g278_reg/NET0131 ,
		_w220_,
		_w221_,
		_w222_
	);
	LUT3 #(
		.INIT('h56)
	) name75 (
		\g478_reg/NET0131 ,
		_w219_,
		_w222_,
		_w223_
	);
	LUT4 #(
		.INIT('h4448)
	) name76 (
		\g478_reg/NET0131 ,
		_w216_,
		_w219_,
		_w222_,
		_w224_
	);
	LUT4 #(
		.INIT('h2d69)
	) name77 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		\g478_reg/NET0131 ,
		_w213_,
		_w225_
	);
	LUT4 #(
		.INIT('h2460)
	) name78 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		\g478_reg/NET0131 ,
		_w213_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\g282_reg/NET0131 ,
		\g283_reg/NET0131 ,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w226_,
		_w227_,
		_w228_
	);
	LUT4 #(
		.INIT('h4c44)
	) name81 (
		\g282_reg/NET0131 ,
		_w214_,
		_w224_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\g283_reg/NET0131 ,
		_w229_,
		_w230_
	);
	LUT4 #(
		.INIT('h8884)
	) name83 (
		\g478_reg/NET0131 ,
		_w216_,
		_w219_,
		_w222_,
		_w231_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\g282_reg/NET0131 ,
		\g283_reg/NET0131 ,
		_w232_
	);
	LUT4 #(
		.INIT('h8d8f)
	) name85 (
		_w216_,
		_w223_,
		_w228_,
		_w232_,
		_w233_
	);
	LUT4 #(
		.INIT('h8000)
	) name86 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w213_,
		_w232_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		_w231_,
		_w234_,
		_w235_
	);
	LUT3 #(
		.INIT('h0e)
	) name88 (
		_w214_,
		_w233_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('hb)
	) name89 (
		_w230_,
		_w236_,
		_w237_
	);
	LUT4 #(
		.INIT('h1b11)
	) name90 (
		\g269_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w230_,
		_w236_,
		_w238_
	);
	LUT4 #(
		.INIT('he4ee)
	) name91 (
		\g269_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w230_,
		_w236_,
		_w239_
	);
	LUT4 #(
		.INIT('h2000)
	) name92 (
		\g685_reg/NET0131 ,
		\g688_reg/NET0131 ,
		\g689_reg/NET0131 ,
		\g698_reg/NET0131 ,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		\g683_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w241_
	);
	LUT3 #(
		.INIT('h40)
	) name94 (
		\g681_reg/NET0131 ,
		\g683_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w242_
	);
	LUT3 #(
		.INIT('h40)
	) name95 (
		\g682_reg/NET0131 ,
		_w240_,
		_w242_,
		_w243_
	);
	LUT4 #(
		.INIT('h8000)
	) name96 (
		\g500_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w175_,
		_w243_,
		_w244_
	);
	LUT3 #(
		.INIT('h80)
	) name97 (
		\g688_reg/NET0131 ,
		\g689_reg/NET0131 ,
		\g698_reg/NET0131 ,
		_w245_
	);
	LUT4 #(
		.INIT('h4000)
	) name98 (
		\g680_reg/NET0131 ,
		_w173_,
		_w174_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		\g679_reg/NET0131 ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w248_
	);
	LUT3 #(
		.INIT('h10)
	) name101 (
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w249_
	);
	LUT4 #(
		.INIT('h8000)
	) name102 (
		_w173_,
		_w174_,
		_w245_,
		_w249_,
		_w250_
	);
	LUT4 #(
		.INIT('h8000)
	) name103 (
		\g684_reg/NET0131 ,
		_w173_,
		_w174_,
		_w240_,
		_w251_
	);
	LUT4 #(
		.INIT('h0007)
	) name104 (
		_w176_,
		_w177_,
		_w250_,
		_w251_,
		_w252_
	);
	LUT4 #(
		.INIT('h1000)
	) name105 (
		\g685_reg/NET0131 ,
		\g688_reg/NET0131 ,
		\g689_reg/NET0131 ,
		\g698_reg/NET0131 ,
		_w253_
	);
	LUT4 #(
		.INIT('h8000)
	) name106 (
		\g676_reg/NET0131 ,
		_w173_,
		_w174_,
		_w253_,
		_w254_
	);
	LUT3 #(
		.INIT('h07)
	) name107 (
		\g689_reg/NET0131 ,
		_w176_,
		_w254_,
		_w255_
	);
	LUT3 #(
		.INIT('h80)
	) name108 (
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w246_,
		_w256_
	);
	LUT4 #(
		.INIT('h0200)
	) name109 (
		_w255_,
		_w247_,
		_w256_,
		_w252_,
		_w257_
	);
	LUT4 #(
		.INIT('h8000)
	) name110 (
		\g557_pad ,
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w246_,
		_w258_
	);
	LUT4 #(
		.INIT('haa80)
	) name111 (
		\g684_reg/NET0131 ,
		\g689_reg/NET0131 ,
		_w176_,
		_w254_,
		_w259_
	);
	LUT3 #(
		.INIT('h80)
	) name112 (
		_w173_,
		_w174_,
		_w241_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\g682_reg/NET0131 ,
		_w240_,
		_w261_
	);
	LUT4 #(
		.INIT('h2000)
	) name114 (
		\g434_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w262_
	);
	LUT4 #(
		.INIT('h8000)
	) name115 (
		\g430_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w263_
	);
	LUT4 #(
		.INIT('h0001)
	) name116 (
		_w259_,
		_w262_,
		_w263_,
		_w258_,
		_w264_
	);
	LUT3 #(
		.INIT('h10)
	) name117 (
		_w244_,
		_w257_,
		_w264_,
		_w265_
	);
	LUT3 #(
		.INIT('hd0)
	) name118 (
		_w212_,
		_w238_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('hb)
	) name119 (
		_w211_,
		_w266_,
		_w267_
	);
	LUT3 #(
		.INIT('h8a)
	) name120 (
		\g210_reg/NET0131 ,
		\g211_reg/NET0131 ,
		_w184_,
		_w268_
	);
	LUT4 #(
		.INIT('h0444)
	) name121 (
		_w193_,
		_w201_,
		_w206_,
		_w268_,
		_w269_
	);
	LUT4 #(
		.INIT('hfbbb)
	) name122 (
		_w193_,
		_w201_,
		_w206_,
		_w268_,
		_w270_
	);
	LUT4 #(
		.INIT('h1b11)
	) name123 (
		\g197_reg/NET0131 ,
		\g683_reg/NET0131 ,
		_w203_,
		_w269_,
		_w271_
	);
	LUT4 #(
		.INIT('he4ee)
	) name124 (
		\g197_reg/NET0131 ,
		\g683_reg/NET0131 ,
		_w203_,
		_w269_,
		_w272_
	);
	LUT3 #(
		.INIT('h06)
	) name125 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		\g283_reg/NET0131 ,
		_w273_
	);
	LUT3 #(
		.INIT('h8a)
	) name126 (
		\g282_reg/NET0131 ,
		_w225_,
		_w273_,
		_w274_
	);
	LUT3 #(
		.INIT('h01)
	) name127 (
		\g282_reg/NET0131 ,
		\g283_reg/NET0131 ,
		\g478_reg/NET0131 ,
		_w275_
	);
	LUT4 #(
		.INIT('hd900)
	) name128 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w213_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		\g282_reg/NET0131 ,
		\g283_reg/NET0131 ,
		_w277_
	);
	LUT4 #(
		.INIT('h8000)
	) name130 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w213_,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w276_,
		_w278_,
		_w279_
	);
	LUT4 #(
		.INIT('h1d00)
	) name132 (
		_w214_,
		_w233_,
		_w274_,
		_w279_,
		_w280_
	);
	LUT4 #(
		.INIT('he2ff)
	) name133 (
		_w214_,
		_w233_,
		_w274_,
		_w279_,
		_w281_
	);
	LUT3 #(
		.INIT('h4e)
	) name134 (
		\g269_reg/NET0131 ,
		\g683_reg/NET0131 ,
		_w280_,
		_w282_
	);
	LUT4 #(
		.INIT('h40e0)
	) name135 (
		\g269_reg/NET0131 ,
		\g683_reg/NET0131 ,
		_w212_,
		_w280_,
		_w283_
	);
	LUT4 #(
		.INIT('h8000)
	) name136 (
		\g558_pad ,
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w246_,
		_w284_
	);
	LUT4 #(
		.INIT('haa80)
	) name137 (
		\g683_reg/NET0131 ,
		\g689_reg/NET0131 ,
		_w176_,
		_w254_,
		_w285_
	);
	LUT4 #(
		.INIT('h8000)
	) name138 (
		\g426_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w286_
	);
	LUT4 #(
		.INIT('h2000)
	) name139 (
		\g437_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w287_
	);
	LUT4 #(
		.INIT('h0001)
	) name140 (
		_w285_,
		_w286_,
		_w287_,
		_w284_,
		_w288_
	);
	LUT3 #(
		.INIT('h10)
	) name141 (
		_w244_,
		_w257_,
		_w288_,
		_w289_
	);
	LUT4 #(
		.INIT('hf2ff)
	) name142 (
		_w179_,
		_w271_,
		_w283_,
		_w289_,
		_w290_
	);
	LUT3 #(
		.INIT('h80)
	) name143 (
		\g567_pad ,
		\g598_reg/NET0131 ,
		\g634_reg/NET0131 ,
		_w291_
	);
	LUT4 #(
		.INIT('h8000)
	) name144 (
		\g567_pad ,
		\g598_reg/NET0131 ,
		\g634_reg/NET0131 ,
		\g642_reg/NET0131 ,
		_w292_
	);
	LUT3 #(
		.INIT('h80)
	) name145 (
		\g606_reg/NET0131 ,
		\g646_reg/NET0131 ,
		_w292_,
		_w293_
	);
	LUT4 #(
		.INIT('h8000)
	) name146 (
		\g606_reg/NET0131 ,
		\g646_reg/NET0131 ,
		\g650_reg/NET0131 ,
		_w292_,
		_w294_
	);
	LUT4 #(
		.INIT('h4888)
	) name147 (
		\g571_reg/NET0131 ,
		\g638_reg/NET0131 ,
		\g654_reg/NET0131 ,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		\g197_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w296_
	);
	LUT4 #(
		.INIT('ha680)
	) name149 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w180_,
		_w198_,
		_w297_
	);
	LUT3 #(
		.INIT('h78)
	) name150 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		\g206_reg/NET0131 ,
		_w298_
	);
	LUT4 #(
		.INIT('h0200)
	) name151 (
		\g197_reg/NET0131 ,
		_w199_,
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('he)
	) name152 (
		_w296_,
		_w299_,
		_w300_
	);
	LUT3 #(
		.INIT('ha8)
	) name153 (
		_w179_,
		_w296_,
		_w299_,
		_w301_
	);
	LUT4 #(
		.INIT('h007f)
	) name154 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w213_,
		_w275_,
		_w302_
	);
	LUT3 #(
		.INIT('h78)
	) name155 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		\g278_reg/NET0131 ,
		_w303_
	);
	LUT4 #(
		.INIT('h1bbb)
	) name156 (
		\g269_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w302_,
		_w303_,
		_w304_
	);
	LUT4 #(
		.INIT('he444)
	) name157 (
		\g269_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w302_,
		_w303_,
		_w305_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		_w212_,
		_w304_,
		_w306_
	);
	LUT4 #(
		.INIT('h8000)
	) name159 (
		\g410_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w307_
	);
	LUT3 #(
		.INIT('h20)
	) name160 (
		\g681_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w240_,
		_w308_
	);
	LUT3 #(
		.INIT('h80)
	) name161 (
		\g551_reg/NET0131 ,
		_w260_,
		_w308_,
		_w309_
	);
	LUT3 #(
		.INIT('h40)
	) name162 (
		\g683_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w240_,
		_w310_
	);
	LUT3 #(
		.INIT('h80)
	) name163 (
		\g293_reg/NET0131 ,
		_w175_,
		_w310_,
		_w311_
	);
	LUT4 #(
		.INIT('h2000)
	) name164 (
		\g453_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w312_
	);
	LUT4 #(
		.INIT('h0001)
	) name165 (
		_w307_,
		_w309_,
		_w311_,
		_w312_,
		_w313_
	);
	LUT4 #(
		.INIT('h2000)
	) name166 (
		\g536_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w175_,
		_w243_,
		_w314_
	);
	LUT4 #(
		.INIT('h8000)
	) name167 (
		\g508_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w175_,
		_w243_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT3 #(
		.INIT('h80)
	) name169 (
		\g562_pad ,
		\g678_reg/NET0131 ,
		_w246_,
		_w317_
	);
	LUT3 #(
		.INIT('ha2)
	) name170 (
		\g679_reg/NET0131 ,
		_w255_,
		_w317_,
		_w318_
	);
	LUT4 #(
		.INIT('h1000)
	) name171 (
		_w257_,
		_w318_,
		_w313_,
		_w316_,
		_w319_
	);
	LUT3 #(
		.INIT('hef)
	) name172 (
		_w306_,
		_w301_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		\g269_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w321_
	);
	LUT4 #(
		.INIT('h7f80)
	) name174 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		\g278_reg/NET0131 ,
		\g279_reg/NET0131 ,
		_w322_
	);
	LUT4 #(
		.INIT('h597f)
	) name175 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w213_,
		_w275_,
		_w323_
	);
	LUT4 #(
		.INIT('h2022)
	) name176 (
		\g269_reg/NET0131 ,
		_w276_,
		_w322_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('he)
	) name177 (
		_w321_,
		_w324_,
		_w325_
	);
	LUT3 #(
		.INIT('ha8)
	) name178 (
		_w212_,
		_w321_,
		_w324_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		\g197_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w327_
	);
	LUT4 #(
		.INIT('h7f80)
	) name180 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		\g206_reg/NET0131 ,
		\g207_reg/NET0131 ,
		_w328_
	);
	LUT4 #(
		.INIT('h2220)
	) name181 (
		\g197_reg/NET0131 ,
		_w199_,
		_w297_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('he)
	) name182 (
		_w327_,
		_w329_,
		_w330_
	);
	LUT3 #(
		.INIT('ha8)
	) name183 (
		_w179_,
		_w327_,
		_w329_,
		_w331_
	);
	LUT4 #(
		.INIT('h8000)
	) name184 (
		\g512_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w175_,
		_w243_,
		_w332_
	);
	LUT4 #(
		.INIT('haa80)
	) name185 (
		\g680_reg/NET0131 ,
		\g689_reg/NET0131 ,
		_w176_,
		_w254_,
		_w333_
	);
	LUT4 #(
		.INIT('h2000)
	) name186 (
		\g541_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w175_,
		_w243_,
		_w334_
	);
	LUT4 #(
		.INIT('h8000)
	) name187 (
		\g561_pad ,
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w246_,
		_w335_
	);
	LUT4 #(
		.INIT('h0001)
	) name188 (
		_w332_,
		_w333_,
		_w334_,
		_w335_,
		_w336_
	);
	LUT4 #(
		.INIT('h8000)
	) name189 (
		\g414_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w337_
	);
	LUT4 #(
		.INIT('h2000)
	) name190 (
		\g449_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w338_
	);
	LUT3 #(
		.INIT('h80)
	) name191 (
		\g554_reg/NET0131 ,
		_w260_,
		_w308_,
		_w339_
	);
	LUT3 #(
		.INIT('h80)
	) name192 (
		\g297_reg/NET0131 ,
		_w175_,
		_w310_,
		_w340_
	);
	LUT4 #(
		.INIT('h0001)
	) name193 (
		_w337_,
		_w338_,
		_w339_,
		_w340_,
		_w341_
	);
	LUT4 #(
		.INIT('h1000)
	) name194 (
		_w257_,
		_w331_,
		_w341_,
		_w336_,
		_w342_
	);
	LUT2 #(
		.INIT('hb)
	) name195 (
		_w326_,
		_w342_,
		_w343_
	);
	LUT4 #(
		.INIT('h596c)
	) name196 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w213_,
		_w275_,
		_w344_
	);
	LUT3 #(
		.INIT('he4)
	) name197 (
		\g269_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w212_,
		_w345_,
		_w346_
	);
	LUT4 #(
		.INIT('h0293)
	) name199 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w180_,
		_w198_,
		_w347_
	);
	LUT4 #(
		.INIT('hbbb1)
	) name200 (
		\g197_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w297_,
		_w347_,
		_w348_
	);
	LUT4 #(
		.INIT('h444e)
	) name201 (
		\g197_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w297_,
		_w347_,
		_w349_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		_w179_,
		_w348_,
		_w350_
	);
	LUT4 #(
		.INIT('h8000)
	) name203 (
		\g559_pad ,
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w246_,
		_w351_
	);
	LUT4 #(
		.INIT('haa80)
	) name204 (
		\g682_reg/NET0131 ,
		\g689_reg/NET0131 ,
		_w176_,
		_w254_,
		_w352_
	);
	LUT4 #(
		.INIT('h8000)
	) name205 (
		\g422_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w353_
	);
	LUT4 #(
		.INIT('h2000)
	) name206 (
		\g441_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w354_
	);
	LUT4 #(
		.INIT('h0001)
	) name207 (
		_w352_,
		_w353_,
		_w354_,
		_w351_,
		_w355_
	);
	LUT4 #(
		.INIT('hfeff)
	) name208 (
		_w257_,
		_w350_,
		_w346_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		\g197_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w357_
	);
	LUT2 #(
		.INIT('h6)
	) name210 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		_w358_
	);
	LUT4 #(
		.INIT('h0200)
	) name211 (
		\g197_reg/NET0131 ,
		_w199_,
		_w297_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('he)
	) name212 (
		_w357_,
		_w359_,
		_w360_
	);
	LUT3 #(
		.INIT('ha8)
	) name213 (
		_w179_,
		_w357_,
		_w359_,
		_w361_
	);
	LUT3 #(
		.INIT('h10)
	) name214 (
		\g489_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w246_,
		_w362_
	);
	LUT3 #(
		.INIT('ha2)
	) name215 (
		\g678_reg/NET0131 ,
		_w255_,
		_w362_,
		_w363_
	);
	LUT4 #(
		.INIT('h2000)
	) name216 (
		\g457_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w364_
	);
	LUT4 #(
		.INIT('h8000)
	) name217 (
		\g406_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w365_
	);
	LUT3 #(
		.INIT('h80)
	) name218 (
		\g269_reg/NET0131 ,
		_w175_,
		_w310_,
		_w366_
	);
	LUT3 #(
		.INIT('h80)
	) name219 (
		\g492_reg/NET0131 ,
		_w248_,
		_w246_,
		_w367_
	);
	LUT4 #(
		.INIT('h0001)
	) name220 (
		_w364_,
		_w365_,
		_w366_,
		_w367_,
		_w368_
	);
	LUT3 #(
		.INIT('h10)
	) name221 (
		_w257_,
		_w363_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h6)
	) name222 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		_w370_
	);
	LUT4 #(
		.INIT('h1bbb)
	) name223 (
		\g269_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w302_,
		_w370_,
		_w371_
	);
	LUT4 #(
		.INIT('he444)
	) name224 (
		\g269_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w302_,
		_w370_,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name225 (
		_w212_,
		_w371_,
		_w373_
	);
	LUT4 #(
		.INIT('h2000)
	) name226 (
		\g465_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w175_,
		_w243_,
		_w374_
	);
	LUT3 #(
		.INIT('h80)
	) name227 (
		\g548_reg/NET0131 ,
		_w260_,
		_w308_,
		_w375_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		\g672_reg/NET0131 ,
		_w250_,
		_w376_
	);
	LUT3 #(
		.INIT('h01)
	) name229 (
		_w375_,
		_w374_,
		_w376_,
		_w377_
	);
	LUT4 #(
		.INIT('h8000)
	) name230 (
		\g563_pad ,
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w246_,
		_w378_
	);
	LUT4 #(
		.INIT('h8000)
	) name231 (
		\g504_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w175_,
		_w243_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT3 #(
		.INIT('h40)
	) name233 (
		_w373_,
		_w377_,
		_w380_,
		_w381_
	);
	LUT3 #(
		.INIT('hbf)
	) name234 (
		_w361_,
		_w369_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		\g197_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w383_
	);
	LUT4 #(
		.INIT('h0002)
	) name236 (
		\g197_reg/NET0131 ,
		\g204_reg/NET0131 ,
		_w199_,
		_w297_,
		_w384_
	);
	LUT2 #(
		.INIT('he)
	) name237 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT3 #(
		.INIT('ha8)
	) name238 (
		_w179_,
		_w383_,
		_w384_,
		_w386_
	);
	LUT4 #(
		.INIT('h2000)
	) name239 (
		\g461_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w387_
	);
	LUT3 #(
		.INIT('h80)
	) name240 (
		\g197_reg/NET0131 ,
		_w175_,
		_w310_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\g486_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w389_
	);
	LUT3 #(
		.INIT('h80)
	) name242 (
		\g678_reg/NET0131 ,
		_w246_,
		_w389_,
		_w390_
	);
	LUT3 #(
		.INIT('h01)
	) name243 (
		_w388_,
		_w390_,
		_w387_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		\g669_reg/NET0131 ,
		_w250_,
		_w392_
	);
	LUT3 #(
		.INIT('h80)
	) name245 (
		\g545_reg/NET0131 ,
		_w260_,
		_w308_,
		_w393_
	);
	LUT4 #(
		.INIT('h8000)
	) name246 (
		\g402_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w394_
	);
	LUT3 #(
		.INIT('h80)
	) name247 (
		\g496_reg/NET0131 ,
		_w248_,
		_w246_,
		_w395_
	);
	LUT4 #(
		.INIT('h0001)
	) name248 (
		_w392_,
		_w393_,
		_w394_,
		_w395_,
		_w396_
	);
	LUT3 #(
		.INIT('h40)
	) name249 (
		_w257_,
		_w391_,
		_w396_,
		_w397_
	);
	LUT4 #(
		.INIT('h8daf)
	) name250 (
		\g269_reg/NET0131 ,
		\g276_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w302_,
		_w398_
	);
	LUT4 #(
		.INIT('h7250)
	) name251 (
		\g269_reg/NET0131 ,
		\g276_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w302_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		_w212_,
		_w398_,
		_w400_
	);
	LUT4 #(
		.INIT('h8000)
	) name253 (
		\g4422_pad ,
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w246_,
		_w401_
	);
	LUT4 #(
		.INIT('haa80)
	) name254 (
		\g677_reg/NET0131 ,
		\g689_reg/NET0131 ,
		_w176_,
		_w254_,
		_w402_
	);
	LUT3 #(
		.INIT('h01)
	) name255 (
		_w244_,
		_w402_,
		_w401_,
		_w403_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		_w400_,
		_w403_,
		_w404_
	);
	LUT3 #(
		.INIT('hbf)
	) name257 (
		_w386_,
		_w397_,
		_w404_,
		_w405_
	);
	LUT4 #(
		.INIT('haa80)
	) name258 (
		\g681_reg/NET0131 ,
		\g689_reg/NET0131 ,
		_w176_,
		_w254_,
		_w406_
	);
	LUT4 #(
		.INIT('h8000)
	) name259 (
		\g560_pad ,
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w246_,
		_w407_
	);
	LUT4 #(
		.INIT('h2000)
	) name260 (
		\g445_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w408_
	);
	LUT4 #(
		.INIT('h8000)
	) name261 (
		\g418_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w260_,
		_w261_,
		_w409_
	);
	LUT4 #(
		.INIT('h0001)
	) name262 (
		_w407_,
		_w408_,
		_w406_,
		_w409_,
		_w410_
	);
	LUT4 #(
		.INIT('h0025)
	) name263 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w213_,
		_w275_,
		_w411_
	);
	LUT3 #(
		.INIT('hb1)
	) name264 (
		\g269_reg/NET0131 ,
		\g681_reg/NET0131 ,
		_w411_,
		_w412_
	);
	LUT3 #(
		.INIT('h4e)
	) name265 (
		\g269_reg/NET0131 ,
		\g681_reg/NET0131 ,
		_w411_,
		_w413_
	);
	LUT4 #(
		.INIT('h0025)
	) name266 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w180_,
		_w198_,
		_w414_
	);
	LUT3 #(
		.INIT('hb1)
	) name267 (
		\g197_reg/NET0131 ,
		\g681_reg/NET0131 ,
		_w414_,
		_w415_
	);
	LUT3 #(
		.INIT('h4e)
	) name268 (
		\g197_reg/NET0131 ,
		\g681_reg/NET0131 ,
		_w414_,
		_w416_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name269 (
		\g687_reg/NET0131 ,
		_w178_,
		_w412_,
		_w415_,
		_w417_
	);
	LUT3 #(
		.INIT('hbf)
	) name270 (
		_w257_,
		_w410_,
		_w417_,
		_w418_
	);
	LUT4 #(
		.INIT('h60c0)
	) name271 (
		\g628_reg/NET0131 ,
		\g631_reg/NET0131 ,
		\g639_pad ,
		_w155_,
		_w419_
	);
	LUT3 #(
		.INIT('h28)
	) name272 (
		\g638_reg/NET0131 ,
		\g654_reg/NET0131 ,
		_w294_,
		_w420_
	);
	LUT3 #(
		.INIT('h48)
	) name273 (
		\g628_reg/NET0131 ,
		\g639_pad ,
		_w155_,
		_w421_
	);
	LUT3 #(
		.INIT('hf4)
	) name274 (
		_w202_,
		_w207_,
		_w269_,
		_w422_
	);
	LUT3 #(
		.INIT('hf4)
	) name275 (
		_w230_,
		_w236_,
		_w280_,
		_w423_
	);
	LUT3 #(
		.INIT('h28)
	) name276 (
		\g638_reg/NET0131 ,
		\g650_reg/NET0131 ,
		_w293_,
		_w424_
	);
	LUT4 #(
		.INIT('h6996)
	) name277 (
		\g10_reg/NET0131 ,
		\g18_reg/NET0131 ,
		\g1_reg/NET0131 ,
		\g28_reg/NET0131 ,
		_w425_
	);
	LUT3 #(
		.INIT('h96)
	) name278 (
		\g14_reg/NET0131 ,
		\g2_reg/NET0131 ,
		\g48_reg/NET0131 ,
		_w426_
	);
	LUT2 #(
		.INIT('h9)
	) name279 (
		\g24_reg/NET0131 ,
		\g6_reg/NET0131 ,
		_w427_
	);
	LUT3 #(
		.INIT('h69)
	) name280 (
		_w425_,
		_w426_,
		_w427_,
		_w428_
	);
	LUT4 #(
		.INIT('h4114)
	) name281 (
		\g4110_pad ,
		_w425_,
		_w426_,
		_w427_,
		_w429_
	);
	LUT3 #(
		.INIT('h20)
	) name282 (
		\g1293_pad ,
		\g4110_pad ,
		\g702_pad ,
		_w430_
	);
	LUT4 #(
		.INIT('h0800)
	) name283 (
		\g676_reg/NET0131 ,
		_w243_,
		_w429_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		\g677_reg/NET0131 ,
		_w431_,
		_w432_
	);
	LUT3 #(
		.INIT('h2a)
	) name285 (
		\g465_reg/NET0131 ,
		_w213_,
		_w215_,
		_w433_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name286 (
		\g212_reg/NET0131 ,
		\g248_reg/NET0131 ,
		\g254_reg/NET0131 ,
		\g500_reg/NET0131 ,
		_w434_
	);
	LUT2 #(
		.INIT('h6)
	) name287 (
		\g218_reg/NET0131 ,
		\g504_reg/NET0131 ,
		_w435_
	);
	LUT3 #(
		.INIT('h01)
	) name288 (
		\g236_reg/NET0131 ,
		\g242_reg/NET0131 ,
		\g260_reg/NET0131 ,
		_w436_
	);
	LUT4 #(
		.INIT('h8421)
	) name289 (
		\g224_reg/NET0131 ,
		\g230_reg/NET0131 ,
		\g508_reg/NET0131 ,
		\g512_reg/NET0131 ,
		_w437_
	);
	LUT4 #(
		.INIT('h1000)
	) name290 (
		_w435_,
		_w434_,
		_w436_,
		_w437_,
		_w438_
	);
	LUT3 #(
		.INIT('h15)
	) name291 (
		\g465_reg/NET0131 ,
		_w180_,
		_w182_,
		_w439_
	);
	LUT4 #(
		.INIT('haaa2)
	) name292 (
		\g536_reg/NET0131 ,
		_w438_,
		_w439_,
		_w433_,
		_w440_
	);
	LUT4 #(
		.INIT('hef40)
	) name293 (
		\g677_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w431_,
		_w440_,
		_w441_
	);
	LUT3 #(
		.INIT('h48)
	) name294 (
		\g625_reg/NET0131 ,
		\g639_pad ,
		_w154_,
		_w442_
	);
	LUT4 #(
		.INIT('h48c0)
	) name295 (
		\g606_reg/NET0131 ,
		\g638_reg/NET0131 ,
		\g646_reg/NET0131 ,
		_w292_,
		_w443_
	);
	LUT3 #(
		.INIT('hba)
	) name296 (
		\g492_reg/NET0131 ,
		_w224_,
		_w228_,
		_w444_
	);
	LUT4 #(
		.INIT('hfeaa)
	) name297 (
		\g496_reg/NET0131 ,
		_w184_,
		_w191_,
		_w192_,
		_w445_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		\g677_reg/NET0131 ,
		_w431_,
		_w446_
	);
	LUT4 #(
		.INIT('h60c0)
	) name299 (
		\g619_reg/NET0131 ,
		\g622_reg/NET0131 ,
		\g639_pad ,
		_w153_,
		_w447_
	);
	LUT4 #(
		.INIT('h0800)
	) name300 (
		\g676_reg/NET0131 ,
		_w310_,
		_w429_,
		_w430_,
		_w448_
	);
	LUT3 #(
		.INIT('h48)
	) name301 (
		\g606_reg/NET0131 ,
		\g638_reg/NET0131 ,
		_w292_,
		_w449_
	);
	LUT4 #(
		.INIT('h6996)
	) name302 (
		\g4099_pad ,
		\g4101_pad ,
		\g4103_pad ,
		\g4105_pad ,
		_w450_
	);
	LUT2 #(
		.INIT('h6)
	) name303 (
		\g4100_pad ,
		\g4102_pad ,
		_w451_
	);
	LUT4 #(
		.INIT('h6996)
	) name304 (
		_w425_,
		_w426_,
		_w427_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h9)
	) name305 (
		_w450_,
		_w452_,
		_w453_
	);
	LUT4 #(
		.INIT('hcddc)
	) name306 (
		\g4104_pad ,
		\g669_reg/NET0131 ,
		_w450_,
		_w452_,
		_w454_
	);
	LUT3 #(
		.INIT('h48)
	) name307 (
		\g619_reg/NET0131 ,
		\g639_pad ,
		_w153_,
		_w455_
	);
	LUT3 #(
		.INIT('h28)
	) name308 (
		\g638_reg/NET0131 ,
		\g642_reg/NET0131 ,
		_w291_,
		_w456_
	);
	LUT3 #(
		.INIT('hdc)
	) name309 (
		\g4104_pad ,
		\g672_reg/NET0131 ,
		_w429_,
		_w457_
	);
	LUT3 #(
		.INIT('h10)
	) name310 (
		\g536_reg/NET0131 ,
		\g541_reg/NET0131 ,
		_w438_,
		_w458_
	);
	LUT4 #(
		.INIT('h084c)
	) name311 (
		\g578_reg/NET0131 ,
		\g582_reg/NET0131 ,
		\g681_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w459_
	);
	LUT4 #(
		.INIT('h0213)
	) name312 (
		\g578_reg/NET0131 ,
		\g582_reg/NET0131 ,
		\g683_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w460_
	);
	LUT3 #(
		.INIT('h54)
	) name313 (
		\g586_reg/NET0131 ,
		_w459_,
		_w460_,
		_w461_
	);
	LUT4 #(
		.INIT('h0213)
	) name314 (
		\g578_reg/NET0131 ,
		\g582_reg/NET0131 ,
		\g679_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w462_
	);
	LUT4 #(
		.INIT('h084c)
	) name315 (
		\g578_reg/NET0131 ,
		\g582_reg/NET0131 ,
		\g677_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w463_
	);
	LUT3 #(
		.INIT('ha8)
	) name316 (
		\g586_reg/NET0131 ,
		_w462_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		\g590_reg/NET0131 ,
		\g594_reg/NET0131 ,
		_w465_
	);
	LUT2 #(
		.INIT('h9)
	) name318 (
		\g590_reg/NET0131 ,
		\g594_reg/NET0131 ,
		_w466_
	);
	LUT4 #(
		.INIT('h8000)
	) name319 (
		\g574_reg/NET0131 ,
		\g578_reg/NET0131 ,
		\g582_reg/NET0131 ,
		\g586_reg/NET0131 ,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w465_,
		_w467_,
		_w468_
	);
	LUT4 #(
		.INIT('h001f)
	) name321 (
		_w461_,
		_w464_,
		_w466_,
		_w468_,
		_w469_
	);
	LUT3 #(
		.INIT('h48)
	) name322 (
		\g616_reg/NET0131 ,
		\g639_pad ,
		_w152_,
		_w470_
	);
	LUT4 #(
		.INIT('h7800)
	) name323 (
		\g567_pad ,
		\g598_reg/NET0131 ,
		\g634_reg/NET0131 ,
		\g638_reg/NET0131 ,
		_w471_
	);
	LUT4 #(
		.INIT('h78ff)
	) name324 (
		\g602_reg/NET0131 ,
		\g610_reg/NET0131 ,
		\g613_reg/NET0131 ,
		\g639_pad ,
		_w472_
	);
	LUT3 #(
		.INIT('he4)
	) name325 (
		\g465_reg/NET0131 ,
		\g471_reg/NET0131 ,
		\g478_reg/NET0131 ,
		_w473_
	);
	LUT3 #(
		.INIT('h60)
	) name326 (
		\g567_pad ,
		\g598_reg/NET0131 ,
		\g638_reg/NET0131 ,
		_w474_
	);
	LUT3 #(
		.INIT('h60)
	) name327 (
		\g602_reg/NET0131 ,
		\g610_reg/NET0131 ,
		\g639_pad ,
		_w475_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		\g266_reg/NET0131 ,
		\g4108_pad ,
		_w476_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		\g602_reg/NET0131 ,
		\g639_pad ,
		_w477_
	);
	LUT3 #(
		.INIT('h10)
	) name330 (
		\g677_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w431_,
		_w478_
	);
	LUT4 #(
		.INIT('h70f0)
	) name331 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		\g465_reg/NET0131 ,
		_w213_,
		_w479_
	);
	LUT4 #(
		.INIT('h070f)
	) name332 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g465_reg/NET0131 ,
		_w180_,
		_w480_
	);
	LUT4 #(
		.INIT('h0004)
	) name333 (
		\g536_reg/NET0131 ,
		_w438_,
		_w480_,
		_w479_,
		_w481_
	);
	LUT4 #(
		.INIT('h0045)
	) name334 (
		\g541_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w431_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w478_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		\g102_pad ,
		\g89_pad ,
		_w484_
	);
	LUT2 #(
		.INIT('h7)
	) name337 (
		\g567_pad ,
		\g638_reg/NET0131 ,
		_w485_
	);
	LUT4 #(
		.INIT('h8acf)
	) name338 (
		\g486_reg/NET0131 ,
		\g489_reg/NET0131 ,
		\g492_reg/NET0131 ,
		\g496_reg/NET0131 ,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name339 (
		\g4104_pad ,
		\g675_reg/NET0131 ,
		_w487_
	);
	LUT3 #(
		.INIT('hdf)
	) name340 (
		\g676_reg/NET0131 ,
		_w429_,
		_w487_,
		_w488_
	);
	LUT4 #(
		.INIT('h8800)
	) name341 (
		\g4110_pad ,
		\g676_reg/NET0131 ,
		_w428_,
		_w487_,
		_w489_
	);
	LUT2 #(
		.INIT('hb)
	) name342 (
		_w172_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('hb)
	) name343 (
		\g25_reg/NET0131 ,
		_w489_,
		_w491_
	);
	LUT2 #(
		.INIT('hb)
	) name344 (
		\g29_reg/NET0131 ,
		_w489_,
		_w492_
	);
	LUT2 #(
		.INIT('hb)
	) name345 (
		\g3_reg/NET0131 ,
		_w489_,
		_w493_
	);
	LUT2 #(
		.INIT('hb)
	) name346 (
		\g33_reg/NET0131 ,
		_w489_,
		_w494_
	);
	LUT2 #(
		.INIT('hb)
	) name347 (
		\g7_reg/NET0131 ,
		_w489_,
		_w495_
	);
	LUT2 #(
		.INIT('hb)
	) name348 (
		\g11_reg/NET0131 ,
		_w489_,
		_w496_
	);
	LUT2 #(
		.INIT('hb)
	) name349 (
		\g15_reg/NET0131 ,
		_w489_,
		_w497_
	);
	LUT2 #(
		.INIT('hb)
	) name350 (
		\g19_reg/NET0131 ,
		_w489_,
		_w498_
	);
	assign \_al_n1  = 1'b1;
	assign \g10560/_0_  = _w159_ ;
	assign \g10562/_1_  = _w161_ ;
	assign \g10564/_1_  = _w163_ ;
	assign \g10566/_1_  = _w164_ ;
	assign \g10567/_0_  = _w166_ ;
	assign \g10569/_1_  = _w168_ ;
	assign \g10580/_0_  = _w172_ ;
	assign \g10616/_2_  = _w267_ ;
	assign \g10627/_2_  = _w290_ ;
	assign \g10628/_0_  = _w295_ ;
	assign \g10629/_2_  = _w320_ ;
	assign \g10630/_2_  = _w343_ ;
	assign \g10633/_2_  = _w356_ ;
	assign \g10635/_2_  = _w382_ ;
	assign \g10636/_2_  = _w405_ ;
	assign \g10637/_2_  = _w418_ ;
	assign \g10641/_0_  = _w419_ ;
	assign \g10649/_0_  = _w420_ ;
	assign \g10672/_0_  = _w239_ ;
	assign \g10673/_0_  = _w210_ ;
	assign \g10680/_0_  = _w421_ ;
	assign \g10683/_0_  = _w422_ ;
	assign \g10686/_0_  = _w423_ ;
	assign \g10695/_0_  = _w282_ ;
	assign \g10700/_0_  = _w424_ ;
	assign \g10703/_0_  = _w208_ ;
	assign \g10704/_0_  = _w441_ ;
	assign \g10748/_0_  = _w442_ ;
	assign \g10750/_2_  = _w270_ ;
	assign \g10757/_0_  = _w345_ ;
	assign \g10758/_0_  = _w349_ ;
	assign \g10782/_0_  = _w443_ ;
	assign \g10826/_0_  = _w444_ ;
	assign \g10827/_0_  = _w445_ ;
	assign \g10828/_1_  = _w446_ ;
	assign \g10832/_2_  = _w416_ ;
	assign \g10834/_2_  = _w413_ ;
	assign \g10836/_0_  = _w447_ ;
	assign \g10837/_1__syn_2  = _w448_ ;
	assign \g10868/_0_  = _w449_ ;
	assign \g10904/_0_  = _w454_ ;
	assign \g10913/_0_  = _w325_ ;
	assign \g10915/_0_  = _w330_ ;
	assign \g10922/_0_  = _w455_ ;
	assign \g10938/_0_  = _w399_ ;
	assign \g10939/_0_  = _w372_ ;
	assign \g10940/_0_  = _w385_ ;
	assign \g10941/_0_  = _w360_ ;
	assign \g10942/_0_  = _w305_ ;
	assign \g10944/_2_  = _w300_ ;
	assign \g10977/_0_  = _w456_ ;
	assign \g10980/_0_  = _w457_ ;
	assign \g11020/_0_  = _w453_ ;
	assign \g11028/_0_  = _w458_ ;
	assign \g11051/_0_  = _w469_ ;
	assign \g11057/_0_  = _w470_ ;
	assign \g11109/_0_  = _w471_ ;
	assign \g11113/_2_  = _w438_ ;
	assign \g11156/_0_  = _w472_ ;
	assign \g11172/_3_  = _w473_ ;
	assign \g11193/_0_  = _w474_ ;
	assign \g11219/_0_  = _w475_ ;
	assign \g11355/_0_  = _w136_ ;
	assign \g11384/_0_  = _w134_ ;
	assign \g11442/_0_  = _w476_ ;
	assign \g11448/_0_  = _w477_ ;
	assign \g11558/_0_  = _w32_ ;
	assign \g11559/_0_  = _w62_ ;
	assign \g11824/_1_  = _w272_ ;
	assign \g11853/_0_  = _w483_ ;
	assign \g11854/_0_  = _w432_ ;
	assign \g11977/_0_  = _w237_ ;
	assign \g11981/_0_  = _w281_ ;
	assign \g2584_pad  = _w484_ ;
	assign \g4121_pad  = _w485_ ;
	assign \g4809_pad  = _w486_ ;
	assign \g5692_pad  = 1'b0;
	assign \g6282_pad  = _w488_ ;
	assign \g6284_pad  = _w490_ ;
	assign \g6360_pad  = _w491_ ;
	assign \g6362_pad  = _w492_ ;
	assign \g6364_pad  = _w493_ ;
	assign \g6366_pad  = _w494_ ;
	assign \g6368_pad  = _w495_ ;
	assign \g6370_pad  = _w496_ ;
	assign \g6372_pad  = _w497_ ;
	assign \g6374_pad  = _w498_ ;
endmodule;